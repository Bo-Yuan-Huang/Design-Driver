
module oc8051_gm_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pc, property_invalid_acc, property_invalid_iram);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire _25005_;
  wire _25006_;
  wire _25007_;
  wire _25008_;
  wire _25009_;
  wire _25010_;
  wire _25011_;
  wire _25012_;
  wire _25013_;
  wire _25014_;
  wire _25015_;
  wire _25016_;
  wire _25017_;
  wire _25018_;
  wire _25019_;
  wire _25020_;
  wire _25021_;
  wire _25022_;
  wire _25023_;
  wire _25024_;
  wire _25025_;
  wire _25026_;
  wire _25027_;
  wire _25028_;
  wire _25029_;
  wire _25030_;
  wire _25031_;
  wire _25032_;
  wire _25033_;
  wire _25034_;
  wire _25035_;
  wire _25036_;
  wire _25037_;
  wire _25038_;
  wire _25039_;
  wire _25040_;
  wire _25041_;
  wire _25042_;
  wire _25043_;
  wire _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire _25454_;
  wire _25455_;
  wire _25456_;
  wire _25457_;
  wire _25458_;
  wire _25459_;
  wire _25460_;
  wire _25461_;
  wire _25462_;
  wire _25463_;
  wire _25464_;
  wire _25465_;
  wire _25466_;
  wire _25467_;
  wire _25468_;
  wire _25469_;
  wire _25470_;
  wire _25471_;
  wire _25472_;
  wire _25473_;
  wire _25474_;
  wire _25475_;
  wire _25476_;
  wire _25477_;
  wire _25478_;
  wire _25479_;
  wire _25480_;
  wire _25481_;
  wire _25482_;
  wire _25483_;
  wire _25484_;
  wire _25485_;
  wire _25486_;
  wire _25487_;
  wire _25488_;
  wire _25489_;
  wire _25490_;
  wire _25491_;
  wire _25492_;
  wire _25493_;
  wire _25494_;
  wire _25495_;
  wire _25496_;
  wire _25497_;
  wire _25498_;
  wire _25499_;
  wire _25500_;
  wire _25501_;
  wire _25502_;
  wire _25503_;
  wire _25504_;
  wire _25505_;
  wire _25506_;
  wire _25507_;
  wire _25508_;
  wire _25509_;
  wire _25510_;
  wire _25511_;
  wire _25512_;
  wire _25513_;
  wire _25514_;
  wire _25515_;
  wire _25516_;
  wire _25517_;
  wire _25518_;
  wire _25519_;
  wire _25520_;
  wire _25521_;
  wire _25522_;
  wire _25523_;
  wire _25524_;
  wire _25525_;
  wire _25526_;
  wire _25527_;
  wire _25528_;
  wire _25529_;
  wire _25530_;
  wire _25531_;
  wire _25532_;
  wire _25533_;
  wire _25534_;
  wire _25535_;
  wire _25536_;
  wire _25537_;
  wire _25538_;
  wire _25539_;
  wire _25540_;
  wire _25541_;
  wire _25542_;
  wire _25543_;
  wire _25544_;
  wire _25545_;
  wire _25546_;
  wire _25547_;
  wire _25548_;
  wire _25549_;
  wire _25550_;
  wire _25551_;
  wire _25552_;
  wire _25553_;
  wire _25554_;
  wire _25555_;
  wire _25556_;
  wire _25557_;
  wire _25558_;
  wire _25559_;
  wire _25560_;
  wire _25561_;
  wire _25562_;
  wire _25563_;
  wire _25564_;
  wire _25565_;
  wire _25566_;
  wire _25567_;
  wire _25568_;
  wire _25569_;
  wire _25570_;
  wire _25571_;
  wire _25572_;
  wire _25573_;
  wire _25574_;
  wire _25575_;
  wire _25576_;
  wire _25577_;
  wire _25578_;
  wire _25579_;
  wire _25580_;
  wire _25581_;
  wire _25582_;
  wire _25583_;
  wire _25584_;
  wire _25585_;
  wire _25586_;
  wire _25587_;
  wire _25588_;
  wire _25589_;
  wire _25590_;
  wire _25591_;
  wire _25592_;
  wire _25593_;
  wire _25594_;
  wire _25595_;
  wire _25596_;
  wire _25597_;
  wire _25598_;
  wire _25599_;
  wire _25600_;
  wire _25601_;
  wire _25602_;
  wire _25603_;
  wire _25604_;
  wire _25605_;
  wire _25606_;
  wire _25607_;
  wire _25608_;
  wire _25609_;
  wire _25610_;
  wire _25611_;
  wire _25612_;
  wire _25613_;
  wire _25614_;
  wire _25615_;
  wire _25616_;
  wire _25617_;
  wire _25618_;
  wire _25619_;
  wire _25620_;
  wire _25621_;
  wire _25622_;
  wire _25623_;
  wire _25624_;
  wire _25625_;
  wire _25626_;
  wire _25627_;
  wire _25628_;
  wire _25629_;
  wire _25630_;
  wire _25631_;
  wire _25632_;
  wire _25633_;
  wire _25634_;
  wire _25635_;
  wire _25636_;
  wire _25637_;
  wire _25638_;
  wire _25639_;
  wire _25640_;
  wire _25641_;
  wire _25642_;
  wire _25643_;
  wire _25644_;
  wire _25645_;
  wire _25646_;
  wire _25647_;
  wire _25648_;
  wire _25649_;
  wire _25650_;
  wire _25651_;
  wire _25652_;
  wire _25653_;
  wire _25654_;
  wire _25655_;
  wire _25656_;
  wire _25657_;
  wire _25658_;
  wire _25659_;
  wire _25660_;
  wire _25661_;
  wire _25662_;
  wire _25663_;
  wire _25664_;
  wire _25665_;
  wire _25666_;
  wire _25667_;
  wire _25668_;
  wire _25669_;
  wire _25670_;
  wire _25671_;
  wire _25672_;
  wire _25673_;
  wire _25674_;
  wire _25675_;
  wire _25676_;
  wire _25677_;
  wire _25678_;
  wire _25679_;
  wire _25680_;
  wire _25681_;
  wire _25682_;
  wire _25683_;
  wire _25684_;
  wire _25685_;
  wire _25686_;
  wire _25687_;
  wire _25688_;
  wire _25689_;
  wire _25690_;
  wire _25691_;
  wire _25692_;
  wire _25693_;
  wire _25694_;
  wire _25695_;
  wire _25696_;
  wire _25697_;
  wire _25698_;
  wire _25699_;
  wire _25700_;
  wire _25701_;
  wire _25702_;
  wire _25703_;
  wire _25704_;
  wire _25705_;
  wire _25706_;
  wire _25707_;
  wire _25708_;
  wire _25709_;
  wire _25710_;
  wire _25711_;
  wire _25712_;
  wire _25713_;
  wire _25714_;
  wire _25715_;
  wire _25716_;
  wire _25717_;
  wire _25718_;
  wire _25719_;
  wire _25720_;
  wire _25721_;
  wire _25722_;
  wire _25723_;
  wire _25724_;
  wire _25725_;
  wire _25726_;
  wire _25727_;
  wire _25728_;
  wire _25729_;
  wire _25730_;
  wire _25731_;
  wire _25732_;
  wire _25733_;
  wire _25734_;
  wire _25735_;
  wire _25736_;
  wire _25737_;
  wire _25738_;
  wire _25739_;
  wire _25740_;
  wire _25741_;
  wire _25742_;
  wire _25743_;
  wire _25744_;
  wire _25745_;
  wire _25746_;
  wire _25747_;
  wire _25748_;
  wire _25749_;
  wire _25750_;
  wire _25751_;
  wire _25752_;
  wire _25753_;
  wire _25754_;
  wire _25755_;
  wire _25756_;
  wire _25757_;
  wire _25758_;
  wire _25759_;
  wire _25760_;
  wire _25761_;
  wire _25762_;
  wire _25763_;
  wire _25764_;
  wire _25765_;
  wire _25766_;
  wire _25767_;
  wire _25768_;
  wire _25769_;
  wire _25770_;
  wire _25771_;
  wire _25772_;
  wire _25773_;
  wire _25774_;
  wire _25775_;
  wire _25776_;
  wire _25777_;
  wire _25778_;
  wire _25779_;
  wire _25780_;
  wire _25781_;
  wire _25782_;
  wire _25783_;
  wire _25784_;
  wire _25785_;
  wire _25786_;
  wire _25787_;
  wire _25788_;
  wire _25789_;
  wire _25790_;
  wire _25791_;
  wire _25792_;
  wire _25793_;
  wire _25794_;
  wire _25795_;
  wire _25796_;
  wire _25797_;
  wire _25798_;
  wire _25799_;
  wire _25800_;
  wire _25801_;
  wire _25802_;
  wire _25803_;
  wire _25804_;
  wire _25805_;
  wire _25806_;
  wire _25807_;
  wire _25808_;
  wire _25809_;
  wire _25810_;
  wire _25811_;
  wire _25812_;
  wire _25813_;
  wire _25814_;
  wire _25815_;
  wire _25816_;
  wire _25817_;
  wire _25818_;
  wire _25819_;
  wire _25820_;
  wire _25821_;
  wire _25822_;
  wire _25823_;
  wire _25824_;
  wire _25825_;
  wire _25826_;
  wire _25827_;
  wire _25828_;
  wire _25829_;
  wire _25830_;
  wire _25831_;
  wire _25832_;
  wire _25833_;
  wire _25834_;
  wire _25835_;
  wire _25836_;
  wire _25837_;
  wire _25838_;
  wire _25839_;
  wire _25840_;
  wire _25841_;
  wire _25842_;
  wire _25843_;
  wire _25844_;
  wire _25845_;
  wire _25846_;
  wire _25847_;
  wire _25848_;
  wire _25849_;
  wire _25850_;
  wire _25851_;
  wire _25852_;
  wire _25853_;
  wire _25854_;
  wire _25855_;
  wire _25856_;
  wire _25857_;
  wire _25858_;
  wire _25859_;
  wire _25860_;
  wire _25861_;
  wire _25862_;
  wire _25863_;
  wire _25864_;
  wire _25865_;
  wire _25866_;
  wire _25867_;
  wire _25868_;
  wire _25869_;
  wire _25870_;
  wire _25871_;
  wire _25872_;
  wire _25873_;
  wire _25874_;
  wire _25875_;
  wire _25876_;
  wire _25877_;
  wire _25878_;
  wire _25879_;
  wire _25880_;
  wire _25881_;
  wire _25882_;
  wire _25883_;
  wire _25884_;
  wire _25885_;
  wire _25886_;
  wire _25887_;
  wire _25888_;
  wire _25889_;
  wire _25890_;
  wire _25891_;
  wire _25892_;
  wire _25893_;
  wire _25894_;
  wire _25895_;
  wire _25896_;
  wire _25897_;
  wire _25898_;
  wire _25899_;
  wire _25900_;
  wire _25901_;
  wire _25902_;
  wire _25903_;
  wire _25904_;
  wire _25905_;
  wire _25906_;
  wire _25907_;
  wire _25908_;
  wire _25909_;
  wire _25910_;
  wire _25911_;
  wire _25912_;
  wire _25913_;
  wire _25914_;
  wire _25915_;
  wire _25916_;
  wire _25917_;
  wire _25918_;
  wire _25919_;
  wire _25920_;
  wire _25921_;
  wire _25922_;
  wire _25923_;
  wire _25924_;
  wire _25925_;
  wire _25926_;
  wire _25927_;
  wire _25928_;
  wire _25929_;
  wire _25930_;
  wire _25931_;
  wire _25932_;
  wire _25933_;
  wire _25934_;
  wire _25935_;
  wire _25936_;
  wire _25937_;
  wire _25938_;
  wire _25939_;
  wire _25940_;
  wire _25941_;
  wire _25942_;
  wire _25943_;
  wire _25944_;
  wire _25945_;
  wire _25946_;
  wire _25947_;
  wire _25948_;
  wire _25949_;
  wire _25950_;
  wire _25951_;
  wire _25952_;
  wire _25953_;
  wire _25954_;
  wire _25955_;
  wire _25956_;
  wire _25957_;
  wire _25958_;
  wire _25959_;
  wire _25960_;
  wire _25961_;
  wire _25962_;
  wire _25963_;
  wire _25964_;
  wire _25965_;
  wire _25966_;
  wire _25967_;
  wire _25968_;
  wire _25969_;
  wire _25970_;
  wire _25971_;
  wire _25972_;
  wire _25973_;
  wire _25974_;
  wire _25975_;
  wire _25976_;
  wire _25977_;
  wire _25978_;
  wire _25979_;
  wire _25980_;
  wire _25981_;
  wire _25982_;
  wire _25983_;
  wire _25984_;
  wire _25985_;
  wire _25986_;
  wire _25987_;
  wire _25988_;
  wire _25989_;
  wire _25990_;
  wire _25991_;
  wire _25992_;
  wire _25993_;
  wire _25994_;
  wire _25995_;
  wire _25996_;
  wire _25997_;
  wire _25998_;
  wire _25999_;
  wire _26000_;
  wire _26001_;
  wire _26002_;
  wire _26003_;
  wire _26004_;
  wire _26005_;
  wire _26006_;
  wire _26007_;
  wire _26008_;
  wire _26009_;
  wire _26010_;
  wire _26011_;
  wire _26012_;
  wire _26013_;
  wire _26014_;
  wire _26015_;
  wire _26016_;
  wire _26017_;
  wire _26018_;
  wire _26019_;
  wire _26020_;
  wire _26021_;
  wire _26022_;
  wire _26023_;
  wire _26024_;
  wire _26025_;
  wire _26026_;
  wire _26027_;
  wire _26028_;
  wire _26029_;
  wire _26030_;
  wire _26031_;
  wire _26032_;
  wire _26033_;
  wire _26034_;
  wire _26035_;
  wire _26036_;
  wire _26037_;
  wire _26038_;
  wire _26039_;
  wire _26040_;
  wire _26041_;
  wire _26042_;
  wire _26043_;
  wire _26044_;
  wire _26045_;
  wire _26046_;
  wire _26047_;
  wire _26048_;
  wire _26049_;
  wire _26050_;
  wire _26051_;
  wire _26052_;
  wire _26053_;
  wire _26054_;
  wire _26055_;
  wire _26056_;
  wire _26057_;
  wire _26058_;
  wire _26059_;
  wire _26060_;
  wire _26061_;
  wire _26062_;
  wire _26063_;
  wire _26064_;
  wire _26065_;
  wire _26066_;
  wire _26067_;
  wire _26068_;
  wire _26069_;
  wire _26070_;
  wire _26071_;
  wire _26072_;
  wire _26073_;
  wire _26074_;
  wire _26075_;
  wire _26076_;
  wire _26077_;
  wire _26078_;
  wire _26079_;
  wire _26080_;
  wire _26081_;
  wire _26082_;
  wire _26083_;
  wire _26084_;
  wire _26085_;
  wire _26086_;
  wire _26087_;
  wire _26088_;
  wire _26089_;
  wire _26090_;
  wire _26091_;
  wire _26092_;
  wire _26093_;
  wire _26094_;
  wire _26095_;
  wire _26096_;
  wire _26097_;
  wire _26098_;
  wire _26099_;
  wire _26100_;
  wire _26101_;
  wire _26102_;
  wire _26103_;
  wire _26104_;
  wire _26105_;
  wire _26106_;
  wire _26107_;
  wire _26108_;
  wire _26109_;
  wire _26110_;
  wire _26111_;
  wire _26112_;
  wire _26113_;
  wire _26114_;
  wire _26115_;
  wire _26116_;
  wire _26117_;
  wire _26118_;
  wire _26119_;
  wire _26120_;
  wire _26121_;
  wire _26122_;
  wire _26123_;
  wire _26124_;
  wire _26125_;
  wire _26126_;
  wire _26127_;
  wire _26128_;
  wire _26129_;
  wire _26130_;
  wire _26131_;
  wire _26132_;
  wire _26133_;
  wire _26134_;
  wire _26135_;
  wire _26136_;
  wire _26137_;
  wire _26138_;
  wire _26139_;
  wire _26140_;
  wire _26141_;
  wire _26142_;
  wire _26143_;
  wire _26144_;
  wire _26145_;
  wire _26146_;
  wire _26147_;
  wire _26148_;
  wire _26149_;
  wire _26150_;
  wire _26151_;
  wire _26152_;
  wire _26153_;
  wire _26154_;
  wire _26155_;
  wire _26156_;
  wire _26157_;
  wire _26158_;
  wire _26159_;
  wire _26160_;
  wire _26161_;
  wire _26162_;
  wire _26163_;
  wire _26164_;
  wire _26165_;
  wire _26166_;
  wire _26167_;
  wire _26168_;
  wire _26169_;
  wire _26170_;
  wire _26171_;
  wire _26172_;
  wire _26173_;
  wire _26174_;
  wire _26175_;
  wire _26176_;
  wire _26177_;
  wire _26178_;
  wire _26179_;
  wire _26180_;
  wire _26181_;
  wire _26182_;
  wire _26183_;
  wire _26184_;
  wire _26185_;
  wire _26186_;
  wire _26187_;
  wire _26188_;
  wire _26189_;
  wire _26190_;
  wire _26191_;
  wire _26192_;
  wire _26193_;
  wire _26194_;
  wire _26195_;
  wire _26196_;
  wire _26197_;
  wire _26198_;
  wire _26199_;
  wire _26200_;
  wire _26201_;
  wire _26202_;
  wire _26203_;
  wire _26204_;
  wire _26205_;
  wire _26206_;
  wire _26207_;
  wire _26208_;
  wire _26209_;
  wire _26210_;
  wire _26211_;
  wire _26212_;
  wire _26213_;
  wire _26214_;
  wire _26215_;
  wire _26216_;
  wire _26217_;
  wire _26218_;
  wire _26219_;
  wire _26220_;
  wire _26221_;
  wire _26222_;
  wire _26223_;
  wire _26224_;
  wire _26225_;
  wire _26226_;
  wire _26227_;
  wire _26228_;
  wire _26229_;
  wire _26230_;
  wire _26231_;
  wire _26232_;
  wire _26233_;
  wire _26234_;
  wire _26235_;
  wire _26236_;
  wire _26237_;
  wire _26238_;
  wire _26239_;
  wire _26240_;
  wire _26241_;
  wire _26242_;
  wire _26243_;
  wire _26244_;
  wire _26245_;
  wire _26246_;
  wire _26247_;
  wire _26248_;
  wire _26249_;
  wire _26250_;
  wire _26251_;
  wire _26252_;
  wire _26253_;
  wire _26254_;
  wire _26255_;
  wire _26256_;
  wire _26257_;
  wire _26258_;
  wire _26259_;
  wire _26260_;
  wire _26261_;
  wire _26262_;
  wire _26263_;
  wire _26264_;
  wire _26265_;
  wire _26266_;
  wire _26267_;
  wire _26268_;
  wire _26269_;
  wire _26270_;
  wire _26271_;
  wire _26272_;
  wire _26273_;
  wire _26274_;
  wire _26275_;
  wire _26276_;
  wire _26277_;
  wire _26278_;
  wire _26279_;
  wire _26280_;
  wire _26281_;
  wire _26282_;
  wire _26283_;
  wire _26284_;
  wire _26285_;
  wire _26286_;
  wire _26287_;
  wire _26288_;
  wire _26289_;
  wire _26290_;
  wire _26291_;
  wire _26292_;
  wire _26293_;
  wire _26294_;
  wire _26295_;
  wire _26296_;
  wire _26297_;
  wire _26298_;
  wire _26299_;
  wire _26300_;
  wire _26301_;
  wire _26302_;
  wire _26303_;
  wire _26304_;
  wire _26305_;
  wire _26306_;
  wire _26307_;
  wire _26308_;
  wire _26309_;
  wire _26310_;
  wire _26311_;
  wire _26312_;
  wire _26313_;
  wire _26314_;
  wire _26315_;
  wire _26316_;
  wire _26317_;
  wire _26318_;
  wire _26319_;
  wire _26320_;
  wire _26321_;
  wire _26322_;
  wire _26323_;
  wire _26324_;
  wire _26325_;
  wire _26326_;
  wire _26327_;
  wire _26328_;
  wire _26329_;
  wire _26330_;
  wire _26331_;
  wire _26332_;
  wire _26333_;
  wire _26334_;
  wire _26335_;
  wire _26336_;
  wire _26337_;
  wire _26338_;
  wire _26339_;
  wire _26340_;
  wire _26341_;
  wire _26342_;
  wire _26343_;
  wire _26344_;
  wire _26345_;
  wire _26346_;
  wire _26347_;
  wire _26348_;
  wire _26349_;
  wire _26350_;
  wire _26351_;
  wire _26352_;
  wire _26353_;
  wire _26354_;
  wire _26355_;
  wire _26356_;
  wire _26357_;
  wire _26358_;
  wire _26359_;
  wire _26360_;
  wire _26361_;
  wire _26362_;
  wire _26363_;
  wire _26364_;
  wire _26365_;
  wire _26366_;
  wire _26367_;
  wire _26368_;
  wire _26369_;
  wire _26370_;
  wire _26371_;
  wire _26372_;
  wire _26373_;
  wire _26374_;
  wire _26375_;
  wire _26376_;
  wire _26377_;
  wire _26378_;
  wire _26379_;
  wire _26380_;
  wire _26381_;
  wire _26382_;
  wire _26383_;
  wire _26384_;
  wire _26385_;
  wire _26386_;
  wire _26387_;
  wire _26388_;
  wire _26389_;
  wire _26390_;
  wire _26391_;
  wire _26392_;
  wire _26393_;
  wire _26394_;
  wire _26395_;
  wire _26396_;
  wire _26397_;
  wire _26398_;
  wire _26399_;
  wire _26400_;
  wire _26401_;
  wire _26402_;
  wire _26403_;
  wire _26404_;
  wire _26405_;
  wire _26406_;
  wire _26407_;
  wire _26408_;
  wire _26409_;
  wire _26410_;
  wire _26411_;
  wire _26412_;
  wire _26413_;
  wire _26414_;
  wire _26415_;
  wire _26416_;
  wire _26417_;
  wire _26418_;
  wire _26419_;
  wire _26420_;
  wire _26421_;
  wire _26422_;
  wire _26423_;
  wire _26424_;
  wire _26425_;
  wire _26426_;
  wire _26427_;
  wire _26428_;
  wire _26429_;
  wire _26430_;
  wire _26431_;
  wire _26432_;
  wire _26433_;
  wire _26434_;
  wire _26435_;
  wire _26436_;
  wire _26437_;
  wire _26438_;
  wire _26439_;
  wire _26440_;
  wire _26441_;
  wire _26442_;
  wire _26443_;
  wire _26444_;
  wire _26445_;
  wire _26446_;
  wire _26447_;
  wire _26448_;
  wire _26449_;
  wire _26450_;
  wire _26451_;
  wire _26452_;
  wire _26453_;
  wire _26454_;
  wire _26455_;
  wire _26456_;
  wire _26457_;
  wire _26458_;
  wire _26459_;
  wire _26460_;
  wire _26461_;
  wire _26462_;
  wire _26463_;
  wire _26464_;
  wire _26465_;
  wire _26466_;
  wire _26467_;
  wire _26468_;
  wire _26469_;
  wire _26470_;
  wire _26471_;
  wire _26472_;
  wire _26473_;
  wire _26474_;
  wire _26475_;
  wire _26476_;
  wire _26477_;
  wire _26478_;
  wire _26479_;
  wire _26480_;
  wire _26481_;
  wire _26482_;
  wire _26483_;
  wire _26484_;
  wire _26485_;
  wire _26486_;
  wire _26487_;
  wire _26488_;
  wire _26489_;
  wire _26490_;
  wire _26491_;
  wire _26492_;
  wire _26493_;
  wire _26494_;
  wire _26495_;
  wire _26496_;
  wire _26497_;
  wire _26498_;
  wire _26499_;
  wire _26500_;
  wire _26501_;
  wire _26502_;
  wire _26503_;
  wire _26504_;
  wire _26505_;
  wire _26506_;
  wire _26507_;
  wire _26508_;
  wire _26509_;
  wire _26510_;
  wire _26511_;
  wire _26512_;
  wire _26513_;
  wire _26514_;
  wire _26515_;
  wire _26516_;
  wire _26517_;
  wire _26518_;
  wire _26519_;
  wire _26520_;
  wire _26521_;
  wire _26522_;
  wire _26523_;
  wire _26524_;
  wire _26525_;
  wire _26526_;
  wire _26527_;
  wire _26528_;
  wire _26529_;
  wire _26530_;
  wire _26531_;
  wire _26532_;
  wire _26533_;
  wire _26534_;
  wire _26535_;
  wire _26536_;
  wire _26537_;
  wire _26538_;
  wire _26539_;
  wire _26540_;
  wire _26541_;
  wire _26542_;
  wire _26543_;
  wire _26544_;
  wire _26545_;
  wire _26546_;
  wire _26547_;
  wire _26548_;
  wire _26549_;
  wire _26550_;
  wire _26551_;
  wire _26552_;
  wire _26553_;
  wire _26554_;
  wire _26555_;
  wire _26556_;
  wire _26557_;
  wire _26558_;
  wire _26559_;
  wire _26560_;
  wire _26561_;
  wire _26562_;
  wire _26563_;
  wire _26564_;
  wire _26565_;
  wire _26566_;
  wire _26567_;
  wire _26568_;
  wire _26569_;
  wire _26570_;
  wire _26571_;
  wire _26572_;
  wire _26573_;
  wire _26574_;
  wire _26575_;
  wire _26576_;
  wire _26577_;
  wire _26578_;
  wire _26579_;
  wire _26580_;
  wire _26581_;
  wire _26582_;
  wire _26583_;
  wire _26584_;
  wire _26585_;
  wire _26586_;
  wire _26587_;
  wire _26588_;
  wire _26589_;
  wire _26590_;
  wire _26591_;
  wire _26592_;
  wire _26593_;
  wire _26594_;
  wire _26595_;
  wire _26596_;
  wire _26597_;
  wire _26598_;
  wire _26599_;
  wire _26600_;
  wire _26601_;
  wire _26602_;
  wire _26603_;
  wire _26604_;
  wire _26605_;
  wire _26606_;
  wire _26607_;
  wire _26608_;
  wire _26609_;
  wire _26610_;
  wire _26611_;
  wire _26612_;
  wire _26613_;
  wire _26614_;
  wire _26615_;
  wire _26616_;
  wire _26617_;
  wire _26618_;
  wire _26619_;
  wire _26620_;
  wire _26621_;
  wire _26622_;
  wire _26623_;
  wire _26624_;
  wire _26625_;
  wire _26626_;
  wire _26627_;
  wire _26628_;
  wire _26629_;
  wire _26630_;
  wire _26631_;
  wire _26632_;
  wire _26633_;
  wire _26634_;
  wire _26635_;
  wire _26636_;
  wire _26637_;
  wire _26638_;
  wire _26639_;
  wire _26640_;
  wire _26641_;
  wire _26642_;
  wire _26643_;
  wire _26644_;
  wire _26645_;
  wire _26646_;
  wire _26647_;
  wire _26648_;
  wire _26649_;
  wire _26650_;
  wire _26651_;
  wire _26652_;
  wire _26653_;
  wire _26654_;
  wire _26655_;
  wire _26656_;
  wire _26657_;
  wire _26658_;
  wire _26659_;
  wire _26660_;
  wire _26661_;
  wire _26662_;
  wire _26663_;
  wire _26664_;
  wire _26665_;
  wire _26666_;
  wire _26667_;
  wire _26668_;
  wire _26669_;
  wire _26670_;
  wire _26671_;
  wire _26672_;
  wire _26673_;
  wire _26674_;
  wire _26675_;
  wire _26676_;
  wire _26677_;
  wire _26678_;
  wire _26679_;
  wire _26680_;
  wire _26681_;
  wire _26682_;
  wire _26683_;
  wire _26684_;
  wire _26685_;
  wire _26686_;
  wire _26687_;
  wire _26688_;
  wire _26689_;
  wire _26690_;
  wire _26691_;
  wire _26692_;
  wire _26693_;
  wire _26694_;
  wire _26695_;
  wire _26696_;
  wire _26697_;
  wire _26698_;
  wire _26699_;
  wire _26700_;
  wire _26701_;
  wire _26702_;
  wire _26703_;
  wire _26704_;
  wire _26705_;
  wire _26706_;
  wire _26707_;
  wire _26708_;
  wire _26709_;
  wire _26710_;
  wire _26711_;
  wire _26712_;
  wire _26713_;
  wire _26714_;
  wire _26715_;
  wire _26716_;
  wire _26717_;
  wire _26718_;
  wire _26719_;
  wire _26720_;
  wire _26721_;
  wire _26722_;
  wire _26723_;
  wire _26724_;
  wire _26725_;
  wire _26726_;
  wire _26727_;
  wire _26728_;
  wire _26729_;
  wire _26730_;
  wire _26731_;
  wire _26732_;
  wire _26733_;
  wire _26734_;
  wire _26735_;
  wire _26736_;
  wire _26737_;
  wire _26738_;
  wire _26739_;
  wire _26740_;
  wire _26741_;
  wire _26742_;
  wire _26743_;
  wire _26744_;
  wire _26745_;
  wire _26746_;
  wire _26747_;
  wire _26748_;
  wire _26749_;
  wire _26750_;
  wire _26751_;
  wire _26752_;
  wire _26753_;
  wire _26754_;
  wire _26755_;
  wire _26756_;
  wire _26757_;
  wire _26758_;
  wire _26759_;
  wire _26760_;
  wire _26761_;
  wire _26762_;
  wire _26763_;
  wire _26764_;
  wire _26765_;
  wire _26766_;
  wire _26767_;
  wire _26768_;
  wire _26769_;
  wire _26770_;
  wire _26771_;
  wire _26772_;
  wire _26773_;
  wire _26774_;
  wire _26775_;
  wire _26776_;
  wire _26777_;
  wire _26778_;
  wire _26779_;
  wire _26780_;
  wire _26781_;
  wire _26782_;
  wire _26783_;
  wire _26784_;
  wire _26785_;
  wire _26786_;
  wire _26787_;
  wire _26788_;
  wire _26789_;
  wire _26790_;
  wire _26791_;
  wire _26792_;
  wire _26793_;
  wire _26794_;
  wire _26795_;
  wire _26796_;
  wire _26797_;
  wire _26798_;
  wire _26799_;
  wire _26800_;
  wire _26801_;
  wire _26802_;
  wire _26803_;
  wire _26804_;
  wire _26805_;
  wire _26806_;
  wire _26807_;
  wire _26808_;
  wire _26809_;
  wire _26810_;
  wire _26811_;
  wire _26812_;
  wire _26813_;
  wire _26814_;
  wire _26815_;
  wire _26816_;
  wire _26817_;
  wire _26818_;
  wire _26819_;
  wire _26820_;
  wire _26821_;
  wire _26822_;
  wire _26823_;
  wire _26824_;
  wire _26825_;
  wire _26826_;
  wire _26827_;
  wire _26828_;
  wire _26829_;
  wire _26830_;
  wire _26831_;
  wire _26832_;
  wire _26833_;
  wire _26834_;
  wire _26835_;
  wire _26836_;
  wire _26837_;
  wire _26838_;
  wire _26839_;
  wire _26840_;
  wire _26841_;
  wire _26842_;
  wire _26843_;
  wire _26844_;
  wire _26845_;
  wire _26846_;
  wire _26847_;
  wire _26848_;
  wire _26849_;
  wire _26850_;
  wire _26851_;
  wire _26852_;
  wire _26853_;
  wire _26854_;
  wire _26855_;
  wire _26856_;
  wire _26857_;
  wire _26858_;
  wire _26859_;
  wire _26860_;
  wire _26861_;
  wire _26862_;
  wire _26863_;
  wire _26864_;
  wire _26865_;
  wire _26866_;
  wire _26867_;
  wire _26868_;
  wire _26869_;
  wire _26870_;
  wire _26871_;
  wire _26872_;
  wire _26873_;
  wire _26874_;
  wire _26875_;
  wire _26876_;
  wire _26877_;
  wire _26878_;
  wire _26879_;
  wire _26880_;
  wire _26881_;
  wire _26882_;
  wire _26883_;
  wire _26884_;
  wire _26885_;
  wire _26886_;
  wire _26887_;
  wire _26888_;
  wire _26889_;
  wire _26890_;
  wire _26891_;
  wire _26892_;
  wire _26893_;
  wire _26894_;
  wire _26895_;
  wire _26896_;
  wire _26897_;
  wire _26898_;
  wire _26899_;
  wire _26900_;
  wire _26901_;
  wire _26902_;
  wire _26903_;
  wire _26904_;
  wire _26905_;
  wire _26906_;
  wire _26907_;
  wire _26908_;
  wire _26909_;
  wire _26910_;
  wire _26911_;
  wire _26912_;
  wire _26913_;
  wire _26914_;
  wire _26915_;
  wire _26916_;
  wire _26917_;
  wire _26918_;
  wire _26919_;
  wire _26920_;
  wire _26921_;
  wire _26922_;
  wire _26923_;
  wire _26924_;
  wire _26925_;
  wire _26926_;
  wire _26927_;
  wire _26928_;
  wire _26929_;
  wire _26930_;
  wire _26931_;
  wire _26932_;
  wire _26933_;
  wire _26934_;
  wire _26935_;
  wire _26936_;
  wire _26937_;
  wire _26938_;
  wire _26939_;
  wire _26940_;
  wire _26941_;
  wire _26942_;
  wire _26943_;
  wire _26944_;
  wire _26945_;
  wire _26946_;
  wire _26947_;
  wire _26948_;
  wire _26949_;
  wire _26950_;
  wire _26951_;
  wire _26952_;
  wire _26953_;
  wire _26954_;
  wire _26955_;
  wire _26956_;
  wire _26957_;
  wire _26958_;
  wire _26959_;
  wire _26960_;
  wire _26961_;
  wire _26962_;
  wire _26963_;
  wire _26964_;
  wire _26965_;
  wire _26966_;
  wire _26967_;
  wire _26968_;
  wire _26969_;
  wire _26970_;
  wire _26971_;
  wire _26972_;
  wire _26973_;
  wire _26974_;
  wire _26975_;
  wire _26976_;
  wire _26977_;
  wire _26978_;
  wire _26979_;
  wire _26980_;
  wire _26981_;
  wire _26982_;
  wire _26983_;
  wire _26984_;
  wire _26985_;
  wire _26986_;
  wire _26987_;
  wire _26988_;
  wire _26989_;
  wire _26990_;
  wire _26991_;
  wire _26992_;
  wire _26993_;
  wire _26994_;
  wire _26995_;
  wire _26996_;
  wire _26997_;
  wire _26998_;
  wire _26999_;
  wire _27000_;
  wire _27001_;
  wire _27002_;
  wire _27003_;
  wire _27004_;
  wire _27005_;
  wire _27006_;
  wire _27007_;
  wire _27008_;
  wire _27009_;
  wire _27010_;
  wire _27011_;
  wire _27012_;
  wire _27013_;
  wire _27014_;
  wire _27015_;
  wire _27016_;
  wire _27017_;
  wire _27018_;
  wire _27019_;
  wire _27020_;
  wire _27021_;
  wire _27022_;
  wire _27023_;
  wire _27024_;
  wire _27025_;
  wire _27026_;
  wire _27027_;
  wire _27028_;
  wire _27029_;
  wire _27030_;
  wire _27031_;
  wire _27032_;
  wire _27033_;
  wire _27034_;
  wire _27035_;
  wire _27036_;
  wire _27037_;
  wire _27038_;
  wire _27039_;
  wire _27040_;
  wire _27041_;
  wire _27042_;
  wire _27043_;
  wire _27044_;
  wire _27045_;
  wire _27046_;
  wire _27047_;
  wire _27048_;
  wire _27049_;
  wire _27050_;
  wire _27051_;
  wire _27052_;
  wire _27053_;
  wire _27054_;
  wire _27055_;
  wire _27056_;
  wire _27057_;
  wire _27058_;
  wire _27059_;
  wire _27060_;
  wire _27061_;
  wire _27062_;
  wire _27063_;
  wire _27064_;
  wire _27065_;
  wire _27066_;
  wire _27067_;
  wire _27068_;
  wire _27069_;
  wire _27070_;
  wire _27071_;
  wire _27072_;
  wire _27073_;
  wire _27074_;
  wire _27075_;
  wire _27076_;
  wire _27077_;
  wire _27078_;
  wire _27079_;
  wire _27080_;
  wire _27081_;
  wire _27082_;
  wire _27083_;
  wire _27084_;
  wire _27085_;
  wire _27086_;
  wire _27087_;
  wire _27088_;
  wire _27089_;
  wire _27090_;
  wire _27091_;
  wire _27092_;
  wire _27093_;
  wire _27094_;
  wire _27095_;
  wire _27096_;
  wire _27097_;
  wire _27098_;
  wire _27099_;
  wire _27100_;
  wire _27101_;
  wire _27102_;
  wire _27103_;
  wire _27104_;
  wire _27105_;
  wire _27106_;
  wire _27107_;
  wire _27108_;
  wire _27109_;
  wire _27110_;
  wire _27111_;
  wire _27112_;
  wire _27113_;
  wire _27114_;
  wire _27115_;
  wire _27116_;
  wire _27117_;
  wire _27118_;
  wire _27119_;
  wire _27120_;
  wire _27121_;
  wire _27122_;
  wire _27123_;
  wire _27124_;
  wire _27125_;
  wire _27126_;
  wire _27127_;
  wire _27128_;
  wire _27129_;
  wire _27130_;
  wire _27131_;
  wire _27132_;
  wire _27133_;
  wire _27134_;
  wire _27135_;
  wire _27136_;
  wire _27137_;
  wire _27138_;
  wire _27139_;
  wire _27140_;
  wire _27141_;
  wire _27142_;
  wire _27143_;
  wire _27144_;
  wire _27145_;
  wire _27146_;
  wire _27147_;
  wire _27148_;
  wire _27149_;
  wire _27150_;
  wire _27151_;
  wire _27152_;
  wire _27153_;
  wire _27154_;
  wire _27155_;
  wire _27156_;
  wire _27157_;
  wire _27158_;
  wire _27159_;
  wire _27160_;
  wire _27161_;
  wire _27162_;
  wire _27163_;
  wire _27164_;
  wire _27165_;
  wire _27166_;
  wire _27167_;
  wire _27168_;
  wire _27169_;
  wire _27170_;
  wire _27171_;
  wire _27172_;
  wire _27173_;
  wire _27174_;
  wire _27175_;
  wire _27176_;
  wire _27177_;
  wire _27178_;
  wire _27179_;
  wire _27180_;
  wire _27181_;
  wire _27182_;
  wire _27183_;
  wire _27184_;
  wire _27185_;
  wire _27186_;
  wire _27187_;
  wire _27188_;
  wire _27189_;
  wire _27190_;
  wire _27191_;
  wire _27192_;
  wire _27193_;
  wire _27194_;
  wire _27195_;
  wire _27196_;
  wire _27197_;
  wire _27198_;
  wire _27199_;
  wire _27200_;
  wire _27201_;
  wire _27202_;
  wire _27203_;
  wire _27204_;
  wire _27205_;
  wire _27206_;
  wire _27207_;
  wire _27208_;
  wire _27209_;
  wire _27210_;
  wire _27211_;
  wire _27212_;
  wire _27213_;
  wire _27214_;
  wire _27215_;
  wire _27216_;
  wire _27217_;
  wire _27218_;
  wire _27219_;
  wire _27220_;
  wire _27221_;
  wire _27222_;
  wire _27223_;
  wire _27224_;
  wire _27225_;
  wire _27226_;
  wire _27227_;
  wire _27228_;
  wire _27229_;
  wire _27230_;
  wire _27231_;
  wire _27232_;
  wire _27233_;
  wire _27234_;
  wire _27235_;
  wire _27236_;
  wire _27237_;
  wire _27238_;
  wire _27239_;
  wire _27240_;
  wire _27241_;
  wire _27242_;
  wire _27243_;
  wire _27244_;
  wire _27245_;
  wire _27246_;
  wire _27247_;
  wire _27248_;
  wire _27249_;
  wire _27250_;
  wire _27251_;
  wire _27252_;
  wire _27253_;
  wire _27254_;
  wire _27255_;
  wire _27256_;
  wire _27257_;
  wire _27258_;
  wire _27259_;
  wire _27260_;
  wire _27261_;
  wire _27262_;
  wire _27263_;
  wire _27264_;
  wire _27265_;
  wire _27266_;
  wire _27267_;
  wire _27268_;
  wire _27269_;
  wire _27270_;
  wire _27271_;
  wire _27272_;
  wire _27273_;
  wire _27274_;
  wire _27275_;
  wire _27276_;
  wire _27277_;
  wire _27278_;
  wire _27279_;
  wire _27280_;
  wire _27281_;
  wire _27282_;
  wire _27283_;
  wire _27284_;
  wire _27285_;
  wire _27286_;
  wire _27287_;
  wire _27288_;
  wire _27289_;
  wire _27290_;
  wire _27291_;
  wire _27292_;
  wire _27293_;
  wire _27294_;
  wire _27295_;
  wire _27296_;
  wire _27297_;
  wire _27298_;
  wire _27299_;
  wire _27300_;
  wire _27301_;
  wire _27302_;
  wire _27303_;
  wire _27304_;
  wire _27305_;
  wire _27306_;
  wire _27307_;
  wire _27308_;
  wire _27309_;
  wire _27310_;
  wire _27311_;
  wire _27312_;
  wire _27313_;
  wire _27314_;
  wire _27315_;
  wire _27316_;
  wire _27317_;
  wire _27318_;
  wire _27319_;
  wire _27320_;
  wire _27321_;
  wire _27322_;
  wire _27323_;
  wire _27324_;
  wire _27325_;
  wire _27326_;
  wire _27327_;
  wire _27328_;
  wire _27329_;
  wire _27330_;
  wire _27331_;
  wire _27332_;
  wire _27333_;
  wire _27334_;
  wire _27335_;
  wire _27336_;
  wire _27337_;
  wire _27338_;
  wire _27339_;
  wire _27340_;
  wire _27341_;
  wire _27342_;
  wire _27343_;
  wire _27344_;
  wire _27345_;
  wire _27346_;
  wire _27347_;
  wire _27348_;
  wire _27349_;
  wire _27350_;
  wire _27351_;
  wire _27352_;
  wire _27353_;
  wire _27354_;
  wire _27355_;
  wire _27356_;
  wire _27357_;
  wire _27358_;
  wire _27359_;
  wire _27360_;
  wire _27361_;
  wire _27362_;
  wire _27363_;
  wire _27364_;
  wire _27365_;
  wire _27366_;
  wire _27367_;
  wire _27368_;
  wire _27369_;
  wire _27370_;
  wire _27371_;
  wire _27372_;
  wire _27373_;
  wire _27374_;
  wire _27375_;
  wire _27376_;
  wire _27377_;
  wire _27378_;
  wire _27379_;
  wire _27380_;
  wire _27381_;
  wire _27382_;
  wire _27383_;
  wire _27384_;
  wire _27385_;
  wire _27386_;
  wire _27387_;
  wire _27388_;
  wire _27389_;
  wire _27390_;
  wire _27391_;
  wire _27392_;
  wire _27393_;
  wire _27394_;
  wire _27395_;
  wire _27396_;
  wire _27397_;
  wire _27398_;
  wire _27399_;
  wire _27400_;
  wire _27401_;
  wire _27402_;
  wire _27403_;
  wire _27404_;
  wire _27405_;
  wire _27406_;
  wire _27407_;
  wire _27408_;
  wire _27409_;
  wire _27410_;
  wire _27411_;
  wire _27412_;
  wire _27413_;
  wire _27414_;
  wire _27415_;
  wire _27416_;
  wire _27417_;
  wire _27418_;
  wire _27419_;
  wire _27420_;
  wire _27421_;
  wire _27422_;
  wire _27423_;
  wire _27424_;
  wire _27425_;
  wire _27426_;
  wire _27427_;
  wire _27428_;
  wire _27429_;
  wire _27430_;
  wire _27431_;
  wire _27432_;
  wire _27433_;
  wire _27434_;
  wire _27435_;
  wire _27436_;
  wire _27437_;
  wire _27438_;
  wire _27439_;
  wire _27440_;
  wire _27441_;
  wire _27442_;
  wire _27443_;
  wire _27444_;
  wire _27445_;
  wire _27446_;
  wire _27447_;
  wire _27448_;
  wire _27449_;
  wire _27450_;
  wire _27451_;
  wire _27452_;
  wire _27453_;
  wire _27454_;
  wire _27455_;
  wire _27456_;
  wire _27457_;
  wire _27458_;
  wire _27459_;
  wire _27460_;
  wire _27461_;
  wire _27462_;
  wire _27463_;
  wire _27464_;
  wire _27465_;
  wire _27466_;
  wire _27467_;
  wire _27468_;
  wire _27469_;
  wire _27470_;
  wire _27471_;
  wire _27472_;
  wire _27473_;
  wire _27474_;
  wire _27475_;
  wire _27476_;
  wire _27477_;
  wire _27478_;
  wire _27479_;
  wire _27480_;
  wire _27481_;
  wire _27482_;
  wire _27483_;
  wire _27484_;
  wire _27485_;
  wire _27486_;
  wire _27487_;
  wire _27488_;
  wire _27489_;
  wire _27490_;
  wire _27491_;
  wire _27492_;
  wire _27493_;
  wire _27494_;
  wire _27495_;
  wire _27496_;
  wire _27497_;
  wire _27498_;
  wire _27499_;
  wire _27500_;
  wire _27501_;
  wire _27502_;
  wire _27503_;
  wire _27504_;
  wire _27505_;
  wire _27506_;
  wire _27507_;
  wire _27508_;
  wire _27509_;
  wire _27510_;
  wire _27511_;
  wire _27512_;
  wire _27513_;
  wire _27514_;
  wire _27515_;
  wire _27516_;
  wire _27517_;
  wire _27518_;
  wire _27519_;
  wire _27520_;
  wire _27521_;
  wire _27522_;
  wire _27523_;
  wire _27524_;
  wire _27525_;
  wire _27526_;
  wire _27527_;
  wire _27528_;
  wire _27529_;
  wire _27530_;
  wire _27531_;
  wire _27532_;
  wire _27533_;
  wire _27534_;
  wire _27535_;
  wire _27536_;
  wire _27537_;
  wire _27538_;
  wire _27539_;
  wire _27540_;
  wire _27541_;
  wire _27542_;
  wire _27543_;
  wire _27544_;
  wire _27545_;
  wire _27546_;
  wire _27547_;
  wire _27548_;
  wire _27549_;
  wire _27550_;
  wire _27551_;
  wire _27552_;
  wire _27553_;
  wire _27554_;
  wire _27555_;
  wire _27556_;
  wire _27557_;
  wire _27558_;
  wire _27559_;
  wire _27560_;
  wire _27561_;
  wire _27562_;
  wire _27563_;
  wire _27564_;
  wire _27565_;
  wire _27566_;
  wire _27567_;
  wire _27568_;
  wire _27569_;
  wire _27570_;
  wire _27571_;
  wire _27572_;
  wire _27573_;
  wire _27574_;
  wire _27575_;
  wire _27576_;
  wire _27577_;
  wire _27578_;
  wire _27579_;
  wire _27580_;
  wire _27581_;
  wire _27582_;
  wire _27583_;
  wire _27584_;
  wire _27585_;
  wire _27586_;
  wire _27587_;
  wire _27588_;
  wire _27589_;
  wire _27590_;
  wire _27591_;
  wire _27592_;
  wire _27593_;
  wire _27594_;
  wire _27595_;
  wire _27596_;
  wire _27597_;
  wire _27598_;
  wire _27599_;
  wire _27600_;
  wire _27601_;
  wire _27602_;
  wire _27603_;
  wire _27604_;
  wire _27605_;
  wire _27606_;
  wire _27607_;
  wire _27608_;
  wire _27609_;
  wire _27610_;
  wire _27611_;
  wire _27612_;
  wire _27613_;
  wire _27614_;
  wire _27615_;
  wire _27616_;
  wire _27617_;
  wire _27618_;
  wire _27619_;
  wire _27620_;
  wire _27621_;
  wire _27622_;
  wire _27623_;
  wire _27624_;
  wire _27625_;
  wire _27626_;
  wire _27627_;
  wire _27628_;
  wire _27629_;
  wire _27630_;
  wire _27631_;
  wire _27632_;
  wire _27633_;
  wire _27634_;
  wire _27635_;
  wire _27636_;
  wire _27637_;
  wire _27638_;
  wire _27639_;
  wire _27640_;
  wire _27641_;
  wire _27642_;
  wire _27643_;
  wire _27644_;
  wire _27645_;
  wire _27646_;
  wire _27647_;
  wire _27648_;
  wire _27649_;
  wire _27650_;
  wire _27651_;
  wire _27652_;
  wire _27653_;
  wire _27654_;
  wire _27655_;
  wire _27656_;
  wire _27657_;
  wire _27658_;
  wire _27659_;
  wire _27660_;
  wire _27661_;
  wire _27662_;
  wire _27663_;
  wire _27664_;
  wire _27665_;
  wire _27666_;
  wire _27667_;
  wire _27668_;
  wire _27669_;
  wire _27670_;
  wire _27671_;
  wire _27672_;
  wire _27673_;
  wire _27674_;
  wire _27675_;
  wire _27676_;
  wire _27677_;
  wire _27678_;
  wire _27679_;
  wire _27680_;
  wire _27681_;
  wire _27682_;
  wire _27683_;
  wire _27684_;
  wire _27685_;
  wire _27686_;
  wire _27687_;
  wire _27688_;
  wire _27689_;
  wire _27690_;
  wire _27691_;
  wire _27692_;
  wire _27693_;
  wire _27694_;
  wire _27695_;
  wire _27696_;
  wire _27697_;
  wire _27698_;
  wire _27699_;
  wire _27700_;
  wire _27701_;
  wire _27702_;
  wire _27703_;
  wire _27704_;
  wire _27705_;
  wire _27706_;
  wire _27707_;
  wire _27708_;
  wire _27709_;
  wire _27710_;
  wire _27711_;
  wire _27712_;
  wire _27713_;
  wire _27714_;
  wire _27715_;
  wire _27716_;
  wire _27717_;
  wire _27718_;
  wire _27719_;
  wire _27720_;
  wire _27721_;
  wire _27722_;
  wire _27723_;
  wire _27724_;
  wire _27725_;
  wire _27726_;
  wire _27727_;
  wire _27728_;
  wire _27729_;
  wire _27730_;
  wire _27731_;
  wire _27732_;
  wire _27733_;
  wire _27734_;
  wire _27735_;
  wire _27736_;
  wire _27737_;
  wire _27738_;
  wire _27739_;
  wire _27740_;
  wire _27741_;
  wire _27742_;
  wire _27743_;
  wire _27744_;
  wire _27745_;
  wire _27746_;
  wire _27747_;
  wire _27748_;
  wire _27749_;
  wire _27750_;
  wire _27751_;
  wire _27752_;
  wire _27753_;
  wire _27754_;
  wire _27755_;
  wire _27756_;
  wire _27757_;
  wire _27758_;
  wire _27759_;
  wire _27760_;
  wire _27761_;
  wire _27762_;
  wire _27763_;
  wire _27764_;
  wire _27765_;
  wire _27766_;
  wire _27767_;
  wire _27768_;
  wire _27769_;
  wire _27770_;
  wire _27771_;
  wire _27772_;
  wire _27773_;
  wire _27774_;
  wire _27775_;
  wire _27776_;
  wire _27777_;
  wire _27778_;
  wire _27779_;
  wire _27780_;
  wire _27781_;
  wire _27782_;
  wire _27783_;
  wire _27784_;
  wire _27785_;
  wire _27786_;
  wire _27787_;
  wire _27788_;
  wire _27789_;
  wire _27790_;
  wire _27791_;
  wire _27792_;
  wire _27793_;
  wire _27794_;
  wire _27795_;
  wire _27796_;
  wire _27797_;
  wire _27798_;
  wire _27799_;
  wire _27800_;
  wire _27801_;
  wire _27802_;
  wire _27803_;
  wire _27804_;
  wire _27805_;
  wire _27806_;
  wire _27807_;
  wire _27808_;
  wire _27809_;
  wire _27810_;
  wire _27811_;
  wire _27812_;
  wire _27813_;
  wire _27814_;
  wire _27815_;
  wire _27816_;
  wire _27817_;
  wire _27818_;
  wire _27819_;
  wire _27820_;
  wire _27821_;
  wire _27822_;
  wire _27823_;
  wire _27824_;
  wire _27825_;
  wire _27826_;
  wire _27827_;
  wire _27828_;
  wire _27829_;
  wire _27830_;
  wire _27831_;
  wire _27832_;
  wire _27833_;
  wire _27834_;
  wire _27835_;
  wire _27836_;
  wire _27837_;
  wire _27838_;
  wire _27839_;
  wire _27840_;
  wire _27841_;
  wire _27842_;
  wire _27843_;
  wire _27844_;
  wire _27845_;
  wire _27846_;
  wire _27847_;
  wire _27848_;
  wire _27849_;
  wire _27850_;
  wire _27851_;
  wire _27852_;
  wire _27853_;
  wire _27854_;
  wire _27855_;
  wire _27856_;
  wire _27857_;
  wire _27858_;
  wire _27859_;
  wire _27860_;
  wire _27861_;
  wire _27862_;
  wire _27863_;
  wire _27864_;
  wire _27865_;
  wire _27866_;
  wire _27867_;
  wire _27868_;
  wire _27869_;
  wire _27870_;
  wire _27871_;
  wire _27872_;
  wire _27873_;
  wire _27874_;
  wire _27875_;
  wire _27876_;
  wire _27877_;
  wire _27878_;
  wire _27879_;
  wire _27880_;
  wire _27881_;
  wire _27882_;
  wire _27883_;
  wire _27884_;
  wire _27885_;
  wire _27886_;
  wire _27887_;
  wire _27888_;
  wire _27889_;
  wire _27890_;
  wire _27891_;
  wire _27892_;
  wire _27893_;
  wire _27894_;
  wire _27895_;
  wire _27896_;
  wire _27897_;
  wire _27898_;
  wire _27899_;
  wire _27900_;
  wire _27901_;
  wire _27902_;
  wire _27903_;
  wire _27904_;
  wire _27905_;
  wire _27906_;
  wire _27907_;
  wire _27908_;
  wire _27909_;
  wire _27910_;
  wire _27911_;
  wire _27912_;
  wire _27913_;
  wire _27914_;
  wire _27915_;
  wire _27916_;
  wire _27917_;
  wire _27918_;
  wire _27919_;
  wire _27920_;
  wire _27921_;
  wire _27922_;
  wire _27923_;
  wire _27924_;
  wire _27925_;
  wire _27926_;
  wire _27927_;
  wire _27928_;
  wire _27929_;
  wire _27930_;
  wire _27931_;
  wire _27932_;
  wire _27933_;
  wire _27934_;
  wire _27935_;
  wire _27936_;
  wire _27937_;
  wire _27938_;
  wire _27939_;
  wire _27940_;
  wire _27941_;
  wire _27942_;
  wire _27943_;
  wire _27944_;
  wire _27945_;
  wire _27946_;
  wire _27947_;
  wire _27948_;
  wire _27949_;
  wire _27950_;
  wire _27951_;
  wire _27952_;
  wire _27953_;
  wire _27954_;
  wire _27955_;
  wire _27956_;
  wire _27957_;
  wire _27958_;
  wire _27959_;
  wire _27960_;
  wire _27961_;
  wire _27962_;
  wire _27963_;
  wire _27964_;
  wire _27965_;
  wire _27966_;
  wire _27967_;
  wire _27968_;
  wire _27969_;
  wire _27970_;
  wire _27971_;
  wire _27972_;
  wire _27973_;
  wire _27974_;
  wire _27975_;
  wire _27976_;
  wire _27977_;
  wire _27978_;
  wire _27979_;
  wire _27980_;
  wire _27981_;
  wire _27982_;
  wire _27983_;
  wire _27984_;
  wire _27985_;
  wire _27986_;
  wire _27987_;
  wire _27988_;
  wire _27989_;
  wire _27990_;
  wire _27991_;
  wire _27992_;
  wire _27993_;
  wire _27994_;
  wire _27995_;
  wire _27996_;
  wire _27997_;
  wire _27998_;
  wire _27999_;
  wire _28000_;
  wire _28001_;
  wire _28002_;
  wire _28003_;
  wire _28004_;
  wire _28005_;
  wire _28006_;
  wire _28007_;
  wire _28008_;
  wire _28009_;
  wire _28010_;
  wire _28011_;
  wire _28012_;
  wire _28013_;
  wire _28014_;
  wire _28015_;
  wire _28016_;
  wire _28017_;
  wire _28018_;
  wire _28019_;
  wire _28020_;
  wire _28021_;
  wire _28022_;
  wire _28023_;
  wire _28024_;
  wire _28025_;
  wire _28026_;
  wire _28027_;
  wire _28028_;
  wire _28029_;
  wire _28030_;
  wire _28031_;
  wire _28032_;
  wire _28033_;
  wire _28034_;
  wire _28035_;
  wire _28036_;
  wire _28037_;
  wire _28038_;
  wire _28039_;
  wire _28040_;
  wire _28041_;
  wire _28042_;
  wire _28043_;
  wire _28044_;
  wire _28045_;
  wire _28046_;
  wire _28047_;
  wire _28048_;
  wire _28049_;
  wire _28050_;
  wire _28051_;
  wire _28052_;
  wire _28053_;
  wire _28054_;
  wire _28055_;
  wire _28056_;
  wire _28057_;
  wire _28058_;
  wire _28059_;
  wire _28060_;
  wire _28061_;
  wire _28062_;
  wire _28063_;
  wire _28064_;
  wire _28065_;
  wire _28066_;
  wire _28067_;
  wire _28068_;
  wire _28069_;
  wire _28070_;
  wire _28071_;
  wire _28072_;
  wire _28073_;
  wire _28074_;
  wire _28075_;
  wire _28076_;
  wire _28077_;
  wire _28078_;
  wire _28079_;
  wire _28080_;
  wire _28081_;
  wire _28082_;
  wire _28083_;
  wire _28084_;
  wire _28085_;
  wire _28086_;
  wire _28087_;
  wire _28088_;
  wire _28089_;
  wire _28090_;
  wire _28091_;
  wire _28092_;
  wire _28093_;
  wire _28094_;
  wire _28095_;
  wire _28096_;
  wire _28097_;
  wire _28098_;
  wire _28099_;
  wire _28100_;
  wire _28101_;
  wire _28102_;
  wire _28103_;
  wire _28104_;
  wire _28105_;
  wire _28106_;
  wire _28107_;
  wire _28108_;
  wire _28109_;
  wire _28110_;
  wire _28111_;
  wire _28112_;
  wire _28113_;
  wire _28114_;
  wire _28115_;
  wire _28116_;
  wire _28117_;
  wire _28118_;
  wire _28119_;
  wire _28120_;
  wire _28121_;
  wire _28122_;
  wire _28123_;
  wire _28124_;
  wire _28125_;
  wire _28126_;
  wire _28127_;
  wire _28128_;
  wire _28129_;
  wire _28130_;
  wire _28131_;
  wire _28132_;
  wire _28133_;
  wire _28134_;
  wire _28135_;
  wire _28136_;
  wire _28137_;
  wire _28138_;
  wire _28139_;
  wire _28140_;
  wire _28141_;
  wire _28142_;
  wire _28143_;
  wire _28144_;
  wire _28145_;
  wire _28146_;
  wire _28147_;
  wire _28148_;
  wire _28149_;
  wire _28150_;
  wire _28151_;
  wire _28152_;
  wire _28153_;
  wire _28154_;
  wire _28155_;
  wire _28156_;
  wire _28157_;
  wire _28158_;
  wire _28159_;
  wire _28160_;
  wire _28161_;
  wire _28162_;
  wire _28163_;
  wire _28164_;
  wire _28165_;
  wire _28166_;
  wire _28167_;
  wire _28168_;
  wire _28169_;
  wire _28170_;
  wire _28171_;
  wire _28172_;
  wire _28173_;
  wire _28174_;
  wire _28175_;
  wire _28176_;
  wire _28177_;
  wire _28178_;
  wire _28179_;
  wire _28180_;
  wire _28181_;
  wire _28182_;
  wire _28183_;
  wire _28184_;
  wire _28185_;
  wire _28186_;
  wire _28187_;
  wire _28188_;
  wire _28189_;
  wire _28190_;
  wire _28191_;
  wire _28192_;
  wire _28193_;
  wire _28194_;
  wire _28195_;
  wire _28196_;
  wire _28197_;
  wire _28198_;
  wire _28199_;
  wire _28200_;
  wire _28201_;
  wire _28202_;
  wire _28203_;
  wire _28204_;
  wire _28205_;
  wire _28206_;
  wire _28207_;
  wire _28208_;
  wire _28209_;
  wire _28210_;
  wire _28211_;
  wire _28212_;
  wire _28213_;
  wire _28214_;
  wire _28215_;
  wire _28216_;
  wire _28217_;
  wire _28218_;
  wire _28219_;
  wire _28220_;
  wire _28221_;
  wire _28222_;
  wire _28223_;
  wire _28224_;
  wire _28225_;
  wire _28226_;
  wire _28227_;
  wire _28228_;
  wire _28229_;
  wire _28230_;
  wire _28231_;
  wire _28232_;
  wire _28233_;
  wire _28234_;
  wire _28235_;
  wire _28236_;
  wire _28237_;
  wire _28238_;
  wire _28239_;
  wire _28240_;
  wire _28241_;
  wire _28242_;
  wire _28243_;
  wire _28244_;
  wire _28245_;
  wire _28246_;
  wire _28247_;
  wire _28248_;
  wire _28249_;
  wire _28250_;
  wire _28251_;
  wire _28252_;
  wire _28253_;
  wire _28254_;
  wire _28255_;
  wire _28256_;
  wire _28257_;
  wire _28258_;
  wire _28259_;
  wire _28260_;
  wire _28261_;
  wire _28262_;
  wire _28263_;
  wire _28264_;
  wire _28265_;
  wire _28266_;
  wire _28267_;
  wire _28268_;
  wire _28269_;
  wire _28270_;
  wire _28271_;
  wire _28272_;
  wire _28273_;
  wire _28274_;
  wire _28275_;
  wire _28276_;
  wire _28277_;
  wire _28278_;
  wire _28279_;
  wire _28280_;
  wire _28281_;
  wire _28282_;
  wire _28283_;
  wire _28284_;
  wire _28285_;
  wire _28286_;
  wire _28287_;
  wire _28288_;
  wire _28289_;
  wire _28290_;
  wire _28291_;
  wire _28292_;
  wire _28293_;
  wire _28294_;
  wire _28295_;
  wire _28296_;
  wire _28297_;
  wire _28298_;
  wire _28299_;
  wire _28300_;
  wire _28301_;
  wire _28302_;
  wire _28303_;
  wire _28304_;
  wire _28305_;
  wire _28306_;
  wire _28307_;
  wire _28308_;
  wire _28309_;
  wire _28310_;
  wire _28311_;
  wire _28312_;
  wire _28313_;
  wire _28314_;
  wire _28315_;
  wire _28316_;
  wire _28317_;
  wire _28318_;
  wire _28319_;
  wire _28320_;
  wire _28321_;
  wire _28322_;
  wire _28323_;
  wire _28324_;
  wire _28325_;
  wire _28326_;
  wire _28327_;
  wire _28328_;
  wire _28329_;
  wire _28330_;
  wire _28331_;
  wire _28332_;
  wire _28333_;
  wire _28334_;
  wire _28335_;
  wire _28336_;
  wire _28337_;
  wire _28338_;
  wire _28339_;
  wire _28340_;
  wire _28341_;
  wire _28342_;
  wire _28343_;
  wire _28344_;
  wire _28345_;
  wire _28346_;
  wire _28347_;
  wire _28348_;
  wire _28349_;
  wire _28350_;
  wire _28351_;
  wire _28352_;
  wire _28353_;
  wire _28354_;
  wire _28355_;
  wire _28356_;
  wire _28357_;
  wire _28358_;
  wire _28359_;
  wire _28360_;
  wire _28361_;
  wire _28362_;
  wire _28363_;
  wire _28364_;
  wire _28365_;
  wire _28366_;
  wire _28367_;
  wire _28368_;
  wire _28369_;
  wire _28370_;
  wire _28371_;
  wire _28372_;
  wire _28373_;
  wire _28374_;
  wire _28375_;
  wire _28376_;
  wire _28377_;
  wire _28378_;
  wire _28379_;
  wire _28380_;
  wire _28381_;
  wire _28382_;
  wire _28383_;
  wire _28384_;
  wire _28385_;
  wire _28386_;
  wire _28387_;
  wire _28388_;
  wire _28389_;
  wire _28390_;
  wire _28391_;
  wire _28392_;
  wire _28393_;
  wire _28394_;
  wire _28395_;
  wire _28396_;
  wire _28397_;
  wire _28398_;
  wire _28399_;
  wire _28400_;
  wire _28401_;
  wire _28402_;
  wire _28403_;
  wire _28404_;
  wire _28405_;
  wire _28406_;
  wire _28407_;
  wire _28408_;
  wire _28409_;
  wire _28410_;
  wire _28411_;
  wire _28412_;
  wire _28413_;
  wire _28414_;
  wire _28415_;
  wire _28416_;
  wire _28417_;
  wire _28418_;
  wire _28419_;
  wire _28420_;
  wire _28421_;
  wire _28422_;
  wire _28423_;
  wire _28424_;
  wire _28425_;
  wire _28426_;
  wire _28427_;
  wire _28428_;
  wire _28429_;
  wire _28430_;
  wire _28431_;
  wire _28432_;
  wire _28433_;
  wire _28434_;
  wire _28435_;
  wire _28436_;
  wire _28437_;
  wire _28438_;
  wire _28439_;
  wire _28440_;
  wire _28441_;
  wire _28442_;
  wire _28443_;
  wire _28444_;
  wire _28445_;
  wire _28446_;
  wire _28447_;
  wire _28448_;
  wire _28449_;
  wire _28450_;
  wire _28451_;
  wire _28452_;
  wire _28453_;
  wire _28454_;
  wire _28455_;
  wire _28456_;
  wire _28457_;
  wire _28458_;
  wire _28459_;
  wire _28460_;
  wire _28461_;
  wire _28462_;
  wire _28463_;
  wire _28464_;
  wire _28465_;
  wire _28466_;
  wire _28467_;
  wire _28468_;
  wire _28469_;
  wire _28470_;
  wire _28471_;
  wire _28472_;
  wire _28473_;
  wire _28474_;
  wire _28475_;
  wire _28476_;
  wire _28477_;
  wire _28478_;
  wire _28479_;
  wire _28480_;
  wire _28481_;
  wire _28482_;
  wire _28483_;
  wire _28484_;
  wire _28485_;
  wire _28486_;
  wire _28487_;
  wire _28488_;
  wire _28489_;
  wire _28490_;
  wire _28491_;
  wire _28492_;
  wire _28493_;
  wire _28494_;
  wire _28495_;
  wire _28496_;
  wire _28497_;
  wire _28498_;
  wire _28499_;
  wire _28500_;
  wire _28501_;
  wire _28502_;
  wire _28503_;
  wire _28504_;
  wire _28505_;
  wire _28506_;
  wire _28507_;
  wire _28508_;
  wire _28509_;
  wire _28510_;
  wire _28511_;
  wire _28512_;
  wire _28513_;
  wire _28514_;
  wire _28515_;
  wire _28516_;
  wire _28517_;
  wire _28518_;
  wire _28519_;
  wire _28520_;
  wire _28521_;
  wire _28522_;
  wire _28523_;
  wire _28524_;
  wire _28525_;
  wire _28526_;
  wire _28527_;
  wire _28528_;
  wire _28529_;
  wire _28530_;
  wire _28531_;
  wire _28532_;
  wire _28533_;
  wire _28534_;
  wire _28535_;
  wire _28536_;
  wire _28537_;
  wire _28538_;
  wire _28539_;
  wire _28540_;
  wire _28541_;
  wire _28542_;
  wire _28543_;
  wire _28544_;
  wire _28545_;
  wire _28546_;
  wire _28547_;
  wire _28548_;
  wire _28549_;
  wire _28550_;
  wire _28551_;
  wire _28552_;
  wire _28553_;
  wire _28554_;
  wire _28555_;
  wire _28556_;
  wire _28557_;
  wire _28558_;
  wire _28559_;
  wire _28560_;
  wire _28561_;
  wire _28562_;
  wire _28563_;
  wire _28564_;
  wire _28565_;
  wire _28566_;
  wire _28567_;
  wire _28568_;
  wire _28569_;
  wire _28570_;
  wire _28571_;
  wire _28572_;
  wire _28573_;
  wire _28574_;
  wire _28575_;
  wire _28576_;
  wire _28577_;
  wire _28578_;
  wire _28579_;
  wire _28580_;
  wire _28581_;
  wire _28582_;
  wire _28583_;
  wire _28584_;
  wire _28585_;
  wire _28586_;
  wire _28587_;
  wire _28588_;
  wire _28589_;
  wire _28590_;
  wire _28591_;
  wire _28592_;
  wire _28593_;
  wire _28594_;
  wire _28595_;
  wire _28596_;
  wire _28597_;
  wire _28598_;
  wire _28599_;
  wire _28600_;
  wire _28601_;
  wire _28602_;
  wire _28603_;
  wire _28604_;
  wire _28605_;
  wire _28606_;
  wire _28607_;
  wire _28608_;
  wire _28609_;
  wire _28610_;
  wire _28611_;
  wire _28612_;
  wire _28613_;
  wire _28614_;
  wire _28615_;
  wire _28616_;
  wire _28617_;
  wire _28618_;
  wire _28619_;
  wire _28620_;
  wire _28621_;
  wire _28622_;
  wire _28623_;
  wire _28624_;
  wire _28625_;
  wire _28626_;
  wire _28627_;
  wire _28628_;
  wire _28629_;
  wire _28630_;
  wire _28631_;
  wire _28632_;
  wire _28633_;
  wire _28634_;
  wire _28635_;
  wire _28636_;
  wire _28637_;
  wire _28638_;
  wire _28639_;
  wire _28640_;
  wire _28641_;
  wire _28642_;
  wire _28643_;
  wire _28644_;
  wire _28645_;
  wire _28646_;
  wire _28647_;
  wire _28648_;
  wire _28649_;
  wire _28650_;
  wire _28651_;
  wire _28652_;
  wire _28653_;
  wire _28654_;
  wire _28655_;
  wire _28656_;
  wire _28657_;
  wire _28658_;
  wire _28659_;
  wire _28660_;
  wire _28661_;
  wire _28662_;
  wire _28663_;
  wire _28664_;
  wire _28665_;
  wire _28666_;
  wire _28667_;
  wire _28668_;
  wire _28669_;
  wire _28670_;
  wire _28671_;
  wire _28672_;
  wire _28673_;
  wire _28674_;
  wire _28675_;
  wire _28676_;
  wire _28677_;
  wire _28678_;
  wire _28679_;
  wire _28680_;
  wire _28681_;
  wire _28682_;
  wire _28683_;
  wire _28684_;
  wire _28685_;
  wire _28686_;
  wire _28687_;
  wire _28688_;
  wire _28689_;
  wire _28690_;
  wire _28691_;
  wire _28692_;
  wire _28693_;
  wire _28694_;
  wire _28695_;
  wire _28696_;
  wire _28697_;
  wire _28698_;
  wire _28699_;
  wire _28700_;
  wire _28701_;
  wire _28702_;
  wire _28703_;
  wire _28704_;
  wire _28705_;
  wire _28706_;
  wire _28707_;
  wire _28708_;
  wire _28709_;
  wire _28710_;
  wire _28711_;
  wire _28712_;
  wire _28713_;
  wire _28714_;
  wire _28715_;
  wire _28716_;
  wire _28717_;
  wire _28718_;
  wire _28719_;
  wire _28720_;
  wire _28721_;
  wire _28722_;
  wire _28723_;
  wire _28724_;
  wire _28725_;
  wire _28726_;
  wire _28727_;
  wire _28728_;
  wire _28729_;
  wire _28730_;
  wire _28731_;
  wire _28732_;
  wire _28733_;
  wire _28734_;
  wire _28735_;
  wire _28736_;
  wire _28737_;
  wire _28738_;
  wire _28739_;
  wire _28740_;
  wire _28741_;
  wire _28742_;
  wire _28743_;
  wire _28744_;
  wire _28745_;
  wire _28746_;
  wire _28747_;
  wire _28748_;
  wire _28749_;
  wire _28750_;
  wire _28751_;
  wire _28752_;
  wire _28753_;
  wire _28754_;
  wire _28755_;
  wire _28756_;
  wire _28757_;
  wire _28758_;
  wire _28759_;
  wire _28760_;
  wire _28761_;
  wire _28762_;
  wire _28763_;
  wire _28764_;
  wire _28765_;
  wire _28766_;
  wire _28767_;
  wire _28768_;
  wire _28769_;
  wire _28770_;
  wire _28771_;
  wire _28772_;
  wire _28773_;
  wire _28774_;
  wire _28775_;
  wire _28776_;
  wire _28777_;
  wire _28778_;
  wire _28779_;
  wire _28780_;
  wire _28781_;
  wire _28782_;
  wire _28783_;
  wire _28784_;
  wire _28785_;
  wire _28786_;
  wire _28787_;
  wire _28788_;
  wire _28789_;
  wire _28790_;
  wire _28791_;
  wire _28792_;
  wire _28793_;
  wire _28794_;
  wire _28795_;
  wire _28796_;
  wire _28797_;
  wire _28798_;
  wire _28799_;
  wire _28800_;
  wire _28801_;
  wire _28802_;
  wire _28803_;
  wire _28804_;
  wire _28805_;
  wire _28806_;
  wire _28807_;
  wire _28808_;
  wire _28809_;
  wire _28810_;
  wire _28811_;
  wire _28812_;
  wire _28813_;
  wire _28814_;
  wire _28815_;
  wire _28816_;
  wire _28817_;
  wire _28818_;
  wire _28819_;
  wire _28820_;
  wire _28821_;
  wire _28822_;
  wire _28823_;
  wire _28824_;
  wire _28825_;
  wire _28826_;
  wire _28827_;
  wire _28828_;
  wire _28829_;
  wire _28830_;
  wire _28831_;
  wire _28832_;
  wire _28833_;
  wire _28834_;
  wire _28835_;
  wire _28836_;
  wire _28837_;
  wire _28838_;
  wire _28839_;
  wire _28840_;
  wire _28841_;
  wire _28842_;
  wire _28843_;
  wire _28844_;
  wire _28845_;
  wire _28846_;
  wire _28847_;
  wire _28848_;
  wire _28849_;
  wire _28850_;
  wire _28851_;
  wire _28852_;
  wire _28853_;
  wire _28854_;
  wire _28855_;
  wire _28856_;
  wire _28857_;
  wire _28858_;
  wire _28859_;
  wire _28860_;
  wire _28861_;
  wire _28862_;
  wire _28863_;
  wire _28864_;
  wire _28865_;
  wire _28866_;
  wire _28867_;
  wire _28868_;
  wire _28869_;
  wire _28870_;
  wire _28871_;
  wire _28872_;
  wire _28873_;
  wire _28874_;
  wire _28875_;
  wire _28876_;
  wire _28877_;
  wire _28878_;
  wire _28879_;
  wire _28880_;
  wire _28881_;
  wire _28882_;
  wire _28883_;
  wire _28884_;
  wire _28885_;
  wire _28886_;
  wire _28887_;
  wire _28888_;
  wire _28889_;
  wire _28890_;
  wire _28891_;
  wire _28892_;
  wire _28893_;
  wire _28894_;
  wire _28895_;
  wire _28896_;
  wire _28897_;
  wire _28898_;
  wire _28899_;
  wire _28900_;
  wire _28901_;
  wire _28902_;
  wire _28903_;
  wire _28904_;
  wire _28905_;
  wire _28906_;
  wire _28907_;
  wire _28908_;
  wire _28909_;
  wire _28910_;
  wire _28911_;
  wire _28912_;
  wire _28913_;
  wire _28914_;
  wire _28915_;
  wire _28916_;
  wire _28917_;
  wire _28918_;
  wire _28919_;
  wire _28920_;
  wire _28921_;
  wire _28922_;
  wire _28923_;
  wire _28924_;
  wire _28925_;
  wire _28926_;
  wire _28927_;
  wire _28928_;
  wire _28929_;
  wire _28930_;
  wire _28931_;
  wire _28932_;
  wire _28933_;
  wire _28934_;
  wire _28935_;
  wire _28936_;
  wire _28937_;
  wire _28938_;
  wire _28939_;
  wire _28940_;
  wire _28941_;
  wire _28942_;
  wire _28943_;
  wire _28944_;
  wire _28945_;
  wire _28946_;
  wire _28947_;
  wire _28948_;
  wire _28949_;
  wire _28950_;
  wire _28951_;
  wire _28952_;
  wire _28953_;
  wire _28954_;
  wire _28955_;
  wire _28956_;
  wire _28957_;
  wire _28958_;
  wire _28959_;
  wire _28960_;
  wire _28961_;
  wire _28962_;
  wire _28963_;
  wire _28964_;
  wire _28965_;
  wire _28966_;
  wire _28967_;
  wire _28968_;
  wire _28969_;
  wire _28970_;
  wire _28971_;
  wire _28972_;
  wire _28973_;
  wire _28974_;
  wire _28975_;
  wire _28976_;
  wire _28977_;
  wire _28978_;
  wire _28979_;
  wire _28980_;
  wire _28981_;
  wire _28982_;
  wire _28983_;
  wire _28984_;
  wire _28985_;
  wire _28986_;
  wire _28987_;
  wire _28988_;
  wire _28989_;
  wire _28990_;
  wire _28991_;
  wire _28992_;
  wire _28993_;
  wire _28994_;
  wire _28995_;
  wire _28996_;
  wire _28997_;
  wire _28998_;
  wire _28999_;
  wire _29000_;
  wire _29001_;
  wire _29002_;
  wire _29003_;
  wire _29004_;
  wire _29005_;
  wire _29006_;
  wire _29007_;
  wire _29008_;
  wire _29009_;
  wire _29010_;
  wire _29011_;
  wire _29012_;
  wire _29013_;
  wire _29014_;
  wire _29015_;
  wire _29016_;
  wire _29017_;
  wire _29018_;
  wire _29019_;
  wire _29020_;
  wire _29021_;
  wire _29022_;
  wire _29023_;
  wire _29024_;
  wire _29025_;
  wire _29026_;
  wire _29027_;
  wire _29028_;
  wire _29029_;
  wire _29030_;
  wire _29031_;
  wire _29032_;
  wire _29033_;
  wire _29034_;
  wire _29035_;
  wire _29036_;
  wire _29037_;
  wire _29038_;
  wire _29039_;
  wire _29040_;
  wire _29041_;
  wire _29042_;
  wire _29043_;
  wire _29044_;
  wire _29045_;
  wire _29046_;
  wire _29047_;
  wire _29048_;
  wire _29049_;
  wire _29050_;
  wire _29051_;
  wire _29052_;
  wire _29053_;
  wire _29054_;
  wire _29055_;
  wire _29056_;
  wire _29057_;
  wire _29058_;
  wire _29059_;
  wire _29060_;
  wire _29061_;
  wire _29062_;
  wire _29063_;
  wire _29064_;
  wire _29065_;
  wire _29066_;
  wire _29067_;
  wire _29068_;
  wire _29069_;
  wire _29070_;
  wire _29071_;
  wire _29072_;
  wire _29073_;
  wire _29074_;
  wire _29075_;
  wire _29076_;
  wire _29077_;
  wire _29078_;
  wire _29079_;
  wire _29080_;
  wire _29081_;
  wire _29082_;
  wire _29083_;
  wire _29084_;
  wire _29085_;
  wire _29086_;
  wire _29087_;
  wire _29088_;
  wire _29089_;
  wire _29090_;
  wire _29091_;
  wire _29092_;
  wire _29093_;
  wire _29094_;
  wire _29095_;
  wire _29096_;
  wire _29097_;
  wire _29098_;
  wire _29099_;
  wire _29100_;
  wire _29101_;
  wire _29102_;
  wire _29103_;
  wire _29104_;
  wire _29105_;
  wire _29106_;
  wire _29107_;
  wire _29108_;
  wire _29109_;
  wire _29110_;
  wire _29111_;
  wire _29112_;
  wire _29113_;
  wire _29114_;
  wire _29115_;
  wire _29116_;
  wire _29117_;
  wire _29118_;
  wire _29119_;
  wire _29120_;
  wire _29121_;
  wire _29122_;
  wire _29123_;
  wire _29124_;
  wire _29125_;
  wire _29126_;
  wire _29127_;
  wire _29128_;
  wire _29129_;
  wire _29130_;
  wire _29131_;
  wire _29132_;
  wire _29133_;
  wire _29134_;
  wire _29135_;
  wire _29136_;
  wire _29137_;
  wire _29138_;
  wire _29139_;
  wire _29140_;
  wire _29141_;
  wire _29142_;
  wire _29143_;
  wire _29144_;
  wire _29145_;
  wire _29146_;
  wire _29147_;
  wire _29148_;
  wire _29149_;
  wire _29150_;
  wire _29151_;
  wire _29152_;
  wire _29153_;
  wire _29154_;
  wire _29155_;
  wire _29156_;
  wire _29157_;
  wire _29158_;
  wire _29159_;
  wire _29160_;
  wire _29161_;
  wire _29162_;
  wire _29163_;
  wire _29164_;
  wire _29165_;
  wire _29166_;
  wire _29167_;
  wire _29168_;
  wire _29169_;
  wire _29170_;
  wire _29171_;
  wire _29172_;
  wire _29173_;
  wire _29174_;
  wire _29175_;
  wire _29176_;
  wire _29177_;
  wire _29178_;
  wire _29179_;
  wire _29180_;
  wire _29181_;
  wire _29182_;
  wire _29183_;
  wire _29184_;
  wire _29185_;
  wire _29186_;
  wire _29187_;
  wire _29188_;
  wire _29189_;
  wire _29190_;
  wire _29191_;
  wire _29192_;
  wire _29193_;
  wire _29194_;
  wire _29195_;
  wire _29196_;
  wire _29197_;
  wire _29198_;
  wire _29199_;
  wire _29200_;
  wire _29201_;
  wire _29202_;
  wire _29203_;
  wire _29204_;
  wire _29205_;
  wire _29206_;
  wire _29207_;
  wire _29208_;
  wire _29209_;
  wire _29210_;
  wire _29211_;
  wire _29212_;
  wire _29213_;
  wire _29214_;
  wire _29215_;
  wire _29216_;
  wire _29217_;
  wire _29218_;
  wire _29219_;
  wire _29220_;
  wire _29221_;
  wire _29222_;
  wire _29223_;
  wire _29224_;
  wire _29225_;
  wire _29226_;
  wire _29227_;
  wire _29228_;
  wire _29229_;
  wire _29230_;
  wire _29231_;
  wire _29232_;
  wire _29233_;
  wire _29234_;
  wire _29235_;
  wire _29236_;
  wire _29237_;
  wire _29238_;
  wire _29239_;
  wire _29240_;
  wire _29241_;
  wire _29242_;
  wire _29243_;
  wire _29244_;
  wire _29245_;
  wire _29246_;
  wire _29247_;
  wire _29248_;
  wire _29249_;
  wire _29250_;
  wire _29251_;
  wire _29252_;
  wire _29253_;
  wire _29254_;
  wire _29255_;
  wire _29256_;
  wire _29257_;
  wire _29258_;
  wire _29259_;
  wire _29260_;
  wire _29261_;
  wire _29262_;
  wire _29263_;
  wire _29264_;
  wire _29265_;
  wire _29266_;
  wire _29267_;
  wire _29268_;
  wire _29269_;
  wire _29270_;
  wire _29271_;
  wire _29272_;
  wire _29273_;
  wire _29274_;
  wire _29275_;
  wire _29276_;
  wire _29277_;
  wire _29278_;
  wire _29279_;
  wire _29280_;
  wire _29281_;
  wire _29282_;
  wire _29283_;
  wire _29284_;
  wire _29285_;
  wire _29286_;
  wire _29287_;
  wire _29288_;
  wire _29289_;
  wire _29290_;
  wire _29291_;
  wire _29292_;
  wire _29293_;
  wire _29294_;
  wire _29295_;
  wire _29296_;
  wire _29297_;
  wire _29298_;
  wire _29299_;
  wire _29300_;
  wire _29301_;
  wire _29302_;
  wire _29303_;
  wire _29304_;
  wire _29305_;
  wire _29306_;
  wire _29307_;
  wire _29308_;
  wire _29309_;
  wire _29310_;
  wire _29311_;
  wire _29312_;
  wire _29313_;
  wire _29314_;
  wire _29315_;
  wire _29316_;
  wire _29317_;
  wire _29318_;
  wire _29319_;
  wire _29320_;
  wire _29321_;
  wire _29322_;
  wire _29323_;
  wire _29324_;
  wire _29325_;
  wire _29326_;
  wire _29327_;
  wire _29328_;
  wire _29329_;
  wire _29330_;
  wire _29331_;
  wire _29332_;
  wire _29333_;
  wire _29334_;
  wire _29335_;
  wire _29336_;
  wire _29337_;
  wire _29338_;
  wire _29339_;
  wire _29340_;
  wire _29341_;
  wire _29342_;
  wire _29343_;
  wire _29344_;
  wire _29345_;
  wire _29346_;
  wire _29347_;
  wire _29348_;
  wire _29349_;
  wire _29350_;
  wire _29351_;
  wire _29352_;
  wire _29353_;
  wire _29354_;
  wire _29355_;
  wire _29356_;
  wire _29357_;
  wire _29358_;
  wire _29359_;
  wire _29360_;
  wire _29361_;
  wire _29362_;
  wire _29363_;
  wire _29364_;
  wire _29365_;
  wire _29366_;
  wire _29367_;
  wire _29368_;
  wire _29369_;
  wire _29370_;
  wire _29371_;
  wire _29372_;
  wire _29373_;
  wire _29374_;
  wire _29375_;
  wire _29376_;
  wire _29377_;
  wire _29378_;
  wire _29379_;
  wire _29380_;
  wire _29381_;
  wire _29382_;
  wire _29383_;
  wire _29384_;
  wire _29385_;
  wire _29386_;
  wire _29387_;
  wire _29388_;
  wire _29389_;
  wire _29390_;
  wire _29391_;
  wire _29392_;
  wire _29393_;
  wire _29394_;
  wire _29395_;
  wire _29396_;
  wire _29397_;
  wire _29398_;
  wire _29399_;
  wire _29400_;
  wire _29401_;
  wire _29402_;
  wire _29403_;
  wire _29404_;
  wire _29405_;
  wire _29406_;
  wire _29407_;
  wire _29408_;
  wire _29409_;
  wire _29410_;
  wire _29411_;
  wire _29412_;
  wire _29413_;
  wire _29414_;
  wire _29415_;
  wire _29416_;
  wire _29417_;
  wire _29418_;
  wire _29419_;
  wire _29420_;
  wire _29421_;
  wire _29422_;
  wire _29423_;
  wire _29424_;
  wire _29425_;
  wire _29426_;
  wire _29427_;
  wire _29428_;
  wire _29429_;
  wire _29430_;
  wire _29431_;
  wire _29432_;
  wire _29433_;
  wire _29434_;
  wire _29435_;
  wire _29436_;
  wire _29437_;
  wire _29438_;
  wire _29439_;
  wire _29440_;
  wire _29441_;
  wire _29442_;
  wire _29443_;
  wire _29444_;
  wire _29445_;
  wire _29446_;
  wire _29447_;
  wire _29448_;
  wire _29449_;
  wire _29450_;
  wire _29451_;
  wire _29452_;
  wire _29453_;
  wire _29454_;
  wire _29455_;
  wire _29456_;
  wire _29457_;
  wire _29458_;
  wire _29459_;
  wire _29460_;
  wire _29461_;
  wire _29462_;
  wire _29463_;
  wire _29464_;
  wire _29465_;
  wire _29466_;
  wire _29467_;
  wire _29468_;
  wire _29469_;
  wire _29470_;
  wire _29471_;
  wire _29472_;
  wire _29473_;
  wire _29474_;
  wire _29475_;
  wire _29476_;
  wire _29477_;
  wire _29478_;
  wire _29479_;
  wire _29480_;
  wire _29481_;
  wire _29482_;
  wire _29483_;
  wire _29484_;
  wire _29485_;
  wire _29486_;
  wire _29487_;
  wire _29488_;
  wire _29489_;
  wire _29490_;
  wire _29491_;
  wire _29492_;
  wire _29493_;
  wire _29494_;
  wire _29495_;
  wire _29496_;
  wire _29497_;
  wire _29498_;
  wire _29499_;
  wire _29500_;
  wire _29501_;
  wire _29502_;
  wire _29503_;
  wire _29504_;
  wire _29505_;
  wire _29506_;
  wire _29507_;
  wire _29508_;
  wire _29509_;
  wire _29510_;
  wire _29511_;
  wire _29512_;
  wire _29513_;
  wire _29514_;
  wire _29515_;
  wire _29516_;
  wire _29517_;
  wire _29518_;
  wire _29519_;
  wire _29520_;
  wire _29521_;
  wire _29522_;
  wire _29523_;
  wire _29524_;
  wire _29525_;
  wire _29526_;
  wire _29527_;
  wire _29528_;
  wire _29529_;
  wire _29530_;
  wire _29531_;
  wire _29532_;
  wire _29533_;
  wire _29534_;
  wire _29535_;
  wire _29536_;
  wire _29537_;
  wire _29538_;
  wire _29539_;
  wire _29540_;
  wire _29541_;
  wire _29542_;
  wire _29543_;
  wire _29544_;
  wire _29545_;
  wire _29546_;
  wire _29547_;
  wire _29548_;
  wire _29549_;
  wire _29550_;
  wire _29551_;
  wire _29552_;
  wire _29553_;
  wire _29554_;
  wire _29555_;
  wire _29556_;
  wire _29557_;
  wire _29558_;
  wire _29559_;
  wire _29560_;
  wire _29561_;
  wire _29562_;
  wire _29563_;
  wire _29564_;
  wire _29565_;
  wire _29566_;
  wire _29567_;
  wire _29568_;
  wire _29569_;
  wire _29570_;
  wire _29571_;
  wire _29572_;
  wire _29573_;
  wire _29574_;
  wire _29575_;
  wire _29576_;
  wire _29577_;
  wire _29578_;
  wire _29579_;
  wire _29580_;
  wire _29581_;
  wire _29582_;
  wire _29583_;
  wire _29584_;
  wire _29585_;
  wire _29586_;
  wire _29587_;
  wire _29588_;
  wire _29589_;
  wire _29590_;
  wire _29591_;
  wire _29592_;
  wire _29593_;
  wire _29594_;
  wire _29595_;
  wire _29596_;
  wire _29597_;
  wire _29598_;
  wire _29599_;
  wire _29600_;
  wire _29601_;
  wire _29602_;
  wire _29603_;
  wire _29604_;
  wire _29605_;
  wire _29606_;
  wire _29607_;
  wire _29608_;
  wire _29609_;
  wire _29610_;
  wire _29611_;
  wire _29612_;
  wire _29613_;
  wire _29614_;
  wire _29615_;
  wire _29616_;
  wire _29617_;
  wire _29618_;
  wire _29619_;
  wire _29620_;
  wire _29621_;
  wire _29622_;
  wire _29623_;
  wire _29624_;
  wire _29625_;
  wire _29626_;
  wire _29627_;
  wire _29628_;
  wire _29629_;
  wire _29630_;
  wire _29631_;
  wire _29632_;
  wire _29633_;
  wire _29634_;
  wire _29635_;
  wire _29636_;
  wire _29637_;
  wire _29638_;
  wire _29639_;
  wire _29640_;
  wire _29641_;
  wire _29642_;
  wire _29643_;
  wire _29644_;
  wire _29645_;
  wire _29646_;
  wire _29647_;
  wire _29648_;
  wire _29649_;
  wire _29650_;
  wire _29651_;
  wire _29652_;
  wire _29653_;
  wire _29654_;
  wire _29655_;
  wire _29656_;
  wire _29657_;
  wire _29658_;
  wire _29659_;
  wire _29660_;
  wire _29661_;
  wire _29662_;
  wire _29663_;
  wire _29664_;
  wire _29665_;
  wire _29666_;
  wire _29667_;
  wire _29668_;
  wire _29669_;
  wire _29670_;
  wire _29671_;
  wire _29672_;
  wire _29673_;
  wire _29674_;
  wire _29675_;
  wire _29676_;
  wire _29677_;
  wire _29678_;
  wire _29679_;
  wire _29680_;
  wire _29681_;
  wire _29682_;
  wire _29683_;
  wire _29684_;
  wire _29685_;
  wire _29686_;
  wire _29687_;
  wire _29688_;
  wire _29689_;
  wire _29690_;
  wire _29691_;
  wire _29692_;
  wire _29693_;
  wire _29694_;
  wire _29695_;
  wire _29696_;
  wire _29697_;
  wire _29698_;
  wire _29699_;
  wire _29700_;
  wire _29701_;
  wire _29702_;
  wire _29703_;
  wire _29704_;
  wire _29705_;
  wire _29706_;
  wire _29707_;
  wire _29708_;
  wire _29709_;
  wire _29710_;
  wire _29711_;
  wire _29712_;
  wire _29713_;
  wire _29714_;
  wire _29715_;
  wire _29716_;
  wire _29717_;
  wire _29718_;
  wire _29719_;
  wire _29720_;
  wire _29721_;
  wire _29722_;
  wire _29723_;
  wire _29724_;
  wire _29725_;
  wire _29726_;
  wire _29727_;
  wire _29728_;
  wire _29729_;
  wire _29730_;
  wire _29731_;
  wire _29732_;
  wire _29733_;
  wire _29734_;
  wire _29735_;
  wire _29736_;
  wire _29737_;
  wire _29738_;
  wire _29739_;
  wire _29740_;
  wire _29741_;
  wire _29742_;
  wire _29743_;
  wire _29744_;
  wire _29745_;
  wire _29746_;
  wire _29747_;
  wire _29748_;
  wire _29749_;
  wire _29750_;
  wire _29751_;
  wire _29752_;
  wire _29753_;
  wire _29754_;
  wire _29755_;
  wire _29756_;
  wire _29757_;
  wire _29758_;
  wire _29759_;
  wire _29760_;
  wire _29761_;
  wire _29762_;
  wire _29763_;
  wire _29764_;
  wire _29765_;
  wire _29766_;
  wire _29767_;
  wire _29768_;
  wire _29769_;
  wire _29770_;
  wire _29771_;
  wire _29772_;
  wire _29773_;
  wire _29774_;
  wire _29775_;
  wire _29776_;
  wire _29777_;
  wire _29778_;
  wire _29779_;
  wire _29780_;
  wire _29781_;
  wire _29782_;
  wire _29783_;
  wire _29784_;
  wire _29785_;
  wire _29786_;
  wire _29787_;
  wire _29788_;
  wire _29789_;
  wire _29790_;
  wire _29791_;
  wire _29792_;
  wire _29793_;
  wire _29794_;
  wire _29795_;
  wire _29796_;
  wire _29797_;
  wire _29798_;
  wire _29799_;
  wire _29800_;
  wire _29801_;
  wire _29802_;
  wire _29803_;
  wire _29804_;
  wire _29805_;
  wire _29806_;
  wire _29807_;
  wire _29808_;
  wire _29809_;
  wire _29810_;
  wire _29811_;
  wire _29812_;
  wire _29813_;
  wire _29814_;
  wire _29815_;
  wire _29816_;
  wire _29817_;
  wire _29818_;
  wire _29819_;
  wire _29820_;
  wire _29821_;
  wire _29822_;
  wire _29823_;
  wire _29824_;
  wire _29825_;
  wire _29826_;
  wire _29827_;
  wire _29828_;
  wire _29829_;
  wire _29830_;
  wire _29831_;
  wire _29832_;
  wire _29833_;
  wire _29834_;
  wire _29835_;
  wire _29836_;
  wire _29837_;
  wire _29838_;
  wire _29839_;
  wire _29840_;
  wire _29841_;
  wire _29842_;
  wire _29843_;
  wire _29844_;
  wire _29845_;
  wire _29846_;
  wire _29847_;
  wire _29848_;
  wire _29849_;
  wire _29850_;
  wire _29851_;
  wire _29852_;
  wire _29853_;
  wire _29854_;
  wire _29855_;
  wire _29856_;
  wire _29857_;
  wire _29858_;
  wire _29859_;
  wire _29860_;
  wire _29861_;
  wire _29862_;
  wire _29863_;
  wire _29864_;
  wire _29865_;
  wire _29866_;
  wire _29867_;
  wire _29868_;
  wire _29869_;
  wire _29870_;
  wire _29871_;
  wire _29872_;
  wire _29873_;
  wire _29874_;
  wire _29875_;
  wire _29876_;
  wire _29877_;
  wire _29878_;
  wire _29879_;
  wire _29880_;
  wire _29881_;
  wire _29882_;
  wire _29883_;
  wire _29884_;
  wire _29885_;
  wire _29886_;
  wire _29887_;
  wire _29888_;
  wire _29889_;
  wire _29890_;
  wire _29891_;
  wire _29892_;
  wire _29893_;
  wire _29894_;
  wire _29895_;
  wire _29896_;
  wire _29897_;
  wire _29898_;
  wire _29899_;
  wire _29900_;
  wire _29901_;
  wire _29902_;
  wire _29903_;
  wire _29904_;
  wire _29905_;
  wire _29906_;
  wire _29907_;
  wire _29908_;
  wire _29909_;
  wire _29910_;
  wire _29911_;
  wire _29912_;
  wire _29913_;
  wire _29914_;
  wire _29915_;
  wire _29916_;
  wire _29917_;
  wire _29918_;
  wire _29919_;
  wire _29920_;
  wire _29921_;
  wire _29922_;
  wire _29923_;
  wire _29924_;
  wire _29925_;
  wire _29926_;
  wire _29927_;
  wire _29928_;
  wire _29929_;
  wire _29930_;
  wire _29931_;
  wire _29932_;
  wire _29933_;
  wire _29934_;
  wire _29935_;
  wire _29936_;
  wire _29937_;
  wire _29938_;
  wire _29939_;
  wire _29940_;
  wire _29941_;
  wire _29942_;
  wire _29943_;
  wire _29944_;
  wire _29945_;
  wire _29946_;
  wire _29947_;
  wire _29948_;
  wire _29949_;
  wire _29950_;
  wire _29951_;
  wire _29952_;
  wire _29953_;
  wire _29954_;
  wire _29955_;
  wire _29956_;
  wire _29957_;
  wire _29958_;
  wire _29959_;
  wire _29960_;
  wire _29961_;
  wire _29962_;
  wire _29963_;
  wire _29964_;
  wire _29965_;
  wire _29966_;
  wire _29967_;
  wire _29968_;
  wire _29969_;
  wire _29970_;
  wire _29971_;
  wire _29972_;
  wire _29973_;
  wire _29974_;
  wire _29975_;
  wire _29976_;
  wire _29977_;
  wire _29978_;
  wire _29979_;
  wire _29980_;
  wire _29981_;
  wire _29982_;
  wire _29983_;
  wire _29984_;
  wire _29985_;
  wire _29986_;
  wire _29987_;
  wire _29988_;
  wire _29989_;
  wire _29990_;
  wire _29991_;
  wire _29992_;
  wire _29993_;
  wire _29994_;
  wire _29995_;
  wire _29996_;
  wire _29997_;
  wire _29998_;
  wire _29999_;
  wire _30000_;
  wire _30001_;
  wire _30002_;
  wire _30003_;
  wire _30004_;
  wire _30005_;
  wire _30006_;
  wire _30007_;
  wire _30008_;
  wire _30009_;
  wire _30010_;
  wire _30011_;
  wire _30012_;
  wire _30013_;
  wire _30014_;
  wire _30015_;
  wire _30016_;
  wire _30017_;
  wire _30018_;
  wire _30019_;
  wire _30020_;
  wire _30021_;
  wire _30022_;
  wire _30023_;
  wire _30024_;
  wire _30025_;
  wire _30026_;
  wire _30027_;
  wire _30028_;
  wire _30029_;
  wire _30030_;
  wire _30031_;
  wire _30032_;
  wire _30033_;
  wire _30034_;
  wire _30035_;
  wire _30036_;
  wire _30037_;
  wire _30038_;
  wire _30039_;
  wire _30040_;
  wire _30041_;
  wire _30042_;
  wire _30043_;
  wire _30044_;
  wire _30045_;
  wire _30046_;
  wire _30047_;
  wire _30048_;
  wire _30049_;
  wire _30050_;
  wire _30051_;
  wire _30052_;
  wire _30053_;
  wire _30054_;
  wire _30055_;
  wire _30056_;
  wire _30057_;
  wire _30058_;
  wire _30059_;
  wire _30060_;
  wire _30061_;
  wire _30062_;
  wire _30063_;
  wire _30064_;
  wire _30065_;
  wire _30066_;
  wire _30067_;
  wire _30068_;
  wire _30069_;
  wire _30070_;
  wire _30071_;
  wire _30072_;
  wire _30073_;
  wire _30074_;
  wire _30075_;
  wire _30076_;
  wire _30077_;
  wire _30078_;
  wire _30079_;
  wire _30080_;
  wire _30081_;
  wire _30082_;
  wire _30083_;
  wire _30084_;
  wire _30085_;
  wire _30086_;
  wire _30087_;
  wire _30088_;
  wire _30089_;
  wire _30090_;
  wire _30091_;
  wire _30092_;
  wire _30093_;
  wire _30094_;
  wire _30095_;
  wire _30096_;
  wire _30097_;
  wire _30098_;
  wire _30099_;
  wire _30100_;
  wire _30101_;
  wire _30102_;
  wire _30103_;
  wire _30104_;
  wire _30105_;
  wire _30106_;
  wire _30107_;
  wire _30108_;
  wire _30109_;
  wire _30110_;
  wire _30111_;
  wire _30112_;
  wire _30113_;
  wire _30114_;
  wire _30115_;
  wire _30116_;
  wire _30117_;
  wire _30118_;
  wire _30119_;
  wire _30120_;
  wire _30121_;
  wire _30122_;
  wire _30123_;
  wire _30124_;
  wire _30125_;
  wire _30126_;
  wire _30127_;
  wire _30128_;
  wire _30129_;
  wire _30130_;
  wire _30131_;
  wire _30132_;
  wire _30133_;
  wire _30134_;
  wire _30135_;
  wire _30136_;
  wire _30137_;
  wire _30138_;
  wire _30139_;
  wire _30140_;
  wire _30141_;
  wire _30142_;
  wire _30143_;
  wire _30144_;
  wire _30145_;
  wire _30146_;
  wire _30147_;
  wire _30148_;
  wire _30149_;
  wire _30150_;
  wire _30151_;
  wire _30152_;
  wire _30153_;
  wire _30154_;
  wire _30155_;
  wire _30156_;
  wire _30157_;
  wire _30158_;
  wire _30159_;
  wire _30160_;
  wire _30161_;
  wire _30162_;
  wire _30163_;
  wire _30164_;
  wire _30165_;
  wire _30166_;
  wire _30167_;
  wire _30168_;
  wire _30169_;
  wire _30170_;
  wire _30171_;
  wire _30172_;
  wire _30173_;
  wire _30174_;
  wire _30175_;
  wire _30176_;
  wire _30177_;
  wire _30178_;
  wire _30179_;
  wire _30180_;
  wire _30181_;
  wire _30182_;
  wire _30183_;
  wire _30184_;
  wire _30185_;
  wire _30186_;
  wire _30187_;
  wire _30188_;
  wire _30189_;
  wire _30190_;
  wire _30191_;
  wire _30192_;
  wire _30193_;
  wire _30194_;
  wire _30195_;
  wire _30196_;
  wire _30197_;
  wire _30198_;
  wire _30199_;
  wire _30200_;
  wire _30201_;
  wire _30202_;
  wire _30203_;
  wire _30204_;
  wire _30205_;
  wire _30206_;
  wire _30207_;
  wire _30208_;
  wire _30209_;
  wire _30210_;
  wire _30211_;
  wire _30212_;
  wire _30213_;
  wire _30214_;
  wire _30215_;
  wire _30216_;
  wire _30217_;
  wire _30218_;
  wire _30219_;
  wire _30220_;
  wire _30221_;
  wire _30222_;
  wire _30223_;
  wire _30224_;
  wire _30225_;
  wire _30226_;
  wire _30227_;
  wire _30228_;
  wire _30229_;
  wire _30230_;
  wire _30231_;
  wire _30232_;
  wire _30233_;
  wire _30234_;
  wire _30235_;
  wire _30236_;
  wire _30237_;
  wire _30238_;
  wire _30239_;
  wire _30240_;
  wire _30241_;
  wire _30242_;
  wire _30243_;
  wire _30244_;
  wire _30245_;
  wire _30246_;
  wire _30247_;
  wire _30248_;
  wire _30249_;
  wire _30250_;
  wire _30251_;
  wire _30252_;
  wire _30253_;
  wire _30254_;
  wire _30255_;
  wire _30256_;
  wire _30257_;
  wire _30258_;
  wire _30259_;
  wire _30260_;
  wire _30261_;
  wire _30262_;
  wire _30263_;
  wire _30264_;
  wire _30265_;
  wire _30266_;
  wire _30267_;
  wire _30268_;
  wire _30269_;
  wire _30270_;
  wire _30271_;
  wire _30272_;
  wire _30273_;
  wire _30274_;
  wire _30275_;
  wire _30276_;
  wire _30277_;
  wire _30278_;
  wire _30279_;
  wire _30280_;
  wire _30281_;
  wire _30282_;
  wire _30283_;
  wire _30284_;
  wire _30285_;
  wire _30286_;
  wire _30287_;
  wire _30288_;
  wire _30289_;
  wire _30290_;
  wire _30291_;
  wire _30292_;
  wire _30293_;
  wire _30294_;
  wire _30295_;
  wire _30296_;
  wire _30297_;
  wire _30298_;
  wire _30299_;
  wire _30300_;
  wire _30301_;
  wire _30302_;
  wire _30303_;
  wire _30304_;
  wire _30305_;
  wire _30306_;
  wire _30307_;
  wire _30308_;
  wire _30309_;
  wire _30310_;
  wire _30311_;
  wire _30312_;
  wire _30313_;
  wire _30314_;
  wire _30315_;
  wire _30316_;
  wire _30317_;
  wire _30318_;
  wire _30319_;
  wire _30320_;
  wire _30321_;
  wire _30322_;
  wire _30323_;
  wire _30324_;
  wire _30325_;
  wire _30326_;
  wire _30327_;
  wire _30328_;
  wire _30329_;
  wire _30330_;
  wire _30331_;
  wire _30332_;
  wire _30333_;
  wire _30334_;
  wire _30335_;
  wire _30336_;
  wire _30337_;
  wire _30338_;
  wire _30339_;
  wire _30340_;
  wire _30341_;
  wire _30342_;
  wire _30343_;
  wire _30344_;
  wire _30345_;
  wire _30346_;
  wire _30347_;
  wire _30348_;
  wire _30349_;
  wire _30350_;
  wire _30351_;
  wire _30352_;
  wire _30353_;
  wire _30354_;
  wire _30355_;
  wire _30356_;
  wire _30357_;
  wire _30358_;
  wire _30359_;
  wire _30360_;
  wire _30361_;
  wire _30362_;
  wire _30363_;
  wire _30364_;
  wire _30365_;
  wire _30366_;
  wire _30367_;
  wire _30368_;
  wire _30369_;
  wire _30370_;
  wire _30371_;
  wire _30372_;
  wire _30373_;
  wire _30374_;
  wire _30375_;
  wire _30376_;
  wire _30377_;
  wire _30378_;
  wire _30379_;
  wire _30380_;
  wire _30381_;
  wire _30382_;
  wire _30383_;
  wire _30384_;
  wire _30385_;
  wire _30386_;
  wire _30387_;
  wire _30388_;
  wire _30389_;
  wire _30390_;
  wire _30391_;
  wire _30392_;
  wire _30393_;
  wire _30394_;
  wire _30395_;
  wire _30396_;
  wire _30397_;
  wire _30398_;
  wire _30399_;
  wire _30400_;
  wire _30401_;
  wire _30402_;
  wire _30403_;
  wire _30404_;
  wire _30405_;
  wire _30406_;
  wire _30407_;
  wire _30408_;
  wire _30409_;
  wire _30410_;
  wire _30411_;
  wire _30412_;
  wire _30413_;
  wire _30414_;
  wire _30415_;
  wire _30416_;
  wire _30417_;
  wire _30418_;
  wire _30419_;
  wire _30420_;
  wire _30421_;
  wire _30422_;
  wire _30423_;
  wire _30424_;
  wire _30425_;
  wire _30426_;
  wire _30427_;
  wire _30428_;
  wire _30429_;
  wire _30430_;
  wire _30431_;
  wire _30432_;
  wire _30433_;
  wire _30434_;
  wire _30435_;
  wire _30436_;
  wire _30437_;
  wire _30438_;
  wire _30439_;
  wire _30440_;
  wire _30441_;
  wire _30442_;
  wire _30443_;
  wire _30444_;
  wire _30445_;
  wire _30446_;
  wire _30447_;
  wire _30448_;
  wire _30449_;
  wire _30450_;
  wire _30451_;
  wire _30452_;
  wire _30453_;
  wire _30454_;
  wire _30455_;
  wire _30456_;
  wire _30457_;
  wire _30458_;
  wire _30459_;
  wire _30460_;
  wire _30461_;
  wire _30462_;
  wire _30463_;
  wire _30464_;
  wire _30465_;
  wire _30466_;
  wire _30467_;
  wire _30468_;
  wire _30469_;
  wire _30470_;
  wire _30471_;
  wire _30472_;
  wire _30473_;
  wire _30474_;
  wire _30475_;
  wire _30476_;
  wire _30477_;
  wire _30478_;
  wire _30479_;
  wire _30480_;
  wire _30481_;
  wire _30482_;
  wire _30483_;
  wire _30484_;
  wire _30485_;
  wire _30486_;
  wire _30487_;
  wire _30488_;
  wire _30489_;
  wire _30490_;
  wire _30491_;
  wire _30492_;
  wire _30493_;
  wire _30494_;
  wire _30495_;
  wire _30496_;
  wire _30497_;
  wire _30498_;
  wire _30499_;
  wire _30500_;
  wire _30501_;
  wire _30502_;
  wire _30503_;
  wire _30504_;
  wire _30505_;
  wire _30506_;
  wire _30507_;
  wire _30508_;
  wire _30509_;
  wire _30510_;
  wire _30511_;
  wire _30512_;
  wire _30513_;
  wire _30514_;
  wire _30515_;
  wire _30516_;
  wire _30517_;
  wire _30518_;
  wire _30519_;
  wire _30520_;
  wire _30521_;
  wire _30522_;
  wire _30523_;
  wire _30524_;
  wire _30525_;
  wire _30526_;
  wire _30527_;
  wire _30528_;
  wire _30529_;
  wire _30530_;
  wire _30531_;
  wire _30532_;
  wire _30533_;
  wire _30534_;
  wire _30535_;
  wire _30536_;
  wire _30537_;
  wire _30538_;
  wire _30539_;
  wire _30540_;
  wire _30541_;
  wire _30542_;
  wire _30543_;
  wire _30544_;
  wire _30545_;
  wire _30546_;
  wire _30547_;
  wire _30548_;
  wire _30549_;
  wire _30550_;
  wire _30551_;
  wire _30552_;
  wire _30553_;
  wire _30554_;
  wire _30555_;
  wire _30556_;
  wire _30557_;
  wire _30558_;
  wire _30559_;
  wire _30560_;
  wire _30561_;
  wire _30562_;
  wire _30563_;
  wire _30564_;
  wire _30565_;
  wire _30566_;
  wire _30567_;
  wire _30568_;
  wire _30569_;
  wire _30570_;
  wire _30571_;
  wire _30572_;
  wire _30573_;
  wire _30574_;
  wire _30575_;
  wire _30576_;
  wire _30577_;
  wire _30578_;
  wire _30579_;
  wire _30580_;
  wire _30581_;
  wire _30582_;
  wire _30583_;
  wire _30584_;
  wire _30585_;
  wire _30586_;
  wire _30587_;
  wire _30588_;
  wire _30589_;
  wire _30590_;
  wire _30591_;
  wire _30592_;
  wire _30593_;
  wire _30594_;
  wire _30595_;
  wire _30596_;
  wire _30597_;
  wire _30598_;
  wire _30599_;
  wire _30600_;
  wire _30601_;
  wire _30602_;
  wire _30603_;
  wire _30604_;
  wire _30605_;
  wire _30606_;
  wire _30607_;
  wire _30608_;
  wire _30609_;
  wire _30610_;
  wire _30611_;
  wire _30612_;
  wire _30613_;
  wire _30614_;
  wire _30615_;
  wire _30616_;
  wire _30617_;
  wire _30618_;
  wire _30619_;
  wire _30620_;
  wire _30621_;
  wire _30622_;
  wire _30623_;
  wire _30624_;
  wire _30625_;
  wire _30626_;
  wire _30627_;
  wire _30628_;
  wire _30629_;
  wire _30630_;
  wire _30631_;
  wire _30632_;
  wire _30633_;
  wire _30634_;
  wire _30635_;
  wire _30636_;
  wire _30637_;
  wire _30638_;
  wire _30639_;
  wire _30640_;
  wire _30641_;
  wire _30642_;
  wire _30643_;
  wire _30644_;
  wire _30645_;
  wire _30646_;
  wire _30647_;
  wire _30648_;
  wire _30649_;
  wire _30650_;
  wire _30651_;
  wire _30652_;
  wire _30653_;
  wire _30654_;
  wire _30655_;
  wire _30656_;
  wire _30657_;
  wire _30658_;
  wire _30659_;
  wire _30660_;
  wire _30661_;
  wire _30662_;
  wire _30663_;
  wire _30664_;
  wire _30665_;
  wire _30666_;
  wire _30667_;
  wire _30668_;
  wire _30669_;
  wire _30670_;
  wire _30671_;
  wire _30672_;
  wire _30673_;
  wire _30674_;
  wire _30675_;
  wire _30676_;
  wire _30677_;
  wire _30678_;
  wire _30679_;
  wire _30680_;
  wire _30681_;
  wire _30682_;
  wire _30683_;
  wire _30684_;
  wire _30685_;
  wire _30686_;
  wire _30687_;
  wire _30688_;
  wire _30689_;
  wire _30690_;
  wire _30691_;
  wire _30692_;
  wire _30693_;
  wire _30694_;
  wire _30695_;
  wire _30696_;
  wire _30697_;
  wire _30698_;
  wire _30699_;
  wire _30700_;
  wire _30701_;
  wire _30702_;
  wire _30703_;
  wire _30704_;
  wire _30705_;
  wire _30706_;
  wire _30707_;
  wire _30708_;
  wire _30709_;
  wire _30710_;
  wire _30711_;
  wire _30712_;
  wire _30713_;
  wire _30714_;
  wire _30715_;
  wire _30716_;
  wire _30717_;
  wire _30718_;
  wire _30719_;
  wire _30720_;
  wire _30721_;
  wire _30722_;
  wire _30723_;
  wire _30724_;
  wire _30725_;
  wire _30726_;
  wire _30727_;
  wire _30728_;
  wire _30729_;
  wire _30730_;
  wire _30731_;
  wire _30732_;
  wire _30733_;
  wire _30734_;
  wire _30735_;
  wire _30736_;
  wire _30737_;
  wire _30738_;
  wire _30739_;
  wire _30740_;
  wire _30741_;
  wire _30742_;
  wire _30743_;
  wire _30744_;
  wire _30745_;
  wire _30746_;
  wire _30747_;
  wire _30748_;
  wire _30749_;
  wire _30750_;
  wire _30751_;
  wire _30752_;
  wire _30753_;
  wire _30754_;
  wire _30755_;
  wire _30756_;
  wire _30757_;
  wire _30758_;
  wire _30759_;
  wire _30760_;
  wire _30761_;
  wire _30762_;
  wire _30763_;
  wire _30764_;
  wire _30765_;
  wire _30766_;
  wire _30767_;
  wire _30768_;
  wire _30769_;
  wire _30770_;
  wire _30771_;
  wire _30772_;
  wire _30773_;
  wire _30774_;
  wire _30775_;
  wire _30776_;
  wire _30777_;
  wire _30778_;
  wire _30779_;
  wire _30780_;
  wire _30781_;
  wire _30782_;
  wire _30783_;
  wire _30784_;
  wire _30785_;
  wire _30786_;
  wire _30787_;
  wire _30788_;
  wire _30789_;
  wire _30790_;
  wire _30791_;
  wire _30792_;
  wire _30793_;
  wire _30794_;
  wire _30795_;
  wire _30796_;
  wire _30797_;
  wire _30798_;
  wire _30799_;
  wire _30800_;
  wire _30801_;
  wire _30802_;
  wire _30803_;
  wire _30804_;
  wire _30805_;
  wire _30806_;
  wire _30807_;
  wire _30808_;
  wire _30809_;
  wire _30810_;
  wire _30811_;
  wire _30812_;
  wire _30813_;
  wire _30814_;
  wire _30815_;
  wire _30816_;
  wire _30817_;
  wire _30818_;
  wire _30819_;
  wire _30820_;
  wire _30821_;
  wire _30822_;
  wire _30823_;
  wire _30824_;
  wire _30825_;
  wire _30826_;
  wire _30827_;
  wire _30828_;
  wire _30829_;
  wire _30830_;
  wire _30831_;
  wire _30832_;
  wire _30833_;
  wire _30834_;
  wire _30835_;
  wire _30836_;
  wire _30837_;
  wire _30838_;
  wire _30839_;
  wire _30840_;
  wire _30841_;
  wire _30842_;
  wire _30843_;
  wire _30844_;
  wire _30845_;
  wire _30846_;
  wire _30847_;
  wire _30848_;
  wire _30849_;
  wire _30850_;
  wire _30851_;
  wire _30852_;
  wire _30853_;
  wire _30854_;
  wire _30855_;
  wire _30856_;
  wire _30857_;
  wire _30858_;
  wire _30859_;
  wire _30860_;
  wire _30861_;
  wire _30862_;
  wire _30863_;
  wire _30864_;
  wire _30865_;
  wire _30866_;
  wire _30867_;
  wire _30868_;
  wire _30869_;
  wire _30870_;
  wire _30871_;
  wire _30872_;
  wire _30873_;
  wire _30874_;
  wire _30875_;
  wire _30876_;
  wire _30877_;
  wire _30878_;
  wire _30879_;
  wire _30880_;
  wire _30881_;
  wire _30882_;
  wire _30883_;
  wire _30884_;
  wire _30885_;
  wire _30886_;
  wire _30887_;
  wire _30888_;
  wire _30889_;
  wire _30890_;
  wire _30891_;
  wire _30892_;
  wire _30893_;
  wire _30894_;
  wire _30895_;
  wire _30896_;
  wire _30897_;
  wire _30898_;
  wire _30899_;
  wire _30900_;
  wire _30901_;
  wire _30902_;
  wire _30903_;
  wire _30904_;
  wire _30905_;
  wire _30906_;
  wire _30907_;
  wire _30908_;
  wire _30909_;
  wire _30910_;
  wire _30911_;
  wire _30912_;
  wire _30913_;
  wire _30914_;
  wire _30915_;
  wire _30916_;
  wire _30917_;
  wire _30918_;
  wire _30919_;
  wire _30920_;
  wire _30921_;
  wire _30922_;
  wire _30923_;
  wire _30924_;
  wire _30925_;
  wire _30926_;
  wire _30927_;
  wire _30928_;
  wire _30929_;
  wire _30930_;
  wire _30931_;
  wire _30932_;
  wire _30933_;
  wire _30934_;
  wire _30935_;
  wire _30936_;
  wire _30937_;
  wire _30938_;
  wire _30939_;
  wire _30940_;
  wire _30941_;
  wire _30942_;
  wire _30943_;
  wire _30944_;
  wire _30945_;
  wire _30946_;
  wire _30947_;
  wire _30948_;
  wire _30949_;
  wire _30950_;
  wire _30951_;
  wire _30952_;
  wire _30953_;
  wire _30954_;
  wire _30955_;
  wire _30956_;
  wire _30957_;
  wire _30958_;
  wire _30959_;
  wire _30960_;
  wire _30961_;
  wire _30962_;
  wire _30963_;
  wire _30964_;
  wire _30965_;
  wire _30966_;
  wire _30967_;
  wire _30968_;
  wire _30969_;
  wire _30970_;
  wire _30971_;
  wire _30972_;
  wire _30973_;
  wire _30974_;
  wire _30975_;
  wire _30976_;
  wire _30977_;
  wire _30978_;
  wire _30979_;
  wire _30980_;
  wire _30981_;
  wire _30982_;
  wire _30983_;
  wire _30984_;
  wire _30985_;
  wire _30986_;
  wire _30987_;
  wire _30988_;
  wire _30989_;
  wire _30990_;
  wire _30991_;
  wire _30992_;
  wire _30993_;
  wire _30994_;
  wire _30995_;
  wire _30996_;
  wire _30997_;
  wire _30998_;
  wire _30999_;
  wire _31000_;
  wire _31001_;
  wire _31002_;
  wire _31003_;
  wire _31004_;
  wire _31005_;
  wire _31006_;
  wire _31007_;
  wire _31008_;
  wire _31009_;
  wire _31010_;
  wire _31011_;
  wire _31012_;
  wire _31013_;
  wire _31014_;
  wire _31015_;
  wire _31016_;
  wire _31017_;
  wire _31018_;
  wire _31019_;
  wire _31020_;
  wire _31021_;
  wire _31022_;
  wire _31023_;
  wire _31024_;
  wire _31025_;
  wire _31026_;
  wire _31027_;
  wire _31028_;
  wire _31029_;
  wire _31030_;
  wire _31031_;
  wire _31032_;
  wire _31033_;
  wire _31034_;
  wire _31035_;
  wire _31036_;
  wire _31037_;
  wire _31038_;
  wire _31039_;
  wire _31040_;
  wire _31041_;
  wire _31042_;
  wire _31043_;
  wire _31044_;
  wire _31045_;
  wire _31046_;
  wire _31047_;
  wire _31048_;
  wire _31049_;
  wire _31050_;
  wire _31051_;
  wire _31052_;
  wire _31053_;
  wire _31054_;
  wire _31055_;
  wire _31056_;
  wire _31057_;
  wire _31058_;
  wire _31059_;
  wire _31060_;
  wire _31061_;
  wire _31062_;
  wire _31063_;
  wire _31064_;
  wire _31065_;
  wire _31066_;
  wire _31067_;
  wire _31068_;
  wire _31069_;
  wire _31070_;
  wire _31071_;
  wire _31072_;
  wire _31073_;
  wire _31074_;
  wire _31075_;
  wire _31076_;
  wire _31077_;
  wire _31078_;
  wire _31079_;
  wire _31080_;
  wire _31081_;
  wire _31082_;
  wire _31083_;
  wire _31084_;
  wire _31085_;
  wire _31086_;
  wire _31087_;
  wire _31088_;
  wire _31089_;
  wire _31090_;
  wire _31091_;
  wire _31092_;
  wire _31093_;
  wire _31094_;
  wire _31095_;
  wire _31096_;
  wire _31097_;
  wire _31098_;
  wire _31099_;
  wire _31100_;
  wire _31101_;
  wire _31102_;
  wire _31103_;
  wire _31104_;
  wire _31105_;
  wire _31106_;
  wire _31107_;
  wire _31108_;
  wire _31109_;
  wire _31110_;
  wire _31111_;
  wire _31112_;
  wire _31113_;
  wire _31114_;
  wire _31115_;
  wire _31116_;
  wire _31117_;
  wire _31118_;
  wire _31119_;
  wire _31120_;
  wire _31121_;
  wire _31122_;
  wire _31123_;
  wire _31124_;
  wire _31125_;
  wire _31126_;
  wire _31127_;
  wire _31128_;
  wire _31129_;
  wire _31130_;
  wire _31131_;
  wire _31132_;
  wire _31133_;
  wire _31134_;
  wire _31135_;
  wire _31136_;
  wire _31137_;
  wire _31138_;
  wire _31139_;
  wire _31140_;
  wire _31141_;
  wire _31142_;
  wire _31143_;
  wire _31144_;
  wire _31145_;
  wire _31146_;
  wire _31147_;
  wire _31148_;
  wire _31149_;
  wire _31150_;
  wire _31151_;
  wire _31152_;
  wire _31153_;
  wire _31154_;
  wire _31155_;
  wire _31156_;
  wire _31157_;
  wire _31158_;
  wire _31159_;
  wire _31160_;
  wire _31161_;
  wire _31162_;
  wire _31163_;
  wire _31164_;
  wire _31165_;
  wire _31166_;
  wire _31167_;
  wire _31168_;
  wire _31169_;
  wire _31170_;
  wire _31171_;
  wire _31172_;
  wire _31173_;
  wire _31174_;
  wire _31175_;
  wire _31176_;
  wire _31177_;
  wire _31178_;
  wire _31179_;
  wire _31180_;
  wire _31181_;
  wire _31182_;
  wire _31183_;
  wire _31184_;
  wire _31185_;
  wire _31186_;
  wire _31187_;
  wire _31188_;
  wire _31189_;
  wire _31190_;
  wire _31191_;
  wire _31192_;
  wire _31193_;
  wire _31194_;
  wire _31195_;
  wire _31196_;
  wire _31197_;
  wire _31198_;
  wire _31199_;
  wire _31200_;
  wire _31201_;
  wire _31202_;
  wire _31203_;
  wire _31204_;
  wire _31205_;
  wire _31206_;
  wire _31207_;
  wire _31208_;
  wire _31209_;
  wire _31210_;
  wire _31211_;
  wire _31212_;
  wire _31213_;
  wire _31214_;
  wire _31215_;
  wire _31216_;
  wire _31217_;
  wire _31218_;
  wire _31219_;
  wire _31220_;
  wire _31221_;
  wire _31222_;
  wire _31223_;
  wire _31224_;
  wire _31225_;
  wire _31226_;
  wire _31227_;
  wire _31228_;
  wire _31229_;
  wire _31230_;
  wire _31231_;
  wire _31232_;
  wire _31233_;
  wire _31234_;
  wire _31235_;
  wire _31236_;
  wire _31237_;
  wire _31238_;
  wire _31239_;
  wire _31240_;
  wire _31241_;
  wire _31242_;
  wire _31243_;
  wire _31244_;
  wire _31245_;
  wire _31246_;
  wire _31247_;
  wire _31248_;
  wire _31249_;
  wire _31250_;
  wire _31251_;
  wire _31252_;
  wire _31253_;
  wire _31254_;
  wire _31255_;
  wire _31256_;
  wire _31257_;
  wire _31258_;
  wire _31259_;
  wire _31260_;
  wire _31261_;
  wire _31262_;
  wire _31263_;
  wire _31264_;
  wire _31265_;
  wire _31266_;
  wire _31267_;
  wire _31268_;
  wire _31269_;
  wire _31270_;
  wire _31271_;
  wire _31272_;
  wire _31273_;
  wire _31274_;
  wire _31275_;
  wire _31276_;
  wire _31277_;
  wire _31278_;
  wire _31279_;
  wire _31280_;
  wire _31281_;
  wire _31282_;
  wire _31283_;
  wire _31284_;
  wire _31285_;
  wire _31286_;
  wire _31287_;
  wire _31288_;
  wire _31289_;
  wire _31290_;
  wire _31291_;
  wire _31292_;
  wire _31293_;
  wire _31294_;
  wire _31295_;
  wire _31296_;
  wire _31297_;
  wire _31298_;
  wire _31299_;
  wire _31300_;
  wire _31301_;
  wire _31302_;
  wire _31303_;
  wire _31304_;
  wire _31305_;
  wire _31306_;
  wire _31307_;
  wire _31308_;
  wire _31309_;
  wire _31310_;
  wire _31311_;
  wire _31312_;
  wire _31313_;
  wire _31314_;
  wire _31315_;
  wire _31316_;
  wire _31317_;
  wire _31318_;
  wire _31319_;
  wire _31320_;
  wire _31321_;
  wire _31322_;
  wire _31323_;
  wire _31324_;
  wire _31325_;
  wire _31326_;
  wire _31327_;
  wire _31328_;
  wire _31329_;
  wire _31330_;
  wire _31331_;
  wire _31332_;
  wire _31333_;
  wire _31334_;
  wire _31335_;
  wire _31336_;
  wire _31337_;
  wire _31338_;
  wire _31339_;
  wire _31340_;
  wire _31341_;
  wire _31342_;
  wire _31343_;
  wire _31344_;
  wire _31345_;
  wire _31346_;
  wire _31347_;
  wire _31348_;
  wire _31349_;
  wire _31350_;
  wire _31351_;
  wire _31352_;
  wire _31353_;
  wire _31354_;
  wire _31355_;
  wire _31356_;
  wire _31357_;
  wire _31358_;
  wire _31359_;
  wire _31360_;
  wire _31361_;
  wire _31362_;
  wire _31363_;
  wire _31364_;
  wire _31365_;
  wire _31366_;
  wire _31367_;
  wire _31368_;
  wire _31369_;
  wire _31370_;
  wire _31371_;
  wire _31372_;
  wire _31373_;
  wire _31374_;
  wire _31375_;
  wire _31376_;
  wire _31377_;
  wire _31378_;
  wire _31379_;
  wire _31380_;
  wire _31381_;
  wire _31382_;
  wire _31383_;
  wire _31384_;
  wire _31385_;
  wire _31386_;
  wire _31387_;
  wire _31388_;
  wire _31389_;
  wire _31390_;
  wire _31391_;
  wire _31392_;
  wire _31393_;
  wire _31394_;
  wire _31395_;
  wire _31396_;
  wire _31397_;
  wire _31398_;
  wire _31399_;
  wire _31400_;
  wire _31401_;
  wire _31402_;
  wire _31403_;
  wire _31404_;
  wire _31405_;
  wire _31406_;
  wire _31407_;
  wire _31408_;
  wire _31409_;
  wire _31410_;
  wire _31411_;
  wire _31412_;
  wire _31413_;
  wire _31414_;
  wire _31415_;
  wire _31416_;
  wire _31417_;
  wire _31418_;
  wire _31419_;
  wire _31420_;
  wire _31421_;
  wire _31422_;
  wire _31423_;
  wire _31424_;
  wire _31425_;
  wire _31426_;
  wire _31427_;
  wire _31428_;
  wire _31429_;
  wire _31430_;
  wire _31431_;
  wire _31432_;
  wire _31433_;
  wire _31434_;
  wire _31435_;
  wire _31436_;
  wire _31437_;
  wire _31438_;
  wire _31439_;
  wire _31440_;
  wire _31441_;
  wire _31442_;
  wire _31443_;
  wire _31444_;
  wire _31445_;
  wire _31446_;
  wire _31447_;
  wire _31448_;
  wire _31449_;
  wire _31450_;
  wire _31451_;
  wire _31452_;
  wire _31453_;
  wire _31454_;
  wire _31455_;
  wire _31456_;
  wire _31457_;
  wire _31458_;
  wire _31459_;
  wire _31460_;
  wire _31461_;
  wire _31462_;
  wire _31463_;
  wire _31464_;
  wire _31465_;
  wire _31466_;
  wire _31467_;
  wire _31468_;
  wire _31469_;
  wire _31470_;
  wire _31471_;
  wire _31472_;
  wire _31473_;
  wire _31474_;
  wire _31475_;
  wire _31476_;
  wire _31477_;
  wire _31478_;
  wire _31479_;
  wire _31480_;
  wire _31481_;
  wire _31482_;
  wire _31483_;
  wire _31484_;
  wire _31485_;
  wire _31486_;
  wire _31487_;
  wire _31488_;
  wire _31489_;
  wire _31490_;
  wire _31491_;
  wire _31492_;
  wire _31493_;
  wire _31494_;
  wire _31495_;
  wire _31496_;
  wire _31497_;
  wire _31498_;
  wire _31499_;
  wire _31500_;
  wire _31501_;
  wire _31502_;
  wire _31503_;
  wire _31504_;
  wire _31505_;
  wire _31506_;
  wire _31507_;
  wire _31508_;
  wire _31509_;
  wire _31510_;
  wire _31511_;
  wire _31512_;
  wire _31513_;
  wire _31514_;
  wire _31515_;
  wire _31516_;
  wire _31517_;
  wire _31518_;
  wire _31519_;
  wire _31520_;
  wire _31521_;
  wire _31522_;
  wire _31523_;
  wire _31524_;
  wire _31525_;
  wire _31526_;
  wire _31527_;
  wire _31528_;
  wire _31529_;
  wire _31530_;
  wire _31531_;
  wire _31532_;
  wire _31533_;
  wire _31534_;
  wire _31535_;
  wire _31536_;
  wire _31537_;
  wire _31538_;
  wire _31539_;
  wire _31540_;
  wire _31541_;
  wire _31542_;
  wire _31543_;
  wire _31544_;
  wire _31545_;
  wire _31546_;
  wire _31547_;
  wire _31548_;
  wire _31549_;
  wire _31550_;
  wire _31551_;
  wire _31552_;
  wire _31553_;
  wire _31554_;
  wire _31555_;
  wire _31556_;
  wire _31557_;
  wire _31558_;
  wire _31559_;
  wire _31560_;
  wire _31561_;
  wire _31562_;
  wire _31563_;
  wire _31564_;
  wire _31565_;
  wire _31566_;
  wire _31567_;
  wire _31568_;
  wire _31569_;
  wire _31570_;
  wire _31571_;
  wire _31572_;
  wire _31573_;
  wire _31574_;
  wire _31575_;
  wire _31576_;
  wire _31577_;
  wire _31578_;
  wire _31579_;
  wire _31580_;
  wire _31581_;
  wire _31582_;
  wire _31583_;
  wire _31584_;
  wire _31585_;
  wire _31586_;
  wire _31587_;
  wire _31588_;
  wire _31589_;
  wire _31590_;
  wire _31591_;
  wire _31592_;
  wire _31593_;
  wire _31594_;
  wire _31595_;
  wire _31596_;
  wire _31597_;
  wire _31598_;
  wire _31599_;
  wire _31600_;
  wire _31601_;
  wire _31602_;
  wire _31603_;
  wire _31604_;
  wire _31605_;
  wire _31606_;
  wire _31607_;
  wire _31608_;
  wire _31609_;
  wire _31610_;
  wire _31611_;
  wire _31612_;
  wire _31613_;
  wire _31614_;
  wire _31615_;
  wire _31616_;
  wire _31617_;
  wire _31618_;
  wire _31619_;
  wire _31620_;
  wire _31621_;
  wire _31622_;
  wire _31623_;
  wire _31624_;
  wire _31625_;
  wire _31626_;
  wire _31627_;
  wire _31628_;
  wire _31629_;
  wire _31630_;
  wire _31631_;
  wire _31632_;
  wire _31633_;
  wire _31634_;
  wire _31635_;
  wire _31636_;
  wire _31637_;
  wire _31638_;
  wire _31639_;
  wire _31640_;
  wire _31641_;
  wire _31642_;
  wire _31643_;
  wire _31644_;
  wire _31645_;
  wire _31646_;
  wire _31647_;
  wire _31648_;
  wire _31649_;
  wire _31650_;
  wire _31651_;
  wire _31652_;
  wire _31653_;
  wire _31654_;
  wire _31655_;
  wire _31656_;
  wire _31657_;
  wire _31658_;
  wire _31659_;
  wire _31660_;
  wire _31661_;
  wire _31662_;
  wire _31663_;
  wire _31664_;
  wire _31665_;
  wire _31666_;
  wire _31667_;
  wire _31668_;
  wire _31669_;
  wire _31670_;
  wire _31671_;
  wire _31672_;
  wire _31673_;
  wire _31674_;
  wire _31675_;
  wire _31676_;
  wire _31677_;
  wire _31678_;
  wire _31679_;
  wire _31680_;
  wire _31681_;
  wire _31682_;
  wire _31683_;
  wire _31684_;
  wire _31685_;
  wire _31686_;
  wire _31687_;
  wire _31688_;
  wire _31689_;
  wire _31690_;
  wire _31691_;
  wire _31692_;
  wire _31693_;
  wire _31694_;
  wire _31695_;
  wire _31696_;
  wire _31697_;
  wire _31698_;
  wire _31699_;
  wire _31700_;
  wire _31701_;
  wire _31702_;
  wire _31703_;
  wire _31704_;
  wire _31705_;
  wire _31706_;
  wire _31707_;
  wire _31708_;
  wire _31709_;
  wire _31710_;
  wire _31711_;
  wire _31712_;
  wire _31713_;
  wire _31714_;
  wire _31715_;
  wire _31716_;
  wire _31717_;
  wire _31718_;
  wire _31719_;
  wire _31720_;
  wire _31721_;
  wire _31722_;
  wire _31723_;
  wire _31724_;
  wire _31725_;
  wire _31726_;
  wire _31727_;
  wire _31728_;
  wire _31729_;
  wire _31730_;
  wire _31731_;
  wire _31732_;
  wire _31733_;
  wire _31734_;
  wire _31735_;
  wire _31736_;
  wire _31737_;
  wire _31738_;
  wire _31739_;
  wire _31740_;
  wire _31741_;
  wire _31742_;
  wire _31743_;
  wire _31744_;
  wire _31745_;
  wire _31746_;
  wire _31747_;
  wire _31748_;
  wire _31749_;
  wire _31750_;
  wire _31751_;
  wire _31752_;
  wire _31753_;
  wire _31754_;
  wire _31755_;
  wire _31756_;
  wire _31757_;
  wire _31758_;
  wire _31759_;
  wire _31760_;
  wire _31761_;
  wire _31762_;
  wire _31763_;
  wire _31764_;
  wire _31765_;
  wire _31766_;
  wire _31767_;
  wire _31768_;
  wire _31769_;
  wire _31770_;
  wire _31771_;
  wire _31772_;
  wire _31773_;
  wire _31774_;
  wire _31775_;
  wire _31776_;
  wire _31777_;
  wire _31778_;
  wire _31779_;
  wire _31780_;
  wire _31781_;
  wire _31782_;
  wire _31783_;
  wire _31784_;
  wire _31785_;
  wire _31786_;
  wire _31787_;
  wire _31788_;
  wire _31789_;
  wire _31790_;
  wire _31791_;
  wire _31792_;
  wire _31793_;
  wire _31794_;
  wire _31795_;
  wire _31796_;
  wire _31797_;
  wire _31798_;
  wire _31799_;
  wire _31800_;
  wire _31801_;
  wire _31802_;
  wire _31803_;
  wire _31804_;
  wire _31805_;
  wire _31806_;
  wire _31807_;
  wire _31808_;
  wire _31809_;
  wire _31810_;
  wire _31811_;
  wire _31812_;
  wire _31813_;
  wire _31814_;
  wire _31815_;
  wire _31816_;
  wire _31817_;
  wire _31818_;
  wire _31819_;
  wire _31820_;
  wire _31821_;
  wire _31822_;
  wire _31823_;
  wire _31824_;
  wire _31825_;
  wire _31826_;
  wire _31827_;
  wire _31828_;
  wire _31829_;
  wire _31830_;
  wire _31831_;
  wire _31832_;
  wire _31833_;
  wire _31834_;
  wire _31835_;
  wire _31836_;
  wire _31837_;
  wire _31838_;
  wire _31839_;
  wire _31840_;
  wire _31841_;
  wire _31842_;
  wire _31843_;
  wire _31844_;
  wire _31845_;
  wire _31846_;
  wire _31847_;
  wire _31848_;
  wire _31849_;
  wire _31850_;
  wire _31851_;
  wire _31852_;
  wire _31853_;
  wire _31854_;
  wire _31855_;
  wire _31856_;
  wire _31857_;
  wire _31858_;
  wire _31859_;
  wire _31860_;
  wire _31861_;
  wire _31862_;
  wire _31863_;
  wire _31864_;
  wire _31865_;
  wire _31866_;
  wire _31867_;
  wire _31868_;
  wire _31869_;
  wire _31870_;
  wire _31871_;
  wire _31872_;
  wire _31873_;
  wire _31874_;
  wire _31875_;
  wire _31876_;
  wire _31877_;
  wire _31878_;
  wire _31879_;
  wire _31880_;
  wire _31881_;
  wire _31882_;
  wire _31883_;
  wire _31884_;
  wire _31885_;
  wire _31886_;
  wire _31887_;
  wire _31888_;
  wire _31889_;
  wire _31890_;
  wire _31891_;
  wire _31892_;
  wire _31893_;
  wire _31894_;
  wire _31895_;
  wire _31896_;
  wire _31897_;
  wire _31898_;
  wire _31899_;
  wire _31900_;
  wire _31901_;
  wire _31902_;
  wire _31903_;
  wire _31904_;
  wire _31905_;
  wire _31906_;
  wire _31907_;
  wire _31908_;
  wire _31909_;
  wire _31910_;
  wire _31911_;
  wire _31912_;
  wire _31913_;
  wire _31914_;
  wire _31915_;
  wire _31916_;
  wire _31917_;
  wire _31918_;
  wire _31919_;
  wire _31920_;
  wire _31921_;
  wire _31922_;
  wire _31923_;
  wire _31924_;
  wire _31925_;
  wire _31926_;
  wire _31927_;
  wire _31928_;
  wire _31929_;
  wire _31930_;
  wire _31931_;
  wire _31932_;
  wire _31933_;
  wire _31934_;
  wire _31935_;
  wire _31936_;
  wire _31937_;
  wire _31938_;
  wire _31939_;
  wire _31940_;
  wire _31941_;
  wire _31942_;
  wire _31943_;
  wire _31944_;
  wire _31945_;
  wire _31946_;
  wire _31947_;
  wire _31948_;
  wire _31949_;
  wire _31950_;
  wire _31951_;
  wire _31952_;
  wire _31953_;
  wire _31954_;
  wire _31955_;
  wire _31956_;
  wire _31957_;
  wire _31958_;
  wire _31959_;
  wire _31960_;
  wire _31961_;
  wire _31962_;
  wire _31963_;
  wire _31964_;
  wire _31965_;
  wire _31966_;
  wire _31967_;
  wire _31968_;
  wire _31969_;
  wire _31970_;
  wire _31971_;
  wire _31972_;
  wire _31973_;
  wire _31974_;
  wire _31975_;
  wire _31976_;
  wire _31977_;
  wire _31978_;
  wire _31979_;
  wire _31980_;
  wire _31981_;
  wire _31982_;
  wire _31983_;
  wire _31984_;
  wire _31985_;
  wire _31986_;
  wire _31987_;
  wire _31988_;
  wire _31989_;
  wire _31990_;
  wire _31991_;
  wire _31992_;
  wire _31993_;
  wire _31994_;
  wire _31995_;
  wire _31996_;
  wire _31997_;
  wire _31998_;
  wire _31999_;
  wire _32000_;
  wire _32001_;
  wire _32002_;
  wire _32003_;
  wire _32004_;
  wire _32005_;
  wire _32006_;
  wire _32007_;
  wire _32008_;
  wire _32009_;
  wire _32010_;
  wire _32011_;
  wire _32012_;
  wire _32013_;
  wire _32014_;
  wire _32015_;
  wire _32016_;
  wire _32017_;
  wire _32018_;
  wire _32019_;
  wire _32020_;
  wire _32021_;
  wire _32022_;
  wire _32023_;
  wire _32024_;
  wire _32025_;
  wire _32026_;
  wire _32027_;
  wire _32028_;
  wire _32029_;
  wire _32030_;
  wire _32031_;
  wire _32032_;
  wire _32033_;
  wire _32034_;
  wire _32035_;
  wire _32036_;
  wire _32037_;
  wire _32038_;
  wire _32039_;
  wire _32040_;
  wire _32041_;
  wire _32042_;
  wire _32043_;
  wire _32044_;
  wire _32045_;
  wire _32046_;
  wire _32047_;
  wire _32048_;
  wire _32049_;
  wire _32050_;
  wire _32051_;
  wire _32052_;
  wire _32053_;
  wire _32054_;
  wire _32055_;
  wire _32056_;
  wire _32057_;
  wire _32058_;
  wire _32059_;
  wire _32060_;
  wire _32061_;
  wire _32062_;
  wire _32063_;
  wire _32064_;
  wire _32065_;
  wire _32066_;
  wire _32067_;
  wire _32068_;
  wire _32069_;
  wire _32070_;
  wire _32071_;
  wire _32072_;
  wire _32073_;
  wire _32074_;
  wire _32075_;
  wire _32076_;
  wire _32077_;
  wire _32078_;
  wire _32079_;
  wire _32080_;
  wire _32081_;
  wire _32082_;
  wire _32083_;
  wire _32084_;
  wire _32085_;
  wire _32086_;
  wire _32087_;
  wire _32088_;
  wire _32089_;
  wire _32090_;
  wire _32091_;
  wire _32092_;
  wire _32093_;
  wire _32094_;
  wire _32095_;
  wire _32096_;
  wire _32097_;
  wire _32098_;
  wire _32099_;
  wire _32100_;
  wire _32101_;
  wire _32102_;
  wire _32103_;
  wire _32104_;
  wire _32105_;
  wire _32106_;
  wire _32107_;
  wire _32108_;
  wire _32109_;
  wire _32110_;
  wire _32111_;
  wire _32112_;
  wire _32113_;
  wire _32114_;
  wire _32115_;
  wire _32116_;
  wire _32117_;
  wire _32118_;
  wire _32119_;
  wire _32120_;
  wire _32121_;
  wire _32122_;
  wire _32123_;
  wire _32124_;
  wire _32125_;
  wire _32126_;
  wire _32127_;
  wire _32128_;
  wire _32129_;
  wire _32130_;
  wire _32131_;
  wire _32132_;
  wire _32133_;
  wire _32134_;
  wire _32135_;
  wire _32136_;
  wire _32137_;
  wire _32138_;
  wire _32139_;
  wire _32140_;
  wire _32141_;
  wire _32142_;
  wire _32143_;
  wire _32144_;
  wire _32145_;
  wire _32146_;
  wire _32147_;
  wire _32148_;
  wire _32149_;
  wire _32150_;
  wire _32151_;
  wire _32152_;
  wire _32153_;
  wire _32154_;
  wire _32155_;
  wire _32156_;
  wire _32157_;
  wire _32158_;
  wire _32159_;
  wire _32160_;
  wire _32161_;
  wire _32162_;
  wire _32163_;
  wire _32164_;
  wire _32165_;
  wire _32166_;
  wire _32167_;
  wire _32168_;
  wire _32169_;
  wire _32170_;
  wire _32171_;
  wire _32172_;
  wire _32173_;
  wire _32174_;
  wire _32175_;
  wire _32176_;
  wire _32177_;
  wire _32178_;
  wire _32179_;
  wire _32180_;
  wire _32181_;
  wire _32182_;
  wire _32183_;
  wire _32184_;
  wire _32185_;
  wire _32186_;
  wire _32187_;
  wire _32188_;
  wire _32189_;
  wire _32190_;
  wire _32191_;
  wire _32192_;
  wire _32193_;
  wire _32194_;
  wire _32195_;
  wire _32196_;
  wire _32197_;
  wire _32198_;
  wire _32199_;
  wire _32200_;
  wire _32201_;
  wire _32202_;
  wire _32203_;
  wire _32204_;
  wire _32205_;
  wire _32206_;
  wire _32207_;
  wire _32208_;
  wire _32209_;
  wire _32210_;
  wire _32211_;
  wire _32212_;
  wire _32213_;
  wire _32214_;
  wire _32215_;
  wire _32216_;
  wire _32217_;
  wire _32218_;
  wire _32219_;
  wire _32220_;
  wire _32221_;
  wire _32222_;
  wire _32223_;
  wire _32224_;
  wire _32225_;
  wire _32226_;
  wire _32227_;
  wire _32228_;
  wire _32229_;
  wire _32230_;
  wire _32231_;
  wire _32232_;
  wire _32233_;
  wire _32234_;
  wire _32235_;
  wire _32236_;
  wire _32237_;
  wire _32238_;
  wire _32239_;
  wire _32240_;
  wire _32241_;
  wire _32242_;
  wire _32243_;
  wire _32244_;
  wire _32245_;
  wire _32246_;
  wire _32247_;
  wire _32248_;
  wire _32249_;
  wire _32250_;
  wire _32251_;
  wire _32252_;
  wire _32253_;
  wire _32254_;
  wire _32255_;
  wire _32256_;
  wire _32257_;
  wire _32258_;
  wire _32259_;
  wire _32260_;
  wire _32261_;
  wire _32262_;
  wire _32263_;
  wire _32264_;
  wire _32265_;
  wire _32266_;
  wire _32267_;
  wire _32268_;
  wire _32269_;
  wire _32270_;
  wire _32271_;
  wire _32272_;
  wire _32273_;
  wire _32274_;
  wire _32275_;
  wire _32276_;
  wire _32277_;
  wire _32278_;
  wire _32279_;
  wire _32280_;
  wire _32281_;
  wire _32282_;
  wire _32283_;
  wire _32284_;
  wire _32285_;
  wire _32286_;
  wire _32287_;
  wire _32288_;
  wire _32289_;
  wire _32290_;
  wire _32291_;
  wire _32292_;
  wire _32293_;
  wire _32294_;
  wire _32295_;
  wire _32296_;
  wire _32297_;
  wire _32298_;
  wire _32299_;
  wire _32300_;
  wire _32301_;
  wire _32302_;
  wire _32303_;
  wire _32304_;
  wire _32305_;
  wire _32306_;
  wire _32307_;
  wire _32308_;
  wire _32309_;
  wire _32310_;
  wire _32311_;
  wire _32312_;
  wire _32313_;
  wire _32314_;
  wire _32315_;
  wire _32316_;
  wire _32317_;
  wire _32318_;
  wire _32319_;
  wire _32320_;
  wire _32321_;
  wire _32322_;
  wire _32323_;
  wire _32324_;
  wire _32325_;
  wire _32326_;
  wire _32327_;
  wire _32328_;
  wire _32329_;
  wire _32330_;
  wire _32331_;
  wire _32332_;
  wire _32333_;
  wire _32334_;
  wire _32335_;
  wire _32336_;
  wire _32337_;
  wire _32338_;
  wire _32339_;
  wire _32340_;
  wire _32341_;
  wire _32342_;
  wire _32343_;
  wire _32344_;
  wire _32345_;
  wire _32346_;
  wire _32347_;
  wire _32348_;
  wire _32349_;
  wire _32350_;
  wire _32351_;
  wire _32352_;
  wire _32353_;
  wire _32354_;
  wire _32355_;
  wire _32356_;
  wire _32357_;
  wire _32358_;
  wire _32359_;
  wire _32360_;
  wire _32361_;
  wire _32362_;
  wire _32363_;
  wire _32364_;
  wire _32365_;
  wire _32366_;
  wire _32367_;
  wire _32368_;
  wire _32369_;
  wire _32370_;
  wire _32371_;
  wire _32372_;
  wire _32373_;
  wire _32374_;
  wire _32375_;
  wire _32376_;
  wire _32377_;
  wire _32378_;
  wire _32379_;
  wire _32380_;
  wire _32381_;
  wire _32382_;
  wire _32383_;
  wire _32384_;
  wire _32385_;
  wire _32386_;
  wire _32387_;
  wire _32388_;
  wire _32389_;
  wire _32390_;
  wire _32391_;
  wire _32392_;
  wire _32393_;
  wire _32394_;
  wire _32395_;
  wire _32396_;
  wire _32397_;
  wire _32398_;
  wire _32399_;
  wire _32400_;
  wire _32401_;
  wire _32402_;
  wire _32403_;
  wire _32404_;
  wire _32405_;
  wire _32406_;
  wire _32407_;
  wire _32408_;
  wire _32409_;
  wire _32410_;
  wire _32411_;
  wire _32412_;
  wire _32413_;
  wire _32414_;
  wire _32415_;
  wire _32416_;
  wire _32417_;
  wire _32418_;
  wire _32419_;
  wire _32420_;
  wire _32421_;
  wire _32422_;
  wire _32423_;
  wire _32424_;
  wire _32425_;
  wire _32426_;
  wire _32427_;
  wire _32428_;
  wire _32429_;
  wire _32430_;
  wire _32431_;
  wire _32432_;
  wire _32433_;
  wire _32434_;
  wire _32435_;
  wire _32436_;
  wire _32437_;
  wire _32438_;
  wire _32439_;
  wire _32440_;
  wire _32441_;
  wire _32442_;
  wire _32443_;
  wire _32444_;
  wire _32445_;
  wire _32446_;
  wire _32447_;
  wire _32448_;
  wire _32449_;
  wire _32450_;
  wire _32451_;
  wire _32452_;
  wire _32453_;
  wire _32454_;
  wire _32455_;
  wire _32456_;
  wire _32457_;
  wire _32458_;
  wire _32459_;
  wire _32460_;
  wire _32461_;
  wire _32462_;
  wire _32463_;
  wire _32464_;
  wire _32465_;
  wire _32466_;
  wire _32467_;
  wire _32468_;
  wire _32469_;
  wire _32470_;
  wire _32471_;
  wire _32472_;
  wire _32473_;
  wire _32474_;
  wire _32475_;
  wire _32476_;
  wire _32477_;
  wire _32478_;
  wire _32479_;
  wire _32480_;
  wire _32481_;
  wire _32482_;
  wire _32483_;
  wire _32484_;
  wire _32485_;
  wire _32486_;
  wire _32487_;
  wire _32488_;
  wire _32489_;
  wire _32490_;
  wire _32491_;
  wire _32492_;
  wire _32493_;
  wire _32494_;
  wire _32495_;
  wire _32496_;
  wire _32497_;
  wire _32498_;
  wire _32499_;
  wire _32500_;
  wire _32501_;
  wire _32502_;
  wire _32503_;
  wire _32504_;
  wire _32505_;
  wire _32506_;
  wire _32507_;
  wire _32508_;
  wire _32509_;
  wire _32510_;
  wire _32511_;
  wire _32512_;
  wire _32513_;
  wire _32514_;
  wire _32515_;
  wire _32516_;
  wire _32517_;
  wire _32518_;
  wire _32519_;
  wire _32520_;
  wire _32521_;
  wire _32522_;
  wire _32523_;
  wire _32524_;
  wire _32525_;
  wire _32526_;
  wire _32527_;
  wire _32528_;
  wire _32529_;
  wire _32530_;
  wire _32531_;
  wire _32532_;
  wire _32533_;
  wire _32534_;
  wire _32535_;
  wire _32536_;
  wire _32537_;
  wire _32538_;
  wire _32539_;
  wire _32540_;
  wire _32541_;
  wire _32542_;
  wire _32543_;
  wire _32544_;
  wire _32545_;
  wire _32546_;
  wire _32547_;
  wire _32548_;
  wire _32549_;
  wire _32550_;
  wire _32551_;
  wire _32552_;
  wire _32553_;
  wire _32554_;
  wire _32555_;
  wire _32556_;
  wire _32557_;
  wire _32558_;
  wire _32559_;
  wire _32560_;
  wire _32561_;
  wire _32562_;
  wire _32563_;
  wire _32564_;
  wire _32565_;
  wire _32566_;
  wire _32567_;
  wire _32568_;
  wire _32569_;
  wire _32570_;
  wire _32571_;
  wire _32572_;
  wire _32573_;
  wire _32574_;
  wire _32575_;
  wire _32576_;
  wire _32577_;
  wire _32578_;
  wire _32579_;
  wire _32580_;
  wire _32581_;
  wire _32582_;
  wire _32583_;
  wire _32584_;
  wire _32585_;
  wire _32586_;
  wire _32587_;
  wire _32588_;
  wire _32589_;
  wire _32590_;
  wire _32591_;
  wire _32592_;
  wire _32593_;
  wire _32594_;
  wire _32595_;
  wire _32596_;
  wire _32597_;
  wire _32598_;
  wire _32599_;
  wire _32600_;
  wire _32601_;
  wire _32602_;
  wire _32603_;
  wire _32604_;
  wire _32605_;
  wire _32606_;
  wire _32607_;
  wire _32608_;
  wire _32609_;
  wire _32610_;
  wire _32611_;
  wire _32612_;
  wire _32613_;
  wire _32614_;
  wire _32615_;
  wire _32616_;
  wire _32617_;
  wire _32618_;
  wire _32619_;
  wire _32620_;
  wire _32621_;
  wire _32622_;
  wire _32623_;
  wire _32624_;
  wire _32625_;
  wire _32626_;
  wire _32627_;
  wire _32628_;
  wire _32629_;
  wire _32630_;
  wire _32631_;
  wire _32632_;
  wire _32633_;
  wire _32634_;
  wire _32635_;
  wire _32636_;
  wire _32637_;
  wire _32638_;
  wire _32639_;
  wire _32640_;
  wire _32641_;
  wire _32642_;
  wire _32643_;
  wire _32644_;
  wire _32645_;
  wire _32646_;
  wire _32647_;
  wire _32648_;
  wire _32649_;
  wire _32650_;
  wire _32651_;
  wire _32652_;
  wire _32653_;
  wire _32654_;
  wire _32655_;
  wire _32656_;
  wire _32657_;
  wire _32658_;
  wire _32659_;
  wire _32660_;
  wire _32661_;
  wire _32662_;
  wire _32663_;
  wire _32664_;
  wire _32665_;
  wire _32666_;
  wire _32667_;
  wire _32668_;
  wire _32669_;
  wire _32670_;
  wire _32671_;
  wire _32672_;
  wire _32673_;
  wire _32674_;
  wire _32675_;
  wire _32676_;
  wire _32677_;
  wire _32678_;
  wire _32679_;
  wire _32680_;
  wire _32681_;
  wire _32682_;
  wire _32683_;
  wire _32684_;
  wire _32685_;
  wire _32686_;
  wire _32687_;
  wire _32688_;
  wire _32689_;
  wire _32690_;
  wire _32691_;
  wire _32692_;
  wire _32693_;
  wire _32694_;
  wire _32695_;
  wire _32696_;
  wire _32697_;
  wire _32698_;
  wire _32699_;
  wire _32700_;
  wire _32701_;
  wire _32702_;
  wire _32703_;
  wire _32704_;
  wire _32705_;
  wire _32706_;
  wire _32707_;
  wire _32708_;
  wire _32709_;
  wire _32710_;
  wire _32711_;
  wire _32712_;
  wire _32713_;
  wire _32714_;
  wire _32715_;
  wire _32716_;
  wire _32717_;
  wire _32718_;
  wire _32719_;
  wire _32720_;
  wire _32721_;
  wire _32722_;
  wire _32723_;
  wire _32724_;
  wire _32725_;
  wire _32726_;
  wire _32727_;
  wire _32728_;
  wire _32729_;
  wire _32730_;
  wire _32731_;
  wire _32732_;
  wire _32733_;
  wire _32734_;
  wire _32735_;
  wire _32736_;
  wire _32737_;
  wire _32738_;
  wire _32739_;
  wire _32740_;
  wire _32741_;
  wire _32742_;
  wire _32743_;
  wire _32744_;
  wire _32745_;
  wire _32746_;
  wire _32747_;
  wire _32748_;
  wire _32749_;
  wire _32750_;
  wire _32751_;
  wire _32752_;
  wire _32753_;
  wire _32754_;
  wire _32755_;
  wire _32756_;
  wire _32757_;
  wire _32758_;
  wire _32759_;
  wire _32760_;
  wire _32761_;
  wire _32762_;
  wire _32763_;
  wire _32764_;
  wire _32765_;
  wire _32766_;
  wire _32767_;
  wire _32768_;
  wire _32769_;
  wire _32770_;
  wire _32771_;
  wire _32772_;
  wire _32773_;
  wire _32774_;
  wire _32775_;
  wire _32776_;
  wire _32777_;
  wire _32778_;
  wire _32779_;
  wire _32780_;
  wire _32781_;
  wire _32782_;
  wire _32783_;
  wire _32784_;
  wire _32785_;
  wire _32786_;
  wire _32787_;
  wire _32788_;
  wire _32789_;
  wire _32790_;
  wire _32791_;
  wire _32792_;
  wire _32793_;
  wire _32794_;
  wire _32795_;
  wire _32796_;
  wire _32797_;
  wire _32798_;
  wire _32799_;
  wire _32800_;
  wire _32801_;
  wire _32802_;
  wire _32803_;
  wire _32804_;
  wire _32805_;
  wire _32806_;
  wire _32807_;
  wire _32808_;
  wire _32809_;
  wire _32810_;
  wire _32811_;
  wire _32812_;
  wire _32813_;
  wire _32814_;
  wire _32815_;
  wire _32816_;
  wire _32817_;
  wire _32818_;
  wire _32819_;
  wire _32820_;
  wire _32821_;
  wire _32822_;
  wire _32823_;
  wire _32824_;
  wire _32825_;
  wire _32826_;
  wire _32827_;
  wire _32828_;
  wire _32829_;
  wire _32830_;
  wire _32831_;
  wire _32832_;
  wire _32833_;
  wire _32834_;
  wire _32835_;
  wire _32836_;
  wire _32837_;
  wire _32838_;
  wire _32839_;
  wire _32840_;
  wire _32841_;
  wire _32842_;
  wire _32843_;
  wire _32844_;
  wire _32845_;
  wire _32846_;
  wire _32847_;
  wire _32848_;
  wire _32849_;
  wire _32850_;
  wire _32851_;
  wire _32852_;
  wire _32853_;
  wire _32854_;
  wire _32855_;
  wire _32856_;
  wire _32857_;
  wire _32858_;
  wire _32859_;
  wire _32860_;
  wire _32861_;
  wire _32862_;
  wire _32863_;
  wire _32864_;
  wire _32865_;
  wire _32866_;
  wire _32867_;
  wire _32868_;
  wire _32869_;
  wire _32870_;
  wire _32871_;
  wire _32872_;
  wire _32873_;
  wire _32874_;
  wire _32875_;
  wire _32876_;
  wire _32877_;
  wire _32878_;
  wire _32879_;
  wire _32880_;
  wire _32881_;
  wire _32882_;
  wire _32883_;
  wire _32884_;
  wire _32885_;
  wire _32886_;
  wire _32887_;
  wire _32888_;
  wire _32889_;
  wire _32890_;
  wire _32891_;
  wire _32892_;
  wire _32893_;
  wire _32894_;
  wire _32895_;
  wire _32896_;
  wire _32897_;
  wire _32898_;
  wire _32899_;
  wire _32900_;
  wire _32901_;
  wire _32902_;
  wire _32903_;
  wire _32904_;
  wire _32905_;
  wire _32906_;
  wire _32907_;
  wire _32908_;
  wire _32909_;
  wire _32910_;
  wire _32911_;
  wire _32912_;
  wire _32913_;
  wire _32914_;
  wire _32915_;
  wire _32916_;
  wire _32917_;
  wire _32918_;
  wire _32919_;
  wire _32920_;
  wire _32921_;
  wire _32922_;
  wire _32923_;
  wire _32924_;
  wire _32925_;
  wire _32926_;
  wire _32927_;
  wire _32928_;
  wire _32929_;
  wire _32930_;
  wire _32931_;
  wire _32932_;
  wire _32933_;
  wire _32934_;
  wire _32935_;
  wire _32936_;
  wire _32937_;
  wire _32938_;
  wire _32939_;
  wire _32940_;
  wire _32941_;
  wire _32942_;
  wire _32943_;
  wire _32944_;
  wire _32945_;
  wire _32946_;
  wire _32947_;
  wire _32948_;
  wire _32949_;
  wire _32950_;
  wire _32951_;
  wire _32952_;
  wire _32953_;
  wire _32954_;
  wire _32955_;
  wire _32956_;
  wire _32957_;
  wire _32958_;
  wire _32959_;
  wire _32960_;
  wire _32961_;
  wire _32962_;
  wire _32963_;
  wire _32964_;
  wire _32965_;
  wire _32966_;
  wire _32967_;
  wire _32968_;
  wire _32969_;
  wire _32970_;
  wire _32971_;
  wire _32972_;
  wire _32973_;
  wire _32974_;
  wire _32975_;
  wire _32976_;
  wire _32977_;
  wire _32978_;
  wire _32979_;
  wire _32980_;
  wire _32981_;
  wire _32982_;
  wire _32983_;
  wire _32984_;
  wire _32985_;
  wire _32986_;
  wire _32987_;
  wire _32988_;
  wire _32989_;
  wire _32990_;
  wire _32991_;
  wire _32992_;
  wire _32993_;
  wire _32994_;
  wire _32995_;
  wire _32996_;
  wire _32997_;
  wire _32998_;
  wire _32999_;
  wire _33000_;
  wire _33001_;
  wire _33002_;
  wire _33003_;
  wire _33004_;
  wire _33005_;
  wire _33006_;
  wire _33007_;
  wire _33008_;
  wire _33009_;
  wire _33010_;
  wire _33011_;
  wire _33012_;
  wire _33013_;
  wire _33014_;
  wire _33015_;
  wire _33016_;
  wire _33017_;
  wire _33018_;
  wire _33019_;
  wire _33020_;
  wire _33021_;
  wire _33022_;
  wire _33023_;
  wire _33024_;
  wire _33025_;
  wire _33026_;
  wire _33027_;
  wire _33028_;
  wire _33029_;
  wire _33030_;
  wire _33031_;
  wire _33032_;
  wire _33033_;
  wire _33034_;
  wire _33035_;
  wire _33036_;
  wire _33037_;
  wire _33038_;
  wire _33039_;
  wire _33040_;
  wire _33041_;
  wire _33042_;
  wire _33043_;
  wire _33044_;
  wire _33045_;
  wire _33046_;
  wire _33047_;
  wire _33048_;
  wire _33049_;
  wire _33050_;
  wire _33051_;
  wire _33052_;
  wire _33053_;
  wire _33054_;
  wire _33055_;
  wire _33056_;
  wire _33057_;
  wire _33058_;
  wire _33059_;
  wire _33060_;
  wire _33061_;
  wire _33062_;
  wire _33063_;
  wire _33064_;
  wire _33065_;
  wire _33066_;
  wire _33067_;
  wire _33068_;
  wire _33069_;
  wire _33070_;
  wire _33071_;
  wire _33072_;
  wire _33073_;
  wire _33074_;
  wire _33075_;
  wire _33076_;
  wire _33077_;
  wire _33078_;
  wire _33079_;
  wire _33080_;
  wire _33081_;
  wire _33082_;
  wire _33083_;
  wire _33084_;
  wire _33085_;
  wire _33086_;
  wire _33087_;
  wire _33088_;
  wire _33089_;
  wire _33090_;
  wire _33091_;
  wire _33092_;
  wire _33093_;
  wire _33094_;
  wire _33095_;
  wire _33096_;
  wire _33097_;
  wire _33098_;
  wire _33099_;
  wire _33100_;
  wire _33101_;
  wire _33102_;
  wire _33103_;
  wire _33104_;
  wire _33105_;
  wire _33106_;
  wire _33107_;
  wire _33108_;
  wire _33109_;
  wire _33110_;
  wire _33111_;
  wire _33112_;
  wire _33113_;
  wire _33114_;
  wire _33115_;
  wire _33116_;
  wire _33117_;
  wire _33118_;
  wire _33119_;
  wire _33120_;
  wire _33121_;
  wire _33122_;
  wire _33123_;
  wire _33124_;
  wire _33125_;
  wire _33126_;
  wire _33127_;
  wire _33128_;
  wire _33129_;
  wire _33130_;
  wire _33131_;
  wire _33132_;
  wire _33133_;
  wire _33134_;
  wire _33135_;
  wire _33136_;
  wire _33137_;
  wire _33138_;
  wire _33139_;
  wire _33140_;
  wire _33141_;
  wire _33142_;
  wire _33143_;
  wire _33144_;
  wire _33145_;
  wire _33146_;
  wire _33147_;
  wire _33148_;
  wire _33149_;
  wire _33150_;
  wire _33151_;
  wire _33152_;
  wire _33153_;
  wire _33154_;
  wire _33155_;
  wire _33156_;
  wire _33157_;
  wire _33158_;
  wire _33159_;
  wire _33160_;
  wire _33161_;
  wire _33162_;
  wire _33163_;
  wire _33164_;
  wire _33165_;
  wire _33166_;
  wire _33167_;
  wire _33168_;
  wire _33169_;
  wire _33170_;
  wire _33171_;
  wire _33172_;
  wire _33173_;
  wire _33174_;
  wire _33175_;
  wire _33176_;
  wire _33177_;
  wire _33178_;
  wire _33179_;
  wire _33180_;
  wire _33181_;
  wire _33182_;
  wire _33183_;
  wire _33184_;
  wire _33185_;
  wire _33186_;
  wire _33187_;
  wire _33188_;
  wire _33189_;
  wire _33190_;
  wire _33191_;
  wire _33192_;
  wire _33193_;
  wire _33194_;
  wire _33195_;
  wire _33196_;
  wire _33197_;
  wire _33198_;
  wire _33199_;
  wire _33200_;
  wire _33201_;
  wire _33202_;
  wire _33203_;
  wire _33204_;
  wire _33205_;
  wire _33206_;
  wire _33207_;
  wire _33208_;
  wire _33209_;
  wire _33210_;
  wire _33211_;
  wire _33212_;
  wire _33213_;
  wire _33214_;
  wire _33215_;
  wire _33216_;
  wire _33217_;
  wire _33218_;
  wire _33219_;
  wire _33220_;
  wire _33221_;
  wire _33222_;
  wire _33223_;
  wire _33224_;
  wire _33225_;
  wire _33226_;
  wire _33227_;
  wire _33228_;
  wire _33229_;
  wire _33230_;
  wire _33231_;
  wire _33232_;
  wire _33233_;
  wire _33234_;
  wire _33235_;
  wire _33236_;
  wire _33237_;
  wire _33238_;
  wire _33239_;
  wire _33240_;
  wire _33241_;
  wire _33242_;
  wire _33243_;
  wire _33244_;
  wire _33245_;
  wire _33246_;
  wire _33247_;
  wire _33248_;
  wire _33249_;
  wire _33250_;
  wire _33251_;
  wire _33252_;
  wire _33253_;
  wire _33254_;
  wire _33255_;
  wire _33256_;
  wire _33257_;
  wire _33258_;
  wire _33259_;
  wire _33260_;
  wire _33261_;
  wire _33262_;
  wire _33263_;
  wire _33264_;
  wire _33265_;
  wire _33266_;
  wire _33267_;
  wire _33268_;
  wire _33269_;
  wire _33270_;
  wire _33271_;
  wire _33272_;
  wire _33273_;
  wire _33274_;
  wire _33275_;
  wire _33276_;
  wire _33277_;
  wire _33278_;
  wire _33279_;
  wire _33280_;
  wire _33281_;
  wire _33282_;
  wire _33283_;
  wire _33284_;
  wire _33285_;
  wire _33286_;
  wire _33287_;
  wire _33288_;
  wire _33289_;
  wire _33290_;
  wire _33291_;
  wire _33292_;
  wire _33293_;
  wire _33294_;
  wire _33295_;
  wire _33296_;
  wire _33297_;
  wire _33298_;
  wire _33299_;
  wire _33300_;
  wire _33301_;
  wire _33302_;
  wire _33303_;
  wire _33304_;
  wire _33305_;
  wire _33306_;
  wire _33307_;
  wire _33308_;
  wire _33309_;
  wire _33310_;
  wire _33311_;
  wire _33312_;
  wire _33313_;
  wire _33314_;
  wire _33315_;
  wire _33316_;
  wire _33317_;
  wire _33318_;
  wire _33319_;
  wire _33320_;
  wire _33321_;
  wire _33322_;
  wire _33323_;
  wire _33324_;
  wire _33325_;
  wire _33326_;
  wire _33327_;
  wire _33328_;
  wire _33329_;
  wire _33330_;
  wire _33331_;
  wire _33332_;
  wire _33333_;
  wire _33334_;
  wire _33335_;
  wire _33336_;
  wire _33337_;
  wire _33338_;
  wire _33339_;
  wire _33340_;
  wire _33341_;
  wire _33342_;
  wire _33343_;
  wire _33344_;
  wire _33345_;
  wire _33346_;
  wire _33347_;
  wire _33348_;
  wire _33349_;
  wire _33350_;
  wire _33351_;
  wire _33352_;
  wire _33353_;
  wire _33354_;
  wire _33355_;
  wire _33356_;
  wire _33357_;
  wire _33358_;
  wire _33359_;
  wire _33360_;
  wire _33361_;
  wire _33362_;
  wire _33363_;
  wire _33364_;
  wire _33365_;
  wire _33366_;
  wire _33367_;
  wire _33368_;
  wire _33369_;
  wire _33370_;
  wire _33371_;
  wire _33372_;
  wire _33373_;
  wire _33374_;
  wire _33375_;
  wire _33376_;
  wire _33377_;
  wire _33378_;
  wire _33379_;
  wire _33380_;
  wire _33381_;
  wire _33382_;
  wire _33383_;
  wire _33384_;
  wire _33385_;
  wire _33386_;
  wire _33387_;
  wire _33388_;
  wire _33389_;
  wire _33390_;
  wire _33391_;
  wire _33392_;
  wire _33393_;
  wire _33394_;
  wire _33395_;
  wire _33396_;
  wire _33397_;
  wire _33398_;
  wire _33399_;
  wire _33400_;
  wire _33401_;
  wire _33402_;
  wire _33403_;
  wire _33404_;
  wire _33405_;
  wire _33406_;
  wire _33407_;
  wire _33408_;
  wire _33409_;
  wire _33410_;
  wire _33411_;
  wire _33412_;
  wire _33413_;
  wire _33414_;
  wire _33415_;
  wire _33416_;
  wire _33417_;
  wire _33418_;
  wire _33419_;
  wire _33420_;
  wire _33421_;
  wire _33422_;
  wire _33423_;
  wire _33424_;
  wire _33425_;
  wire _33426_;
  wire _33427_;
  wire _33428_;
  wire _33429_;
  wire _33430_;
  wire _33431_;
  wire _33432_;
  wire _33433_;
  wire _33434_;
  wire _33435_;
  wire _33436_;
  wire _33437_;
  wire _33438_;
  wire _33439_;
  wire _33440_;
  wire _33441_;
  wire _33442_;
  wire _33443_;
  wire _33444_;
  wire _33445_;
  wire _33446_;
  wire _33447_;
  wire _33448_;
  wire _33449_;
  wire _33450_;
  wire _33451_;
  wire _33452_;
  wire _33453_;
  wire _33454_;
  wire _33455_;
  wire _33456_;
  wire _33457_;
  wire _33458_;
  wire _33459_;
  wire _33460_;
  wire _33461_;
  wire _33462_;
  wire _33463_;
  wire _33464_;
  wire _33465_;
  wire _33466_;
  wire _33467_;
  wire _33468_;
  wire _33469_;
  wire _33470_;
  wire _33471_;
  wire _33472_;
  wire _33473_;
  wire _33474_;
  wire _33475_;
  wire _33476_;
  wire _33477_;
  wire _33478_;
  wire _33479_;
  wire _33480_;
  wire _33481_;
  wire _33482_;
  wire _33483_;
  wire _33484_;
  wire _33485_;
  wire _33486_;
  wire _33487_;
  wire _33488_;
  wire _33489_;
  wire _33490_;
  wire _33491_;
  wire _33492_;
  wire _33493_;
  wire _33494_;
  wire _33495_;
  wire _33496_;
  wire _33497_;
  wire _33498_;
  wire _33499_;
  wire _33500_;
  wire _33501_;
  wire _33502_;
  wire _33503_;
  wire _33504_;
  wire _33505_;
  wire _33506_;
  wire _33507_;
  wire _33508_;
  wire _33509_;
  wire _33510_;
  wire _33511_;
  wire _33512_;
  wire _33513_;
  wire _33514_;
  wire _33515_;
  wire _33516_;
  wire _33517_;
  wire _33518_;
  wire _33519_;
  wire _33520_;
  wire _33521_;
  wire _33522_;
  wire _33523_;
  wire _33524_;
  wire _33525_;
  wire _33526_;
  wire _33527_;
  wire _33528_;
  wire _33529_;
  wire _33530_;
  wire _33531_;
  wire _33532_;
  wire _33533_;
  wire _33534_;
  wire _33535_;
  wire _33536_;
  wire _33537_;
  wire _33538_;
  wire _33539_;
  wire _33540_;
  wire _33541_;
  wire _33542_;
  wire _33543_;
  wire _33544_;
  wire _33545_;
  wire _33546_;
  wire _33547_;
  wire _33548_;
  wire _33549_;
  wire _33550_;
  wire _33551_;
  wire _33552_;
  wire _33553_;
  wire _33554_;
  wire _33555_;
  wire _33556_;
  wire _33557_;
  wire _33558_;
  wire _33559_;
  wire _33560_;
  wire _33561_;
  wire _33562_;
  wire _33563_;
  wire _33564_;
  wire _33565_;
  wire _33566_;
  wire _33567_;
  wire _33568_;
  wire _33569_;
  wire _33570_;
  wire _33571_;
  wire _33572_;
  wire _33573_;
  wire _33574_;
  wire _33575_;
  wire _33576_;
  wire _33577_;
  wire _33578_;
  wire _33579_;
  wire _33580_;
  wire _33581_;
  wire _33582_;
  wire _33583_;
  wire _33584_;
  wire _33585_;
  wire _33586_;
  wire _33587_;
  wire _33588_;
  wire _33589_;
  wire _33590_;
  wire _33591_;
  wire _33592_;
  wire _33593_;
  wire _33594_;
  wire _33595_;
  wire _33596_;
  wire _33597_;
  wire _33598_;
  wire _33599_;
  wire _33600_;
  wire _33601_;
  wire _33602_;
  wire _33603_;
  wire _33604_;
  wire _33605_;
  wire _33606_;
  wire _33607_;
  wire _33608_;
  wire _33609_;
  wire _33610_;
  wire _33611_;
  wire _33612_;
  wire _33613_;
  wire _33614_;
  wire _33615_;
  wire _33616_;
  wire _33617_;
  wire _33618_;
  wire _33619_;
  wire _33620_;
  wire _33621_;
  wire _33622_;
  wire _33623_;
  wire _33624_;
  wire _33625_;
  wire _33626_;
  wire _33627_;
  wire _33628_;
  wire _33629_;
  wire _33630_;
  wire _33631_;
  wire _33632_;
  wire _33633_;
  wire _33634_;
  wire _33635_;
  wire _33636_;
  wire _33637_;
  wire _33638_;
  wire _33639_;
  wire _33640_;
  wire _33641_;
  wire _33642_;
  wire _33643_;
  wire _33644_;
  wire _33645_;
  wire _33646_;
  wire _33647_;
  wire _33648_;
  wire _33649_;
  wire _33650_;
  wire _33651_;
  wire _33652_;
  wire _33653_;
  wire _33654_;
  wire _33655_;
  wire _33656_;
  wire _33657_;
  wire _33658_;
  wire _33659_;
  wire _33660_;
  wire _33661_;
  wire _33662_;
  wire _33663_;
  wire _33664_;
  wire _33665_;
  wire _33666_;
  wire _33667_;
  wire _33668_;
  wire _33669_;
  wire _33670_;
  wire _33671_;
  wire _33672_;
  wire _33673_;
  wire _33674_;
  wire _33675_;
  wire _33676_;
  wire _33677_;
  wire _33678_;
  wire _33679_;
  wire _33680_;
  wire _33681_;
  wire _33682_;
  wire _33683_;
  wire _33684_;
  wire _33685_;
  wire _33686_;
  wire _33687_;
  wire _33688_;
  wire _33689_;
  wire _33690_;
  wire _33691_;
  wire _33692_;
  wire _33693_;
  wire _33694_;
  wire _33695_;
  wire _33696_;
  wire _33697_;
  wire _33698_;
  wire _33699_;
  wire _33700_;
  wire _33701_;
  wire _33702_;
  wire _33703_;
  wire _33704_;
  wire _33705_;
  wire _33706_;
  wire _33707_;
  wire _33708_;
  wire _33709_;
  wire _33710_;
  wire _33711_;
  wire _33712_;
  wire _33713_;
  wire _33714_;
  wire _33715_;
  wire _33716_;
  wire _33717_;
  wire _33718_;
  wire _33719_;
  wire _33720_;
  wire _33721_;
  wire _33722_;
  wire _33723_;
  wire _33724_;
  wire _33725_;
  wire _33726_;
  wire _33727_;
  wire _33728_;
  wire _33729_;
  wire _33730_;
  wire _33731_;
  wire _33732_;
  wire _33733_;
  wire _33734_;
  wire _33735_;
  wire _33736_;
  wire _33737_;
  wire _33738_;
  wire _33739_;
  wire _33740_;
  wire _33741_;
  wire _33742_;
  wire _33743_;
  wire _33744_;
  wire _33745_;
  wire _33746_;
  wire _33747_;
  wire _33748_;
  wire _33749_;
  wire _33750_;
  wire _33751_;
  wire _33752_;
  wire _33753_;
  wire _33754_;
  wire _33755_;
  wire _33756_;
  wire _33757_;
  wire _33758_;
  wire _33759_;
  wire _33760_;
  wire _33761_;
  wire _33762_;
  wire _33763_;
  wire _33764_;
  wire _33765_;
  wire _33766_;
  wire _33767_;
  wire _33768_;
  wire _33769_;
  wire _33770_;
  wire _33771_;
  wire _33772_;
  wire _33773_;
  wire _33774_;
  wire _33775_;
  wire _33776_;
  wire _33777_;
  wire _33778_;
  wire _33779_;
  wire _33780_;
  wire _33781_;
  wire _33782_;
  wire _33783_;
  wire _33784_;
  wire _33785_;
  wire _33786_;
  wire _33787_;
  wire _33788_;
  wire _33789_;
  wire _33790_;
  wire _33791_;
  wire _33792_;
  wire _33793_;
  wire _33794_;
  wire _33795_;
  wire _33796_;
  wire _33797_;
  wire _33798_;
  wire _33799_;
  wire _33800_;
  wire _33801_;
  wire _33802_;
  wire _33803_;
  wire _33804_;
  wire _33805_;
  wire _33806_;
  wire _33807_;
  wire _33808_;
  wire _33809_;
  wire _33810_;
  wire _33811_;
  wire _33812_;
  wire _33813_;
  wire _33814_;
  wire _33815_;
  wire _33816_;
  wire _33817_;
  wire _33818_;
  wire _33819_;
  wire _33820_;
  wire _33821_;
  wire _33822_;
  wire _33823_;
  wire _33824_;
  wire _33825_;
  wire _33826_;
  wire _33827_;
  wire _33828_;
  wire _33829_;
  wire _33830_;
  wire _33831_;
  wire _33832_;
  wire _33833_;
  wire _33834_;
  wire _33835_;
  wire _33836_;
  wire _33837_;
  wire _33838_;
  wire _33839_;
  wire _33840_;
  wire _33841_;
  wire _33842_;
  wire _33843_;
  wire _33844_;
  wire _33845_;
  wire _33846_;
  wire _33847_;
  wire _33848_;
  wire _33849_;
  wire _33850_;
  wire _33851_;
  wire _33852_;
  wire _33853_;
  wire _33854_;
  wire _33855_;
  wire _33856_;
  wire _33857_;
  wire _33858_;
  wire _33859_;
  wire _33860_;
  wire _33861_;
  wire _33862_;
  wire _33863_;
  wire _33864_;
  wire _33865_;
  wire _33866_;
  wire _33867_;
  wire _33868_;
  wire _33869_;
  wire _33870_;
  wire _33871_;
  wire _33872_;
  wire _33873_;
  wire _33874_;
  wire _33875_;
  wire _33876_;
  wire _33877_;
  wire _33878_;
  wire _33879_;
  wire _33880_;
  wire _33881_;
  wire _33882_;
  wire _33883_;
  wire _33884_;
  wire _33885_;
  wire _33886_;
  wire _33887_;
  wire _33888_;
  wire _33889_;
  wire _33890_;
  wire _33891_;
  wire _33892_;
  wire _33893_;
  wire _33894_;
  wire _33895_;
  wire _33896_;
  wire _33897_;
  wire _33898_;
  wire _33899_;
  wire _33900_;
  wire _33901_;
  wire _33902_;
  wire _33903_;
  wire _33904_;
  wire _33905_;
  wire _33906_;
  wire _33907_;
  wire _33908_;
  wire _33909_;
  wire _33910_;
  wire _33911_;
  wire _33912_;
  wire _33913_;
  wire _33914_;
  wire _33915_;
  wire _33916_;
  wire _33917_;
  wire _33918_;
  wire _33919_;
  wire _33920_;
  wire _33921_;
  wire _33922_;
  wire _33923_;
  wire _33924_;
  wire _33925_;
  wire _33926_;
  wire _33927_;
  wire _33928_;
  wire _33929_;
  wire _33930_;
  wire _33931_;
  wire _33932_;
  wire _33933_;
  wire _33934_;
  wire _33935_;
  wire _33936_;
  wire _33937_;
  wire _33938_;
  wire _33939_;
  wire _33940_;
  wire _33941_;
  wire _33942_;
  wire _33943_;
  wire _33944_;
  wire _33945_;
  wire _33946_;
  wire _33947_;
  wire _33948_;
  wire _33949_;
  wire _33950_;
  wire _33951_;
  wire _33952_;
  wire _33953_;
  wire _33954_;
  wire _33955_;
  wire _33956_;
  wire _33957_;
  wire _33958_;
  wire _33959_;
  wire _33960_;
  wire _33961_;
  wire _33962_;
  wire _33963_;
  wire _33964_;
  wire _33965_;
  wire _33966_;
  wire _33967_;
  wire _33968_;
  wire _33969_;
  wire _33970_;
  wire _33971_;
  wire _33972_;
  wire _33973_;
  wire _33974_;
  wire _33975_;
  wire _33976_;
  wire _33977_;
  wire _33978_;
  wire _33979_;
  wire _33980_;
  wire _33981_;
  wire _33982_;
  wire _33983_;
  wire _33984_;
  wire _33985_;
  wire _33986_;
  wire _33987_;
  wire _33988_;
  wire _33989_;
  wire _33990_;
  wire _33991_;
  wire _33992_;
  wire _33993_;
  wire _33994_;
  wire _33995_;
  wire _33996_;
  wire _33997_;
  wire _33998_;
  wire _33999_;
  wire _34000_;
  wire _34001_;
  wire _34002_;
  wire _34003_;
  wire _34004_;
  wire _34005_;
  wire _34006_;
  wire _34007_;
  wire _34008_;
  wire _34009_;
  wire _34010_;
  wire _34011_;
  wire _34012_;
  wire _34013_;
  wire _34014_;
  wire _34015_;
  wire _34016_;
  wire _34017_;
  wire _34018_;
  wire _34019_;
  wire _34020_;
  wire _34021_;
  wire _34022_;
  wire _34023_;
  wire _34024_;
  wire _34025_;
  wire _34026_;
  wire _34027_;
  wire _34028_;
  wire _34029_;
  wire _34030_;
  wire _34031_;
  wire _34032_;
  wire _34033_;
  wire _34034_;
  wire _34035_;
  wire _34036_;
  wire _34037_;
  wire _34038_;
  wire _34039_;
  wire _34040_;
  wire _34041_;
  wire _34042_;
  wire _34043_;
  wire _34044_;
  wire _34045_;
  wire _34046_;
  wire _34047_;
  wire _34048_;
  wire _34049_;
  wire _34050_;
  wire _34051_;
  wire _34052_;
  wire _34053_;
  wire _34054_;
  wire _34055_;
  wire _34056_;
  wire _34057_;
  wire _34058_;
  wire _34059_;
  wire _34060_;
  wire _34061_;
  wire _34062_;
  wire _34063_;
  wire _34064_;
  wire _34065_;
  wire _34066_;
  wire _34067_;
  wire _34068_;
  wire _34069_;
  wire _34070_;
  wire _34071_;
  wire _34072_;
  wire _34073_;
  wire _34074_;
  wire _34075_;
  wire _34076_;
  wire _34077_;
  wire _34078_;
  wire _34079_;
  wire _34080_;
  wire _34081_;
  wire _34082_;
  wire _34083_;
  wire _34084_;
  wire _34085_;
  wire _34086_;
  wire _34087_;
  wire _34088_;
  wire _34089_;
  wire _34090_;
  wire _34091_;
  wire _34092_;
  wire _34093_;
  wire _34094_;
  wire _34095_;
  wire _34096_;
  wire _34097_;
  wire _34098_;
  wire _34099_;
  wire _34100_;
  wire _34101_;
  wire _34102_;
  wire _34103_;
  wire _34104_;
  wire _34105_;
  wire _34106_;
  wire _34107_;
  wire _34108_;
  wire _34109_;
  wire _34110_;
  wire _34111_;
  wire _34112_;
  wire _34113_;
  wire _34114_;
  wire _34115_;
  wire _34116_;
  wire _34117_;
  wire _34118_;
  wire _34119_;
  wire _34120_;
  wire _34121_;
  wire _34122_;
  wire _34123_;
  wire _34124_;
  wire _34125_;
  wire _34126_;
  wire _34127_;
  wire _34128_;
  wire _34129_;
  wire _34130_;
  wire _34131_;
  wire _34132_;
  wire _34133_;
  wire _34134_;
  wire _34135_;
  wire _34136_;
  wire _34137_;
  wire _34138_;
  wire _34139_;
  wire _34140_;
  wire _34141_;
  wire _34142_;
  wire _34143_;
  wire _34144_;
  wire _34145_;
  wire _34146_;
  wire _34147_;
  wire _34148_;
  wire _34149_;
  wire _34150_;
  wire _34151_;
  wire _34152_;
  wire _34153_;
  wire _34154_;
  wire _34155_;
  wire _34156_;
  wire _34157_;
  wire _34158_;
  wire _34159_;
  wire _34160_;
  wire _34161_;
  wire _34162_;
  wire _34163_;
  wire _34164_;
  wire _34165_;
  wire _34166_;
  wire _34167_;
  wire _34168_;
  wire _34169_;
  wire _34170_;
  wire _34171_;
  wire _34172_;
  wire _34173_;
  wire _34174_;
  wire _34175_;
  wire _34176_;
  wire _34177_;
  wire _34178_;
  wire _34179_;
  wire _34180_;
  wire _34181_;
  wire _34182_;
  wire _34183_;
  wire _34184_;
  wire _34185_;
  wire _34186_;
  wire _34187_;
  wire _34188_;
  wire _34189_;
  wire _34190_;
  wire _34191_;
  wire _34192_;
  wire _34193_;
  wire _34194_;
  wire _34195_;
  wire _34196_;
  wire _34197_;
  wire _34198_;
  wire _34199_;
  wire _34200_;
  wire _34201_;
  wire _34202_;
  wire _34203_;
  wire _34204_;
  wire _34205_;
  wire _34206_;
  wire _34207_;
  wire _34208_;
  wire _34209_;
  wire _34210_;
  wire _34211_;
  wire _34212_;
  wire _34213_;
  wire _34214_;
  wire _34215_;
  wire _34216_;
  wire _34217_;
  wire _34218_;
  wire _34219_;
  wire _34220_;
  wire _34221_;
  wire _34222_;
  wire _34223_;
  wire _34224_;
  wire _34225_;
  wire _34226_;
  wire _34227_;
  wire _34228_;
  wire _34229_;
  wire _34230_;
  wire _34231_;
  wire _34232_;
  wire _34233_;
  wire _34234_;
  wire _34235_;
  wire _34236_;
  wire _34237_;
  wire _34238_;
  wire _34239_;
  wire _34240_;
  wire _34241_;
  wire _34242_;
  wire _34243_;
  wire _34244_;
  wire _34245_;
  wire _34246_;
  wire _34247_;
  wire _34248_;
  wire _34249_;
  wire _34250_;
  wire _34251_;
  wire _34252_;
  wire _34253_;
  wire _34254_;
  wire _34255_;
  wire _34256_;
  wire _34257_;
  wire _34258_;
  wire _34259_;
  wire _34260_;
  wire _34261_;
  wire _34262_;
  wire _34263_;
  wire _34264_;
  wire _34265_;
  wire _34266_;
  wire _34267_;
  wire _34268_;
  wire _34269_;
  wire _34270_;
  wire _34271_;
  wire _34272_;
  wire _34273_;
  wire _34274_;
  wire _34275_;
  wire _34276_;
  wire _34277_;
  wire _34278_;
  wire _34279_;
  wire _34280_;
  wire _34281_;
  wire _34282_;
  wire _34283_;
  wire _34284_;
  wire _34285_;
  wire _34286_;
  wire _34287_;
  wire _34288_;
  wire _34289_;
  wire _34290_;
  wire _34291_;
  wire _34292_;
  wire _34293_;
  wire _34294_;
  wire _34295_;
  wire _34296_;
  wire _34297_;
  wire _34298_;
  wire _34299_;
  wire _34300_;
  wire _34301_;
  wire _34302_;
  wire _34303_;
  wire _34304_;
  wire _34305_;
  wire _34306_;
  wire _34307_;
  wire _34308_;
  wire _34309_;
  wire _34310_;
  wire _34311_;
  wire _34312_;
  wire _34313_;
  wire _34314_;
  wire _34315_;
  wire _34316_;
  wire _34317_;
  wire _34318_;
  wire _34319_;
  wire _34320_;
  wire _34321_;
  wire _34322_;
  wire _34323_;
  wire _34324_;
  wire _34325_;
  wire _34326_;
  wire _34327_;
  wire _34328_;
  wire _34329_;
  wire _34330_;
  wire _34331_;
  wire _34332_;
  wire _34333_;
  wire _34334_;
  wire _34335_;
  wire _34336_;
  wire _34337_;
  wire _34338_;
  wire _34339_;
  wire _34340_;
  wire _34341_;
  wire _34342_;
  wire _34343_;
  wire _34344_;
  wire _34345_;
  wire _34346_;
  wire _34347_;
  wire _34348_;
  wire _34349_;
  wire _34350_;
  wire _34351_;
  wire _34352_;
  wire _34353_;
  wire _34354_;
  wire _34355_;
  wire _34356_;
  wire _34357_;
  wire _34358_;
  wire _34359_;
  wire _34360_;
  wire _34361_;
  wire _34362_;
  wire _34363_;
  wire _34364_;
  wire _34365_;
  wire _34366_;
  wire _34367_;
  wire _34368_;
  wire _34369_;
  wire _34370_;
  wire _34371_;
  wire _34372_;
  wire _34373_;
  wire _34374_;
  wire _34375_;
  wire _34376_;
  wire _34377_;
  wire _34378_;
  wire _34379_;
  wire _34380_;
  wire _34381_;
  wire _34382_;
  wire _34383_;
  wire _34384_;
  wire _34385_;
  wire _34386_;
  wire _34387_;
  wire _34388_;
  wire _34389_;
  wire _34390_;
  wire _34391_;
  wire _34392_;
  wire _34393_;
  wire _34394_;
  wire _34395_;
  wire _34396_;
  wire _34397_;
  wire _34398_;
  wire _34399_;
  wire _34400_;
  wire _34401_;
  wire _34402_;
  wire _34403_;
  wire _34404_;
  wire _34405_;
  wire _34406_;
  wire _34407_;
  wire _34408_;
  wire _34409_;
  wire _34410_;
  wire _34411_;
  wire _34412_;
  wire _34413_;
  wire _34414_;
  wire _34415_;
  wire _34416_;
  wire _34417_;
  wire _34418_;
  wire _34419_;
  wire _34420_;
  wire _34421_;
  wire _34422_;
  wire _34423_;
  wire _34424_;
  wire _34425_;
  wire _34426_;
  wire _34427_;
  wire _34428_;
  wire _34429_;
  wire _34430_;
  wire _34431_;
  wire _34432_;
  wire _34433_;
  wire _34434_;
  wire _34435_;
  wire _34436_;
  wire _34437_;
  wire _34438_;
  wire _34439_;
  wire _34440_;
  wire _34441_;
  wire _34442_;
  wire _34443_;
  wire _34444_;
  wire _34445_;
  wire _34446_;
  wire _34447_;
  wire _34448_;
  wire _34449_;
  wire _34450_;
  wire _34451_;
  wire _34452_;
  wire _34453_;
  wire _34454_;
  wire _34455_;
  wire _34456_;
  wire _34457_;
  wire _34458_;
  wire _34459_;
  wire _34460_;
  wire _34461_;
  wire _34462_;
  wire _34463_;
  wire _34464_;
  wire _34465_;
  wire _34466_;
  wire _34467_;
  wire _34468_;
  wire _34469_;
  wire _34470_;
  wire _34471_;
  wire _34472_;
  wire _34473_;
  wire _34474_;
  wire _34475_;
  wire _34476_;
  wire _34477_;
  wire _34478_;
  wire _34479_;
  wire _34480_;
  wire _34481_;
  wire _34482_;
  wire _34483_;
  wire _34484_;
  wire _34485_;
  wire _34486_;
  wire _34487_;
  wire _34488_;
  wire _34489_;
  wire _34490_;
  wire _34491_;
  wire _34492_;
  wire _34493_;
  wire _34494_;
  wire _34495_;
  wire _34496_;
  wire _34497_;
  wire _34498_;
  wire _34499_;
  wire _34500_;
  wire _34501_;
  wire _34502_;
  wire _34503_;
  wire _34504_;
  wire _34505_;
  wire _34506_;
  wire _34507_;
  wire _34508_;
  wire _34509_;
  wire _34510_;
  wire _34511_;
  wire _34512_;
  wire _34513_;
  wire _34514_;
  wire _34515_;
  wire _34516_;
  wire _34517_;
  wire _34518_;
  wire _34519_;
  wire _34520_;
  wire _34521_;
  wire _34522_;
  wire _34523_;
  wire _34524_;
  wire _34525_;
  wire _34526_;
  wire _34527_;
  wire _34528_;
  wire _34529_;
  wire _34530_;
  wire _34531_;
  wire _34532_;
  wire _34533_;
  wire _34534_;
  wire _34535_;
  wire _34536_;
  wire _34537_;
  wire _34538_;
  wire _34539_;
  wire _34540_;
  wire _34541_;
  wire _34542_;
  wire _34543_;
  wire _34544_;
  wire _34545_;
  wire _34546_;
  wire _34547_;
  wire _34548_;
  wire _34549_;
  wire _34550_;
  wire _34551_;
  wire _34552_;
  wire _34553_;
  wire _34554_;
  wire _34555_;
  wire _34556_;
  wire _34557_;
  wire _34558_;
  wire _34559_;
  wire _34560_;
  wire _34561_;
  wire _34562_;
  wire _34563_;
  wire _34564_;
  wire _34565_;
  wire _34566_;
  wire _34567_;
  wire _34568_;
  wire _34569_;
  wire _34570_;
  wire _34571_;
  wire _34572_;
  wire _34573_;
  wire _34574_;
  wire _34575_;
  wire _34576_;
  wire _34577_;
  wire _34578_;
  wire _34579_;
  wire _34580_;
  wire _34581_;
  wire _34582_;
  wire _34583_;
  wire _34584_;
  wire _34585_;
  wire _34586_;
  wire _34587_;
  wire _34588_;
  wire _34589_;
  wire _34590_;
  wire _34591_;
  wire _34592_;
  wire _34593_;
  wire _34594_;
  wire _34595_;
  wire _34596_;
  wire _34597_;
  wire _34598_;
  wire _34599_;
  wire _34600_;
  wire _34601_;
  wire _34602_;
  wire _34603_;
  wire _34604_;
  wire _34605_;
  wire _34606_;
  wire _34607_;
  wire _34608_;
  wire _34609_;
  wire _34610_;
  wire _34611_;
  wire _34612_;
  wire _34613_;
  wire _34614_;
  wire _34615_;
  wire _34616_;
  wire _34617_;
  wire _34618_;
  wire _34619_;
  wire _34620_;
  wire _34621_;
  wire _34622_;
  wire _34623_;
  wire _34624_;
  wire _34625_;
  wire _34626_;
  wire _34627_;
  wire _34628_;
  wire _34629_;
  wire _34630_;
  wire _34631_;
  wire _34632_;
  wire _34633_;
  wire _34634_;
  wire _34635_;
  wire _34636_;
  wire _34637_;
  wire _34638_;
  wire _34639_;
  wire _34640_;
  wire _34641_;
  wire _34642_;
  wire _34643_;
  wire _34644_;
  wire _34645_;
  wire _34646_;
  wire _34647_;
  wire _34648_;
  wire _34649_;
  wire _34650_;
  wire _34651_;
  wire _34652_;
  wire _34653_;
  wire _34654_;
  wire _34655_;
  wire _34656_;
  wire _34657_;
  wire _34658_;
  wire _34659_;
  wire _34660_;
  wire _34661_;
  wire _34662_;
  wire _34663_;
  wire _34664_;
  wire _34665_;
  wire _34666_;
  wire _34667_;
  wire _34668_;
  wire _34669_;
  wire _34670_;
  wire _34671_;
  wire _34672_;
  wire _34673_;
  wire _34674_;
  wire _34675_;
  wire _34676_;
  wire _34677_;
  wire _34678_;
  wire _34679_;
  wire _34680_;
  wire _34681_;
  wire _34682_;
  wire _34683_;
  wire _34684_;
  wire _34685_;
  wire _34686_;
  wire _34687_;
  wire _34688_;
  wire _34689_;
  wire _34690_;
  wire _34691_;
  wire _34692_;
  wire _34693_;
  wire _34694_;
  wire _34695_;
  wire _34696_;
  wire _34697_;
  wire _34698_;
  wire _34699_;
  wire _34700_;
  wire _34701_;
  wire _34702_;
  wire _34703_;
  wire _34704_;
  wire _34705_;
  wire _34706_;
  wire _34707_;
  wire _34708_;
  wire _34709_;
  wire _34710_;
  wire _34711_;
  wire _34712_;
  wire _34713_;
  wire _34714_;
  wire _34715_;
  wire _34716_;
  wire _34717_;
  wire _34718_;
  wire _34719_;
  wire _34720_;
  wire _34721_;
  wire _34722_;
  wire _34723_;
  wire _34724_;
  wire _34725_;
  wire _34726_;
  wire _34727_;
  wire _34728_;
  wire _34729_;
  wire _34730_;
  wire _34731_;
  wire _34732_;
  wire _34733_;
  wire _34734_;
  wire _34735_;
  wire _34736_;
  wire _34737_;
  wire _34738_;
  wire _34739_;
  wire _34740_;
  wire _34741_;
  wire _34742_;
  wire _34743_;
  wire _34744_;
  wire _34745_;
  wire _34746_;
  wire _34747_;
  wire _34748_;
  wire _34749_;
  wire _34750_;
  wire _34751_;
  wire _34752_;
  wire _34753_;
  wire _34754_;
  wire _34755_;
  wire _34756_;
  wire _34757_;
  wire _34758_;
  wire _34759_;
  wire _34760_;
  wire _34761_;
  wire _34762_;
  wire _34763_;
  wire _34764_;
  wire _34765_;
  wire _34766_;
  wire _34767_;
  wire _34768_;
  wire _34769_;
  wire _34770_;
  wire _34771_;
  wire _34772_;
  wire _34773_;
  wire _34774_;
  wire _34775_;
  wire _34776_;
  wire _34777_;
  wire _34778_;
  wire _34779_;
  wire _34780_;
  wire _34781_;
  wire _34782_;
  wire _34783_;
  wire _34784_;
  wire _34785_;
  wire _34786_;
  wire _34787_;
  wire _34788_;
  wire _34789_;
  wire _34790_;
  wire _34791_;
  wire _34792_;
  wire _34793_;
  wire _34794_;
  wire _34795_;
  wire _34796_;
  wire _34797_;
  wire _34798_;
  wire _34799_;
  wire _34800_;
  wire _34801_;
  wire _34802_;
  wire _34803_;
  wire _34804_;
  wire _34805_;
  wire _34806_;
  wire _34807_;
  wire _34808_;
  wire _34809_;
  wire _34810_;
  wire _34811_;
  wire _34812_;
  wire _34813_;
  wire _34814_;
  wire _34815_;
  wire _34816_;
  wire _34817_;
  wire _34818_;
  wire _34819_;
  wire _34820_;
  wire _34821_;
  wire _34822_;
  wire _34823_;
  wire _34824_;
  wire _34825_;
  wire _34826_;
  wire _34827_;
  wire _34828_;
  wire _34829_;
  wire _34830_;
  wire _34831_;
  wire _34832_;
  wire _34833_;
  wire _34834_;
  wire _34835_;
  wire _34836_;
  wire _34837_;
  wire _34838_;
  wire _34839_;
  wire _34840_;
  wire _34841_;
  wire _34842_;
  wire _34843_;
  wire _34844_;
  wire _34845_;
  wire _34846_;
  wire _34847_;
  wire _34848_;
  wire _34849_;
  wire _34850_;
  wire _34851_;
  wire _34852_;
  wire _34853_;
  wire _34854_;
  wire _34855_;
  wire _34856_;
  wire _34857_;
  wire _34858_;
  wire _34859_;
  wire _34860_;
  wire _34861_;
  wire _34862_;
  wire _34863_;
  wire _34864_;
  wire _34865_;
  wire _34866_;
  wire _34867_;
  wire _34868_;
  wire _34869_;
  wire _34870_;
  wire _34871_;
  wire _34872_;
  wire _34873_;
  wire _34874_;
  wire _34875_;
  wire _34876_;
  wire _34877_;
  wire _34878_;
  wire _34879_;
  wire _34880_;
  wire _34881_;
  wire _34882_;
  wire _34883_;
  wire _34884_;
  wire _34885_;
  wire _34886_;
  wire _34887_;
  wire _34888_;
  wire _34889_;
  wire _34890_;
  wire _34891_;
  wire _34892_;
  wire _34893_;
  wire _34894_;
  wire _34895_;
  wire _34896_;
  wire _34897_;
  wire _34898_;
  wire _34899_;
  wire _34900_;
  wire _34901_;
  wire _34902_;
  wire _34903_;
  wire _34904_;
  wire _34905_;
  wire _34906_;
  wire _34907_;
  wire _34908_;
  wire _34909_;
  wire _34910_;
  wire _34911_;
  wire _34912_;
  wire _34913_;
  wire _34914_;
  wire _34915_;
  wire _34916_;
  wire _34917_;
  wire _34918_;
  wire _34919_;
  wire _34920_;
  wire _34921_;
  wire _34922_;
  wire _34923_;
  wire _34924_;
  wire _34925_;
  wire _34926_;
  wire _34927_;
  wire _34928_;
  wire _34929_;
  wire _34930_;
  wire _34931_;
  wire _34932_;
  wire _34933_;
  wire _34934_;
  wire _34935_;
  wire _34936_;
  wire _34937_;
  wire _34938_;
  wire _34939_;
  wire _34940_;
  wire _34941_;
  wire _34942_;
  wire _34943_;
  wire _34944_;
  wire _34945_;
  wire _34946_;
  wire _34947_;
  wire _34948_;
  wire _34949_;
  wire _34950_;
  wire _34951_;
  wire _34952_;
  wire _34953_;
  wire _34954_;
  wire _34955_;
  wire _34956_;
  wire _34957_;
  wire _34958_;
  wire _34959_;
  wire _34960_;
  wire _34961_;
  wire _34962_;
  wire _34963_;
  wire _34964_;
  wire _34965_;
  wire _34966_;
  wire _34967_;
  wire _34968_;
  wire _34969_;
  wire _34970_;
  wire _34971_;
  wire _34972_;
  wire _34973_;
  wire _34974_;
  wire _34975_;
  wire _34976_;
  wire _34977_;
  wire _34978_;
  wire _34979_;
  wire _34980_;
  wire _34981_;
  wire _34982_;
  wire _34983_;
  wire _34984_;
  wire _34985_;
  wire _34986_;
  wire _34987_;
  wire _34988_;
  wire _34989_;
  wire _34990_;
  wire _34991_;
  wire _34992_;
  wire _34993_;
  wire _34994_;
  wire _34995_;
  wire _34996_;
  wire _34997_;
  wire _34998_;
  wire _34999_;
  wire _35000_;
  wire _35001_;
  wire _35002_;
  wire _35003_;
  wire _35004_;
  wire _35005_;
  wire _35006_;
  wire _35007_;
  wire _35008_;
  wire _35009_;
  wire _35010_;
  wire _35011_;
  wire _35012_;
  wire _35013_;
  wire _35014_;
  wire _35015_;
  wire _35016_;
  wire _35017_;
  wire _35018_;
  wire _35019_;
  wire _35020_;
  wire _35021_;
  wire _35022_;
  wire _35023_;
  wire _35024_;
  wire _35025_;
  wire _35026_;
  wire _35027_;
  wire _35028_;
  wire _35029_;
  wire _35030_;
  wire _35031_;
  wire _35032_;
  wire _35033_;
  wire _35034_;
  wire _35035_;
  wire _35036_;
  wire _35037_;
  wire _35038_;
  wire _35039_;
  wire _35040_;
  wire _35041_;
  wire _35042_;
  wire _35043_;
  wire _35044_;
  wire _35045_;
  wire _35046_;
  wire _35047_;
  wire _35048_;
  wire _35049_;
  wire _35050_;
  wire _35051_;
  wire _35052_;
  wire _35053_;
  wire _35054_;
  wire _35055_;
  wire _35056_;
  wire _35057_;
  wire _35058_;
  wire _35059_;
  wire _35060_;
  wire _35061_;
  wire _35062_;
  wire _35063_;
  wire _35064_;
  wire _35065_;
  wire _35066_;
  wire _35067_;
  wire _35068_;
  wire _35069_;
  wire _35070_;
  wire _35071_;
  wire _35072_;
  wire _35073_;
  wire _35074_;
  wire _35075_;
  wire _35076_;
  wire _35077_;
  wire _35078_;
  wire _35079_;
  wire _35080_;
  wire _35081_;
  wire _35082_;
  wire _35083_;
  wire _35084_;
  wire _35085_;
  wire _35086_;
  wire _35087_;
  wire _35088_;
  wire _35089_;
  wire _35090_;
  wire _35091_;
  wire _35092_;
  wire _35093_;
  wire _35094_;
  wire _35095_;
  wire _35096_;
  wire _35097_;
  wire _35098_;
  wire _35099_;
  wire _35100_;
  wire _35101_;
  wire _35102_;
  wire _35103_;
  wire _35104_;
  wire _35105_;
  wire _35106_;
  wire _35107_;
  wire _35108_;
  wire _35109_;
  wire _35110_;
  wire _35111_;
  wire _35112_;
  wire _35113_;
  wire _35114_;
  wire _35115_;
  wire _35116_;
  wire _35117_;
  wire _35118_;
  wire _35119_;
  wire _35120_;
  wire _35121_;
  wire _35122_;
  wire _35123_;
  wire _35124_;
  wire _35125_;
  wire _35126_;
  wire _35127_;
  wire _35128_;
  wire _35129_;
  wire _35130_;
  wire _35131_;
  wire _35132_;
  wire _35133_;
  wire _35134_;
  wire _35135_;
  wire _35136_;
  wire _35137_;
  wire _35138_;
  wire _35139_;
  wire _35140_;
  wire _35141_;
  wire _35142_;
  wire _35143_;
  wire _35144_;
  wire _35145_;
  wire _35146_;
  wire _35147_;
  wire _35148_;
  wire _35149_;
  wire _35150_;
  wire _35151_;
  wire _35152_;
  wire _35153_;
  wire _35154_;
  wire _35155_;
  wire _35156_;
  wire _35157_;
  wire _35158_;
  wire _35159_;
  wire _35160_;
  wire _35161_;
  wire _35162_;
  wire _35163_;
  wire _35164_;
  wire _35165_;
  wire _35166_;
  wire _35167_;
  wire _35168_;
  wire _35169_;
  wire _35170_;
  wire _35171_;
  wire _35172_;
  wire _35173_;
  wire _35174_;
  wire _35175_;
  wire _35176_;
  wire _35177_;
  wire _35178_;
  wire _35179_;
  wire _35180_;
  wire _35181_;
  wire _35182_;
  wire _35183_;
  wire _35184_;
  wire _35185_;
  wire _35186_;
  wire _35187_;
  wire _35188_;
  wire _35189_;
  wire _35190_;
  wire _35191_;
  wire _35192_;
  wire _35193_;
  wire _35194_;
  wire _35195_;
  wire _35196_;
  wire _35197_;
  wire _35198_;
  wire _35199_;
  wire _35200_;
  wire _35201_;
  wire _35202_;
  wire _35203_;
  wire _35204_;
  wire _35205_;
  wire _35206_;
  wire _35207_;
  wire _35208_;
  wire _35209_;
  wire _35210_;
  wire _35211_;
  wire _35212_;
  wire _35213_;
  wire _35214_;
  wire _35215_;
  wire _35216_;
  wire _35217_;
  wire _35218_;
  wire _35219_;
  wire _35220_;
  wire _35221_;
  wire _35222_;
  wire _35223_;
  wire _35224_;
  wire _35225_;
  wire _35226_;
  wire _35227_;
  wire _35228_;
  wire _35229_;
  wire _35230_;
  wire _35231_;
  wire _35232_;
  wire _35233_;
  wire _35234_;
  wire _35235_;
  wire _35236_;
  wire _35237_;
  wire _35238_;
  wire _35239_;
  wire _35240_;
  wire _35241_;
  wire _35242_;
  wire _35243_;
  wire _35244_;
  wire _35245_;
  wire _35246_;
  wire _35247_;
  wire _35248_;
  wire _35249_;
  wire _35250_;
  wire _35251_;
  wire _35252_;
  wire _35253_;
  wire _35254_;
  wire _35255_;
  wire _35256_;
  wire _35257_;
  wire _35258_;
  wire _35259_;
  wire _35260_;
  wire _35261_;
  wire _35262_;
  wire _35263_;
  wire _35264_;
  wire _35265_;
  wire _35266_;
  wire _35267_;
  wire _35268_;
  wire _35269_;
  wire _35270_;
  wire _35271_;
  wire _35272_;
  wire _35273_;
  wire _35274_;
  wire _35275_;
  wire _35276_;
  wire _35277_;
  wire _35278_;
  wire _35279_;
  wire _35280_;
  wire _35281_;
  wire _35282_;
  wire _35283_;
  wire _35284_;
  wire _35285_;
  wire _35286_;
  wire _35287_;
  wire _35288_;
  wire _35289_;
  wire _35290_;
  wire _35291_;
  wire _35292_;
  wire _35293_;
  wire _35294_;
  wire _35295_;
  wire _35296_;
  wire _35297_;
  wire _35298_;
  wire _35299_;
  wire _35300_;
  wire _35301_;
  wire _35302_;
  wire _35303_;
  wire _35304_;
  wire _35305_;
  wire _35306_;
  wire _35307_;
  wire _35308_;
  wire _35309_;
  wire _35310_;
  wire _35311_;
  wire _35312_;
  wire _35313_;
  wire _35314_;
  wire _35315_;
  wire _35316_;
  wire _35317_;
  wire _35318_;
  wire _35319_;
  wire _35320_;
  wire _35321_;
  wire _35322_;
  wire _35323_;
  wire _35324_;
  wire _35325_;
  wire _35326_;
  wire _35327_;
  wire _35328_;
  wire _35329_;
  wire _35330_;
  wire _35331_;
  wire _35332_;
  wire _35333_;
  wire _35334_;
  wire _35335_;
  wire _35336_;
  wire _35337_;
  wire _35338_;
  wire _35339_;
  wire _35340_;
  wire _35341_;
  wire _35342_;
  wire _35343_;
  wire _35344_;
  wire _35345_;
  wire _35346_;
  wire _35347_;
  wire _35348_;
  wire _35349_;
  wire _35350_;
  wire _35351_;
  wire _35352_;
  wire _35353_;
  wire _35354_;
  wire _35355_;
  wire _35356_;
  wire _35357_;
  wire _35358_;
  wire _35359_;
  wire _35360_;
  wire _35361_;
  wire _35362_;
  wire _35363_;
  wire _35364_;
  wire _35365_;
  wire _35366_;
  wire _35367_;
  wire _35368_;
  wire _35369_;
  wire _35370_;
  wire _35371_;
  wire _35372_;
  wire _35373_;
  wire _35374_;
  wire _35375_;
  wire _35376_;
  wire _35377_;
  wire _35378_;
  wire _35379_;
  wire _35380_;
  wire _35381_;
  wire _35382_;
  wire _35383_;
  wire _35384_;
  wire _35385_;
  wire _35386_;
  wire _35387_;
  wire _35388_;
  wire _35389_;
  wire _35390_;
  wire _35391_;
  wire _35392_;
  wire _35393_;
  wire _35394_;
  wire _35395_;
  wire _35396_;
  wire _35397_;
  wire _35398_;
  wire _35399_;
  wire _35400_;
  wire _35401_;
  wire _35402_;
  wire _35403_;
  wire _35404_;
  wire _35405_;
  wire _35406_;
  wire _35407_;
  wire _35408_;
  wire _35409_;
  wire _35410_;
  wire _35411_;
  wire _35412_;
  wire _35413_;
  wire _35414_;
  wire _35415_;
  wire _35416_;
  wire _35417_;
  wire _35418_;
  wire _35419_;
  wire _35420_;
  wire _35421_;
  wire _35422_;
  wire _35423_;
  wire _35424_;
  wire _35425_;
  wire _35426_;
  wire _35427_;
  wire _35428_;
  wire _35429_;
  wire _35430_;
  wire _35431_;
  wire _35432_;
  wire _35433_;
  wire _35434_;
  wire _35435_;
  wire _35436_;
  wire _35437_;
  wire _35438_;
  wire _35439_;
  wire _35440_;
  wire _35441_;
  wire _35442_;
  wire _35443_;
  wire _35444_;
  wire _35445_;
  wire _35446_;
  wire _35447_;
  wire _35448_;
  wire _35449_;
  wire _35450_;
  wire _35451_;
  wire _35452_;
  wire _35453_;
  wire _35454_;
  wire _35455_;
  wire _35456_;
  wire _35457_;
  wire _35458_;
  wire _35459_;
  wire _35460_;
  wire _35461_;
  wire _35462_;
  wire _35463_;
  wire _35464_;
  wire _35465_;
  wire _35466_;
  wire _35467_;
  wire _35468_;
  wire _35469_;
  wire _35470_;
  wire _35471_;
  wire _35472_;
  wire _35473_;
  wire _35474_;
  wire _35475_;
  wire _35476_;
  wire _35477_;
  wire _35478_;
  wire _35479_;
  wire _35480_;
  wire _35481_;
  wire _35482_;
  wire _35483_;
  wire _35484_;
  wire _35485_;
  wire _35486_;
  wire _35487_;
  wire _35488_;
  wire _35489_;
  wire _35490_;
  wire _35491_;
  wire _35492_;
  wire _35493_;
  wire _35494_;
  wire _35495_;
  wire _35496_;
  wire _35497_;
  wire _35498_;
  wire _35499_;
  wire _35500_;
  wire _35501_;
  wire _35502_;
  wire _35503_;
  wire _35504_;
  wire _35505_;
  wire _35506_;
  wire _35507_;
  wire _35508_;
  wire _35509_;
  wire _35510_;
  wire _35511_;
  wire _35512_;
  wire _35513_;
  wire _35514_;
  wire _35515_;
  wire _35516_;
  wire _35517_;
  wire _35518_;
  wire _35519_;
  wire _35520_;
  wire _35521_;
  wire _35522_;
  wire _35523_;
  wire _35524_;
  wire _35525_;
  wire _35526_;
  wire _35527_;
  wire _35528_;
  wire _35529_;
  wire _35530_;
  wire _35531_;
  wire _35532_;
  wire _35533_;
  wire _35534_;
  wire _35535_;
  wire _35536_;
  wire _35537_;
  wire _35538_;
  wire _35539_;
  wire _35540_;
  wire _35541_;
  wire _35542_;
  wire _35543_;
  wire _35544_;
  wire _35545_;
  wire _35546_;
  wire _35547_;
  wire _35548_;
  wire _35549_;
  wire _35550_;
  wire _35551_;
  wire _35552_;
  wire _35553_;
  wire _35554_;
  wire _35555_;
  wire _35556_;
  wire _35557_;
  wire _35558_;
  wire _35559_;
  wire _35560_;
  wire _35561_;
  wire _35562_;
  wire _35563_;
  wire _35564_;
  wire _35565_;
  wire _35566_;
  wire _35567_;
  wire _35568_;
  wire _35569_;
  wire _35570_;
  wire _35571_;
  wire _35572_;
  wire _35573_;
  wire _35574_;
  wire _35575_;
  wire _35576_;
  wire _35577_;
  wire _35578_;
  wire _35579_;
  wire _35580_;
  wire _35581_;
  wire _35582_;
  wire _35583_;
  wire _35584_;
  wire _35585_;
  wire _35586_;
  wire _35587_;
  wire _35588_;
  wire _35589_;
  wire _35590_;
  wire _35591_;
  wire _35592_;
  wire _35593_;
  wire _35594_;
  wire _35595_;
  wire _35596_;
  wire _35597_;
  wire _35598_;
  wire _35599_;
  wire _35600_;
  wire _35601_;
  wire _35602_;
  wire _35603_;
  wire _35604_;
  wire _35605_;
  wire _35606_;
  wire _35607_;
  wire _35608_;
  wire _35609_;
  wire _35610_;
  wire _35611_;
  wire _35612_;
  wire _35613_;
  wire _35614_;
  wire _35615_;
  wire _35616_;
  wire _35617_;
  wire _35618_;
  wire _35619_;
  wire _35620_;
  wire _35621_;
  wire _35622_;
  wire _35623_;
  wire _35624_;
  wire _35625_;
  wire _35626_;
  wire _35627_;
  wire _35628_;
  wire _35629_;
  wire _35630_;
  wire _35631_;
  wire _35632_;
  wire _35633_;
  wire _35634_;
  wire _35635_;
  wire _35636_;
  wire _35637_;
  wire _35638_;
  wire _35639_;
  wire _35640_;
  wire _35641_;
  wire _35642_;
  wire _35643_;
  wire _35644_;
  wire _35645_;
  wire _35646_;
  wire _35647_;
  wire _35648_;
  wire _35649_;
  wire _35650_;
  wire _35651_;
  wire _35652_;
  wire _35653_;
  wire _35654_;
  wire _35655_;
  wire _35656_;
  wire _35657_;
  wire _35658_;
  wire _35659_;
  wire _35660_;
  wire _35661_;
  wire _35662_;
  wire _35663_;
  wire _35664_;
  wire _35665_;
  wire _35666_;
  wire _35667_;
  wire _35668_;
  wire _35669_;
  wire _35670_;
  wire _35671_;
  wire _35672_;
  wire _35673_;
  wire _35674_;
  wire _35675_;
  wire _35676_;
  wire _35677_;
  wire _35678_;
  wire _35679_;
  wire _35680_;
  wire _35681_;
  wire _35682_;
  wire _35683_;
  wire _35684_;
  wire _35685_;
  wire _35686_;
  wire _35687_;
  wire _35688_;
  wire _35689_;
  wire _35690_;
  wire _35691_;
  wire _35692_;
  wire _35693_;
  wire _35694_;
  wire _35695_;
  wire _35696_;
  wire _35697_;
  wire _35698_;
  wire _35699_;
  wire _35700_;
  wire _35701_;
  wire _35702_;
  wire _35703_;
  wire _35704_;
  wire _35705_;
  wire _35706_;
  wire _35707_;
  wire _35708_;
  wire _35709_;
  wire _35710_;
  wire _35711_;
  wire _35712_;
  wire _35713_;
  wire _35714_;
  wire _35715_;
  wire _35716_;
  wire _35717_;
  wire _35718_;
  wire _35719_;
  wire _35720_;
  wire _35721_;
  wire _35722_;
  wire _35723_;
  wire _35724_;
  wire _35725_;
  wire _35726_;
  wire _35727_;
  wire _35728_;
  wire _35729_;
  wire _35730_;
  wire _35731_;
  wire _35732_;
  wire _35733_;
  wire _35734_;
  wire _35735_;
  wire _35736_;
  wire _35737_;
  wire _35738_;
  wire _35739_;
  wire _35740_;
  wire _35741_;
  wire _35742_;
  wire _35743_;
  wire _35744_;
  wire _35745_;
  wire _35746_;
  wire _35747_;
  wire _35748_;
  wire _35749_;
  wire _35750_;
  wire _35751_;
  wire _35752_;
  wire _35753_;
  wire _35754_;
  wire _35755_;
  wire _35756_;
  wire _35757_;
  wire _35758_;
  wire _35759_;
  wire _35760_;
  wire _35761_;
  wire _35762_;
  wire _35763_;
  wire _35764_;
  wire _35765_;
  wire _35766_;
  wire _35767_;
  wire _35768_;
  wire _35769_;
  wire _35770_;
  wire _35771_;
  wire _35772_;
  wire _35773_;
  wire _35774_;
  wire _35775_;
  wire _35776_;
  wire _35777_;
  wire _35778_;
  wire _35779_;
  wire _35780_;
  wire _35781_;
  wire _35782_;
  wire _35783_;
  wire _35784_;
  wire _35785_;
  wire _35786_;
  wire _35787_;
  wire _35788_;
  wire _35789_;
  wire _35790_;
  wire _35791_;
  wire _35792_;
  wire _35793_;
  wire _35794_;
  wire _35795_;
  wire _35796_;
  wire _35797_;
  wire _35798_;
  wire _35799_;
  wire _35800_;
  wire _35801_;
  wire _35802_;
  wire _35803_;
  wire _35804_;
  wire _35805_;
  wire _35806_;
  wire _35807_;
  wire _35808_;
  wire _35809_;
  wire _35810_;
  wire _35811_;
  wire _35812_;
  wire _35813_;
  wire _35814_;
  wire _35815_;
  wire _35816_;
  wire _35817_;
  wire _35818_;
  wire _35819_;
  wire _35820_;
  wire _35821_;
  wire _35822_;
  wire _35823_;
  wire _35824_;
  wire _35825_;
  wire _35826_;
  wire _35827_;
  wire _35828_;
  wire _35829_;
  wire _35830_;
  wire _35831_;
  wire _35832_;
  wire _35833_;
  wire _35834_;
  wire _35835_;
  wire _35836_;
  wire _35837_;
  wire _35838_;
  wire _35839_;
  wire _35840_;
  wire _35841_;
  wire _35842_;
  wire _35843_;
  wire _35844_;
  wire _35845_;
  wire _35846_;
  wire _35847_;
  wire _35848_;
  wire _35849_;
  wire _35850_;
  wire _35851_;
  wire _35852_;
  wire _35853_;
  wire _35854_;
  wire _35855_;
  wire _35856_;
  wire _35857_;
  wire _35858_;
  wire _35859_;
  wire _35860_;
  wire _35861_;
  wire _35862_;
  wire _35863_;
  wire _35864_;
  wire _35865_;
  wire _35866_;
  wire _35867_;
  wire _35868_;
  wire _35869_;
  wire _35870_;
  wire _35871_;
  wire _35872_;
  wire _35873_;
  wire _35874_;
  wire _35875_;
  wire _35876_;
  wire _35877_;
  wire _35878_;
  wire _35879_;
  wire _35880_;
  wire _35881_;
  wire _35882_;
  wire _35883_;
  wire _35884_;
  wire _35885_;
  wire _35886_;
  wire _35887_;
  wire _35888_;
  wire _35889_;
  wire _35890_;
  wire _35891_;
  wire _35892_;
  wire _35893_;
  wire _35894_;
  wire _35895_;
  wire _35896_;
  wire _35897_;
  wire _35898_;
  wire _35899_;
  wire _35900_;
  wire _35901_;
  wire _35902_;
  wire _35903_;
  wire _35904_;
  wire _35905_;
  wire _35906_;
  wire _35907_;
  wire _35908_;
  wire _35909_;
  wire _35910_;
  wire _35911_;
  wire _35912_;
  wire _35913_;
  wire _35914_;
  wire _35915_;
  wire _35916_;
  wire _35917_;
  wire _35918_;
  wire _35919_;
  wire _35920_;
  wire _35921_;
  wire _35922_;
  wire _35923_;
  wire _35924_;
  wire _35925_;
  wire _35926_;
  wire _35927_;
  wire _35928_;
  wire _35929_;
  wire _35930_;
  wire _35931_;
  wire _35932_;
  wire _35933_;
  wire _35934_;
  wire _35935_;
  wire _35936_;
  wire _35937_;
  wire _35938_;
  wire _35939_;
  wire _35940_;
  wire _35941_;
  wire _35942_;
  wire _35943_;
  wire _35944_;
  wire _35945_;
  wire _35946_;
  wire _35947_;
  wire _35948_;
  wire _35949_;
  wire _35950_;
  wire _35951_;
  wire _35952_;
  wire _35953_;
  wire _35954_;
  wire _35955_;
  wire _35956_;
  wire _35957_;
  wire _35958_;
  wire _35959_;
  wire _35960_;
  wire _35961_;
  wire _35962_;
  wire _35963_;
  wire _35964_;
  wire _35965_;
  wire _35966_;
  wire _35967_;
  wire _35968_;
  wire _35969_;
  wire _35970_;
  wire _35971_;
  wire _35972_;
  wire _35973_;
  wire _35974_;
  wire _35975_;
  wire _35976_;
  wire _35977_;
  wire _35978_;
  wire _35979_;
  wire _35980_;
  wire _35981_;
  wire _35982_;
  wire _35983_;
  wire _35984_;
  wire _35985_;
  wire _35986_;
  wire _35987_;
  wire _35988_;
  wire _35989_;
  wire _35990_;
  wire _35991_;
  wire _35992_;
  wire _35993_;
  wire _35994_;
  wire _35995_;
  wire _35996_;
  wire _35997_;
  wire _35998_;
  wire _35999_;
  wire _36000_;
  wire _36001_;
  wire _36002_;
  wire _36003_;
  wire _36004_;
  wire _36005_;
  wire _36006_;
  wire _36007_;
  wire _36008_;
  wire _36009_;
  wire _36010_;
  wire _36011_;
  wire _36012_;
  wire _36013_;
  wire _36014_;
  wire _36015_;
  wire _36016_;
  wire _36017_;
  wire _36018_;
  wire _36019_;
  wire _36020_;
  wire _36021_;
  wire _36022_;
  wire _36023_;
  wire _36024_;
  wire _36025_;
  wire _36026_;
  wire _36027_;
  wire _36028_;
  wire _36029_;
  wire _36030_;
  wire _36031_;
  wire _36032_;
  wire _36033_;
  wire _36034_;
  wire _36035_;
  wire _36036_;
  wire _36037_;
  wire _36038_;
  wire _36039_;
  wire _36040_;
  wire _36041_;
  wire _36042_;
  wire _36043_;
  wire _36044_;
  wire _36045_;
  wire _36046_;
  wire _36047_;
  wire _36048_;
  wire _36049_;
  wire _36050_;
  wire _36051_;
  wire _36052_;
  wire _36053_;
  wire _36054_;
  wire _36055_;
  wire _36056_;
  wire _36057_;
  wire _36058_;
  wire _36059_;
  wire _36060_;
  wire _36061_;
  wire _36062_;
  wire _36063_;
  wire _36064_;
  wire _36065_;
  wire _36066_;
  wire _36067_;
  wire _36068_;
  wire _36069_;
  wire _36070_;
  wire _36071_;
  wire _36072_;
  wire _36073_;
  wire _36074_;
  wire _36075_;
  wire _36076_;
  wire _36077_;
  wire _36078_;
  wire _36079_;
  wire _36080_;
  wire _36081_;
  wire _36082_;
  wire _36083_;
  wire _36084_;
  wire _36085_;
  wire _36086_;
  wire _36087_;
  wire _36088_;
  wire _36089_;
  wire _36090_;
  wire _36091_;
  wire _36092_;
  wire _36093_;
  wire _36094_;
  wire _36095_;
  wire _36096_;
  wire _36097_;
  wire _36098_;
  wire _36099_;
  wire _36100_;
  wire _36101_;
  wire _36102_;
  wire _36103_;
  wire _36104_;
  wire _36105_;
  wire _36106_;
  wire _36107_;
  wire _36108_;
  wire _36109_;
  wire _36110_;
  wire _36111_;
  wire _36112_;
  wire _36113_;
  wire _36114_;
  wire _36115_;
  wire _36116_;
  wire _36117_;
  wire _36118_;
  wire _36119_;
  wire _36120_;
  wire _36121_;
  wire _36122_;
  wire _36123_;
  wire _36124_;
  wire _36125_;
  wire _36126_;
  wire _36127_;
  wire _36128_;
  wire _36129_;
  wire _36130_;
  wire _36131_;
  wire _36132_;
  wire _36133_;
  wire _36134_;
  wire _36135_;
  wire _36136_;
  wire _36137_;
  wire _36138_;
  wire _36139_;
  wire _36140_;
  wire _36141_;
  wire _36142_;
  wire _36143_;
  wire _36144_;
  wire _36145_;
  wire _36146_;
  wire _36147_;
  wire _36148_;
  wire _36149_;
  wire _36150_;
  wire _36151_;
  wire _36152_;
  wire _36153_;
  wire _36154_;
  wire _36155_;
  wire _36156_;
  wire _36157_;
  wire _36158_;
  wire _36159_;
  wire _36160_;
  wire _36161_;
  wire _36162_;
  wire _36163_;
  wire _36164_;
  wire _36165_;
  wire _36166_;
  wire _36167_;
  wire _36168_;
  wire _36169_;
  wire _36170_;
  wire _36171_;
  wire _36172_;
  wire _36173_;
  wire _36174_;
  wire _36175_;
  wire _36176_;
  wire _36177_;
  wire _36178_;
  wire _36179_;
  wire _36180_;
  wire _36181_;
  wire _36182_;
  wire _36183_;
  wire _36184_;
  wire _36185_;
  wire _36186_;
  wire _36187_;
  wire _36188_;
  wire _36189_;
  wire _36190_;
  wire _36191_;
  wire _36192_;
  wire _36193_;
  wire _36194_;
  wire _36195_;
  wire _36196_;
  wire _36197_;
  wire _36198_;
  wire _36199_;
  wire _36200_;
  wire _36201_;
  wire _36202_;
  wire _36203_;
  wire _36204_;
  wire _36205_;
  wire _36206_;
  wire _36207_;
  wire _36208_;
  wire _36209_;
  wire _36210_;
  wire _36211_;
  wire _36212_;
  wire _36213_;
  wire _36214_;
  wire _36215_;
  wire _36216_;
  wire _36217_;
  wire _36218_;
  wire _36219_;
  wire _36220_;
  wire _36221_;
  wire _36222_;
  wire _36223_;
  wire _36224_;
  wire _36225_;
  wire _36226_;
  wire _36227_;
  wire _36228_;
  wire _36229_;
  wire _36230_;
  wire _36231_;
  wire _36232_;
  wire _36233_;
  wire _36234_;
  wire _36235_;
  wire _36236_;
  wire _36237_;
  wire _36238_;
  wire _36239_;
  wire _36240_;
  wire _36241_;
  wire _36242_;
  wire _36243_;
  wire _36244_;
  wire _36245_;
  wire _36246_;
  wire _36247_;
  wire _36248_;
  wire _36249_;
  wire _36250_;
  wire _36251_;
  wire _36252_;
  wire _36253_;
  wire _36254_;
  wire _36255_;
  wire _36256_;
  wire _36257_;
  wire _36258_;
  wire _36259_;
  wire _36260_;
  wire _36261_;
  wire _36262_;
  wire _36263_;
  wire _36264_;
  wire _36265_;
  wire _36266_;
  wire _36267_;
  wire _36268_;
  wire _36269_;
  wire _36270_;
  wire _36271_;
  wire _36272_;
  wire _36273_;
  wire _36274_;
  wire _36275_;
  wire _36276_;
  wire _36277_;
  wire _36278_;
  wire _36279_;
  wire _36280_;
  wire _36281_;
  wire _36282_;
  wire _36283_;
  wire _36284_;
  wire _36285_;
  wire _36286_;
  wire _36287_;
  wire _36288_;
  wire _36289_;
  wire _36290_;
  wire _36291_;
  wire _36292_;
  wire _36293_;
  wire _36294_;
  wire _36295_;
  wire _36296_;
  wire _36297_;
  wire _36298_;
  wire _36299_;
  wire _36300_;
  wire _36301_;
  wire _36302_;
  wire _36303_;
  wire _36304_;
  wire _36305_;
  wire _36306_;
  wire _36307_;
  wire _36308_;
  wire _36309_;
  wire _36310_;
  wire _36311_;
  wire _36312_;
  wire _36313_;
  wire _36314_;
  wire _36315_;
  wire _36316_;
  wire _36317_;
  wire _36318_;
  wire _36319_;
  wire _36320_;
  wire _36321_;
  wire _36322_;
  wire _36323_;
  wire _36324_;
  wire _36325_;
  wire _36326_;
  wire _36327_;
  wire _36328_;
  wire _36329_;
  wire _36330_;
  wire _36331_;
  wire _36332_;
  wire _36333_;
  wire _36334_;
  wire _36335_;
  wire _36336_;
  wire _36337_;
  wire _36338_;
  wire _36339_;
  wire _36340_;
  wire _36341_;
  wire _36342_;
  wire _36343_;
  wire _36344_;
  wire _36345_;
  wire _36346_;
  wire _36347_;
  wire _36348_;
  wire _36349_;
  wire _36350_;
  wire _36351_;
  wire _36352_;
  wire _36353_;
  wire _36354_;
  wire _36355_;
  wire _36356_;
  wire _36357_;
  wire _36358_;
  wire _36359_;
  wire _36360_;
  wire _36361_;
  wire _36362_;
  wire _36363_;
  wire _36364_;
  wire _36365_;
  wire _36366_;
  wire _36367_;
  wire _36368_;
  wire _36369_;
  wire _36370_;
  wire _36371_;
  wire _36372_;
  wire _36373_;
  wire _36374_;
  wire _36375_;
  wire _36376_;
  wire _36377_;
  wire _36378_;
  wire _36379_;
  wire _36380_;
  wire _36381_;
  wire _36382_;
  wire _36383_;
  wire _36384_;
  wire _36385_;
  wire _36386_;
  wire _36387_;
  wire _36388_;
  wire _36389_;
  wire _36390_;
  wire _36391_;
  wire _36392_;
  wire _36393_;
  wire _36394_;
  wire _36395_;
  wire _36396_;
  wire _36397_;
  wire _36398_;
  wire _36399_;
  wire _36400_;
  wire _36401_;
  wire _36402_;
  wire _36403_;
  wire _36404_;
  wire _36405_;
  wire _36406_;
  wire _36407_;
  wire _36408_;
  wire _36409_;
  wire _36410_;
  wire _36411_;
  wire _36412_;
  wire _36413_;
  wire _36414_;
  wire _36415_;
  wire _36416_;
  wire _36417_;
  wire _36418_;
  wire _36419_;
  wire _36420_;
  wire _36421_;
  wire _36422_;
  wire _36423_;
  wire _36424_;
  wire _36425_;
  wire _36426_;
  wire _36427_;
  wire _36428_;
  wire _36429_;
  wire _36430_;
  wire _36431_;
  wire _36432_;
  wire _36433_;
  wire _36434_;
  wire _36435_;
  wire _36436_;
  wire _36437_;
  wire _36438_;
  wire _36439_;
  wire _36440_;
  wire _36441_;
  wire _36442_;
  wire _36443_;
  wire _36444_;
  wire _36445_;
  wire _36446_;
  wire _36447_;
  wire _36448_;
  wire _36449_;
  wire _36450_;
  wire _36451_;
  wire _36452_;
  wire _36453_;
  wire _36454_;
  wire _36455_;
  wire _36456_;
  wire _36457_;
  wire _36458_;
  wire _36459_;
  wire _36460_;
  wire _36461_;
  wire _36462_;
  wire _36463_;
  wire _36464_;
  wire _36465_;
  wire _36466_;
  wire _36467_;
  wire _36468_;
  wire _36469_;
  wire _36470_;
  wire _36471_;
  wire _36472_;
  wire _36473_;
  wire _36474_;
  wire _36475_;
  wire _36476_;
  wire _36477_;
  wire _36478_;
  wire _36479_;
  wire _36480_;
  wire _36481_;
  wire _36482_;
  wire _36483_;
  wire _36484_;
  wire _36485_;
  wire _36486_;
  wire _36487_;
  wire _36488_;
  wire _36489_;
  wire _36490_;
  wire _36491_;
  wire _36492_;
  wire _36493_;
  wire _36494_;
  wire _36495_;
  wire _36496_;
  wire _36497_;
  wire _36498_;
  wire _36499_;
  wire _36500_;
  wire _36501_;
  wire _36502_;
  wire _36503_;
  wire _36504_;
  wire _36505_;
  wire _36506_;
  wire _36507_;
  wire _36508_;
  wire _36509_;
  wire _36510_;
  wire _36511_;
  wire _36512_;
  wire _36513_;
  wire _36514_;
  wire _36515_;
  wire _36516_;
  wire _36517_;
  wire _36518_;
  wire _36519_;
  wire _36520_;
  wire _36521_;
  wire _36522_;
  wire _36523_;
  wire _36524_;
  wire _36525_;
  wire _36526_;
  wire _36527_;
  wire _36528_;
  wire _36529_;
  wire _36530_;
  wire _36531_;
  wire _36532_;
  wire _36533_;
  wire _36534_;
  wire _36535_;
  wire _36536_;
  wire _36537_;
  wire _36538_;
  wire _36539_;
  wire _36540_;
  wire _36541_;
  wire _36542_;
  wire _36543_;
  wire _36544_;
  wire _36545_;
  wire _36546_;
  wire _36547_;
  wire _36548_;
  wire _36549_;
  wire _36550_;
  wire _36551_;
  wire _36552_;
  wire _36553_;
  wire _36554_;
  wire _36555_;
  wire _36556_;
  wire _36557_;
  wire _36558_;
  wire _36559_;
  wire _36560_;
  wire _36561_;
  wire _36562_;
  wire _36563_;
  wire _36564_;
  wire _36565_;
  wire _36566_;
  wire _36567_;
  wire _36568_;
  wire _36569_;
  wire _36570_;
  wire _36571_;
  wire _36572_;
  wire _36573_;
  wire _36574_;
  wire _36575_;
  wire _36576_;
  wire _36577_;
  wire _36578_;
  wire _36579_;
  wire _36580_;
  wire _36581_;
  wire _36582_;
  wire _36583_;
  wire _36584_;
  wire _36585_;
  wire _36586_;
  wire _36587_;
  wire _36588_;
  wire _36589_;
  wire _36590_;
  wire _36591_;
  wire _36592_;
  wire _36593_;
  wire _36594_;
  wire _36595_;
  wire _36596_;
  wire _36597_;
  wire _36598_;
  wire _36599_;
  wire _36600_;
  wire _36601_;
  wire _36602_;
  wire _36603_;
  wire _36604_;
  wire _36605_;
  wire _36606_;
  wire _36607_;
  wire _36608_;
  wire _36609_;
  wire _36610_;
  wire _36611_;
  wire _36612_;
  wire _36613_;
  wire _36614_;
  wire _36615_;
  wire _36616_;
  wire _36617_;
  wire _36618_;
  wire _36619_;
  wire _36620_;
  wire _36621_;
  wire _36622_;
  wire _36623_;
  wire _36624_;
  wire _36625_;
  wire _36626_;
  wire _36627_;
  wire _36628_;
  wire _36629_;
  wire _36630_;
  wire _36631_;
  wire _36632_;
  wire _36633_;
  wire _36634_;
  wire _36635_;
  wire _36636_;
  wire _36637_;
  wire _36638_;
  wire _36639_;
  wire _36640_;
  wire _36641_;
  wire _36642_;
  wire _36643_;
  wire _36644_;
  wire _36645_;
  wire _36646_;
  wire _36647_;
  wire _36648_;
  wire _36649_;
  wire _36650_;
  wire _36651_;
  wire _36652_;
  wire _36653_;
  wire _36654_;
  wire _36655_;
  wire _36656_;
  wire _36657_;
  wire _36658_;
  wire _36659_;
  wire _36660_;
  wire _36661_;
  wire _36662_;
  wire _36663_;
  wire _36664_;
  wire _36665_;
  wire _36666_;
  wire _36667_;
  wire _36668_;
  wire _36669_;
  wire _36670_;
  wire _36671_;
  wire _36672_;
  wire _36673_;
  wire _36674_;
  wire _36675_;
  wire _36676_;
  wire _36677_;
  wire _36678_;
  wire _36679_;
  wire _36680_;
  wire _36681_;
  wire _36682_;
  wire _36683_;
  wire _36684_;
  wire _36685_;
  wire _36686_;
  wire _36687_;
  wire _36688_;
  wire _36689_;
  wire _36690_;
  wire _36691_;
  wire _36692_;
  wire _36693_;
  wire _36694_;
  wire _36695_;
  wire _36696_;
  wire _36697_;
  wire _36698_;
  wire _36699_;
  wire _36700_;
  wire _36701_;
  wire _36702_;
  wire _36703_;
  wire _36704_;
  wire _36705_;
  wire _36706_;
  wire _36707_;
  wire _36708_;
  wire _36709_;
  wire _36710_;
  wire _36711_;
  wire _36712_;
  wire _36713_;
  wire _36714_;
  wire _36715_;
  wire _36716_;
  wire _36717_;
  wire _36718_;
  wire _36719_;
  wire _36720_;
  wire _36721_;
  wire _36722_;
  wire _36723_;
  wire _36724_;
  wire _36725_;
  wire _36726_;
  wire _36727_;
  wire _36728_;
  wire _36729_;
  wire _36730_;
  wire _36731_;
  wire _36732_;
  wire _36733_;
  wire _36734_;
  wire _36735_;
  wire _36736_;
  wire _36737_;
  wire _36738_;
  wire _36739_;
  wire _36740_;
  wire _36741_;
  wire _36742_;
  wire _36743_;
  wire _36744_;
  wire _36745_;
  wire _36746_;
  wire _36747_;
  wire _36748_;
  wire _36749_;
  wire _36750_;
  wire _36751_;
  wire _36752_;
  wire _36753_;
  wire _36754_;
  wire _36755_;
  wire _36756_;
  wire _36757_;
  wire _36758_;
  wire _36759_;
  wire _36760_;
  wire _36761_;
  wire _36762_;
  wire _36763_;
  wire _36764_;
  wire _36765_;
  wire _36766_;
  wire _36767_;
  wire _36768_;
  wire _36769_;
  wire _36770_;
  wire _36771_;
  wire _36772_;
  wire _36773_;
  wire _36774_;
  wire _36775_;
  wire _36776_;
  wire _36777_;
  wire _36778_;
  wire _36779_;
  wire _36780_;
  wire _36781_;
  wire _36782_;
  wire _36783_;
  wire _36784_;
  wire _36785_;
  wire _36786_;
  wire _36787_;
  wire _36788_;
  wire _36789_;
  wire _36790_;
  wire _36791_;
  wire _36792_;
  wire _36793_;
  wire _36794_;
  wire _36795_;
  wire _36796_;
  wire _36797_;
  wire _36798_;
  wire _36799_;
  wire _36800_;
  wire _36801_;
  wire _36802_;
  wire _36803_;
  wire _36804_;
  wire _36805_;
  wire _36806_;
  wire _36807_;
  wire _36808_;
  wire _36809_;
  wire _36810_;
  wire _36811_;
  wire _36812_;
  wire _36813_;
  wire _36814_;
  wire _36815_;
  wire _36816_;
  wire _36817_;
  wire _36818_;
  wire _36819_;
  wire _36820_;
  wire _36821_;
  wire _36822_;
  wire _36823_;
  wire _36824_;
  wire _36825_;
  wire _36826_;
  wire _36827_;
  wire _36828_;
  wire _36829_;
  wire _36830_;
  wire _36831_;
  wire _36832_;
  wire _36833_;
  wire _36834_;
  wire _36835_;
  wire _36836_;
  wire _36837_;
  wire _36838_;
  wire _36839_;
  wire _36840_;
  wire _36841_;
  wire _36842_;
  wire _36843_;
  wire _36844_;
  wire _36845_;
  wire _36846_;
  wire _36847_;
  wire _36848_;
  wire _36849_;
  wire _36850_;
  wire _36851_;
  wire _36852_;
  wire _36853_;
  wire _36854_;
  wire _36855_;
  wire _36856_;
  wire _36857_;
  wire _36858_;
  wire _36859_;
  wire _36860_;
  wire _36861_;
  wire _36862_;
  wire _36863_;
  wire _36864_;
  wire _36865_;
  wire _36866_;
  wire _36867_;
  wire _36868_;
  wire _36869_;
  wire _36870_;
  wire _36871_;
  wire _36872_;
  wire _36873_;
  wire _36874_;
  wire _36875_;
  wire _36876_;
  wire _36877_;
  wire _36878_;
  wire _36879_;
  wire _36880_;
  wire _36881_;
  wire _36882_;
  wire _36883_;
  wire _36884_;
  wire _36885_;
  wire _36886_;
  wire _36887_;
  wire _36888_;
  wire _36889_;
  wire _36890_;
  wire _36891_;
  wire _36892_;
  wire _36893_;
  wire _36894_;
  wire _36895_;
  wire _36896_;
  wire _36897_;
  wire _36898_;
  wire _36899_;
  wire _36900_;
  wire _36901_;
  wire _36902_;
  wire _36903_;
  wire _36904_;
  wire _36905_;
  wire _36906_;
  wire _36907_;
  wire _36908_;
  wire _36909_;
  wire _36910_;
  wire _36911_;
  wire _36912_;
  wire _36913_;
  wire _36914_;
  wire _36915_;
  wire _36916_;
  wire _36917_;
  wire _36918_;
  wire _36919_;
  wire _36920_;
  wire _36921_;
  wire _36922_;
  wire _36923_;
  wire _36924_;
  wire _36925_;
  wire _36926_;
  wire _36927_;
  wire _36928_;
  wire _36929_;
  wire _36930_;
  wire _36931_;
  wire _36932_;
  wire _36933_;
  wire _36934_;
  wire _36935_;
  wire _36936_;
  wire _36937_;
  wire _36938_;
  wire _36939_;
  wire _36940_;
  wire _36941_;
  wire _36942_;
  wire _36943_;
  wire _36944_;
  wire _36945_;
  wire _36946_;
  wire _36947_;
  wire _36948_;
  wire _36949_;
  wire _36950_;
  wire _36951_;
  wire _36952_;
  wire _36953_;
  wire _36954_;
  wire _36955_;
  wire _36956_;
  wire _36957_;
  wire _36958_;
  wire _36959_;
  wire _36960_;
  wire _36961_;
  wire _36962_;
  wire _36963_;
  wire _36964_;
  wire _36965_;
  wire _36966_;
  wire _36967_;
  wire _36968_;
  wire _36969_;
  wire _36970_;
  wire _36971_;
  wire _36972_;
  wire _36973_;
  wire _36974_;
  wire _36975_;
  wire _36976_;
  wire _36977_;
  wire _36978_;
  wire _36979_;
  wire _36980_;
  wire _36981_;
  wire _36982_;
  wire _36983_;
  wire _36984_;
  wire _36985_;
  wire _36986_;
  wire _36987_;
  wire _36988_;
  wire _36989_;
  wire _36990_;
  wire _36991_;
  wire _36992_;
  wire _36993_;
  wire _36994_;
  wire _36995_;
  wire _36996_;
  wire _36997_;
  wire _36998_;
  wire _36999_;
  wire _37000_;
  wire _37001_;
  wire _37002_;
  wire _37003_;
  wire _37004_;
  wire _37005_;
  wire _37006_;
  wire _37007_;
  wire _37008_;
  wire _37009_;
  wire _37010_;
  wire _37011_;
  wire _37012_;
  wire _37013_;
  wire _37014_;
  wire _37015_;
  wire _37016_;
  wire _37017_;
  wire _37018_;
  wire _37019_;
  wire _37020_;
  wire _37021_;
  wire _37022_;
  wire _37023_;
  wire _37024_;
  wire _37025_;
  wire _37026_;
  wire _37027_;
  wire _37028_;
  wire _37029_;
  wire _37030_;
  wire _37031_;
  wire _37032_;
  wire _37033_;
  wire _37034_;
  wire _37035_;
  wire _37036_;
  wire _37037_;
  wire _37038_;
  wire _37039_;
  wire _37040_;
  wire _37041_;
  wire _37042_;
  wire _37043_;
  wire _37044_;
  wire _37045_;
  wire _37046_;
  wire _37047_;
  wire _37048_;
  wire _37049_;
  wire _37050_;
  wire _37051_;
  wire _37052_;
  wire _37053_;
  wire _37054_;
  wire _37055_;
  wire _37056_;
  wire _37057_;
  wire _37058_;
  wire _37059_;
  wire _37060_;
  wire _37061_;
  wire _37062_;
  wire _37063_;
  wire _37064_;
  wire _37065_;
  wire _37066_;
  wire _37067_;
  wire _37068_;
  wire _37069_;
  wire _37070_;
  wire _37071_;
  wire _37072_;
  wire _37073_;
  wire _37074_;
  wire _37075_;
  wire _37076_;
  wire _37077_;
  wire _37078_;
  wire _37079_;
  wire _37080_;
  wire _37081_;
  wire _37082_;
  wire _37083_;
  wire _37084_;
  wire _37085_;
  wire _37086_;
  wire _37087_;
  wire _37088_;
  wire _37089_;
  wire _37090_;
  wire _37091_;
  wire _37092_;
  wire _37093_;
  wire _37094_;
  wire _37095_;
  wire _37096_;
  wire _37097_;
  wire _37098_;
  wire _37099_;
  wire _37100_;
  wire _37101_;
  wire _37102_;
  wire _37103_;
  wire _37104_;
  wire _37105_;
  wire _37106_;
  wire _37107_;
  wire _37108_;
  wire _37109_;
  wire _37110_;
  wire _37111_;
  wire _37112_;
  wire _37113_;
  wire _37114_;
  wire _37115_;
  wire _37116_;
  wire _37117_;
  wire _37118_;
  wire _37119_;
  wire _37120_;
  wire _37121_;
  wire _37122_;
  wire _37123_;
  wire _37124_;
  wire _37125_;
  wire _37126_;
  wire _37127_;
  wire _37128_;
  wire _37129_;
  wire _37130_;
  wire _37131_;
  wire _37132_;
  wire _37133_;
  wire _37134_;
  wire _37135_;
  wire _37136_;
  wire _37137_;
  wire _37138_;
  wire _37139_;
  wire _37140_;
  wire _37141_;
  wire _37142_;
  wire _37143_;
  wire _37144_;
  wire _37145_;
  wire _37146_;
  wire _37147_;
  wire _37148_;
  wire _37149_;
  wire _37150_;
  wire _37151_;
  wire _37152_;
  wire _37153_;
  wire _37154_;
  wire _37155_;
  wire _37156_;
  wire _37157_;
  wire _37158_;
  wire _37159_;
  wire _37160_;
  wire _37161_;
  wire _37162_;
  wire _37163_;
  wire _37164_;
  wire _37165_;
  wire _37166_;
  wire _37167_;
  wire _37168_;
  wire _37169_;
  wire _37170_;
  wire _37171_;
  wire _37172_;
  wire _37173_;
  wire _37174_;
  wire _37175_;
  wire _37176_;
  wire _37177_;
  wire _37178_;
  wire _37179_;
  wire _37180_;
  wire _37181_;
  wire _37182_;
  wire _37183_;
  wire _37184_;
  wire _37185_;
  wire _37186_;
  wire _37187_;
  wire _37188_;
  wire _37189_;
  wire _37190_;
  wire _37191_;
  wire _37192_;
  wire _37193_;
  wire _37194_;
  wire _37195_;
  wire _37196_;
  wire _37197_;
  wire _37198_;
  wire _37199_;
  wire _37200_;
  wire _37201_;
  wire _37202_;
  wire _37203_;
  wire _37204_;
  wire _37205_;
  wire _37206_;
  wire _37207_;
  wire _37208_;
  wire _37209_;
  wire _37210_;
  wire _37211_;
  wire _37212_;
  wire _37213_;
  wire _37214_;
  wire _37215_;
  wire _37216_;
  wire _37217_;
  wire _37218_;
  wire _37219_;
  wire _37220_;
  wire _37221_;
  wire _37222_;
  wire _37223_;
  wire _37224_;
  wire _37225_;
  wire _37226_;
  wire _37227_;
  wire _37228_;
  wire _37229_;
  wire _37230_;
  wire _37231_;
  wire _37232_;
  wire _37233_;
  wire _37234_;
  wire _37235_;
  wire _37236_;
  wire _37237_;
  wire _37238_;
  wire _37239_;
  wire _37240_;
  wire _37241_;
  wire _37242_;
  wire _37243_;
  wire _37244_;
  wire _37245_;
  wire _37246_;
  wire _37247_;
  wire _37248_;
  wire _37249_;
  wire _37250_;
  wire _37251_;
  wire _37252_;
  wire _37253_;
  wire _37254_;
  wire _37255_;
  wire _37256_;
  wire _37257_;
  wire _37258_;
  wire _37259_;
  wire _37260_;
  wire _37261_;
  wire _37262_;
  wire _37263_;
  wire _37264_;
  wire _37265_;
  wire _37266_;
  wire _37267_;
  wire _37268_;
  wire _37269_;
  wire _37270_;
  wire _37271_;
  wire _37272_;
  wire _37273_;
  wire _37274_;
  wire _37275_;
  wire _37276_;
  wire _37277_;
  wire _37278_;
  wire _37279_;
  wire _37280_;
  wire _37281_;
  wire _37282_;
  wire _37283_;
  wire _37284_;
  wire _37285_;
  wire _37286_;
  wire _37287_;
  wire _37288_;
  wire _37289_;
  wire _37290_;
  wire _37291_;
  wire _37292_;
  wire _37293_;
  wire _37294_;
  wire _37295_;
  wire _37296_;
  wire _37297_;
  wire _37298_;
  wire _37299_;
  wire _37300_;
  wire _37301_;
  wire _37302_;
  wire _37303_;
  wire _37304_;
  wire _37305_;
  wire _37306_;
  wire _37307_;
  wire _37308_;
  wire _37309_;
  wire _37310_;
  wire _37311_;
  wire _37312_;
  wire _37313_;
  wire _37314_;
  wire _37315_;
  wire _37316_;
  wire _37317_;
  wire _37318_;
  wire _37319_;
  wire _37320_;
  wire _37321_;
  wire _37322_;
  wire _37323_;
  wire _37324_;
  wire _37325_;
  wire _37326_;
  wire _37327_;
  wire _37328_;
  wire _37329_;
  wire _37330_;
  wire _37331_;
  wire _37332_;
  wire _37333_;
  wire _37334_;
  wire _37335_;
  wire _37336_;
  wire _37337_;
  wire _37338_;
  wire _37339_;
  wire _37340_;
  wire _37341_;
  wire _37342_;
  wire _37343_;
  wire _37344_;
  wire _37345_;
  wire _37346_;
  wire _37347_;
  wire _37348_;
  wire _37349_;
  wire _37350_;
  wire _37351_;
  wire _37352_;
  wire _37353_;
  wire _37354_;
  wire _37355_;
  wire _37356_;
  wire _37357_;
  wire _37358_;
  wire _37359_;
  wire _37360_;
  wire _37361_;
  wire _37362_;
  wire _37363_;
  wire _37364_;
  wire _37365_;
  wire _37366_;
  wire _37367_;
  wire _37368_;
  wire _37369_;
  wire _37370_;
  wire _37371_;
  wire _37372_;
  wire _37373_;
  wire _37374_;
  wire _37375_;
  wire _37376_;
  wire _37377_;
  wire _37378_;
  wire _37379_;
  wire _37380_;
  wire _37381_;
  wire _37382_;
  wire _37383_;
  wire _37384_;
  wire _37385_;
  wire _37386_;
  wire _37387_;
  wire _37388_;
  wire _37389_;
  wire _37390_;
  wire _37391_;
  wire _37392_;
  wire _37393_;
  wire _37394_;
  wire _37395_;
  wire _37396_;
  wire _37397_;
  wire _37398_;
  wire _37399_;
  wire _37400_;
  wire _37401_;
  wire _37402_;
  wire _37403_;
  wire _37404_;
  wire _37405_;
  wire _37406_;
  wire _37407_;
  wire _37408_;
  wire _37409_;
  wire _37410_;
  wire _37411_;
  wire _37412_;
  wire _37413_;
  wire _37414_;
  wire _37415_;
  wire _37416_;
  wire _37417_;
  wire _37418_;
  wire _37419_;
  wire _37420_;
  wire _37421_;
  wire _37422_;
  wire _37423_;
  wire _37424_;
  wire _37425_;
  wire _37426_;
  wire _37427_;
  wire _37428_;
  wire _37429_;
  wire _37430_;
  wire _37431_;
  wire _37432_;
  wire _37433_;
  wire _37434_;
  wire _37435_;
  wire _37436_;
  wire _37437_;
  wire _37438_;
  wire _37439_;
  wire _37440_;
  wire _37441_;
  wire _37442_;
  wire _37443_;
  wire _37444_;
  wire _37445_;
  wire _37446_;
  wire _37447_;
  wire _37448_;
  wire _37449_;
  wire _37450_;
  wire _37451_;
  wire _37452_;
  wire _37453_;
  wire _37454_;
  wire _37455_;
  wire _37456_;
  wire _37457_;
  wire _37458_;
  wire _37459_;
  wire _37460_;
  wire _37461_;
  wire _37462_;
  wire _37463_;
  wire _37464_;
  wire _37465_;
  wire _37466_;
  wire _37467_;
  wire _37468_;
  wire _37469_;
  wire _37470_;
  wire _37471_;
  wire _37472_;
  wire _37473_;
  wire _37474_;
  wire _37475_;
  wire _37476_;
  wire _37477_;
  wire _37478_;
  wire _37479_;
  wire _37480_;
  wire _37481_;
  wire _37482_;
  wire _37483_;
  wire _37484_;
  wire _37485_;
  wire _37486_;
  wire _37487_;
  wire _37488_;
  wire _37489_;
  wire _37490_;
  wire _37491_;
  wire _37492_;
  wire _37493_;
  wire _37494_;
  wire _37495_;
  wire _37496_;
  wire _37497_;
  wire _37498_;
  wire _37499_;
  wire _37500_;
  wire _37501_;
  wire _37502_;
  wire _37503_;
  wire _37504_;
  wire _37505_;
  wire _37506_;
  wire _37507_;
  wire _37508_;
  wire _37509_;
  wire _37510_;
  wire _37511_;
  wire _37512_;
  wire _37513_;
  wire _37514_;
  wire _37515_;
  wire _37516_;
  wire _37517_;
  wire _37518_;
  wire _37519_;
  wire _37520_;
  wire _37521_;
  wire _37522_;
  wire _37523_;
  wire _37524_;
  wire _37525_;
  wire _37526_;
  wire _37527_;
  wire _37528_;
  wire _37529_;
  wire _37530_;
  wire _37531_;
  wire _37532_;
  wire _37533_;
  wire _37534_;
  wire _37535_;
  wire _37536_;
  wire _37537_;
  wire _37538_;
  wire _37539_;
  wire _37540_;
  wire _37541_;
  wire _37542_;
  wire _37543_;
  wire _37544_;
  wire _37545_;
  wire _37546_;
  wire _37547_;
  wire _37548_;
  wire _37549_;
  wire _37550_;
  wire _37551_;
  wire _37552_;
  wire _37553_;
  wire _37554_;
  wire _37555_;
  wire _37556_;
  wire _37557_;
  wire _37558_;
  wire _37559_;
  wire _37560_;
  wire _37561_;
  wire _37562_;
  wire _37563_;
  wire _37564_;
  wire _37565_;
  wire _37566_;
  wire _37567_;
  wire _37568_;
  wire _37569_;
  wire _37570_;
  wire _37571_;
  wire _37572_;
  wire _37573_;
  wire _37574_;
  wire _37575_;
  wire _37576_;
  wire _37577_;
  wire _37578_;
  wire _37579_;
  wire _37580_;
  wire _37581_;
  wire _37582_;
  wire _37583_;
  wire _37584_;
  wire _37585_;
  wire _37586_;
  wire _37587_;
  wire _37588_;
  wire _37589_;
  wire _37590_;
  wire _37591_;
  wire _37592_;
  wire _37593_;
  wire _37594_;
  wire _37595_;
  wire _37596_;
  wire _37597_;
  wire _37598_;
  wire _37599_;
  wire _37600_;
  wire _37601_;
  wire _37602_;
  wire _37603_;
  wire _37604_;
  wire _37605_;
  wire _37606_;
  wire _37607_;
  wire _37608_;
  wire _37609_;
  wire _37610_;
  wire _37611_;
  wire _37612_;
  wire _37613_;
  wire _37614_;
  wire _37615_;
  wire _37616_;
  wire _37617_;
  wire _37618_;
  wire _37619_;
  wire _37620_;
  wire _37621_;
  wire _37622_;
  wire _37623_;
  wire _37624_;
  wire _37625_;
  wire _37626_;
  wire _37627_;
  wire _37628_;
  wire _37629_;
  wire _37630_;
  wire _37631_;
  wire _37632_;
  wire _37633_;
  wire _37634_;
  wire _37635_;
  wire _37636_;
  wire _37637_;
  wire _37638_;
  wire _37639_;
  wire _37640_;
  wire _37641_;
  wire _37642_;
  wire _37643_;
  wire _37644_;
  wire _37645_;
  wire _37646_;
  wire _37647_;
  wire _37648_;
  wire _37649_;
  wire _37650_;
  wire _37651_;
  wire _37652_;
  wire _37653_;
  wire _37654_;
  wire _37655_;
  wire _37656_;
  wire _37657_;
  wire _37658_;
  wire _37659_;
  wire _37660_;
  wire _37661_;
  wire _37662_;
  wire _37663_;
  wire _37664_;
  wire _37665_;
  wire _37666_;
  wire _37667_;
  wire _37668_;
  wire _37669_;
  wire _37670_;
  wire _37671_;
  wire _37672_;
  wire _37673_;
  wire _37674_;
  wire _37675_;
  wire _37676_;
  wire _37677_;
  wire _37678_;
  wire _37679_;
  wire _37680_;
  wire _37681_;
  wire _37682_;
  wire _37683_;
  wire _37684_;
  wire _37685_;
  wire _37686_;
  wire _37687_;
  wire _37688_;
  wire _37689_;
  wire _37690_;
  wire _37691_;
  wire _37692_;
  wire _37693_;
  wire _37694_;
  wire _37695_;
  wire _37696_;
  wire _37697_;
  wire _37698_;
  wire _37699_;
  wire _37700_;
  wire _37701_;
  wire _37702_;
  wire _37703_;
  wire _37704_;
  wire _37705_;
  wire _37706_;
  wire _37707_;
  wire _37708_;
  wire _37709_;
  wire _37710_;
  wire _37711_;
  wire _37712_;
  wire _37713_;
  wire _37714_;
  wire _37715_;
  wire _37716_;
  wire _37717_;
  wire _37718_;
  wire _37719_;
  wire _37720_;
  wire _37721_;
  wire _37722_;
  wire _37723_;
  wire _37724_;
  wire _37725_;
  wire _37726_;
  wire _37727_;
  wire _37728_;
  wire _37729_;
  wire _37730_;
  wire _37731_;
  wire _37732_;
  wire _37733_;
  wire _37734_;
  wire _37735_;
  wire _37736_;
  wire _37737_;
  wire _37738_;
  wire _37739_;
  wire _37740_;
  wire _37741_;
  wire _37742_;
  wire _37743_;
  wire _37744_;
  wire _37745_;
  wire _37746_;
  wire _37747_;
  wire _37748_;
  wire _37749_;
  wire _37750_;
  wire _37751_;
  wire _37752_;
  wire _37753_;
  wire _37754_;
  wire _37755_;
  wire _37756_;
  wire _37757_;
  wire _37758_;
  wire _37759_;
  wire _37760_;
  wire _37761_;
  wire _37762_;
  wire _37763_;
  wire _37764_;
  wire _37765_;
  wire _37766_;
  wire _37767_;
  wire _37768_;
  wire _37769_;
  wire _37770_;
  wire _37771_;
  wire _37772_;
  wire _37773_;
  wire _37774_;
  wire _37775_;
  wire _37776_;
  wire _37777_;
  wire _37778_;
  wire _37779_;
  wire _37780_;
  wire _37781_;
  wire _37782_;
  wire _37783_;
  wire _37784_;
  wire _37785_;
  wire _37786_;
  wire _37787_;
  wire _37788_;
  wire _37789_;
  wire _37790_;
  wire _37791_;
  wire _37792_;
  wire _37793_;
  wire _37794_;
  wire _37795_;
  wire _37796_;
  wire _37797_;
  wire _37798_;
  wire _37799_;
  wire _37800_;
  wire _37801_;
  wire _37802_;
  wire _37803_;
  wire _37804_;
  wire _37805_;
  wire _37806_;
  wire _37807_;
  wire _37808_;
  wire _37809_;
  wire _37810_;
  wire _37811_;
  wire _37812_;
  wire _37813_;
  wire _37814_;
  wire _37815_;
  wire _37816_;
  wire _37817_;
  wire _37818_;
  wire _37819_;
  wire _37820_;
  wire _37821_;
  wire _37822_;
  wire _37823_;
  wire _37824_;
  wire _37825_;
  wire _37826_;
  wire _37827_;
  wire _37828_;
  wire _37829_;
  wire _37830_;
  wire _37831_;
  wire _37832_;
  wire _37833_;
  wire _37834_;
  wire _37835_;
  wire _37836_;
  wire _37837_;
  wire _37838_;
  wire _37839_;
  wire _37840_;
  wire _37841_;
  wire _37842_;
  wire _37843_;
  wire _37844_;
  wire _37845_;
  wire _37846_;
  wire _37847_;
  wire _37848_;
  wire _37849_;
  wire _37850_;
  wire _37851_;
  wire _37852_;
  wire _37853_;
  wire _37854_;
  wire _37855_;
  wire _37856_;
  wire _37857_;
  wire _37858_;
  wire _37859_;
  wire _37860_;
  wire _37861_;
  wire _37862_;
  wire _37863_;
  wire _37864_;
  wire _37865_;
  wire _37866_;
  wire _37867_;
  wire _37868_;
  wire _37869_;
  wire _37870_;
  wire _37871_;
  wire _37872_;
  wire _37873_;
  wire _37874_;
  wire _37875_;
  wire _37876_;
  wire _37877_;
  wire _37878_;
  wire _37879_;
  wire _37880_;
  wire _37881_;
  wire _37882_;
  wire _37883_;
  wire _37884_;
  wire _37885_;
  wire _37886_;
  wire _37887_;
  wire _37888_;
  wire _37889_;
  wire _37890_;
  wire _37891_;
  wire _37892_;
  wire _37893_;
  wire _37894_;
  wire _37895_;
  wire _37896_;
  wire _37897_;
  wire _37898_;
  wire _37899_;
  wire _37900_;
  wire _37901_;
  wire _37902_;
  wire _37903_;
  wire _37904_;
  wire _37905_;
  wire _37906_;
  wire _37907_;
  wire _37908_;
  wire _37909_;
  wire _37910_;
  wire _37911_;
  wire _37912_;
  wire _37913_;
  wire _37914_;
  wire _37915_;
  wire _37916_;
  wire _37917_;
  wire _37918_;
  wire _37919_;
  wire _37920_;
  wire _37921_;
  wire _37922_;
  wire _37923_;
  wire _37924_;
  wire _37925_;
  wire _37926_;
  wire _37927_;
  wire _37928_;
  wire _37929_;
  wire _37930_;
  wire _37931_;
  wire _37932_;
  wire _37933_;
  wire _37934_;
  wire _37935_;
  wire _37936_;
  wire _37937_;
  wire _37938_;
  wire _37939_;
  wire _37940_;
  wire _37941_;
  wire _37942_;
  wire _37943_;
  wire _37944_;
  wire _37945_;
  wire _37946_;
  wire _37947_;
  wire _37948_;
  wire _37949_;
  wire _37950_;
  wire _37951_;
  wire _37952_;
  wire _37953_;
  wire _37954_;
  wire _37955_;
  wire _37956_;
  wire _37957_;
  wire _37958_;
  wire _37959_;
  wire _37960_;
  wire _37961_;
  wire _37962_;
  wire _37963_;
  wire _37964_;
  wire _37965_;
  wire _37966_;
  wire _37967_;
  wire _37968_;
  wire _37969_;
  wire _37970_;
  wire _37971_;
  wire _37972_;
  wire _37973_;
  wire _37974_;
  wire _37975_;
  wire _37976_;
  wire _37977_;
  wire _37978_;
  wire _37979_;
  wire _37980_;
  wire _37981_;
  wire _37982_;
  wire _37983_;
  wire _37984_;
  wire _37985_;
  wire _37986_;
  wire _37987_;
  wire _37988_;
  wire _37989_;
  wire _37990_;
  wire _37991_;
  wire _37992_;
  wire _37993_;
  wire _37994_;
  wire _37995_;
  wire _37996_;
  wire _37997_;
  wire _37998_;
  wire _37999_;
  wire _38000_;
  wire _38001_;
  wire _38002_;
  wire _38003_;
  wire _38004_;
  wire _38005_;
  wire _38006_;
  wire _38007_;
  wire _38008_;
  wire _38009_;
  wire _38010_;
  wire _38011_;
  wire _38012_;
  wire _38013_;
  wire _38014_;
  wire _38015_;
  wire _38016_;
  wire _38017_;
  wire _38018_;
  wire _38019_;
  wire _38020_;
  wire _38021_;
  wire _38022_;
  wire _38023_;
  wire _38024_;
  wire _38025_;
  wire _38026_;
  wire _38027_;
  wire _38028_;
  wire _38029_;
  wire _38030_;
  wire _38031_;
  wire _38032_;
  wire _38033_;
  wire _38034_;
  wire _38035_;
  wire _38036_;
  wire _38037_;
  wire _38038_;
  wire _38039_;
  wire _38040_;
  wire _38041_;
  wire _38042_;
  wire _38043_;
  wire _38044_;
  wire _38045_;
  wire _38046_;
  wire _38047_;
  wire _38048_;
  wire _38049_;
  wire _38050_;
  wire _38051_;
  wire _38052_;
  wire _38053_;
  wire _38054_;
  wire _38055_;
  wire _38056_;
  wire _38057_;
  wire _38058_;
  wire _38059_;
  wire _38060_;
  wire _38061_;
  wire _38062_;
  wire _38063_;
  wire _38064_;
  wire _38065_;
  wire _38066_;
  wire _38067_;
  wire _38068_;
  wire _38069_;
  wire _38070_;
  wire _38071_;
  wire _38072_;
  wire _38073_;
  wire _38074_;
  wire _38075_;
  wire _38076_;
  wire _38077_;
  wire _38078_;
  wire _38079_;
  wire _38080_;
  wire _38081_;
  wire _38082_;
  wire _38083_;
  wire _38084_;
  wire _38085_;
  wire _38086_;
  wire _38087_;
  wire _38088_;
  wire _38089_;
  wire _38090_;
  wire _38091_;
  wire _38092_;
  wire _38093_;
  wire _38094_;
  wire _38095_;
  wire _38096_;
  wire _38097_;
  wire _38098_;
  wire _38099_;
  wire _38100_;
  wire _38101_;
  wire _38102_;
  wire _38103_;
  wire _38104_;
  wire _38105_;
  wire _38106_;
  wire _38107_;
  wire _38108_;
  wire _38109_;
  wire _38110_;
  wire _38111_;
  wire _38112_;
  wire _38113_;
  wire _38114_;
  wire _38115_;
  wire _38116_;
  wire _38117_;
  wire _38118_;
  wire _38119_;
  wire _38120_;
  wire _38121_;
  wire _38122_;
  wire _38123_;
  wire _38124_;
  wire _38125_;
  wire _38126_;
  wire _38127_;
  wire _38128_;
  wire _38129_;
  wire _38130_;
  wire _38131_;
  wire _38132_;
  wire _38133_;
  wire _38134_;
  wire _38135_;
  wire _38136_;
  wire _38137_;
  wire _38138_;
  wire _38139_;
  wire _38140_;
  wire _38141_;
  wire _38142_;
  wire _38143_;
  wire _38144_;
  wire _38145_;
  wire _38146_;
  wire _38147_;
  wire _38148_;
  wire _38149_;
  wire _38150_;
  wire _38151_;
  wire _38152_;
  wire _38153_;
  wire _38154_;
  wire _38155_;
  wire _38156_;
  wire _38157_;
  wire _38158_;
  wire _38159_;
  wire _38160_;
  wire _38161_;
  wire _38162_;
  wire _38163_;
  wire _38164_;
  wire _38165_;
  wire _38166_;
  wire _38167_;
  wire _38168_;
  wire _38169_;
  wire _38170_;
  wire _38171_;
  wire _38172_;
  wire _38173_;
  wire _38174_;
  wire _38175_;
  wire _38176_;
  wire _38177_;
  wire _38178_;
  wire _38179_;
  wire _38180_;
  wire _38181_;
  wire _38182_;
  wire _38183_;
  wire _38184_;
  wire _38185_;
  wire _38186_;
  wire _38187_;
  wire _38188_;
  wire _38189_;
  wire _38190_;
  wire _38191_;
  wire _38192_;
  wire _38193_;
  wire _38194_;
  wire _38195_;
  wire _38196_;
  wire _38197_;
  wire _38198_;
  wire _38199_;
  wire _38200_;
  wire _38201_;
  wire _38202_;
  wire _38203_;
  wire _38204_;
  wire _38205_;
  wire _38206_;
  wire _38207_;
  wire _38208_;
  wire _38209_;
  wire _38210_;
  wire _38211_;
  wire _38212_;
  wire _38213_;
  wire _38214_;
  wire _38215_;
  wire _38216_;
  wire _38217_;
  wire _38218_;
  wire _38219_;
  wire _38220_;
  wire _38221_;
  wire _38222_;
  wire _38223_;
  wire _38224_;
  wire _38225_;
  wire _38226_;
  wire _38227_;
  wire _38228_;
  wire _38229_;
  wire _38230_;
  wire _38231_;
  wire _38232_;
  wire _38233_;
  wire _38234_;
  wire _38235_;
  wire _38236_;
  wire _38237_;
  wire _38238_;
  wire _38239_;
  wire _38240_;
  wire _38241_;
  wire _38242_;
  wire _38243_;
  wire _38244_;
  wire _38245_;
  wire _38246_;
  wire _38247_;
  wire _38248_;
  wire _38249_;
  wire _38250_;
  wire _38251_;
  wire _38252_;
  wire _38253_;
  wire _38254_;
  wire _38255_;
  wire _38256_;
  wire _38257_;
  wire _38258_;
  wire _38259_;
  wire _38260_;
  wire _38261_;
  wire _38262_;
  wire _38263_;
  wire _38264_;
  wire _38265_;
  wire _38266_;
  wire _38267_;
  wire _38268_;
  wire _38269_;
  wire _38270_;
  wire _38271_;
  wire _38272_;
  wire _38273_;
  wire _38274_;
  wire _38275_;
  wire _38276_;
  wire _38277_;
  wire _38278_;
  wire _38279_;
  wire _38280_;
  wire _38281_;
  wire _38282_;
  wire _38283_;
  wire _38284_;
  wire _38285_;
  wire _38286_;
  wire _38287_;
  wire _38288_;
  wire _38289_;
  wire _38290_;
  wire _38291_;
  wire _38292_;
  wire _38293_;
  wire _38294_;
  wire _38295_;
  wire _38296_;
  wire _38297_;
  wire _38298_;
  wire _38299_;
  wire _38300_;
  wire _38301_;
  wire _38302_;
  wire _38303_;
  wire _38304_;
  wire _38305_;
  wire _38306_;
  wire _38307_;
  wire _38308_;
  wire _38309_;
  wire _38310_;
  wire _38311_;
  wire _38312_;
  wire _38313_;
  wire _38314_;
  wire _38315_;
  wire _38316_;
  wire _38317_;
  wire _38318_;
  wire _38319_;
  wire _38320_;
  wire _38321_;
  wire _38322_;
  wire _38323_;
  wire _38324_;
  wire _38325_;
  wire _38326_;
  wire _38327_;
  wire _38328_;
  wire _38329_;
  wire _38330_;
  wire _38331_;
  wire _38332_;
  wire _38333_;
  wire _38334_;
  wire _38335_;
  wire _38336_;
  wire _38337_;
  wire _38338_;
  wire _38339_;
  wire _38340_;
  wire _38341_;
  wire _38342_;
  wire _38343_;
  wire _38344_;
  wire _38345_;
  wire _38346_;
  wire _38347_;
  wire _38348_;
  wire _38349_;
  wire _38350_;
  wire _38351_;
  wire _38352_;
  wire _38353_;
  wire _38354_;
  wire _38355_;
  wire _38356_;
  wire _38357_;
  wire _38358_;
  wire _38359_;
  wire _38360_;
  wire _38361_;
  wire _38362_;
  wire _38363_;
  wire _38364_;
  wire _38365_;
  wire _38366_;
  wire _38367_;
  wire _38368_;
  wire _38369_;
  wire _38370_;
  wire _38371_;
  wire _38372_;
  wire _38373_;
  wire _38374_;
  wire _38375_;
  wire _38376_;
  wire _38377_;
  wire _38378_;
  wire _38379_;
  wire _38380_;
  wire _38381_;
  wire _38382_;
  wire _38383_;
  wire _38384_;
  wire _38385_;
  wire _38386_;
  wire _38387_;
  wire _38388_;
  wire _38389_;
  wire _38390_;
  wire _38391_;
  wire _38392_;
  wire _38393_;
  wire _38394_;
  wire _38395_;
  wire _38396_;
  wire _38397_;
  wire _38398_;
  wire _38399_;
  wire _38400_;
  wire _38401_;
  wire _38402_;
  wire _38403_;
  wire _38404_;
  wire _38405_;
  wire _38406_;
  wire _38407_;
  wire _38408_;
  wire _38409_;
  wire _38410_;
  wire _38411_;
  wire _38412_;
  wire _38413_;
  wire _38414_;
  wire _38415_;
  wire _38416_;
  wire _38417_;
  wire _38418_;
  wire _38419_;
  wire _38420_;
  wire _38421_;
  wire _38422_;
  wire _38423_;
  wire _38424_;
  wire _38425_;
  wire _38426_;
  wire _38427_;
  wire _38428_;
  wire _38429_;
  wire _38430_;
  wire _38431_;
  wire _38432_;
  wire _38433_;
  wire _38434_;
  wire _38435_;
  wire _38436_;
  wire _38437_;
  wire _38438_;
  wire _38439_;
  wire _38440_;
  wire _38441_;
  wire _38442_;
  wire _38443_;
  wire _38444_;
  wire _38445_;
  wire _38446_;
  wire _38447_;
  wire _38448_;
  wire _38449_;
  wire _38450_;
  wire _38451_;
  wire _38452_;
  wire _38453_;
  wire _38454_;
  wire _38455_;
  wire _38456_;
  wire _38457_;
  wire _38458_;
  wire _38459_;
  wire _38460_;
  wire _38461_;
  wire _38462_;
  wire _38463_;
  wire _38464_;
  wire _38465_;
  wire _38466_;
  wire _38467_;
  wire _38468_;
  wire _38469_;
  wire _38470_;
  wire _38471_;
  wire _38472_;
  wire _38473_;
  wire _38474_;
  wire _38475_;
  wire _38476_;
  wire _38477_;
  wire _38478_;
  wire _38479_;
  wire _38480_;
  wire _38481_;
  wire _38482_;
  wire _38483_;
  wire _38484_;
  wire _38485_;
  wire _38486_;
  wire _38487_;
  wire _38488_;
  wire _38489_;
  wire _38490_;
  wire _38491_;
  wire _38492_;
  wire _38493_;
  wire _38494_;
  wire _38495_;
  wire _38496_;
  wire _38497_;
  wire _38498_;
  wire _38499_;
  wire _38500_;
  wire _38501_;
  wire _38502_;
  wire _38503_;
  wire _38504_;
  wire _38505_;
  wire _38506_;
  wire _38507_;
  wire _38508_;
  wire _38509_;
  wire _38510_;
  wire _38511_;
  wire _38512_;
  wire _38513_;
  wire _38514_;
  wire _38515_;
  wire _38516_;
  wire _38517_;
  wire _38518_;
  wire _38519_;
  wire _38520_;
  wire _38521_;
  wire _38522_;
  wire _38523_;
  wire _38524_;
  wire _38525_;
  wire _38526_;
  wire _38527_;
  wire _38528_;
  wire _38529_;
  wire _38530_;
  wire _38531_;
  wire _38532_;
  wire _38533_;
  wire _38534_;
  wire _38535_;
  wire _38536_;
  wire _38537_;
  wire _38538_;
  wire _38539_;
  wire _38540_;
  wire _38541_;
  wire _38542_;
  wire _38543_;
  wire _38544_;
  wire _38545_;
  wire _38546_;
  wire _38547_;
  wire _38548_;
  wire _38549_;
  wire _38550_;
  wire _38551_;
  wire _38552_;
  wire _38553_;
  wire _38554_;
  wire _38555_;
  wire _38556_;
  wire _38557_;
  wire _38558_;
  wire _38559_;
  wire _38560_;
  wire _38561_;
  wire _38562_;
  wire _38563_;
  wire _38564_;
  wire _38565_;
  wire _38566_;
  wire _38567_;
  wire _38568_;
  wire _38569_;
  wire _38570_;
  wire _38571_;
  wire _38572_;
  wire _38573_;
  wire _38574_;
  wire _38575_;
  wire _38576_;
  wire _38577_;
  wire _38578_;
  wire _38579_;
  wire _38580_;
  wire _38581_;
  wire _38582_;
  wire _38583_;
  wire _38584_;
  wire _38585_;
  wire _38586_;
  wire _38587_;
  wire _38588_;
  wire _38589_;
  wire _38590_;
  wire _38591_;
  wire _38592_;
  wire _38593_;
  wire _38594_;
  wire _38595_;
  wire _38596_;
  wire _38597_;
  wire _38598_;
  wire _38599_;
  wire _38600_;
  wire _38601_;
  wire _38602_;
  wire _38603_;
  wire _38604_;
  wire _38605_;
  wire _38606_;
  wire _38607_;
  wire _38608_;
  wire _38609_;
  wire _38610_;
  wire _38611_;
  wire _38612_;
  wire _38613_;
  wire _38614_;
  wire _38615_;
  wire _38616_;
  wire _38617_;
  wire _38618_;
  wire _38619_;
  wire _38620_;
  wire _38621_;
  wire _38622_;
  wire _38623_;
  wire _38624_;
  wire _38625_;
  wire _38626_;
  wire _38627_;
  wire _38628_;
  wire _38629_;
  wire _38630_;
  wire _38631_;
  wire _38632_;
  wire _38633_;
  wire _38634_;
  wire _38635_;
  wire _38636_;
  wire _38637_;
  wire _38638_;
  wire _38639_;
  wire _38640_;
  wire _38641_;
  wire _38642_;
  wire _38643_;
  wire _38644_;
  wire _38645_;
  wire _38646_;
  wire _38647_;
  wire _38648_;
  wire _38649_;
  wire _38650_;
  wire _38651_;
  wire _38652_;
  wire _38653_;
  wire _38654_;
  wire _38655_;
  wire _38656_;
  wire _38657_;
  wire _38658_;
  wire _38659_;
  wire _38660_;
  wire _38661_;
  wire _38662_;
  wire _38663_;
  wire _38664_;
  wire _38665_;
  wire _38666_;
  wire _38667_;
  wire _38668_;
  wire _38669_;
  wire _38670_;
  wire _38671_;
  wire _38672_;
  wire _38673_;
  wire _38674_;
  wire _38675_;
  wire _38676_;
  wire _38677_;
  wire _38678_;
  wire _38679_;
  wire _38680_;
  wire _38681_;
  wire _38682_;
  wire _38683_;
  wire _38684_;
  wire _38685_;
  wire _38686_;
  wire _38687_;
  wire _38688_;
  wire _38689_;
  wire _38690_;
  wire _38691_;
  wire _38692_;
  wire _38693_;
  wire _38694_;
  wire _38695_;
  wire _38696_;
  wire _38697_;
  wire _38698_;
  wire _38699_;
  wire _38700_;
  wire _38701_;
  wire _38702_;
  wire _38703_;
  wire _38704_;
  wire _38705_;
  wire _38706_;
  wire _38707_;
  wire _38708_;
  wire _38709_;
  wire _38710_;
  wire _38711_;
  wire _38712_;
  wire _38713_;
  wire _38714_;
  wire _38715_;
  wire _38716_;
  wire _38717_;
  wire _38718_;
  wire _38719_;
  wire _38720_;
  wire _38721_;
  wire _38722_;
  wire _38723_;
  wire _38724_;
  wire _38725_;
  wire _38726_;
  wire _38727_;
  wire _38728_;
  wire _38729_;
  wire _38730_;
  wire _38731_;
  wire _38732_;
  wire _38733_;
  wire _38734_;
  wire _38735_;
  wire _38736_;
  wire _38737_;
  wire _38738_;
  wire _38739_;
  wire _38740_;
  wire _38741_;
  wire _38742_;
  wire _38743_;
  wire _38744_;
  wire _38745_;
  wire _38746_;
  wire _38747_;
  wire _38748_;
  wire _38749_;
  wire _38750_;
  wire _38751_;
  wire _38752_;
  wire _38753_;
  wire _38754_;
  wire _38755_;
  wire _38756_;
  wire _38757_;
  wire _38758_;
  wire _38759_;
  wire _38760_;
  wire _38761_;
  wire _38762_;
  wire _38763_;
  wire _38764_;
  wire _38765_;
  wire _38766_;
  wire _38767_;
  wire _38768_;
  wire _38769_;
  wire _38770_;
  wire _38771_;
  wire _38772_;
  wire _38773_;
  wire _38774_;
  wire _38775_;
  wire _38776_;
  wire _38777_;
  wire _38778_;
  wire _38779_;
  wire _38780_;
  wire _38781_;
  wire _38782_;
  wire _38783_;
  wire _38784_;
  wire _38785_;
  wire _38786_;
  wire _38787_;
  wire _38788_;
  wire _38789_;
  wire _38790_;
  wire _38791_;
  wire _38792_;
  wire _38793_;
  wire _38794_;
  wire _38795_;
  wire _38796_;
  wire _38797_;
  wire _38798_;
  wire _38799_;
  wire _38800_;
  wire _38801_;
  wire _38802_;
  wire _38803_;
  wire _38804_;
  wire _38805_;
  wire _38806_;
  wire _38807_;
  wire _38808_;
  wire _38809_;
  wire _38810_;
  wire _38811_;
  wire _38812_;
  wire _38813_;
  wire _38814_;
  wire _38815_;
  wire _38816_;
  wire _38817_;
  wire _38818_;
  wire _38819_;
  wire _38820_;
  wire _38821_;
  wire _38822_;
  wire _38823_;
  wire _38824_;
  wire _38825_;
  wire _38826_;
  wire _38827_;
  wire _38828_;
  wire _38829_;
  wire _38830_;
  wire _38831_;
  wire _38832_;
  wire _38833_;
  wire _38834_;
  wire _38835_;
  wire _38836_;
  wire _38837_;
  wire _38838_;
  wire _38839_;
  wire _38840_;
  wire _38841_;
  wire _38842_;
  wire _38843_;
  wire _38844_;
  wire _38845_;
  wire _38846_;
  wire _38847_;
  wire _38848_;
  wire _38849_;
  wire _38850_;
  wire _38851_;
  wire _38852_;
  wire _38853_;
  wire _38854_;
  wire _38855_;
  wire _38856_;
  wire _38857_;
  wire _38858_;
  wire _38859_;
  wire _38860_;
  wire _38861_;
  wire _38862_;
  wire _38863_;
  wire _38864_;
  wire _38865_;
  wire _38866_;
  wire _38867_;
  wire _38868_;
  wire _38869_;
  wire _38870_;
  wire _38871_;
  wire _38872_;
  wire _38873_;
  wire _38874_;
  wire _38875_;
  wire _38876_;
  wire _38877_;
  wire _38878_;
  wire _38879_;
  wire _38880_;
  wire _38881_;
  wire _38882_;
  wire _38883_;
  wire _38884_;
  wire _38885_;
  wire _38886_;
  wire _38887_;
  wire _38888_;
  wire _38889_;
  wire _38890_;
  wire _38891_;
  wire _38892_;
  wire _38893_;
  wire _38894_;
  wire _38895_;
  wire _38896_;
  wire _38897_;
  wire _38898_;
  wire _38899_;
  wire _38900_;
  wire _38901_;
  wire _38902_;
  wire _38903_;
  wire _38904_;
  wire _38905_;
  wire _38906_;
  wire _38907_;
  wire _38908_;
  wire _38909_;
  wire _38910_;
  wire _38911_;
  wire _38912_;
  wire _38913_;
  wire _38914_;
  wire _38915_;
  wire _38916_;
  wire _38917_;
  wire _38918_;
  wire _38919_;
  wire _38920_;
  wire _38921_;
  wire _38922_;
  wire _38923_;
  wire _38924_;
  wire _38925_;
  wire _38926_;
  wire _38927_;
  wire _38928_;
  wire _38929_;
  wire _38930_;
  wire _38931_;
  wire _38932_;
  wire _38933_;
  wire _38934_;
  wire _38935_;
  wire _38936_;
  wire _38937_;
  wire _38938_;
  wire _38939_;
  wire _38940_;
  wire _38941_;
  wire _38942_;
  wire _38943_;
  wire _38944_;
  wire _38945_;
  wire _38946_;
  wire _38947_;
  wire _38948_;
  wire _38949_;
  wire _38950_;
  wire _38951_;
  wire _38952_;
  wire _38953_;
  wire _38954_;
  wire _38955_;
  wire _38956_;
  wire _38957_;
  wire _38958_;
  wire _38959_;
  wire _38960_;
  wire _38961_;
  wire _38962_;
  wire _38963_;
  wire _38964_;
  wire _38965_;
  wire _38966_;
  wire _38967_;
  wire _38968_;
  wire _38969_;
  wire _38970_;
  wire _38971_;
  wire _38972_;
  wire _38973_;
  wire _38974_;
  wire _38975_;
  wire _38976_;
  wire _38977_;
  wire _38978_;
  wire _38979_;
  wire _38980_;
  wire _38981_;
  wire _38982_;
  wire _38983_;
  wire _38984_;
  wire _38985_;
  wire _38986_;
  wire _38987_;
  wire _38988_;
  wire _38989_;
  wire _38990_;
  wire _38991_;
  wire _38992_;
  wire _38993_;
  wire _38994_;
  wire _38995_;
  wire _38996_;
  wire _38997_;
  wire _38998_;
  wire _38999_;
  wire _39000_;
  wire _39001_;
  wire _39002_;
  wire _39003_;
  wire _39004_;
  wire _39005_;
  wire _39006_;
  wire _39007_;
  wire _39008_;
  wire _39009_;
  wire _39010_;
  wire _39011_;
  wire _39012_;
  wire _39013_;
  wire _39014_;
  wire _39015_;
  wire _39016_;
  wire _39017_;
  wire _39018_;
  wire _39019_;
  wire _39020_;
  wire _39021_;
  wire _39022_;
  wire _39023_;
  wire _39024_;
  wire _39025_;
  wire _39026_;
  wire _39027_;
  wire _39028_;
  wire _39029_;
  wire _39030_;
  wire _39031_;
  wire _39032_;
  wire _39033_;
  wire _39034_;
  wire _39035_;
  wire _39036_;
  wire _39037_;
  wire _39038_;
  wire _39039_;
  wire _39040_;
  wire _39041_;
  wire _39042_;
  wire _39043_;
  wire _39044_;
  wire _39045_;
  wire _39046_;
  wire _39047_;
  wire _39048_;
  wire _39049_;
  wire _39050_;
  wire _39051_;
  wire _39052_;
  wire _39053_;
  wire _39054_;
  wire _39055_;
  wire _39056_;
  wire _39057_;
  wire _39058_;
  wire _39059_;
  wire _39060_;
  wire _39061_;
  wire _39062_;
  wire _39063_;
  wire _39064_;
  wire _39065_;
  wire _39066_;
  wire _39067_;
  wire _39068_;
  wire _39069_;
  wire _39070_;
  wire _39071_;
  wire _39072_;
  wire _39073_;
  wire _39074_;
  wire _39075_;
  wire _39076_;
  wire _39077_;
  wire _39078_;
  wire _39079_;
  wire _39080_;
  wire _39081_;
  wire _39082_;
  wire _39083_;
  wire _39084_;
  wire _39085_;
  wire _39086_;
  wire _39087_;
  wire _39088_;
  wire _39089_;
  wire _39090_;
  wire _39091_;
  wire _39092_;
  wire _39093_;
  wire _39094_;
  wire _39095_;
  wire _39096_;
  wire _39097_;
  wire _39098_;
  wire _39099_;
  wire _39100_;
  wire _39101_;
  wire _39102_;
  wire _39103_;
  wire _39104_;
  wire _39105_;
  wire _39106_;
  wire _39107_;
  wire _39108_;
  wire _39109_;
  wire _39110_;
  wire _39111_;
  wire _39112_;
  wire _39113_;
  wire _39114_;
  wire _39115_;
  wire _39116_;
  wire _39117_;
  wire _39118_;
  wire _39119_;
  wire _39120_;
  wire _39121_;
  wire _39122_;
  wire _39123_;
  wire _39124_;
  wire _39125_;
  wire _39126_;
  wire _39127_;
  wire _39128_;
  wire _39129_;
  wire _39130_;
  wire _39131_;
  wire _39132_;
  wire _39133_;
  wire _39134_;
  wire _39135_;
  wire _39136_;
  wire _39137_;
  wire _39138_;
  wire _39139_;
  wire _39140_;
  wire _39141_;
  wire _39142_;
  wire _39143_;
  wire _39144_;
  wire _39145_;
  wire _39146_;
  wire _39147_;
  wire _39148_;
  wire _39149_;
  wire _39150_;
  wire _39151_;
  wire _39152_;
  wire _39153_;
  wire _39154_;
  wire _39155_;
  wire _39156_;
  wire _39157_;
  wire _39158_;
  wire _39159_;
  wire _39160_;
  wire _39161_;
  wire _39162_;
  wire _39163_;
  wire _39164_;
  wire _39165_;
  wire _39166_;
  wire _39167_;
  wire _39168_;
  wire _39169_;
  wire _39170_;
  wire _39171_;
  wire _39172_;
  wire _39173_;
  wire _39174_;
  wire _39175_;
  wire _39176_;
  wire _39177_;
  wire _39178_;
  wire _39179_;
  wire _39180_;
  wire _39181_;
  wire _39182_;
  wire _39183_;
  wire _39184_;
  wire _39185_;
  wire _39186_;
  wire _39187_;
  wire _39188_;
  wire _39189_;
  wire _39190_;
  wire _39191_;
  wire _39192_;
  wire _39193_;
  wire _39194_;
  wire _39195_;
  wire _39196_;
  wire _39197_;
  wire _39198_;
  wire _39199_;
  wire _39200_;
  wire _39201_;
  wire _39202_;
  wire _39203_;
  wire _39204_;
  wire _39205_;
  wire _39206_;
  wire _39207_;
  wire _39208_;
  wire _39209_;
  wire _39210_;
  wire _39211_;
  wire _39212_;
  wire _39213_;
  wire _39214_;
  wire _39215_;
  wire _39216_;
  wire _39217_;
  wire _39218_;
  wire _39219_;
  wire _39220_;
  wire _39221_;
  wire _39222_;
  wire _39223_;
  wire _39224_;
  wire _39225_;
  wire _39226_;
  wire _39227_;
  wire _39228_;
  wire _39229_;
  wire _39230_;
  wire _39231_;
  wire _39232_;
  wire _39233_;
  wire _39234_;
  wire _39235_;
  wire _39236_;
  wire _39237_;
  wire _39238_;
  wire _39239_;
  wire _39240_;
  wire _39241_;
  wire _39242_;
  wire _39243_;
  wire _39244_;
  wire _39245_;
  wire _39246_;
  wire _39247_;
  wire _39248_;
  wire _39249_;
  wire _39250_;
  wire _39251_;
  wire _39252_;
  wire _39253_;
  wire _39254_;
  wire _39255_;
  wire _39256_;
  wire _39257_;
  wire _39258_;
  wire _39259_;
  wire _39260_;
  wire _39261_;
  wire _39262_;
  wire _39263_;
  wire _39264_;
  wire _39265_;
  wire _39266_;
  wire _39267_;
  wire _39268_;
  wire _39269_;
  wire _39270_;
  wire _39271_;
  wire _39272_;
  wire _39273_;
  wire _39274_;
  wire _39275_;
  wire _39276_;
  wire _39277_;
  wire _39278_;
  wire _39279_;
  wire _39280_;
  wire _39281_;
  wire _39282_;
  wire _39283_;
  wire _39284_;
  wire _39285_;
  wire _39286_;
  wire _39287_;
  wire _39288_;
  wire _39289_;
  wire _39290_;
  wire _39291_;
  wire _39292_;
  wire _39293_;
  wire _39294_;
  wire _39295_;
  wire _39296_;
  wire _39297_;
  wire _39298_;
  wire _39299_;
  wire _39300_;
  wire _39301_;
  wire _39302_;
  wire _39303_;
  wire _39304_;
  wire _39305_;
  wire _39306_;
  wire _39307_;
  wire _39308_;
  wire _39309_;
  wire _39310_;
  wire _39311_;
  wire _39312_;
  wire _39313_;
  wire _39314_;
  wire _39315_;
  wire _39316_;
  wire _39317_;
  wire _39318_;
  wire _39319_;
  wire _39320_;
  wire _39321_;
  wire _39322_;
  wire _39323_;
  wire _39324_;
  wire _39325_;
  wire _39326_;
  wire _39327_;
  wire _39328_;
  wire _39329_;
  wire _39330_;
  wire _39331_;
  wire _39332_;
  wire _39333_;
  wire _39334_;
  wire _39335_;
  wire _39336_;
  wire _39337_;
  wire _39338_;
  wire _39339_;
  wire _39340_;
  wire _39341_;
  wire _39342_;
  wire _39343_;
  wire _39344_;
  wire _39345_;
  wire _39346_;
  wire _39347_;
  wire _39348_;
  wire _39349_;
  wire _39350_;
  wire _39351_;
  wire _39352_;
  wire _39353_;
  wire _39354_;
  wire _39355_;
  wire _39356_;
  wire _39357_;
  wire _39358_;
  wire _39359_;
  wire _39360_;
  wire _39361_;
  wire _39362_;
  wire _39363_;
  wire _39364_;
  wire _39365_;
  wire _39366_;
  wire _39367_;
  wire _39368_;
  wire _39369_;
  wire _39370_;
  wire _39371_;
  wire _39372_;
  wire _39373_;
  wire _39374_;
  wire _39375_;
  wire _39376_;
  wire _39377_;
  wire _39378_;
  wire _39379_;
  wire _39380_;
  wire _39381_;
  wire _39382_;
  wire _39383_;
  wire _39384_;
  wire _39385_;
  wire _39386_;
  wire _39387_;
  wire _39388_;
  wire _39389_;
  wire _39390_;
  wire _39391_;
  wire _39392_;
  wire _39393_;
  wire _39394_;
  wire _39395_;
  wire _39396_;
  wire _39397_;
  wire _39398_;
  wire _39399_;
  wire _39400_;
  wire _39401_;
  wire _39402_;
  wire _39403_;
  wire _39404_;
  wire _39405_;
  wire _39406_;
  wire _39407_;
  wire _39408_;
  wire _39409_;
  wire _39410_;
  wire _39411_;
  wire _39412_;
  wire _39413_;
  wire _39414_;
  wire _39415_;
  wire _39416_;
  wire _39417_;
  wire _39418_;
  wire _39419_;
  wire _39420_;
  wire _39421_;
  wire _39422_;
  wire _39423_;
  wire _39424_;
  wire _39425_;
  wire _39426_;
  wire _39427_;
  wire _39428_;
  wire _39429_;
  wire _39430_;
  wire _39431_;
  wire _39432_;
  wire _39433_;
  wire _39434_;
  wire _39435_;
  wire _39436_;
  wire _39437_;
  wire _39438_;
  wire _39439_;
  wire _39440_;
  wire _39441_;
  wire _39442_;
  wire _39443_;
  wire _39444_;
  wire _39445_;
  wire _39446_;
  wire _39447_;
  wire _39448_;
  wire _39449_;
  wire _39450_;
  wire _39451_;
  wire _39452_;
  wire _39453_;
  wire _39454_;
  wire _39455_;
  wire _39456_;
  wire _39457_;
  wire _39458_;
  wire _39459_;
  wire _39460_;
  wire _39461_;
  wire _39462_;
  wire _39463_;
  wire _39464_;
  wire _39465_;
  wire _39466_;
  wire _39467_;
  wire _39468_;
  wire _39469_;
  wire _39470_;
  wire _39471_;
  wire _39472_;
  wire _39473_;
  wire _39474_;
  wire _39475_;
  wire _39476_;
  wire _39477_;
  wire _39478_;
  wire _39479_;
  wire _39480_;
  wire _39481_;
  wire _39482_;
  wire _39483_;
  wire _39484_;
  wire _39485_;
  wire _39486_;
  wire _39487_;
  wire _39488_;
  wire _39489_;
  wire _39490_;
  wire _39491_;
  wire _39492_;
  wire _39493_;
  wire _39494_;
  wire _39495_;
  wire _39496_;
  wire _39497_;
  wire _39498_;
  wire _39499_;
  wire _39500_;
  wire _39501_;
  wire _39502_;
  wire _39503_;
  wire _39504_;
  wire _39505_;
  wire _39506_;
  wire _39507_;
  wire _39508_;
  wire _39509_;
  wire _39510_;
  wire _39511_;
  wire _39512_;
  wire _39513_;
  wire _39514_;
  wire _39515_;
  wire _39516_;
  wire _39517_;
  wire _39518_;
  wire _39519_;
  wire _39520_;
  wire _39521_;
  wire _39522_;
  wire _39523_;
  wire _39524_;
  wire _39525_;
  wire _39526_;
  wire _39527_;
  wire _39528_;
  wire _39529_;
  wire _39530_;
  wire _39531_;
  wire _39532_;
  wire _39533_;
  wire _39534_;
  wire _39535_;
  wire _39536_;
  wire _39537_;
  wire _39538_;
  wire _39539_;
  wire _39540_;
  wire _39541_;
  wire _39542_;
  wire _39543_;
  wire _39544_;
  wire _39545_;
  wire _39546_;
  wire _39547_;
  wire _39548_;
  wire _39549_;
  wire _39550_;
  wire _39551_;
  wire _39552_;
  wire _39553_;
  wire _39554_;
  wire _39555_;
  wire _39556_;
  wire _39557_;
  wire _39558_;
  wire _39559_;
  wire _39560_;
  wire _39561_;
  wire _39562_;
  wire _39563_;
  wire _39564_;
  wire _39565_;
  wire _39566_;
  wire _39567_;
  wire _39568_;
  wire _39569_;
  wire _39570_;
  wire _39571_;
  wire _39572_;
  wire _39573_;
  wire _39574_;
  wire _39575_;
  wire _39576_;
  wire _39577_;
  wire _39578_;
  wire _39579_;
  wire _39580_;
  wire _39581_;
  wire _39582_;
  wire _39583_;
  wire _39584_;
  wire _39585_;
  wire _39586_;
  wire _39587_;
  wire _39588_;
  wire _39589_;
  wire _39590_;
  wire _39591_;
  wire _39592_;
  wire _39593_;
  wire _39594_;
  wire _39595_;
  wire _39596_;
  wire _39597_;
  wire _39598_;
  wire _39599_;
  wire _39600_;
  wire _39601_;
  wire _39602_;
  wire _39603_;
  wire _39604_;
  wire _39605_;
  wire _39606_;
  wire _39607_;
  wire _39608_;
  wire _39609_;
  wire _39610_;
  wire _39611_;
  wire _39612_;
  wire _39613_;
  wire _39614_;
  wire _39615_;
  wire _39616_;
  wire _39617_;
  wire _39618_;
  wire _39619_;
  wire _39620_;
  wire _39621_;
  wire _39622_;
  wire _39623_;
  wire _39624_;
  wire _39625_;
  wire _39626_;
  wire _39627_;
  wire _39628_;
  wire _39629_;
  wire _39630_;
  wire _39631_;
  wire _39632_;
  wire _39633_;
  wire _39634_;
  wire _39635_;
  wire _39636_;
  wire _39637_;
  wire _39638_;
  wire _39639_;
  wire _39640_;
  wire _39641_;
  wire _39642_;
  wire _39643_;
  wire _39644_;
  wire _39645_;
  wire _39646_;
  wire _39647_;
  wire _39648_;
  wire _39649_;
  wire _39650_;
  wire _39651_;
  wire _39652_;
  wire _39653_;
  wire _39654_;
  wire _39655_;
  wire _39656_;
  wire _39657_;
  wire _39658_;
  wire _39659_;
  wire _39660_;
  wire _39661_;
  wire _39662_;
  wire _39663_;
  wire _39664_;
  wire _39665_;
  wire _39666_;
  wire _39667_;
  wire _39668_;
  wire _39669_;
  wire _39670_;
  wire _39671_;
  wire _39672_;
  wire _39673_;
  wire _39674_;
  wire _39675_;
  wire _39676_;
  wire _39677_;
  wire _39678_;
  wire _39679_;
  wire _39680_;
  wire _39681_;
  wire _39682_;
  wire _39683_;
  wire _39684_;
  wire _39685_;
  wire _39686_;
  wire _39687_;
  wire _39688_;
  wire _39689_;
  wire _39690_;
  wire _39691_;
  wire _39692_;
  wire _39693_;
  wire _39694_;
  wire _39695_;
  wire _39696_;
  wire _39697_;
  wire _39698_;
  wire _39699_;
  wire _39700_;
  wire _39701_;
  wire _39702_;
  wire _39703_;
  wire _39704_;
  wire _39705_;
  wire _39706_;
  wire _39707_;
  wire _39708_;
  wire _39709_;
  wire _39710_;
  wire _39711_;
  wire _39712_;
  wire _39713_;
  wire _39714_;
  wire _39715_;
  wire _39716_;
  wire _39717_;
  wire _39718_;
  wire _39719_;
  wire _39720_;
  wire _39721_;
  wire _39722_;
  wire _39723_;
  wire _39724_;
  wire _39725_;
  wire _39726_;
  wire _39727_;
  wire _39728_;
  wire _39729_;
  wire _39730_;
  wire _39731_;
  wire _39732_;
  wire _39733_;
  wire _39734_;
  wire _39735_;
  wire _39736_;
  wire _39737_;
  wire _39738_;
  wire _39739_;
  wire _39740_;
  wire _39741_;
  wire _39742_;
  wire _39743_;
  wire _39744_;
  wire _39745_;
  wire _39746_;
  wire _39747_;
  wire _39748_;
  wire _39749_;
  wire _39750_;
  wire _39751_;
  wire _39752_;
  wire _39753_;
  wire _39754_;
  wire _39755_;
  wire _39756_;
  wire _39757_;
  wire _39758_;
  wire _39759_;
  wire _39760_;
  wire _39761_;
  wire _39762_;
  wire _39763_;
  wire _39764_;
  wire _39765_;
  wire _39766_;
  wire _39767_;
  wire _39768_;
  wire _39769_;
  wire _39770_;
  wire _39771_;
  wire _39772_;
  wire _39773_;
  wire _39774_;
  wire _39775_;
  wire _39776_;
  wire _39777_;
  wire _39778_;
  wire _39779_;
  wire _39780_;
  wire _39781_;
  wire _39782_;
  wire _39783_;
  wire _39784_;
  wire _39785_;
  wire _39786_;
  wire _39787_;
  wire _39788_;
  wire _39789_;
  wire _39790_;
  wire _39791_;
  wire _39792_;
  wire _39793_;
  wire _39794_;
  wire _39795_;
  wire _39796_;
  wire _39797_;
  wire _39798_;
  wire _39799_;
  wire _39800_;
  wire _39801_;
  wire _39802_;
  wire _39803_;
  wire _39804_;
  wire _39805_;
  wire _39806_;
  wire _39807_;
  wire _39808_;
  wire _39809_;
  wire _39810_;
  wire _39811_;
  wire _39812_;
  wire _39813_;
  wire _39814_;
  wire _39815_;
  wire _39816_;
  wire _39817_;
  wire _39818_;
  wire _39819_;
  wire _39820_;
  wire _39821_;
  wire _39822_;
  wire _39823_;
  wire _39824_;
  wire _39825_;
  wire _39826_;
  wire _39827_;
  wire _39828_;
  wire _39829_;
  wire _39830_;
  wire _39831_;
  wire _39832_;
  wire _39833_;
  wire _39834_;
  wire _39835_;
  wire _39836_;
  wire _39837_;
  wire _39838_;
  wire _39839_;
  wire _39840_;
  wire _39841_;
  wire _39842_;
  wire _39843_;
  wire _39844_;
  wire _39845_;
  wire _39846_;
  wire _39847_;
  wire _39848_;
  wire _39849_;
  wire _39850_;
  wire _39851_;
  wire _39852_;
  wire _39853_;
  wire _39854_;
  wire _39855_;
  wire _39856_;
  wire _39857_;
  wire _39858_;
  wire _39859_;
  wire _39860_;
  wire _39861_;
  wire _39862_;
  wire _39863_;
  wire _39864_;
  wire _39865_;
  wire _39866_;
  wire _39867_;
  wire _39868_;
  wire _39869_;
  wire _39870_;
  wire _39871_;
  wire _39872_;
  wire _39873_;
  wire _39874_;
  wire _39875_;
  wire _39876_;
  wire _39877_;
  wire _39878_;
  wire _39879_;
  wire _39880_;
  wire _39881_;
  wire _39882_;
  wire _39883_;
  wire _39884_;
  wire _39885_;
  wire _39886_;
  wire _39887_;
  wire _39888_;
  wire _39889_;
  wire _39890_;
  wire _39891_;
  wire _39892_;
  wire _39893_;
  wire _39894_;
  wire _39895_;
  wire _39896_;
  wire _39897_;
  wire _39898_;
  wire _39899_;
  wire _39900_;
  wire _39901_;
  wire _39902_;
  wire _39903_;
  wire _39904_;
  wire _39905_;
  wire _39906_;
  wire _39907_;
  wire _39908_;
  wire _39909_;
  wire _39910_;
  wire _39911_;
  wire _39912_;
  wire _39913_;
  wire _39914_;
  wire _39915_;
  wire _39916_;
  wire _39917_;
  wire _39918_;
  wire _39919_;
  wire _39920_;
  wire _39921_;
  wire _39922_;
  wire _39923_;
  wire _39924_;
  wire _39925_;
  wire _39926_;
  wire _39927_;
  wire _39928_;
  wire _39929_;
  wire _39930_;
  wire _39931_;
  wire _39932_;
  wire _39933_;
  wire _39934_;
  wire _39935_;
  wire _39936_;
  wire _39937_;
  wire _39938_;
  wire _39939_;
  wire _39940_;
  wire _39941_;
  wire _39942_;
  wire _39943_;
  wire _39944_;
  wire _39945_;
  wire _39946_;
  wire _39947_;
  wire _39948_;
  wire _39949_;
  wire _39950_;
  wire _39951_;
  wire _39952_;
  wire _39953_;
  wire _39954_;
  wire _39955_;
  wire _39956_;
  wire _39957_;
  wire _39958_;
  wire _39959_;
  wire _39960_;
  wire _39961_;
  wire _39962_;
  wire _39963_;
  wire _39964_;
  wire _39965_;
  wire _39966_;
  wire _39967_;
  wire _39968_;
  wire _39969_;
  wire _39970_;
  wire _39971_;
  wire _39972_;
  wire _39973_;
  wire _39974_;
  wire _39975_;
  wire _39976_;
  wire _39977_;
  wire _39978_;
  wire _39979_;
  wire _39980_;
  wire _39981_;
  wire _39982_;
  wire _39983_;
  wire _39984_;
  wire _39985_;
  wire _39986_;
  wire _39987_;
  wire _39988_;
  wire _39989_;
  wire _39990_;
  wire _39991_;
  wire _39992_;
  wire _39993_;
  wire _39994_;
  wire _39995_;
  wire _39996_;
  wire _39997_;
  wire _39998_;
  wire _39999_;
  wire _40000_;
  wire _40001_;
  wire _40002_;
  wire _40003_;
  wire _40004_;
  wire _40005_;
  wire _40006_;
  wire _40007_;
  wire _40008_;
  wire _40009_;
  wire _40010_;
  wire _40011_;
  wire _40012_;
  wire _40013_;
  wire _40014_;
  wire _40015_;
  wire _40016_;
  wire _40017_;
  wire _40018_;
  wire _40019_;
  wire _40020_;
  wire _40021_;
  wire _40022_;
  wire _40023_;
  wire _40024_;
  wire _40025_;
  wire _40026_;
  wire _40027_;
  wire _40028_;
  wire _40029_;
  wire _40030_;
  wire _40031_;
  wire _40032_;
  wire _40033_;
  wire _40034_;
  wire _40035_;
  wire _40036_;
  wire _40037_;
  wire _40038_;
  wire _40039_;
  wire _40040_;
  wire _40041_;
  wire _40042_;
  wire _40043_;
  wire _40044_;
  wire _40045_;
  wire _40046_;
  wire _40047_;
  wire _40048_;
  wire _40049_;
  wire _40050_;
  wire _40051_;
  wire _40052_;
  wire _40053_;
  wire _40054_;
  wire _40055_;
  wire _40056_;
  wire _40057_;
  wire _40058_;
  wire _40059_;
  wire _40060_;
  wire _40061_;
  wire _40062_;
  wire _40063_;
  wire _40064_;
  wire _40065_;
  wire _40066_;
  wire _40067_;
  wire _40068_;
  wire _40069_;
  wire _40070_;
  wire _40071_;
  wire _40072_;
  wire _40073_;
  wire _40074_;
  wire _40075_;
  wire _40076_;
  wire _40077_;
  wire _40078_;
  wire _40079_;
  wire _40080_;
  wire _40081_;
  wire _40082_;
  wire _40083_;
  wire _40084_;
  wire _40085_;
  wire _40086_;
  wire _40087_;
  wire _40088_;
  wire _40089_;
  wire _40090_;
  wire _40091_;
  wire _40092_;
  wire _40093_;
  wire _40094_;
  wire _40095_;
  wire _40096_;
  wire _40097_;
  wire _40098_;
  wire _40099_;
  wire _40100_;
  wire _40101_;
  wire _40102_;
  wire _40103_;
  wire _40104_;
  wire _40105_;
  wire _40106_;
  wire _40107_;
  wire _40108_;
  wire _40109_;
  wire _40110_;
  wire _40111_;
  wire _40112_;
  wire _40113_;
  wire _40114_;
  wire _40115_;
  wire _40116_;
  wire _40117_;
  wire _40118_;
  wire _40119_;
  wire _40120_;
  wire _40121_;
  wire _40122_;
  wire _40123_;
  wire _40124_;
  wire _40125_;
  wire _40126_;
  wire _40127_;
  wire _40128_;
  wire _40129_;
  wire _40130_;
  wire _40131_;
  wire _40132_;
  wire _40133_;
  wire _40134_;
  wire _40135_;
  wire _40136_;
  wire _40137_;
  wire _40138_;
  wire _40139_;
  wire _40140_;
  wire _40141_;
  wire _40142_;
  wire _40143_;
  wire _40144_;
  wire _40145_;
  wire _40146_;
  wire _40147_;
  wire _40148_;
  wire _40149_;
  wire _40150_;
  wire _40151_;
  wire _40152_;
  wire _40153_;
  wire _40154_;
  wire _40155_;
  wire _40156_;
  wire _40157_;
  wire _40158_;
  wire _40159_;
  wire _40160_;
  wire _40161_;
  wire _40162_;
  wire _40163_;
  wire _40164_;
  wire _40165_;
  wire _40166_;
  wire _40167_;
  wire _40168_;
  wire _40169_;
  wire _40170_;
  wire _40171_;
  wire _40172_;
  wire _40173_;
  wire _40174_;
  wire _40175_;
  wire _40176_;
  wire _40177_;
  wire _40178_;
  wire _40179_;
  wire _40180_;
  wire _40181_;
  wire _40182_;
  wire _40183_;
  wire _40184_;
  wire _40185_;
  wire _40186_;
  wire _40187_;
  wire _40188_;
  wire _40189_;
  wire _40190_;
  wire _40191_;
  wire _40192_;
  wire _40193_;
  wire _40194_;
  wire _40195_;
  wire _40196_;
  wire _40197_;
  wire _40198_;
  wire _40199_;
  wire _40200_;
  wire _40201_;
  wire _40202_;
  wire _40203_;
  wire _40204_;
  wire _40205_;
  wire _40206_;
  wire _40207_;
  wire _40208_;
  wire _40209_;
  wire _40210_;
  wire _40211_;
  wire _40212_;
  wire _40213_;
  wire _40214_;
  wire _40215_;
  wire _40216_;
  wire _40217_;
  wire _40218_;
  wire _40219_;
  wire _40220_;
  wire _40221_;
  wire _40222_;
  wire _40223_;
  wire _40224_;
  wire _40225_;
  wire _40226_;
  wire _40227_;
  wire _40228_;
  wire _40229_;
  wire _40230_;
  wire _40231_;
  wire _40232_;
  wire _40233_;
  wire _40234_;
  wire _40235_;
  wire _40236_;
  wire _40237_;
  wire _40238_;
  wire _40239_;
  wire _40240_;
  wire _40241_;
  wire _40242_;
  wire _40243_;
  wire _40244_;
  wire _40245_;
  wire _40246_;
  wire _40247_;
  wire _40248_;
  wire _40249_;
  wire _40250_;
  wire _40251_;
  wire _40252_;
  wire _40253_;
  wire _40254_;
  wire _40255_;
  wire _40256_;
  wire _40257_;
  wire _40258_;
  wire _40259_;
  wire _40260_;
  wire _40261_;
  wire _40262_;
  wire _40263_;
  wire _40264_;
  wire _40265_;
  wire _40266_;
  wire _40267_;
  wire _40268_;
  wire _40269_;
  wire _40270_;
  wire _40271_;
  wire _40272_;
  wire _40273_;
  wire _40274_;
  wire _40275_;
  wire _40276_;
  wire _40277_;
  wire _40278_;
  wire _40279_;
  wire _40280_;
  wire _40281_;
  wire _40282_;
  wire _40283_;
  wire _40284_;
  wire _40285_;
  wire _40286_;
  wire _40287_;
  wire _40288_;
  wire _40289_;
  wire _40290_;
  wire _40291_;
  wire _40292_;
  wire _40293_;
  wire _40294_;
  wire _40295_;
  wire _40296_;
  wire _40297_;
  wire _40298_;
  wire _40299_;
  wire _40300_;
  wire _40301_;
  wire _40302_;
  wire _40303_;
  wire _40304_;
  wire _40305_;
  wire _40306_;
  wire _40307_;
  wire _40308_;
  wire _40309_;
  wire _40310_;
  wire _40311_;
  wire _40312_;
  wire _40313_;
  wire _40314_;
  wire _40315_;
  wire _40316_;
  wire _40317_;
  wire _40318_;
  wire _40319_;
  wire _40320_;
  wire _40321_;
  wire _40322_;
  wire _40323_;
  wire _40324_;
  wire _40325_;
  wire _40326_;
  wire _40327_;
  wire _40328_;
  wire _40329_;
  wire _40330_;
  wire _40331_;
  wire _40332_;
  wire _40333_;
  wire _40334_;
  wire _40335_;
  wire _40336_;
  wire _40337_;
  wire _40338_;
  wire _40339_;
  wire _40340_;
  wire _40341_;
  wire _40342_;
  wire _40343_;
  wire _40344_;
  wire _40345_;
  wire _40346_;
  wire _40347_;
  wire _40348_;
  wire _40349_;
  wire _40350_;
  wire _40351_;
  wire _40352_;
  wire _40353_;
  wire _40354_;
  wire _40355_;
  wire _40356_;
  wire _40357_;
  wire _40358_;
  wire _40359_;
  wire _40360_;
  wire _40361_;
  wire _40362_;
  wire _40363_;
  wire _40364_;
  wire _40365_;
  wire _40366_;
  wire _40367_;
  wire _40368_;
  wire _40369_;
  wire _40370_;
  wire _40371_;
  wire _40372_;
  wire _40373_;
  wire _40374_;
  wire _40375_;
  wire _40376_;
  wire _40377_;
  wire _40378_;
  wire _40379_;
  wire _40380_;
  wire _40381_;
  wire _40382_;
  wire _40383_;
  wire _40384_;
  wire _40385_;
  wire _40386_;
  wire _40387_;
  wire _40388_;
  wire _40389_;
  wire _40390_;
  wire _40391_;
  wire _40392_;
  wire _40393_;
  wire _40394_;
  wire _40395_;
  wire _40396_;
  wire _40397_;
  wire _40398_;
  wire _40399_;
  wire _40400_;
  wire _40401_;
  wire _40402_;
  wire _40403_;
  wire _40404_;
  wire _40405_;
  wire _40406_;
  wire _40407_;
  wire _40408_;
  wire _40409_;
  wire _40410_;
  wire _40411_;
  wire _40412_;
  wire _40413_;
  wire _40414_;
  wire _40415_;
  wire _40416_;
  wire _40417_;
  wire _40418_;
  wire _40419_;
  wire _40420_;
  wire _40421_;
  wire _40422_;
  wire _40423_;
  wire _40424_;
  wire _40425_;
  wire _40426_;
  wire _40427_;
  wire _40428_;
  wire _40429_;
  wire _40430_;
  wire _40431_;
  wire _40432_;
  wire _40433_;
  wire _40434_;
  wire _40435_;
  wire _40436_;
  wire _40437_;
  wire _40438_;
  wire _40439_;
  wire _40440_;
  wire _40441_;
  wire _40442_;
  wire _40443_;
  wire _40444_;
  wire _40445_;
  wire _40446_;
  wire _40447_;
  wire _40448_;
  wire _40449_;
  wire _40450_;
  wire _40451_;
  wire _40452_;
  wire _40453_;
  wire _40454_;
  wire _40455_;
  wire _40456_;
  wire _40457_;
  wire _40458_;
  wire _40459_;
  wire _40460_;
  wire _40461_;
  wire _40462_;
  wire _40463_;
  wire _40464_;
  wire _40465_;
  wire _40466_;
  wire _40467_;
  wire _40468_;
  wire _40469_;
  wire _40470_;
  wire _40471_;
  wire _40472_;
  wire _40473_;
  wire _40474_;
  wire _40475_;
  wire _40476_;
  wire _40477_;
  wire _40478_;
  wire _40479_;
  wire _40480_;
  wire _40481_;
  wire _40482_;
  wire _40483_;
  wire _40484_;
  wire _40485_;
  wire _40486_;
  wire _40487_;
  wire _40488_;
  wire _40489_;
  wire _40490_;
  wire _40491_;
  wire _40492_;
  wire _40493_;
  wire _40494_;
  wire _40495_;
  wire _40496_;
  wire _40497_;
  wire _40498_;
  wire _40499_;
  wire _40500_;
  wire _40501_;
  wire _40502_;
  wire _40503_;
  wire _40504_;
  wire _40505_;
  wire _40506_;
  wire _40507_;
  wire _40508_;
  wire _40509_;
  wire _40510_;
  wire _40511_;
  wire _40512_;
  wire _40513_;
  wire _40514_;
  wire _40515_;
  wire _40516_;
  wire _40517_;
  wire _40518_;
  wire _40519_;
  wire _40520_;
  wire _40521_;
  wire _40522_;
  wire _40523_;
  wire _40524_;
  wire _40525_;
  wire _40526_;
  wire _40527_;
  wire _40528_;
  wire _40529_;
  wire _40530_;
  wire _40531_;
  wire _40532_;
  wire _40533_;
  wire _40534_;
  wire _40535_;
  wire _40536_;
  wire _40537_;
  wire _40538_;
  wire _40539_;
  wire _40540_;
  wire _40541_;
  wire _40542_;
  wire _40543_;
  wire _40544_;
  wire _40545_;
  wire _40546_;
  wire _40547_;
  wire _40548_;
  wire _40549_;
  wire _40550_;
  wire _40551_;
  wire _40552_;
  wire _40553_;
  wire _40554_;
  wire _40555_;
  wire _40556_;
  wire _40557_;
  wire _40558_;
  wire _40559_;
  wire _40560_;
  wire _40561_;
  wire _40562_;
  wire _40563_;
  wire _40564_;
  wire _40565_;
  wire _40566_;
  wire _40567_;
  wire _40568_;
  wire _40569_;
  wire _40570_;
  wire _40571_;
  wire _40572_;
  wire _40573_;
  wire _40574_;
  wire _40575_;
  wire _40576_;
  wire _40577_;
  wire _40578_;
  wire _40579_;
  wire _40580_;
  wire _40581_;
  wire _40582_;
  wire _40583_;
  wire _40584_;
  wire _40585_;
  wire _40586_;
  wire _40587_;
  wire _40588_;
  wire _40589_;
  wire _40590_;
  wire _40591_;
  wire _40592_;
  wire _40593_;
  wire _40594_;
  wire _40595_;
  wire _40596_;
  wire _40597_;
  wire _40598_;
  wire _40599_;
  wire _40600_;
  wire _40601_;
  wire _40602_;
  wire _40603_;
  wire _40604_;
  wire _40605_;
  wire _40606_;
  wire _40607_;
  wire _40608_;
  wire _40609_;
  wire _40610_;
  wire _40611_;
  wire _40612_;
  wire _40613_;
  wire _40614_;
  wire _40615_;
  wire _40616_;
  wire _40617_;
  wire _40618_;
  wire _40619_;
  wire _40620_;
  wire _40621_;
  wire _40622_;
  wire _40623_;
  wire _40624_;
  wire _40625_;
  wire _40626_;
  wire _40627_;
  wire _40628_;
  wire _40629_;
  wire _40630_;
  wire _40631_;
  wire _40632_;
  wire _40633_;
  wire _40634_;
  wire _40635_;
  wire _40636_;
  wire _40637_;
  wire _40638_;
  wire _40639_;
  wire _40640_;
  wire _40641_;
  wire _40642_;
  wire _40643_;
  wire _40644_;
  wire _40645_;
  wire _40646_;
  wire _40647_;
  wire _40648_;
  wire _40649_;
  wire _40650_;
  wire _40651_;
  wire _40652_;
  wire _40653_;
  wire _40654_;
  wire _40655_;
  wire _40656_;
  wire _40657_;
  wire _40658_;
  wire _40659_;
  wire _40660_;
  wire _40661_;
  wire _40662_;
  wire _40663_;
  wire _40664_;
  wire _40665_;
  wire _40666_;
  wire _40667_;
  wire _40668_;
  wire _40669_;
  wire _40670_;
  wire _40671_;
  wire _40672_;
  wire _40673_;
  wire _40674_;
  wire _40675_;
  wire _40676_;
  wire _40677_;
  wire _40678_;
  wire _40679_;
  wire _40680_;
  wire _40681_;
  wire _40682_;
  wire _40683_;
  wire _40684_;
  wire _40685_;
  wire _40686_;
  wire _40687_;
  wire _40688_;
  wire _40689_;
  wire _40690_;
  wire _40691_;
  wire _40692_;
  wire _40693_;
  wire _40694_;
  wire _40695_;
  wire _40696_;
  wire _40697_;
  wire _40698_;
  wire _40699_;
  wire _40700_;
  wire _40701_;
  wire _40702_;
  wire _40703_;
  wire _40704_;
  wire _40705_;
  wire _40706_;
  wire _40707_;
  wire _40708_;
  wire _40709_;
  wire _40710_;
  wire _40711_;
  wire _40712_;
  wire _40713_;
  wire _40714_;
  wire _40715_;
  wire _40716_;
  wire _40717_;
  wire _40718_;
  wire _40719_;
  wire _40720_;
  wire _40721_;
  wire _40722_;
  wire _40723_;
  wire _40724_;
  wire _40725_;
  wire _40726_;
  wire _40727_;
  wire _40728_;
  wire _40729_;
  wire _40730_;
  wire _40731_;
  wire _40732_;
  wire _40733_;
  wire _40734_;
  wire _40735_;
  wire _40736_;
  wire _40737_;
  wire _40738_;
  wire _40739_;
  wire _40740_;
  wire _40741_;
  wire _40742_;
  wire _40743_;
  wire _40744_;
  wire _40745_;
  wire _40746_;
  wire _40747_;
  wire _40748_;
  wire _40749_;
  wire _40750_;
  wire _40751_;
  wire _40752_;
  wire _40753_;
  wire _40754_;
  wire _40755_;
  wire _40756_;
  wire _40757_;
  wire _40758_;
  wire _40759_;
  wire _40760_;
  wire _40761_;
  wire _40762_;
  wire _40763_;
  wire _40764_;
  wire _40765_;
  wire _40766_;
  wire _40767_;
  wire _40768_;
  wire _40769_;
  wire _40770_;
  wire _40771_;
  wire _40772_;
  wire _40773_;
  wire _40774_;
  wire _40775_;
  wire _40776_;
  wire _40777_;
  wire _40778_;
  wire _40779_;
  wire _40780_;
  wire _40781_;
  wire _40782_;
  wire _40783_;
  wire _40784_;
  wire _40785_;
  wire _40786_;
  wire _40787_;
  wire _40788_;
  wire _40789_;
  wire _40790_;
  wire _40791_;
  wire _40792_;
  wire _40793_;
  wire _40794_;
  wire _40795_;
  wire _40796_;
  wire _40797_;
  wire _40798_;
  wire _40799_;
  wire _40800_;
  wire _40801_;
  wire _40802_;
  wire _40803_;
  wire _40804_;
  wire _40805_;
  wire _40806_;
  wire _40807_;
  wire _40808_;
  wire _40809_;
  wire _40810_;
  wire _40811_;
  wire _40812_;
  wire _40813_;
  wire _40814_;
  wire _40815_;
  wire _40816_;
  wire _40817_;
  wire _40818_;
  wire _40819_;
  wire _40820_;
  wire _40821_;
  wire _40822_;
  wire _40823_;
  wire _40824_;
  wire _40825_;
  wire _40826_;
  wire _40827_;
  wire _40828_;
  wire _40829_;
  wire _40830_;
  wire _40831_;
  wire _40832_;
  wire _40833_;
  wire _40834_;
  wire _40835_;
  wire _40836_;
  wire _40837_;
  wire _40838_;
  wire _40839_;
  wire _40840_;
  wire _40841_;
  wire _40842_;
  wire _40843_;
  wire _40844_;
  wire _40845_;
  wire _40846_;
  wire _40847_;
  wire _40848_;
  wire _40849_;
  wire _40850_;
  wire _40851_;
  wire _40852_;
  wire _40853_;
  wire _40854_;
  wire _40855_;
  wire _40856_;
  wire _40857_;
  wire _40858_;
  wire _40859_;
  wire _40860_;
  wire _40861_;
  wire _40862_;
  wire _40863_;
  wire _40864_;
  wire _40865_;
  wire _40866_;
  wire _40867_;
  wire _40868_;
  wire _40869_;
  wire _40870_;
  wire _40871_;
  wire _40872_;
  wire _40873_;
  wire _40874_;
  wire _40875_;
  wire _40876_;
  wire _40877_;
  wire _40878_;
  wire _40879_;
  wire _40880_;
  wire _40881_;
  wire _40882_;
  wire _40883_;
  wire _40884_;
  wire _40885_;
  wire _40886_;
  wire _40887_;
  wire _40888_;
  wire _40889_;
  wire _40890_;
  wire _40891_;
  wire _40892_;
  wire _40893_;
  wire _40894_;
  wire _40895_;
  wire _40896_;
  wire _40897_;
  wire _40898_;
  wire _40899_;
  wire _40900_;
  wire _40901_;
  wire _40902_;
  wire _40903_;
  wire _40904_;
  wire _40905_;
  wire _40906_;
  wire _40907_;
  wire _40908_;
  wire _40909_;
  wire _40910_;
  wire _40911_;
  wire _40912_;
  wire _40913_;
  wire _40914_;
  wire _40915_;
  wire _40916_;
  wire _40917_;
  wire _40918_;
  wire _40919_;
  wire _40920_;
  wire _40921_;
  wire _40922_;
  wire _40923_;
  wire _40924_;
  wire _40925_;
  wire _40926_;
  wire _40927_;
  wire _40928_;
  wire _40929_;
  wire _40930_;
  wire _40931_;
  wire _40932_;
  wire _40933_;
  wire _40934_;
  wire _40935_;
  wire _40936_;
  wire _40937_;
  wire _40938_;
  wire _40939_;
  wire _40940_;
  wire _40941_;
  wire _40942_;
  wire _40943_;
  wire _40944_;
  wire _40945_;
  wire _40946_;
  wire _40947_;
  wire _40948_;
  wire _40949_;
  wire _40950_;
  wire _40951_;
  wire _40952_;
  wire _40953_;
  wire _40954_;
  wire _40955_;
  wire _40956_;
  wire _40957_;
  wire _40958_;
  wire _40959_;
  wire _40960_;
  wire _40961_;
  wire _40962_;
  wire _40963_;
  wire _40964_;
  wire _40965_;
  wire _40966_;
  wire _40967_;
  wire _40968_;
  wire _40969_;
  wire _40970_;
  wire _40971_;
  wire _40972_;
  wire _40973_;
  wire _40974_;
  wire _40975_;
  wire _40976_;
  wire _40977_;
  wire _40978_;
  wire _40979_;
  wire _40980_;
  wire _40981_;
  wire _40982_;
  wire _40983_;
  wire _40984_;
  wire _40985_;
  wire _40986_;
  wire _40987_;
  wire _40988_;
  wire _40989_;
  wire _40990_;
  wire _40991_;
  wire _40992_;
  wire _40993_;
  wire _40994_;
  wire _40995_;
  wire _40996_;
  wire _40997_;
  wire _40998_;
  wire _40999_;
  wire _41000_;
  wire _41001_;
  wire _41002_;
  wire _41003_;
  wire _41004_;
  wire _41005_;
  wire _41006_;
  wire _41007_;
  wire _41008_;
  wire _41009_;
  wire _41010_;
  wire _41011_;
  wire _41012_;
  wire _41013_;
  wire _41014_;
  wire _41015_;
  wire _41016_;
  wire _41017_;
  wire _41018_;
  wire _41019_;
  wire _41020_;
  wire _41021_;
  wire _41022_;
  wire _41023_;
  wire _41024_;
  wire _41025_;
  wire _41026_;
  wire _41027_;
  wire _41028_;
  wire _41029_;
  wire _41030_;
  wire _41031_;
  wire _41032_;
  wire _41033_;
  wire _41034_;
  wire _41035_;
  wire _41036_;
  wire _41037_;
  wire _41038_;
  wire _41039_;
  wire _41040_;
  wire _41041_;
  wire _41042_;
  wire _41043_;
  wire _41044_;
  wire _41045_;
  wire _41046_;
  wire _41047_;
  wire _41048_;
  wire _41049_;
  wire _41050_;
  wire _41051_;
  wire _41052_;
  wire _41053_;
  wire _41054_;
  wire _41055_;
  wire _41056_;
  wire _41057_;
  wire _41058_;
  wire _41059_;
  wire _41060_;
  wire _41061_;
  wire _41062_;
  wire _41063_;
  wire _41064_;
  wire _41065_;
  wire _41066_;
  wire _41067_;
  wire _41068_;
  wire _41069_;
  wire _41070_;
  wire _41071_;
  wire _41072_;
  wire _41073_;
  wire _41074_;
  wire _41075_;
  wire _41076_;
  wire _41077_;
  wire _41078_;
  wire _41079_;
  wire _41080_;
  wire _41081_;
  wire _41082_;
  wire _41083_;
  wire _41084_;
  wire _41085_;
  wire _41086_;
  wire _41087_;
  wire _41088_;
  wire _41089_;
  wire _41090_;
  wire _41091_;
  wire _41092_;
  wire _41093_;
  wire _41094_;
  wire _41095_;
  wire _41096_;
  wire _41097_;
  wire _41098_;
  wire _41099_;
  wire _41100_;
  wire _41101_;
  wire _41102_;
  wire _41103_;
  wire _41104_;
  wire _41105_;
  wire _41106_;
  wire _41107_;
  wire _41108_;
  wire _41109_;
  wire _41110_;
  wire _41111_;
  wire _41112_;
  wire _41113_;
  wire _41114_;
  wire _41115_;
  wire _41116_;
  wire _41117_;
  wire _41118_;
  wire _41119_;
  wire _41120_;
  wire _41121_;
  wire _41122_;
  wire _41123_;
  wire _41124_;
  wire _41125_;
  wire _41126_;
  wire _41127_;
  wire _41128_;
  wire _41129_;
  wire _41130_;
  wire _41131_;
  wire _41132_;
  wire _41133_;
  wire _41134_;
  wire _41135_;
  wire _41136_;
  wire _41137_;
  wire _41138_;
  wire _41139_;
  wire _41140_;
  wire _41141_;
  wire _41142_;
  wire _41143_;
  wire _41144_;
  wire _41145_;
  wire _41146_;
  wire _41147_;
  wire _41148_;
  wire _41149_;
  wire _41150_;
  wire _41151_;
  wire _41152_;
  wire _41153_;
  wire _41154_;
  wire _41155_;
  wire _41156_;
  wire _41157_;
  wire _41158_;
  wire _41159_;
  wire _41160_;
  wire _41161_;
  wire _41162_;
  wire _41163_;
  wire _41164_;
  wire _41165_;
  wire _41166_;
  wire _41167_;
  wire _41168_;
  wire _41169_;
  wire _41170_;
  wire _41171_;
  wire _41172_;
  wire _41173_;
  wire _41174_;
  wire _41175_;
  wire _41176_;
  wire _41177_;
  wire _41178_;
  wire _41179_;
  wire _41180_;
  wire _41181_;
  wire _41182_;
  wire _41183_;
  wire _41184_;
  wire _41185_;
  wire _41186_;
  wire _41187_;
  wire _41188_;
  wire _41189_;
  wire _41190_;
  wire _41191_;
  wire _41192_;
  wire _41193_;
  wire _41194_;
  wire _41195_;
  wire _41196_;
  wire _41197_;
  wire _41198_;
  wire _41199_;
  wire _41200_;
  wire _41201_;
  wire _41202_;
  wire _41203_;
  wire _41204_;
  wire _41205_;
  wire _41206_;
  wire _41207_;
  wire _41208_;
  wire _41209_;
  wire _41210_;
  wire _41211_;
  wire _41212_;
  wire _41213_;
  wire _41214_;
  wire _41215_;
  wire _41216_;
  wire _41217_;
  wire _41218_;
  wire _41219_;
  wire _41220_;
  wire _41221_;
  wire _41222_;
  wire _41223_;
  wire _41224_;
  wire _41225_;
  wire _41226_;
  wire _41227_;
  wire _41228_;
  wire _41229_;
  wire _41230_;
  wire _41231_;
  wire _41232_;
  wire _41233_;
  wire _41234_;
  wire _41235_;
  wire _41236_;
  wire _41237_;
  wire _41238_;
  wire _41239_;
  wire _41240_;
  wire _41241_;
  wire _41242_;
  wire _41243_;
  wire _41244_;
  wire _41245_;
  wire _41246_;
  wire _41247_;
  wire _41248_;
  wire _41249_;
  wire _41250_;
  wire _41251_;
  wire _41252_;
  wire _41253_;
  wire _41254_;
  wire _41255_;
  wire _41256_;
  wire _41257_;
  wire _41258_;
  wire _41259_;
  wire _41260_;
  wire _41261_;
  wire _41262_;
  wire _41263_;
  wire _41264_;
  wire _41265_;
  wire _41266_;
  wire _41267_;
  wire _41268_;
  wire _41269_;
  wire _41270_;
  wire _41271_;
  wire _41272_;
  wire _41273_;
  wire _41274_;
  wire _41275_;
  wire _41276_;
  wire _41277_;
  wire _41278_;
  wire _41279_;
  wire _41280_;
  wire _41281_;
  wire _41282_;
  wire _41283_;
  wire _41284_;
  wire _41285_;
  wire _41286_;
  wire _41287_;
  wire _41288_;
  wire _41289_;
  wire _41290_;
  wire _41291_;
  wire _41292_;
  wire _41293_;
  wire _41294_;
  wire _41295_;
  wire _41296_;
  wire _41297_;
  wire _41298_;
  wire _41299_;
  wire _41300_;
  wire _41301_;
  wire _41302_;
  wire _41303_;
  wire _41304_;
  wire _41305_;
  wire _41306_;
  wire _41307_;
  wire _41308_;
  wire _41309_;
  wire _41310_;
  wire _41311_;
  wire _41312_;
  wire _41313_;
  wire _41314_;
  wire _41315_;
  wire _41316_;
  wire _41317_;
  wire _41318_;
  wire _41319_;
  wire _41320_;
  wire _41321_;
  wire _41322_;
  wire _41323_;
  wire _41324_;
  wire _41325_;
  wire _41326_;
  wire _41327_;
  wire _41328_;
  wire _41329_;
  wire _41330_;
  wire _41331_;
  wire _41332_;
  wire _41333_;
  wire _41334_;
  wire _41335_;
  wire _41336_;
  wire _41337_;
  wire _41338_;
  wire _41339_;
  wire _41340_;
  wire _41341_;
  wire _41342_;
  wire _41343_;
  wire _41344_;
  wire _41345_;
  wire _41346_;
  wire _41347_;
  wire _41348_;
  wire _41349_;
  wire _41350_;
  wire _41351_;
  wire _41352_;
  wire _41353_;
  wire _41354_;
  wire _41355_;
  wire _41356_;
  wire _41357_;
  wire _41358_;
  wire _41359_;
  wire _41360_;
  wire _41361_;
  wire _41362_;
  wire _41363_;
  wire _41364_;
  wire _41365_;
  wire _41366_;
  wire _41367_;
  wire _41368_;
  wire _41369_;
  wire _41370_;
  wire _41371_;
  wire _41372_;
  wire _41373_;
  wire _41374_;
  wire _41375_;
  wire _41376_;
  wire _41377_;
  wire _41378_;
  wire _41379_;
  wire _41380_;
  wire _41381_;
  wire _41382_;
  wire _41383_;
  wire _41384_;
  wire _41385_;
  wire _41386_;
  wire _41387_;
  wire _41388_;
  wire _41389_;
  wire _41390_;
  wire _41391_;
  wire _41392_;
  wire _41393_;
  wire _41394_;
  wire _41395_;
  wire _41396_;
  wire _41397_;
  wire _41398_;
  wire _41399_;
  wire _41400_;
  wire _41401_;
  wire _41402_;
  wire _41403_;
  wire _41404_;
  wire _41405_;
  wire _41406_;
  wire _41407_;
  wire _41408_;
  wire _41409_;
  wire _41410_;
  wire _41411_;
  wire _41412_;
  wire _41413_;
  wire _41414_;
  wire _41415_;
  wire _41416_;
  wire _41417_;
  wire _41418_;
  wire _41419_;
  wire _41420_;
  wire _41421_;
  wire _41422_;
  wire _41423_;
  wire _41424_;
  wire _41425_;
  wire _41426_;
  wire _41427_;
  wire _41428_;
  wire _41429_;
  wire _41430_;
  wire _41431_;
  wire _41432_;
  wire _41433_;
  wire _41434_;
  wire _41435_;
  wire _41436_;
  wire _41437_;
  wire _41438_;
  wire _41439_;
  wire _41440_;
  wire _41441_;
  wire _41442_;
  wire _41443_;
  wire _41444_;
  wire _41445_;
  wire _41446_;
  wire _41447_;
  wire _41448_;
  wire _41449_;
  wire _41450_;
  wire _41451_;
  wire _41452_;
  wire _41453_;
  wire _41454_;
  wire _41455_;
  wire _41456_;
  wire _41457_;
  wire _41458_;
  wire _41459_;
  wire _41460_;
  wire _41461_;
  wire _41462_;
  wire _41463_;
  wire _41464_;
  wire _41465_;
  wire _41466_;
  wire _41467_;
  wire _41468_;
  wire _41469_;
  wire _41470_;
  wire _41471_;
  wire _41472_;
  wire _41473_;
  wire _41474_;
  wire _41475_;
  wire _41476_;
  wire _41477_;
  wire _41478_;
  wire _41479_;
  wire _41480_;
  wire _41481_;
  wire _41482_;
  wire _41483_;
  wire _41484_;
  wire _41485_;
  wire _41486_;
  wire _41487_;
  wire _41488_;
  wire _41489_;
  wire _41490_;
  wire _41491_;
  wire _41492_;
  wire _41493_;
  wire _41494_;
  wire _41495_;
  wire _41496_;
  wire _41497_;
  wire _41498_;
  wire _41499_;
  wire _41500_;
  wire _41501_;
  wire _41502_;
  wire _41503_;
  wire _41504_;
  wire _41505_;
  wire _41506_;
  wire _41507_;
  wire _41508_;
  wire _41509_;
  wire _41510_;
  wire _41511_;
  wire _41512_;
  wire _41513_;
  wire _41514_;
  wire _41515_;
  wire _41516_;
  wire _41517_;
  wire _41518_;
  wire _41519_;
  wire _41520_;
  wire _41521_;
  wire _41522_;
  wire _41523_;
  wire _41524_;
  wire _41525_;
  wire _41526_;
  wire _41527_;
  wire _41528_;
  wire _41529_;
  wire _41530_;
  wire _41531_;
  wire _41532_;
  wire _41533_;
  wire _41534_;
  wire _41535_;
  wire _41536_;
  wire _41537_;
  wire _41538_;
  wire _41539_;
  wire _41540_;
  wire _41541_;
  wire _41542_;
  wire _41543_;
  wire _41544_;
  wire _41545_;
  wire _41546_;
  wire _41547_;
  wire _41548_;
  wire _41549_;
  wire _41550_;
  wire _41551_;
  wire _41552_;
  wire _41553_;
  wire _41554_;
  wire _41555_;
  wire _41556_;
  wire _41557_;
  wire _41558_;
  wire _41559_;
  wire _41560_;
  wire _41561_;
  wire _41562_;
  wire _41563_;
  wire _41564_;
  wire _41565_;
  wire _41566_;
  wire _41567_;
  wire _41568_;
  wire _41569_;
  wire _41570_;
  wire _41571_;
  wire _41572_;
  wire _41573_;
  wire _41574_;
  wire _41575_;
  wire _41576_;
  wire _41577_;
  wire _41578_;
  wire _41579_;
  wire _41580_;
  wire _41581_;
  wire _41582_;
  wire _41583_;
  wire _41584_;
  wire _41585_;
  wire _41586_;
  wire _41587_;
  wire _41588_;
  wire _41589_;
  wire _41590_;
  wire _41591_;
  wire _41592_;
  wire _41593_;
  wire _41594_;
  wire _41595_;
  wire _41596_;
  wire _41597_;
  wire _41598_;
  wire _41599_;
  wire _41600_;
  wire _41601_;
  wire _41602_;
  wire _41603_;
  wire _41604_;
  wire _41605_;
  wire _41606_;
  wire _41607_;
  wire _41608_;
  wire _41609_;
  wire _41610_;
  wire _41611_;
  wire _41612_;
  wire _41613_;
  wire _41614_;
  wire _41615_;
  wire _41616_;
  wire _41617_;
  wire _41618_;
  wire _41619_;
  wire _41620_;
  wire _41621_;
  wire _41622_;
  wire _41623_;
  wire _41624_;
  wire _41625_;
  wire _41626_;
  wire _41627_;
  wire _41628_;
  wire _41629_;
  wire _41630_;
  wire _41631_;
  wire _41632_;
  wire _41633_;
  wire _41634_;
  wire _41635_;
  wire _41636_;
  wire _41637_;
  wire _41638_;
  wire _41639_;
  wire _41640_;
  wire _41641_;
  wire _41642_;
  wire _41643_;
  wire _41644_;
  wire _41645_;
  wire _41646_;
  wire _41647_;
  wire _41648_;
  wire _41649_;
  wire _41650_;
  wire _41651_;
  wire _41652_;
  wire _41653_;
  wire _41654_;
  wire _41655_;
  wire _41656_;
  wire _41657_;
  wire _41658_;
  wire _41659_;
  wire _41660_;
  wire _41661_;
  wire _41662_;
  wire _41663_;
  wire _41664_;
  wire _41665_;
  wire _41666_;
  wire _41667_;
  wire _41668_;
  wire _41669_;
  wire _41670_;
  wire _41671_;
  wire _41672_;
  wire _41673_;
  wire _41674_;
  wire _41675_;
  wire _41676_;
  wire _41677_;
  wire _41678_;
  wire _41679_;
  wire _41680_;
  wire _41681_;
  wire _41682_;
  wire _41683_;
  wire _41684_;
  wire _41685_;
  wire _41686_;
  wire _41687_;
  wire _41688_;
  wire _41689_;
  wire _41690_;
  wire _41691_;
  wire _41692_;
  wire _41693_;
  wire _41694_;
  wire _41695_;
  wire _41696_;
  wire _41697_;
  wire _41698_;
  wire _41699_;
  wire _41700_;
  wire _41701_;
  wire _41702_;
  wire _41703_;
  wire _41704_;
  wire _41705_;
  wire _41706_;
  wire _41707_;
  wire _41708_;
  wire _41709_;
  wire _41710_;
  wire _41711_;
  wire _41712_;
  wire _41713_;
  wire _41714_;
  wire _41715_;
  wire _41716_;
  wire _41717_;
  wire _41718_;
  wire _41719_;
  wire _41720_;
  wire _41721_;
  wire _41722_;
  wire _41723_;
  wire _41724_;
  wire _41725_;
  wire _41726_;
  wire _41727_;
  wire _41728_;
  wire _41729_;
  wire _41730_;
  wire _41731_;
  wire _41732_;
  wire _41733_;
  wire _41734_;
  wire _41735_;
  wire _41736_;
  wire _41737_;
  wire _41738_;
  wire _41739_;
  wire _41740_;
  wire _41741_;
  wire _41742_;
  wire _41743_;
  wire _41744_;
  wire _41745_;
  wire _41746_;
  wire _41747_;
  wire _41748_;
  wire _41749_;
  wire _41750_;
  wire _41751_;
  wire _41752_;
  wire _41753_;
  wire _41754_;
  wire _41755_;
  wire _41756_;
  wire _41757_;
  wire _41758_;
  wire _41759_;
  wire _41760_;
  wire _41761_;
  wire _41762_;
  wire _41763_;
  wire _41764_;
  wire _41765_;
  wire _41766_;
  wire _41767_;
  wire _41768_;
  wire _41769_;
  wire _41770_;
  wire _41771_;
  wire _41772_;
  wire _41773_;
  wire _41774_;
  wire _41775_;
  wire _41776_;
  wire _41777_;
  wire _41778_;
  wire _41779_;
  wire _41780_;
  wire _41781_;
  wire _41782_;
  wire _41783_;
  wire _41784_;
  wire _41785_;
  wire _41786_;
  wire _41787_;
  wire _41788_;
  wire _41789_;
  wire _41790_;
  wire _41791_;
  wire _41792_;
  wire _41793_;
  wire _41794_;
  wire _41795_;
  wire _41796_;
  wire _41797_;
  wire _41798_;
  wire _41799_;
  wire _41800_;
  wire _41801_;
  wire _41802_;
  wire _41803_;
  wire _41804_;
  wire _41805_;
  wire _41806_;
  wire _41807_;
  wire _41808_;
  wire _41809_;
  wire _41810_;
  wire _41811_;
  wire _41812_;
  wire _41813_;
  wire _41814_;
  wire _41815_;
  wire _41816_;
  wire _41817_;
  wire _41818_;
  wire _41819_;
  wire _41820_;
  wire _41821_;
  wire _41822_;
  wire _41823_;
  wire _41824_;
  wire _41825_;
  wire _41826_;
  wire _41827_;
  wire _41828_;
  wire _41829_;
  wire _41830_;
  wire _41831_;
  wire _41832_;
  wire _41833_;
  wire _41834_;
  wire _41835_;
  wire _41836_;
  wire _41837_;
  wire _41838_;
  wire _41839_;
  wire _41840_;
  wire _41841_;
  wire _41842_;
  wire _41843_;
  wire _41844_;
  wire _41845_;
  wire _41846_;
  wire _41847_;
  wire _41848_;
  wire _41849_;
  wire _41850_;
  wire _41851_;
  wire _41852_;
  wire _41853_;
  wire _41854_;
  wire _41855_;
  wire _41856_;
  wire _41857_;
  wire _41858_;
  wire _41859_;
  wire _41860_;
  wire _41861_;
  wire _41862_;
  wire _41863_;
  wire _41864_;
  wire _41865_;
  wire _41866_;
  wire _41867_;
  wire _41868_;
  wire _41869_;
  wire _41870_;
  wire _41871_;
  wire _41872_;
  wire _41873_;
  wire _41874_;
  wire _41875_;
  wire _41876_;
  wire _41877_;
  wire _41878_;
  wire _41879_;
  wire _41880_;
  wire _41881_;
  wire _41882_;
  wire _41883_;
  wire _41884_;
  wire _41885_;
  wire _41886_;
  wire _41887_;
  wire _41888_;
  wire _41889_;
  wire _41890_;
  wire _41891_;
  wire _41892_;
  wire _41893_;
  wire _41894_;
  wire _41895_;
  wire _41896_;
  wire _41897_;
  wire _41898_;
  wire _41899_;
  wire _41900_;
  wire _41901_;
  wire _41902_;
  wire _41903_;
  wire _41904_;
  wire _41905_;
  wire _41906_;
  wire _41907_;
  wire _41908_;
  wire _41909_;
  wire _41910_;
  wire _41911_;
  wire _41912_;
  wire _41913_;
  wire _41914_;
  wire _41915_;
  wire _41916_;
  wire _41917_;
  wire _41918_;
  wire _41919_;
  wire _41920_;
  wire _41921_;
  wire _41922_;
  wire _41923_;
  wire _41924_;
  wire _41925_;
  wire _41926_;
  wire _41927_;
  wire _41928_;
  wire _41929_;
  wire _41930_;
  wire _41931_;
  wire _41932_;
  wire _41933_;
  wire _41934_;
  wire _41935_;
  wire _41936_;
  wire _41937_;
  wire _41938_;
  wire _41939_;
  wire _41940_;
  wire _41941_;
  wire _41942_;
  wire _41943_;
  wire _41944_;
  wire _41945_;
  wire _41946_;
  wire _41947_;
  wire _41948_;
  wire _41949_;
  wire _41950_;
  wire _41951_;
  wire _41952_;
  wire _41953_;
  wire _41954_;
  wire _41955_;
  wire _41956_;
  wire _41957_;
  wire _41958_;
  wire _41959_;
  wire _41960_;
  wire _41961_;
  wire _41962_;
  wire _41963_;
  wire _41964_;
  wire _41965_;
  wire _41966_;
  wire _41967_;
  wire _41968_;
  wire _41969_;
  wire _41970_;
  wire _41971_;
  wire _41972_;
  wire _41973_;
  wire _41974_;
  wire _41975_;
  wire _41976_;
  wire _41977_;
  wire _41978_;
  wire _41979_;
  wire _41980_;
  wire _41981_;
  wire _41982_;
  wire _41983_;
  wire _41984_;
  wire _41985_;
  wire _41986_;
  wire _41987_;
  wire _41988_;
  wire _41989_;
  wire _41990_;
  wire _41991_;
  wire _41992_;
  wire _41993_;
  wire _41994_;
  wire _41995_;
  wire _41996_;
  wire _41997_;
  wire _41998_;
  wire _41999_;
  wire _42000_;
  wire _42001_;
  wire _42002_;
  wire _42003_;
  wire _42004_;
  wire _42005_;
  wire _42006_;
  wire _42007_;
  wire _42008_;
  wire _42009_;
  wire _42010_;
  wire _42011_;
  wire _42012_;
  wire _42013_;
  wire _42014_;
  wire _42015_;
  wire _42016_;
  wire _42017_;
  wire _42018_;
  wire _42019_;
  wire _42020_;
  wire _42021_;
  wire _42022_;
  wire _42023_;
  wire _42024_;
  wire _42025_;
  wire _42026_;
  wire _42027_;
  wire _42028_;
  wire _42029_;
  wire _42030_;
  wire _42031_;
  wire _42032_;
  wire _42033_;
  wire _42034_;
  wire _42035_;
  wire _42036_;
  wire _42037_;
  wire _42038_;
  wire _42039_;
  wire _42040_;
  wire _42041_;
  wire _42042_;
  wire _42043_;
  wire _42044_;
  wire _42045_;
  wire _42046_;
  wire _42047_;
  wire _42048_;
  wire _42049_;
  wire _42050_;
  wire _42051_;
  wire _42052_;
  wire _42053_;
  wire _42054_;
  wire _42055_;
  wire _42056_;
  wire _42057_;
  wire _42058_;
  wire _42059_;
  wire _42060_;
  wire _42061_;
  wire _42062_;
  wire _42063_;
  wire _42064_;
  wire _42065_;
  wire _42066_;
  wire _42067_;
  wire _42068_;
  wire _42069_;
  wire _42070_;
  wire _42071_;
  wire _42072_;
  wire _42073_;
  wire _42074_;
  wire _42075_;
  wire _42076_;
  wire _42077_;
  wire _42078_;
  wire _42079_;
  wire _42080_;
  wire _42081_;
  wire _42082_;
  wire _42083_;
  wire _42084_;
  wire _42085_;
  wire _42086_;
  wire _42087_;
  wire _42088_;
  wire _42089_;
  wire _42090_;
  wire _42091_;
  wire _42092_;
  wire _42093_;
  wire _42094_;
  wire _42095_;
  wire _42096_;
  wire _42097_;
  wire _42098_;
  wire _42099_;
  wire _42100_;
  wire _42101_;
  wire _42102_;
  wire _42103_;
  wire _42104_;
  wire _42105_;
  wire _42106_;
  wire _42107_;
  wire _42108_;
  wire _42109_;
  wire _42110_;
  wire _42111_;
  wire _42112_;
  wire _42113_;
  wire _42114_;
  wire _42115_;
  wire _42116_;
  wire _42117_;
  wire _42118_;
  wire _42119_;
  wire _42120_;
  wire _42121_;
  wire _42122_;
  wire _42123_;
  wire _42124_;
  wire _42125_;
  wire _42126_;
  wire _42127_;
  wire _42128_;
  wire _42129_;
  wire _42130_;
  wire _42131_;
  wire _42132_;
  wire _42133_;
  wire _42134_;
  wire _42135_;
  wire _42136_;
  wire _42137_;
  wire _42138_;
  wire _42139_;
  wire _42140_;
  wire _42141_;
  wire _42142_;
  wire _42143_;
  wire _42144_;
  wire _42145_;
  wire _42146_;
  wire _42147_;
  wire _42148_;
  wire _42149_;
  wire _42150_;
  wire _42151_;
  wire _42152_;
  wire _42153_;
  wire _42154_;
  wire _42155_;
  wire _42156_;
  wire _42157_;
  wire _42158_;
  wire _42159_;
  wire _42160_;
  wire _42161_;
  wire _42162_;
  wire _42163_;
  wire _42164_;
  wire _42165_;
  wire _42166_;
  wire _42167_;
  wire _42168_;
  wire _42169_;
  wire _42170_;
  wire _42171_;
  wire _42172_;
  wire _42173_;
  wire _42174_;
  wire _42175_;
  wire _42176_;
  wire _42177_;
  wire _42178_;
  wire _42179_;
  wire _42180_;
  wire _42181_;
  wire _42182_;
  wire _42183_;
  wire _42184_;
  wire _42185_;
  wire _42186_;
  wire _42187_;
  wire _42188_;
  wire _42189_;
  wire _42190_;
  wire _42191_;
  wire _42192_;
  wire _42193_;
  wire _42194_;
  wire _42195_;
  wire _42196_;
  wire _42197_;
  wire _42198_;
  wire _42199_;
  wire _42200_;
  wire _42201_;
  wire _42202_;
  wire _42203_;
  wire _42204_;
  wire _42205_;
  wire _42206_;
  wire _42207_;
  wire _42208_;
  wire _42209_;
  wire _42210_;
  wire _42211_;
  wire _42212_;
  wire _42213_;
  wire _42214_;
  wire _42215_;
  wire _42216_;
  wire _42217_;
  wire _42218_;
  wire _42219_;
  wire _42220_;
  wire _42221_;
  wire _42222_;
  wire _42223_;
  wire _42224_;
  wire _42225_;
  wire _42226_;
  wire _42227_;
  wire _42228_;
  wire _42229_;
  wire _42230_;
  wire _42231_;
  wire _42232_;
  wire _42233_;
  wire _42234_;
  wire _42235_;
  wire _42236_;
  wire _42237_;
  wire _42238_;
  wire _42239_;
  wire _42240_;
  wire _42241_;
  wire _42242_;
  wire _42243_;
  wire _42244_;
  wire _42245_;
  wire _42246_;
  wire _42247_;
  wire _42248_;
  wire _42249_;
  wire _42250_;
  wire _42251_;
  wire _42252_;
  wire _42253_;
  wire _42254_;
  wire _42255_;
  wire _42256_;
  wire _42257_;
  wire _42258_;
  wire _42259_;
  wire _42260_;
  wire _42261_;
  wire _42262_;
  wire _42263_;
  wire _42264_;
  wire _42265_;
  wire _42266_;
  wire _42267_;
  wire _42268_;
  wire _42269_;
  wire _42270_;
  wire _42271_;
  wire _42272_;
  wire _42273_;
  wire _42274_;
  wire _42275_;
  wire _42276_;
  wire _42277_;
  wire _42278_;
  wire _42279_;
  wire _42280_;
  wire _42281_;
  wire _42282_;
  wire _42283_;
  wire _42284_;
  wire _42285_;
  wire _42286_;
  wire _42287_;
  wire _42288_;
  wire _42289_;
  wire _42290_;
  wire _42291_;
  wire _42292_;
  wire _42293_;
  wire _42294_;
  wire _42295_;
  wire _42296_;
  wire _42297_;
  wire _42298_;
  wire _42299_;
  wire _42300_;
  wire _42301_;
  wire _42302_;
  wire _42303_;
  wire _42304_;
  wire _42305_;
  wire _42306_;
  wire _42307_;
  wire _42308_;
  wire _42309_;
  wire _42310_;
  wire _42311_;
  wire _42312_;
  wire _42313_;
  wire _42314_;
  wire _42315_;
  wire _42316_;
  wire _42317_;
  wire _42318_;
  wire _42319_;
  wire _42320_;
  wire _42321_;
  wire _42322_;
  wire _42323_;
  wire _42324_;
  wire _42325_;
  wire _42326_;
  wire _42327_;
  wire _42328_;
  wire _42329_;
  wire _42330_;
  wire _42331_;
  wire _42332_;
  wire _42333_;
  wire _42334_;
  wire _42335_;
  wire _42336_;
  wire _42337_;
  wire _42338_;
  wire _42339_;
  wire _42340_;
  wire _42341_;
  wire _42342_;
  wire _42343_;
  wire _42344_;
  wire _42345_;
  wire _42346_;
  wire _42347_;
  wire _42348_;
  wire _42349_;
  wire _42350_;
  wire _42351_;
  wire _42352_;
  wire _42353_;
  wire _42354_;
  wire _42355_;
  wire _42356_;
  wire _42357_;
  wire _42358_;
  wire _42359_;
  wire _42360_;
  wire _42361_;
  wire _42362_;
  wire _42363_;
  wire _42364_;
  wire _42365_;
  wire _42366_;
  wire _42367_;
  wire _42368_;
  wire _42369_;
  wire _42370_;
  wire _42371_;
  wire _42372_;
  wire _42373_;
  wire _42374_;
  wire _42375_;
  wire _42376_;
  wire _42377_;
  wire _42378_;
  wire _42379_;
  wire _42380_;
  wire _42381_;
  wire _42382_;
  wire _42383_;
  wire _42384_;
  wire _42385_;
  wire _42386_;
  wire _42387_;
  wire _42388_;
  wire _42389_;
  wire _42390_;
  wire _42391_;
  wire _42392_;
  wire _42393_;
  wire _42394_;
  wire _42395_;
  wire _42396_;
  wire _42397_;
  wire _42398_;
  wire _42399_;
  wire _42400_;
  wire _42401_;
  wire _42402_;
  wire _42403_;
  wire _42404_;
  wire _42405_;
  wire _42406_;
  wire _42407_;
  wire _42408_;
  wire _42409_;
  wire _42410_;
  wire _42411_;
  wire _42412_;
  wire _42413_;
  wire _42414_;
  wire _42415_;
  wire _42416_;
  wire _42417_;
  wire _42418_;
  wire _42419_;
  wire _42420_;
  wire _42421_;
  wire _42422_;
  wire _42423_;
  wire _42424_;
  wire _42425_;
  wire _42426_;
  wire _42427_;
  wire _42428_;
  wire _42429_;
  wire _42430_;
  wire _42431_;
  wire _42432_;
  wire _42433_;
  wire _42434_;
  wire _42435_;
  wire _42436_;
  wire _42437_;
  wire _42438_;
  wire _42439_;
  wire _42440_;
  wire _42441_;
  wire _42442_;
  wire _42443_;
  wire _42444_;
  wire _42445_;
  wire _42446_;
  wire _42447_;
  wire _42448_;
  wire _42449_;
  wire _42450_;
  wire _42451_;
  wire _42452_;
  wire _42453_;
  wire _42454_;
  wire _42455_;
  wire _42456_;
  wire _42457_;
  wire _42458_;
  wire _42459_;
  wire _42460_;
  wire _42461_;
  wire _42462_;
  wire _42463_;
  wire _42464_;
  wire _42465_;
  wire _42466_;
  wire _42467_;
  wire _42468_;
  wire _42469_;
  wire _42470_;
  wire _42471_;
  wire _42472_;
  wire _42473_;
  wire _42474_;
  wire _42475_;
  wire _42476_;
  wire _42477_;
  wire _42478_;
  wire _42479_;
  wire _42480_;
  wire _42481_;
  wire _42482_;
  wire _42483_;
  wire _42484_;
  wire _42485_;
  wire _42486_;
  wire _42487_;
  wire _42488_;
  wire _42489_;
  wire _42490_;
  wire _42491_;
  wire _42492_;
  wire _42493_;
  wire _42494_;
  wire _42495_;
  wire _42496_;
  wire _42497_;
  wire _42498_;
  wire _42499_;
  wire _42500_;
  wire _42501_;
  wire _42502_;
  wire _42503_;
  wire _42504_;
  wire _42505_;
  wire _42506_;
  wire _42507_;
  wire _42508_;
  wire _42509_;
  wire _42510_;
  wire _42511_;
  wire _42512_;
  wire _42513_;
  wire _42514_;
  wire _42515_;
  wire _42516_;
  wire _42517_;
  wire _42518_;
  wire _42519_;
  wire _42520_;
  wire _42521_;
  wire _42522_;
  wire _42523_;
  wire _42524_;
  wire _42525_;
  wire _42526_;
  wire _42527_;
  wire _42528_;
  wire _42529_;
  wire _42530_;
  wire _42531_;
  wire _42532_;
  wire _42533_;
  wire _42534_;
  wire _42535_;
  wire _42536_;
  wire _42537_;
  wire _42538_;
  wire _42539_;
  wire _42540_;
  wire _42541_;
  wire _42542_;
  wire _42543_;
  wire _42544_;
  wire _42545_;
  wire _42546_;
  wire _42547_;
  wire _42548_;
  wire _42549_;
  wire _42550_;
  wire _42551_;
  wire _42552_;
  wire _42553_;
  wire _42554_;
  wire _42555_;
  wire _42556_;
  wire _42557_;
  wire _42558_;
  wire _42559_;
  wire _42560_;
  wire _42561_;
  wire _42562_;
  wire _42563_;
  wire _42564_;
  wire _42565_;
  wire _42566_;
  wire _42567_;
  wire _42568_;
  wire _42569_;
  wire _42570_;
  wire _42571_;
  wire _42572_;
  wire _42573_;
  wire _42574_;
  wire _42575_;
  wire _42576_;
  wire _42577_;
  wire _42578_;
  wire _42579_;
  wire _42580_;
  wire _42581_;
  wire _42582_;
  wire _42583_;
  wire _42584_;
  wire _42585_;
  wire _42586_;
  wire _42587_;
  wire _42588_;
  wire _42589_;
  wire _42590_;
  wire _42591_;
  wire _42592_;
  wire _42593_;
  wire _42594_;
  wire _42595_;
  wire _42596_;
  wire _42597_;
  wire _42598_;
  wire _42599_;
  wire _42600_;
  wire _42601_;
  wire _42602_;
  wire _42603_;
  wire _42604_;
  wire _42605_;
  wire _42606_;
  wire _42607_;
  wire _42608_;
  wire _42609_;
  wire _42610_;
  wire _42611_;
  wire _42612_;
  wire _42613_;
  wire _42614_;
  wire _42615_;
  wire _42616_;
  wire _42617_;
  wire _42618_;
  wire _42619_;
  wire _42620_;
  wire _42621_;
  wire _42622_;
  wire _42623_;
  wire _42624_;
  wire _42625_;
  wire _42626_;
  wire _42627_;
  wire _42628_;
  wire _42629_;
  wire _42630_;
  wire _42631_;
  wire _42632_;
  wire _42633_;
  wire _42634_;
  wire _42635_;
  wire _42636_;
  wire _42637_;
  wire _42638_;
  wire _42639_;
  wire _42640_;
  wire _42641_;
  wire _42642_;
  wire _42643_;
  wire _42644_;
  wire _42645_;
  wire _42646_;
  wire _42647_;
  wire _42648_;
  wire _42649_;
  wire _42650_;
  wire _42651_;
  wire _42652_;
  wire _42653_;
  wire _42654_;
  wire _42655_;
  wire _42656_;
  wire _42657_;
  wire _42658_;
  wire _42659_;
  wire _42660_;
  wire _42661_;
  wire _42662_;
  wire _42663_;
  wire _42664_;
  wire _42665_;
  wire _42666_;
  wire _42667_;
  wire _42668_;
  wire _42669_;
  wire _42670_;
  wire _42671_;
  wire _42672_;
  wire _42673_;
  wire _42674_;
  wire _42675_;
  wire _42676_;
  wire _42677_;
  wire _42678_;
  wire _42679_;
  wire _42680_;
  wire _42681_;
  wire _42682_;
  wire _42683_;
  wire _42684_;
  wire _42685_;
  wire _42686_;
  wire _42687_;
  wire _42688_;
  wire _42689_;
  wire _42690_;
  wire _42691_;
  wire _42692_;
  wire _42693_;
  wire _42694_;
  wire _42695_;
  wire _42696_;
  wire _42697_;
  wire _42698_;
  wire _42699_;
  wire _42700_;
  wire _42701_;
  wire _42702_;
  wire _42703_;
  wire _42704_;
  wire _42705_;
  wire _42706_;
  wire _42707_;
  wire _42708_;
  wire _42709_;
  wire _42710_;
  wire _42711_;
  wire _42712_;
  wire _42713_;
  wire _42714_;
  wire _42715_;
  wire _42716_;
  wire _42717_;
  wire _42718_;
  wire _42719_;
  wire _42720_;
  wire _42721_;
  wire _42722_;
  wire _42723_;
  wire _42724_;
  wire _42725_;
  wire _42726_;
  wire _42727_;
  wire _42728_;
  wire _42729_;
  wire _42730_;
  wire _42731_;
  wire _42732_;
  wire _42733_;
  wire _42734_;
  wire _42735_;
  wire _42736_;
  wire _42737_;
  wire _42738_;
  wire _42739_;
  wire _42740_;
  wire _42741_;
  wire _42742_;
  wire _42743_;
  wire _42744_;
  wire _42745_;
  wire _42746_;
  wire _42747_;
  wire _42748_;
  wire _42749_;
  wire _42750_;
  wire _42751_;
  wire _42752_;
  wire _42753_;
  wire _42754_;
  wire _42755_;
  wire _42756_;
  wire _42757_;
  wire _42758_;
  wire _42759_;
  wire _42760_;
  wire _42761_;
  wire _42762_;
  wire _42763_;
  wire _42764_;
  wire _42765_;
  wire _42766_;
  wire _42767_;
  wire _42768_;
  wire _42769_;
  wire _42770_;
  wire _42771_;
  wire _42772_;
  wire _42773_;
  wire _42774_;
  wire _42775_;
  wire _42776_;
  wire _42777_;
  wire _42778_;
  wire _42779_;
  wire _42780_;
  wire _42781_;
  wire _42782_;
  wire _42783_;
  wire _42784_;
  wire _42785_;
  wire _42786_;
  wire _42787_;
  wire _42788_;
  wire _42789_;
  wire _42790_;
  wire _42791_;
  wire _42792_;
  wire _42793_;
  wire _42794_;
  wire _42795_;
  wire _42796_;
  wire _42797_;
  wire _42798_;
  wire _42799_;
  wire _42800_;
  wire _42801_;
  wire _42802_;
  wire _42803_;
  wire _42804_;
  wire _42805_;
  wire _42806_;
  wire _42807_;
  wire _42808_;
  wire _42809_;
  wire _42810_;
  wire _42811_;
  wire _42812_;
  wire _42813_;
  wire _42814_;
  wire _42815_;
  wire _42816_;
  wire _42817_;
  wire _42818_;
  wire _42819_;
  wire _42820_;
  wire _42821_;
  wire _42822_;
  wire _42823_;
  wire _42824_;
  wire _42825_;
  wire _42826_;
  wire _42827_;
  wire _42828_;
  wire _42829_;
  wire _42830_;
  wire _42831_;
  wire _42832_;
  wire _42833_;
  wire _42834_;
  wire _42835_;
  wire _42836_;
  wire _42837_;
  wire _42838_;
  wire _42839_;
  wire _42840_;
  wire _42841_;
  wire _42842_;
  wire _42843_;
  wire _42844_;
  wire _42845_;
  wire _42846_;
  wire _42847_;
  wire _42848_;
  wire _42849_;
  wire _42850_;
  wire _42851_;
  wire _42852_;
  wire _42853_;
  wire _42854_;
  wire _42855_;
  wire _42856_;
  wire _42857_;
  wire _42858_;
  wire _42859_;
  wire _42860_;
  wire _42861_;
  wire _42862_;
  wire _42863_;
  wire _42864_;
  wire _42865_;
  wire _42866_;
  wire _42867_;
  wire _42868_;
  wire _42869_;
  wire _42870_;
  wire _42871_;
  wire _42872_;
  wire _42873_;
  wire _42874_;
  wire _42875_;
  wire _42876_;
  wire _42877_;
  wire _42878_;
  wire _42879_;
  wire _42880_;
  wire _42881_;
  wire _42882_;
  wire _42883_;
  wire _42884_;
  wire _42885_;
  wire _42886_;
  wire _42887_;
  wire _42888_;
  wire _42889_;
  wire _42890_;
  wire _42891_;
  wire _42892_;
  wire _42893_;
  wire _42894_;
  wire _42895_;
  wire _42896_;
  wire _42897_;
  wire _42898_;
  wire _42899_;
  wire _42900_;
  wire _42901_;
  wire _42902_;
  wire _42903_;
  wire _42904_;
  wire _42905_;
  wire _42906_;
  wire _42907_;
  wire _42908_;
  wire _42909_;
  wire _42910_;
  wire _42911_;
  wire _42912_;
  wire _42913_;
  wire _42914_;
  wire _42915_;
  wire _42916_;
  wire _42917_;
  wire _42918_;
  wire _42919_;
  wire _42920_;
  wire _42921_;
  wire _42922_;
  wire _42923_;
  wire _42924_;
  wire _42925_;
  wire _42926_;
  wire _42927_;
  wire _42928_;
  wire _42929_;
  wire _42930_;
  wire _42931_;
  wire _42932_;
  wire _42933_;
  wire _42934_;
  wire _42935_;
  wire _42936_;
  wire _42937_;
  wire _42938_;
  wire _42939_;
  wire _42940_;
  wire _42941_;
  wire _42942_;
  wire _42943_;
  wire _42944_;
  wire _42945_;
  wire _42946_;
  wire _42947_;
  wire _42948_;
  wire _42949_;
  wire _42950_;
  wire _42951_;
  wire _42952_;
  wire _42953_;
  wire _42954_;
  wire _42955_;
  wire _42956_;
  wire _42957_;
  wire _42958_;
  wire _42959_;
  wire _42960_;
  wire _42961_;
  wire _42962_;
  wire _42963_;
  wire _42964_;
  wire _42965_;
  wire _42966_;
  wire _42967_;
  wire _42968_;
  wire _42969_;
  wire _42970_;
  wire _42971_;
  wire _42972_;
  wire _42973_;
  wire _42974_;
  wire _42975_;
  wire _42976_;
  wire _42977_;
  wire _42978_;
  wire _42979_;
  wire _42980_;
  wire _42981_;
  wire _42982_;
  wire _42983_;
  wire _42984_;
  wire _42985_;
  wire _42986_;
  wire _42987_;
  wire _42988_;
  wire _42989_;
  wire _42990_;
  wire _42991_;
  wire _42992_;
  wire _42993_;
  wire _42994_;
  wire _42995_;
  wire _42996_;
  wire _42997_;
  wire _42998_;
  wire _42999_;
  wire _43000_;
  wire _43001_;
  wire _43002_;
  wire _43003_;
  wire _43004_;
  wire _43005_;
  wire _43006_;
  wire _43007_;
  wire _43008_;
  wire _43009_;
  wire _43010_;
  wire _43011_;
  wire _43012_;
  wire _43013_;
  wire _43014_;
  wire _43015_;
  wire _43016_;
  wire _43017_;
  wire _43018_;
  wire _43019_;
  wire _43020_;
  wire _43021_;
  wire _43022_;
  wire _43023_;
  wire _43024_;
  wire _43025_;
  wire _43026_;
  wire _43027_;
  wire _43028_;
  wire _43029_;
  wire _43030_;
  wire _43031_;
  wire _43032_;
  wire _43033_;
  wire _43034_;
  wire _43035_;
  wire _43036_;
  wire _43037_;
  wire _43038_;
  wire _43039_;
  wire _43040_;
  wire _43041_;
  wire _43042_;
  wire _43043_;
  wire _43044_;
  wire _43045_;
  wire _43046_;
  wire _43047_;
  wire _43048_;
  wire _43049_;
  wire _43050_;
  wire _43051_;
  wire _43052_;
  wire _43053_;
  wire _43054_;
  wire _43055_;
  wire _43056_;
  wire _43057_;
  wire _43058_;
  wire _43059_;
  wire _43060_;
  wire _43061_;
  wire _43062_;
  wire _43063_;
  wire _43064_;
  wire _43065_;
  wire _43066_;
  wire _43067_;
  wire _43068_;
  wire _43069_;
  wire _43070_;
  wire _43071_;
  wire _43072_;
  wire _43073_;
  wire _43074_;
  wire _43075_;
  wire _43076_;
  wire _43077_;
  wire _43078_;
  wire _43079_;
  wire _43080_;
  wire _43081_;
  wire _43082_;
  wire _43083_;
  wire _43084_;
  wire _43085_;
  wire _43086_;
  wire _43087_;
  wire _43088_;
  wire _43089_;
  wire _43090_;
  wire _43091_;
  wire _43092_;
  wire _43093_;
  wire _43094_;
  wire _43095_;
  wire _43096_;
  wire _43097_;
  wire _43098_;
  wire _43099_;
  wire _43100_;
  wire _43101_;
  wire _43102_;
  wire _43103_;
  wire _43104_;
  wire _43105_;
  wire _43106_;
  wire _43107_;
  wire _43108_;
  wire _43109_;
  wire _43110_;
  wire _43111_;
  wire _43112_;
  wire _43113_;
  wire _43114_;
  wire _43115_;
  wire _43116_;
  wire _43117_;
  wire _43118_;
  wire _43119_;
  wire _43120_;
  wire _43121_;
  wire _43122_;
  wire _43123_;
  wire _43124_;
  wire _43125_;
  wire _43126_;
  wire _43127_;
  wire _43128_;
  wire _43129_;
  wire _43130_;
  wire _43131_;
  wire _43132_;
  wire _43133_;
  wire _43134_;
  wire _43135_;
  wire _43136_;
  wire _43137_;
  wire _43138_;
  wire _43139_;
  wire _43140_;
  wire _43141_;
  wire _43142_;
  wire _43143_;
  wire _43144_;
  wire _43145_;
  wire _43146_;
  wire _43147_;
  wire _43148_;
  wire _43149_;
  wire _43150_;
  wire _43151_;
  wire _43152_;
  wire _43153_;
  wire _43154_;
  wire _43155_;
  wire _43156_;
  wire _43157_;
  wire _43158_;
  wire _43159_;
  wire _43160_;
  wire _43161_;
  wire _43162_;
  wire _43163_;
  wire _43164_;
  wire _43165_;
  wire _43166_;
  wire _43167_;
  wire _43168_;
  wire _43169_;
  wire _43170_;
  wire _43171_;
  wire _43172_;
  wire _43173_;
  wire _43174_;
  wire _43175_;
  wire _43176_;
  wire _43177_;
  wire _43178_;
  wire _43179_;
  wire _43180_;
  wire _43181_;
  wire _43182_;
  wire _43183_;
  wire _43184_;
  wire _43185_;
  wire _43186_;
  wire _43187_;
  wire _43188_;
  wire _43189_;
  wire _43190_;
  wire _43191_;
  wire _43192_;
  wire _43193_;
  wire _43194_;
  wire _43195_;
  wire _43196_;
  wire _43197_;
  wire _43198_;
  wire _43199_;
  wire _43200_;
  wire _43201_;
  wire _43202_;
  wire _43203_;
  wire _43204_;
  wire _43205_;
  wire _43206_;
  wire _43207_;
  wire _43208_;
  wire _43209_;
  wire _43210_;
  wire _43211_;
  wire _43212_;
  wire _43213_;
  wire _43214_;
  wire _43215_;
  wire _43216_;
  wire _43217_;
  wire _43218_;
  wire _43219_;
  wire _43220_;
  wire _43221_;
  wire _43222_;
  wire _43223_;
  wire _43224_;
  wire _43225_;
  wire _43226_;
  wire _43227_;
  wire _43228_;
  wire _43229_;
  wire _43230_;
  wire _43231_;
  wire _43232_;
  wire _43233_;
  wire _43234_;
  wire _43235_;
  wire _43236_;
  wire _43237_;
  wire _43238_;
  wire _43239_;
  wire _43240_;
  wire _43241_;
  wire _43242_;
  wire _43243_;
  wire _43244_;
  wire _43245_;
  wire _43246_;
  wire _43247_;
  wire _43248_;
  wire _43249_;
  wire _43250_;
  wire _43251_;
  wire _43252_;
  wire _43253_;
  wire _43254_;
  wire _43255_;
  wire _43256_;
  wire _43257_;
  wire _43258_;
  wire _43259_;
  wire _43260_;
  wire _43261_;
  wire _43262_;
  wire _43263_;
  wire _43264_;
  wire _43265_;
  wire _43266_;
  wire _43267_;
  wire _43268_;
  wire _43269_;
  wire _43270_;
  wire _43271_;
  wire _43272_;
  wire _43273_;
  wire _43274_;
  wire _43275_;
  wire _43276_;
  wire _43277_;
  wire _43278_;
  wire _43279_;
  wire _43280_;
  wire _43281_;
  wire _43282_;
  wire _43283_;
  wire _43284_;
  wire _43285_;
  wire _43286_;
  wire _43287_;
  wire _43288_;
  wire _43289_;
  wire _43290_;
  wire _43291_;
  wire _43292_;
  wire _43293_;
  wire _43294_;
  wire _43295_;
  wire _43296_;
  wire _43297_;
  wire _43298_;
  wire _43299_;
  wire _43300_;
  wire _43301_;
  wire _43302_;
  wire _43303_;
  wire _43304_;
  wire _43305_;
  wire _43306_;
  wire _43307_;
  wire _43308_;
  wire _43309_;
  wire _43310_;
  wire _43311_;
  wire _43312_;
  wire _43313_;
  wire _43314_;
  wire _43315_;
  wire _43316_;
  wire _43317_;
  wire _43318_;
  wire _43319_;
  wire _43320_;
  wire _43321_;
  wire _43322_;
  wire _43323_;
  wire _43324_;
  wire _43325_;
  wire _43326_;
  wire _43327_;
  wire _43328_;
  wire _43329_;
  wire _43330_;
  wire _43331_;
  wire _43332_;
  wire _43333_;
  wire _43334_;
  wire _43335_;
  wire _43336_;
  wire _43337_;
  wire _43338_;
  wire _43339_;
  wire _43340_;
  wire _43341_;
  wire _43342_;
  wire _43343_;
  wire _43344_;
  wire _43345_;
  wire _43346_;
  wire _43347_;
  wire _43348_;
  wire _43349_;
  wire _43350_;
  wire _43351_;
  wire _43352_;
  wire _43353_;
  wire _43354_;
  wire _43355_;
  wire _43356_;
  wire _43357_;
  wire _43358_;
  wire _43359_;
  wire _43360_;
  wire _43361_;
  wire _43362_;
  wire _43363_;
  wire _43364_;
  wire _43365_;
  wire _43366_;
  wire _43367_;
  wire _43368_;
  wire _43369_;
  wire _43370_;
  wire _43371_;
  wire _43372_;
  wire _43373_;
  wire _43374_;
  wire _43375_;
  wire _43376_;
  wire _43377_;
  wire _43378_;
  wire _43379_;
  wire _43380_;
  wire _43381_;
  wire _43382_;
  wire _43383_;
  wire _43384_;
  wire _43385_;
  wire _43386_;
  wire _43387_;
  wire _43388_;
  wire _43389_;
  wire _43390_;
  wire _43391_;
  wire _43392_;
  wire _43393_;
  wire _43394_;
  wire _43395_;
  wire _43396_;
  wire _43397_;
  wire _43398_;
  wire _43399_;
  wire _43400_;
  wire _43401_;
  wire _43402_;
  wire _43403_;
  wire _43404_;
  wire _43405_;
  wire _43406_;
  wire _43407_;
  wire _43408_;
  wire _43409_;
  wire _43410_;
  wire _43411_;
  wire _43412_;
  wire _43413_;
  wire _43414_;
  wire _43415_;
  wire _43416_;
  wire _43417_;
  wire _43418_;
  wire _43419_;
  wire _43420_;
  wire _43421_;
  wire _43422_;
  wire _43423_;
  wire _43424_;
  wire _43425_;
  wire _43426_;
  wire _43427_;
  wire _43428_;
  wire _43429_;
  wire _43430_;
  wire _43431_;
  wire _43432_;
  wire _43433_;
  wire _43434_;
  wire _43435_;
  wire _43436_;
  wire _43437_;
  wire _43438_;
  wire _43439_;
  wire _43440_;
  wire _43441_;
  wire _43442_;
  wire _43443_;
  wire _43444_;
  wire _43445_;
  wire _43446_;
  wire _43447_;
  wire _43448_;
  wire _43449_;
  wire _43450_;
  wire _43451_;
  wire _43452_;
  wire _43453_;
  wire _43454_;
  wire _43455_;
  wire _43456_;
  wire _43457_;
  wire _43458_;
  wire _43459_;
  wire _43460_;
  wire _43461_;
  wire _43462_;
  wire _43463_;
  wire _43464_;
  wire _43465_;
  wire _43466_;
  wire _43467_;
  wire _43468_;
  wire _43469_;
  wire _43470_;
  wire _43471_;
  wire _43472_;
  wire _43473_;
  wire _43474_;
  wire _43475_;
  wire _43476_;
  wire _43477_;
  wire _43478_;
  wire _43479_;
  wire _43480_;
  wire _43481_;
  wire _43482_;
  wire _43483_;
  wire _43484_;
  wire _43485_;
  wire _43486_;
  wire _43487_;
  wire _43488_;
  wire _43489_;
  wire _43490_;
  wire _43491_;
  wire _43492_;
  wire _43493_;
  wire _43494_;
  wire _43495_;
  wire _43496_;
  wire _43497_;
  wire _43498_;
  wire _43499_;
  wire _43500_;
  wire _43501_;
  wire _43502_;
  wire _43503_;
  wire _43504_;
  wire _43505_;
  wire _43506_;
  wire _43507_;
  wire _43508_;
  wire _43509_;
  wire _43510_;
  wire _43511_;
  wire _43512_;
  wire _43513_;
  wire _43514_;
  wire _43515_;
  wire _43516_;
  wire _43517_;
  wire _43518_;
  wire _43519_;
  wire _43520_;
  wire _43521_;
  wire _43522_;
  wire _43523_;
  wire _43524_;
  wire _43525_;
  wire _43526_;
  wire _43527_;
  wire _43528_;
  wire _43529_;
  wire _43530_;
  wire _43531_;
  wire _43532_;
  wire _43533_;
  wire _43534_;
  wire _43535_;
  wire _43536_;
  wire _43537_;
  wire _43538_;
  wire _43539_;
  wire _43540_;
  wire _43541_;
  wire _43542_;
  wire _43543_;
  wire _43544_;
  wire _43545_;
  wire _43546_;
  wire _43547_;
  wire _43548_;
  wire _43549_;
  wire _43550_;
  wire _43551_;
  wire _43552_;
  wire _43553_;
  wire _43554_;
  wire _43555_;
  wire _43556_;
  wire _43557_;
  wire _43558_;
  wire _43559_;
  wire _43560_;
  wire _43561_;
  wire _43562_;
  wire _43563_;
  wire _43564_;
  wire _43565_;
  wire _43566_;
  wire _43567_;
  wire _43568_;
  wire _43569_;
  wire _43570_;
  wire _43571_;
  wire _43572_;
  wire _43573_;
  wire _43574_;
  wire _43575_;
  wire _43576_;
  wire _43577_;
  wire _43578_;
  wire _43579_;
  wire _43580_;
  wire _43581_;
  wire _43582_;
  wire _43583_;
  wire _43584_;
  wire _43585_;
  wire _43586_;
  wire _43587_;
  wire _43588_;
  wire _43589_;
  wire _43590_;
  wire _43591_;
  wire _43592_;
  wire _43593_;
  wire _43594_;
  wire _43595_;
  wire _43596_;
  wire _43597_;
  wire _43598_;
  wire _43599_;
  wire _43600_;
  wire _43601_;
  wire _43602_;
  wire _43603_;
  wire _43604_;
  wire _43605_;
  wire _43606_;
  wire _43607_;
  wire _43608_;
  wire _43609_;
  wire _43610_;
  wire _43611_;
  wire _43612_;
  wire _43613_;
  wire _43614_;
  wire _43615_;
  wire _43616_;
  wire _43617_;
  wire _43618_;
  wire _43619_;
  wire _43620_;
  wire _43621_;
  wire _43622_;
  wire _43623_;
  wire _43624_;
  wire _43625_;
  wire _43626_;
  wire _43627_;
  wire _43628_;
  wire _43629_;
  wire _43630_;
  wire _43631_;
  wire _43632_;
  wire _43633_;
  wire _43634_;
  wire _43635_;
  wire _43636_;
  wire _43637_;
  wire _43638_;
  wire _43639_;
  wire _43640_;
  wire _43641_;
  wire _43642_;
  wire _43643_;
  wire _43644_;
  wire _43645_;
  wire _43646_;
  wire _43647_;
  wire _43648_;
  wire _43649_;
  wire _43650_;
  wire _43651_;
  wire _43652_;
  wire _43653_;
  wire _43654_;
  wire _43655_;
  wire _43656_;
  wire _43657_;
  wire _43658_;
  wire _43659_;
  wire _43660_;
  wire _43661_;
  wire _43662_;
  wire _43663_;
  wire _43664_;
  wire _43665_;
  wire _43666_;
  wire _43667_;
  wire _43668_;
  wire _43669_;
  wire _43670_;
  wire _43671_;
  wire _43672_;
  wire _43673_;
  wire _43674_;
  wire _43675_;
  wire _43676_;
  wire _43677_;
  wire _43678_;
  wire _43679_;
  wire _43680_;
  wire _43681_;
  wire _43682_;
  wire _43683_;
  wire _43684_;
  wire _43685_;
  wire _43686_;
  wire _43687_;
  wire _43688_;
  wire _43689_;
  wire _43690_;
  wire _43691_;
  wire _43692_;
  wire _43693_;
  wire _43694_;
  wire _43695_;
  wire _43696_;
  wire _43697_;
  wire _43698_;
  wire _43699_;
  wire _43700_;
  wire _43701_;
  wire _43702_;
  wire _43703_;
  wire _43704_;
  wire _43705_;
  wire _43706_;
  wire _43707_;
  wire _43708_;
  wire _43709_;
  wire _43710_;
  wire _43711_;
  wire _43712_;
  wire _43713_;
  wire _43714_;
  wire _43715_;
  wire _43716_;
  wire _43717_;
  wire _43718_;
  wire _43719_;
  wire _43720_;
  wire _43721_;
  wire _43722_;
  wire _43723_;
  wire _43724_;
  wire _43725_;
  wire _43726_;
  wire _43727_;
  wire _43728_;
  wire _43729_;
  wire _43730_;
  wire _43731_;
  wire _43732_;
  wire _43733_;
  wire _43734_;
  wire _43735_;
  wire _43736_;
  wire _43737_;
  wire _43738_;
  wire _43739_;
  wire _43740_;
  wire _43741_;
  wire _43742_;
  wire _43743_;
  wire _43744_;
  wire _43745_;
  wire _43746_;
  wire _43747_;
  wire _43748_;
  wire _43749_;
  wire _43750_;
  wire _43751_;
  wire _43752_;
  wire _43753_;
  wire _43754_;
  wire _43755_;
  wire _43756_;
  wire _43757_;
  wire _43758_;
  wire _43759_;
  wire _43760_;
  wire _43761_;
  wire _43762_;
  wire _43763_;
  wire _43764_;
  wire _43765_;
  wire _43766_;
  wire _43767_;
  wire _43768_;
  wire _43769_;
  wire _43770_;
  wire _43771_;
  wire _43772_;
  wire _43773_;
  wire _43774_;
  wire _43775_;
  wire _43776_;
  wire _43777_;
  wire _43778_;
  wire _43779_;
  wire _43780_;
  wire _43781_;
  wire _43782_;
  wire _43783_;
  wire _43784_;
  wire _43785_;
  wire _43786_;
  wire _43787_;
  wire _43788_;
  wire _43789_;
  wire _43790_;
  wire _43791_;
  wire _43792_;
  wire _43793_;
  wire _43794_;
  wire _43795_;
  wire _43796_;
  wire _43797_;
  wire _43798_;
  wire _43799_;
  wire _43800_;
  wire _43801_;
  wire _43802_;
  wire _43803_;
  wire _43804_;
  wire _43805_;
  wire _43806_;
  wire _43807_;
  wire _43808_;
  wire _43809_;
  wire _43810_;
  wire _43811_;
  wire [7:0] ACC_gm;
  wire [7:0] acc;
  input clk;
  wire [31:0] cxrom_data_out;
  wire inst_finished_r;
  wire \oc8051_gm_cxrom_1.cell0.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.data ;
  wire \oc8051_gm_cxrom_1.cell0.rst ;
  wire \oc8051_gm_cxrom_1.cell0.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell0.word ;
  wire \oc8051_gm_cxrom_1.cell1.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.data ;
  wire \oc8051_gm_cxrom_1.cell1.rst ;
  wire \oc8051_gm_cxrom_1.cell1.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell1.word ;
  wire \oc8051_gm_cxrom_1.cell10.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.data ;
  wire \oc8051_gm_cxrom_1.cell10.rst ;
  wire \oc8051_gm_cxrom_1.cell10.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell10.word ;
  wire \oc8051_gm_cxrom_1.cell11.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.data ;
  wire \oc8051_gm_cxrom_1.cell11.rst ;
  wire \oc8051_gm_cxrom_1.cell11.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell11.word ;
  wire \oc8051_gm_cxrom_1.cell12.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.data ;
  wire \oc8051_gm_cxrom_1.cell12.rst ;
  wire \oc8051_gm_cxrom_1.cell12.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell12.word ;
  wire \oc8051_gm_cxrom_1.cell13.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.data ;
  wire \oc8051_gm_cxrom_1.cell13.rst ;
  wire \oc8051_gm_cxrom_1.cell13.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell13.word ;
  wire \oc8051_gm_cxrom_1.cell14.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.data ;
  wire \oc8051_gm_cxrom_1.cell14.rst ;
  wire \oc8051_gm_cxrom_1.cell14.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell14.word ;
  wire \oc8051_gm_cxrom_1.cell15.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.data ;
  wire \oc8051_gm_cxrom_1.cell15.rst ;
  wire \oc8051_gm_cxrom_1.cell15.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell15.word ;
  wire \oc8051_gm_cxrom_1.cell2.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.data ;
  wire \oc8051_gm_cxrom_1.cell2.rst ;
  wire \oc8051_gm_cxrom_1.cell2.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell2.word ;
  wire \oc8051_gm_cxrom_1.cell3.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.data ;
  wire \oc8051_gm_cxrom_1.cell3.rst ;
  wire \oc8051_gm_cxrom_1.cell3.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell3.word ;
  wire \oc8051_gm_cxrom_1.cell4.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.data ;
  wire \oc8051_gm_cxrom_1.cell4.rst ;
  wire \oc8051_gm_cxrom_1.cell4.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell4.word ;
  wire \oc8051_gm_cxrom_1.cell5.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.data ;
  wire \oc8051_gm_cxrom_1.cell5.rst ;
  wire \oc8051_gm_cxrom_1.cell5.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell5.word ;
  wire \oc8051_gm_cxrom_1.cell6.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.data ;
  wire \oc8051_gm_cxrom_1.cell6.rst ;
  wire \oc8051_gm_cxrom_1.cell6.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell6.word ;
  wire \oc8051_gm_cxrom_1.cell7.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.data ;
  wire \oc8051_gm_cxrom_1.cell7.rst ;
  wire \oc8051_gm_cxrom_1.cell7.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell7.word ;
  wire \oc8051_gm_cxrom_1.cell8.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.data ;
  wire \oc8051_gm_cxrom_1.cell8.rst ;
  wire \oc8051_gm_cxrom_1.cell8.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell8.word ;
  wire \oc8051_gm_cxrom_1.cell9.clk ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.data ;
  wire \oc8051_gm_cxrom_1.cell9.rst ;
  wire \oc8051_gm_cxrom_1.cell9.valid ;
  wire [7:0] \oc8051_gm_cxrom_1.cell9.word ;
  wire \oc8051_gm_cxrom_1.clk ;
  wire [31:0] \oc8051_gm_cxrom_1.cxrom_data_out ;
  wire [15:0] \oc8051_gm_cxrom_1.rd_addr_0 ;
  wire \oc8051_gm_cxrom_1.rst ;
  wire [127:0] \oc8051_gm_cxrom_1.word_in ;
  wire [7:0] \oc8051_golden_model_1.ACC ;
  wire [7:0] \oc8051_golden_model_1.ACC_03 ;
  wire [7:0] \oc8051_golden_model_1.ACC_13 ;
  wire [7:0] \oc8051_golden_model_1.ACC_23 ;
  wire [7:0] \oc8051_golden_model_1.ACC_33 ;
  wire [7:0] \oc8051_golden_model_1.ACC_c4 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d6 ;
  wire [7:0] \oc8051_golden_model_1.ACC_d7 ;
  wire [7:0] \oc8051_golden_model_1.ACC_e4 ;
  wire [7:0] \oc8051_golden_model_1.B ;
  wire [7:0] \oc8051_golden_model_1.DPH ;
  wire [7:0] \oc8051_golden_model_1.DPL ;
  wire [7:0] \oc8051_golden_model_1.IE ;
  wire [7:0] \oc8051_golden_model_1.IP ;
  wire [7:0] \oc8051_golden_model_1.IRAM[0] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[10] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[11] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[12] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[13] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[14] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[15] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[1] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[2] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[3] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[4] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[5] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[6] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[7] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[8] ;
  wire [7:0] \oc8051_golden_model_1.IRAM[9] ;
  wire [7:0] \oc8051_golden_model_1.P0 ;
  wire [7:0] \oc8051_golden_model_1.P1 ;
  wire [7:0] \oc8051_golden_model_1.P2 ;
  wire [7:0] \oc8051_golden_model_1.P3 ;
  wire [15:0] \oc8051_golden_model_1.PC ;
  wire [7:0] \oc8051_golden_model_1.PCON ;
  wire [15:0] \oc8051_golden_model_1.PC_22 ;
  wire [15:0] \oc8051_golden_model_1.PC_32 ;
  wire [7:0] \oc8051_golden_model_1.PSW ;
  wire [7:0] \oc8051_golden_model_1.PSW_13 ;
  wire [7:0] \oc8051_golden_model_1.PSW_24 ;
  wire [7:0] \oc8051_golden_model_1.PSW_25 ;
  wire [7:0] \oc8051_golden_model_1.PSW_26 ;
  wire [7:0] \oc8051_golden_model_1.PSW_27 ;
  wire [7:0] \oc8051_golden_model_1.PSW_28 ;
  wire [7:0] \oc8051_golden_model_1.PSW_29 ;
  wire [7:0] \oc8051_golden_model_1.PSW_2a ;
  wire [7:0] \oc8051_golden_model_1.PSW_2b ;
  wire [7:0] \oc8051_golden_model_1.PSW_2c ;
  wire [7:0] \oc8051_golden_model_1.PSW_2d ;
  wire [7:0] \oc8051_golden_model_1.PSW_2e ;
  wire [7:0] \oc8051_golden_model_1.PSW_2f ;
  wire [7:0] \oc8051_golden_model_1.PSW_33 ;
  wire [7:0] \oc8051_golden_model_1.PSW_34 ;
  wire [7:0] \oc8051_golden_model_1.PSW_35 ;
  wire [7:0] \oc8051_golden_model_1.PSW_36 ;
  wire [7:0] \oc8051_golden_model_1.PSW_37 ;
  wire [7:0] \oc8051_golden_model_1.PSW_38 ;
  wire [7:0] \oc8051_golden_model_1.PSW_39 ;
  wire [7:0] \oc8051_golden_model_1.PSW_3a ;
  wire [7:0] \oc8051_golden_model_1.PSW_3b ;
  wire [7:0] \oc8051_golden_model_1.PSW_3c ;
  wire [7:0] \oc8051_golden_model_1.PSW_3d ;
  wire [7:0] \oc8051_golden_model_1.PSW_3e ;
  wire [7:0] \oc8051_golden_model_1.PSW_3f ;
  wire [7:0] \oc8051_golden_model_1.PSW_72 ;
  wire [7:0] \oc8051_golden_model_1.PSW_82 ;
  wire [7:0] \oc8051_golden_model_1.PSW_84 ;
  wire [7:0] \oc8051_golden_model_1.PSW_94 ;
  wire [7:0] \oc8051_golden_model_1.PSW_95 ;
  wire [7:0] \oc8051_golden_model_1.PSW_96 ;
  wire [7:0] \oc8051_golden_model_1.PSW_97 ;
  wire [7:0] \oc8051_golden_model_1.PSW_98 ;
  wire [7:0] \oc8051_golden_model_1.PSW_99 ;
  wire [7:0] \oc8051_golden_model_1.PSW_9a ;
  wire [7:0] \oc8051_golden_model_1.PSW_9b ;
  wire [7:0] \oc8051_golden_model_1.PSW_9c ;
  wire [7:0] \oc8051_golden_model_1.PSW_9d ;
  wire [7:0] \oc8051_golden_model_1.PSW_9e ;
  wire [7:0] \oc8051_golden_model_1.PSW_9f ;
  wire [7:0] \oc8051_golden_model_1.PSW_a0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a2 ;
  wire [7:0] \oc8051_golden_model_1.PSW_a4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b0 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b4 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b5 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b6 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b7 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b8 ;
  wire [7:0] \oc8051_golden_model_1.PSW_b9 ;
  wire [7:0] \oc8051_golden_model_1.PSW_ba ;
  wire [7:0] \oc8051_golden_model_1.PSW_bb ;
  wire [7:0] \oc8051_golden_model_1.PSW_bc ;
  wire [7:0] \oc8051_golden_model_1.PSW_bd ;
  wire [7:0] \oc8051_golden_model_1.PSW_be ;
  wire [7:0] \oc8051_golden_model_1.PSW_bf ;
  wire [7:0] \oc8051_golden_model_1.PSW_c3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d3 ;
  wire [7:0] \oc8051_golden_model_1.PSW_d4 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_0 ;
  wire [7:0] \oc8051_golden_model_1.RD_IRAM_1 ;
  wire [3:0] \oc8051_golden_model_1.RD_IRAM_ADDR ;
  wire [15:0] \oc8051_golden_model_1.RD_ROM_0_ADDR ;
  wire [7:0] \oc8051_golden_model_1.SBUF ;
  wire [7:0] \oc8051_golden_model_1.SCON ;
  wire [7:0] \oc8051_golden_model_1.SP ;
  wire [7:0] \oc8051_golden_model_1.TCON ;
  wire [7:0] \oc8051_golden_model_1.TH0 ;
  wire [7:0] \oc8051_golden_model_1.TH1 ;
  wire [7:0] \oc8051_golden_model_1.TL0 ;
  wire [7:0] \oc8051_golden_model_1.TL1 ;
  wire [7:0] \oc8051_golden_model_1.TMOD ;
  wire \oc8051_golden_model_1.clk ;
  wire [1:0] \oc8051_golden_model_1.n0006 ;
  wire [7:0] \oc8051_golden_model_1.n0007 ;
  wire [7:0] \oc8051_golden_model_1.n0011 ;
  wire [7:0] \oc8051_golden_model_1.n0019 ;
  wire [7:0] \oc8051_golden_model_1.n0023 ;
  wire [7:0] \oc8051_golden_model_1.n0027 ;
  wire [7:0] \oc8051_golden_model_1.n0031 ;
  wire [7:0] \oc8051_golden_model_1.n0035 ;
  wire [7:0] \oc8051_golden_model_1.n0039 ;
  wire [7:0] \oc8051_golden_model_1.n0561 ;
  wire [7:0] \oc8051_golden_model_1.n0594 ;
  wire [15:0] \oc8051_golden_model_1.n0701 ;
  wire [15:0] \oc8051_golden_model_1.n0733 ;
  wire [7:0] \oc8051_golden_model_1.n0994 ;
  wire [3:0] \oc8051_golden_model_1.n1071 ;
  wire [3:0] \oc8051_golden_model_1.n1073 ;
  wire [3:0] \oc8051_golden_model_1.n1075 ;
  wire [3:0] \oc8051_golden_model_1.n1076 ;
  wire [3:0] \oc8051_golden_model_1.n1077 ;
  wire [3:0] \oc8051_golden_model_1.n1078 ;
  wire [3:0] \oc8051_golden_model_1.n1079 ;
  wire [3:0] \oc8051_golden_model_1.n1080 ;
  wire [3:0] \oc8051_golden_model_1.n1081 ;
  wire \oc8051_golden_model_1.n1118 ;
  wire \oc8051_golden_model_1.n1146 ;
  wire [8:0] \oc8051_golden_model_1.n1147 ;
  wire [8:0] \oc8051_golden_model_1.n1148 ;
  wire [7:0] \oc8051_golden_model_1.n1149 ;
  wire \oc8051_golden_model_1.n1150 ;
  wire \oc8051_golden_model_1.n1151 ;
  wire [2:0] \oc8051_golden_model_1.n1152 ;
  wire \oc8051_golden_model_1.n1153 ;
  wire [1:0] \oc8051_golden_model_1.n1154 ;
  wire [7:0] \oc8051_golden_model_1.n1155 ;
  wire [15:0] \oc8051_golden_model_1.n1181 ;
  wire [7:0] \oc8051_golden_model_1.n1183 ;
  wire [8:0] \oc8051_golden_model_1.n1185 ;
  wire [8:0] \oc8051_golden_model_1.n1189 ;
  wire \oc8051_golden_model_1.n1190 ;
  wire [3:0] \oc8051_golden_model_1.n1191 ;
  wire [4:0] \oc8051_golden_model_1.n1192 ;
  wire [4:0] \oc8051_golden_model_1.n1196 ;
  wire \oc8051_golden_model_1.n1197 ;
  wire [8:0] \oc8051_golden_model_1.n1198 ;
  wire \oc8051_golden_model_1.n1206 ;
  wire [7:0] \oc8051_golden_model_1.n1207 ;
  wire [8:0] \oc8051_golden_model_1.n1211 ;
  wire \oc8051_golden_model_1.n1212 ;
  wire [4:0] \oc8051_golden_model_1.n1217 ;
  wire \oc8051_golden_model_1.n1218 ;
  wire \oc8051_golden_model_1.n1226 ;
  wire [7:0] \oc8051_golden_model_1.n1227 ;
  wire [8:0] \oc8051_golden_model_1.n1229 ;
  wire [8:0] \oc8051_golden_model_1.n1231 ;
  wire \oc8051_golden_model_1.n1232 ;
  wire [3:0] \oc8051_golden_model_1.n1233 ;
  wire [4:0] \oc8051_golden_model_1.n1234 ;
  wire [4:0] \oc8051_golden_model_1.n1236 ;
  wire \oc8051_golden_model_1.n1237 ;
  wire [8:0] \oc8051_golden_model_1.n1238 ;
  wire \oc8051_golden_model_1.n1245 ;
  wire [7:0] \oc8051_golden_model_1.n1246 ;
  wire [8:0] \oc8051_golden_model_1.n1249 ;
  wire \oc8051_golden_model_1.n1250 ;
  wire \oc8051_golden_model_1.n1257 ;
  wire [7:0] \oc8051_golden_model_1.n1258 ;
  wire [8:0] \oc8051_golden_model_1.n1260 ;
  wire [8:0] \oc8051_golden_model_1.n1262 ;
  wire \oc8051_golden_model_1.n1263 ;
  wire [4:0] \oc8051_golden_model_1.n1264 ;
  wire [4:0] \oc8051_golden_model_1.n1266 ;
  wire \oc8051_golden_model_1.n1267 ;
  wire [8:0] \oc8051_golden_model_1.n1268 ;
  wire \oc8051_golden_model_1.n1275 ;
  wire [7:0] \oc8051_golden_model_1.n1276 ;
  wire [4:0] \oc8051_golden_model_1.n1278 ;
  wire \oc8051_golden_model_1.n1279 ;
  wire [7:0] \oc8051_golden_model_1.n1280 ;
  wire [8:0] \oc8051_golden_model_1.n1282 ;
  wire \oc8051_golden_model_1.n1283 ;
  wire \oc8051_golden_model_1.n1290 ;
  wire [7:0] \oc8051_golden_model_1.n1291 ;
  wire [7:0] \oc8051_golden_model_1.n1292 ;
  wire [8:0] \oc8051_golden_model_1.n1295 ;
  wire [8:0] \oc8051_golden_model_1.n1296 ;
  wire [7:0] \oc8051_golden_model_1.n1297 ;
  wire \oc8051_golden_model_1.n1298 ;
  wire [7:0] \oc8051_golden_model_1.n1299 ;
  wire [7:0] \oc8051_golden_model_1.n1300 ;
  wire [8:0] \oc8051_golden_model_1.n1303 ;
  wire [8:0] \oc8051_golden_model_1.n1305 ;
  wire \oc8051_golden_model_1.n1306 ;
  wire [4:0] \oc8051_golden_model_1.n1307 ;
  wire [4:0] \oc8051_golden_model_1.n1309 ;
  wire \oc8051_golden_model_1.n1310 ;
  wire \oc8051_golden_model_1.n1317 ;
  wire [7:0] \oc8051_golden_model_1.n1318 ;
  wire [8:0] \oc8051_golden_model_1.n1322 ;
  wire \oc8051_golden_model_1.n1323 ;
  wire [4:0] \oc8051_golden_model_1.n1325 ;
  wire \oc8051_golden_model_1.n1326 ;
  wire \oc8051_golden_model_1.n1333 ;
  wire [7:0] \oc8051_golden_model_1.n1334 ;
  wire [8:0] \oc8051_golden_model_1.n1338 ;
  wire \oc8051_golden_model_1.n1339 ;
  wire [4:0] \oc8051_golden_model_1.n1341 ;
  wire \oc8051_golden_model_1.n1342 ;
  wire \oc8051_golden_model_1.n1349 ;
  wire [7:0] \oc8051_golden_model_1.n1350 ;
  wire [8:0] \oc8051_golden_model_1.n1354 ;
  wire \oc8051_golden_model_1.n1355 ;
  wire [4:0] \oc8051_golden_model_1.n1357 ;
  wire \oc8051_golden_model_1.n1358 ;
  wire \oc8051_golden_model_1.n1365 ;
  wire [7:0] \oc8051_golden_model_1.n1366 ;
  wire \oc8051_golden_model_1.n1520 ;
  wire [6:0] \oc8051_golden_model_1.n1521 ;
  wire [7:0] \oc8051_golden_model_1.n1522 ;
  wire \oc8051_golden_model_1.n1545 ;
  wire [7:0] \oc8051_golden_model_1.n1546 ;
  wire [3:0] \oc8051_golden_model_1.n1553 ;
  wire \oc8051_golden_model_1.n1554 ;
  wire [7:0] \oc8051_golden_model_1.n1555 ;
  wire [7:0] \oc8051_golden_model_1.n1680 ;
  wire \oc8051_golden_model_1.n1683 ;
  wire \oc8051_golden_model_1.n1685 ;
  wire \oc8051_golden_model_1.n1691 ;
  wire [7:0] \oc8051_golden_model_1.n1692 ;
  wire \oc8051_golden_model_1.n1696 ;
  wire \oc8051_golden_model_1.n1698 ;
  wire \oc8051_golden_model_1.n1704 ;
  wire [7:0] \oc8051_golden_model_1.n1705 ;
  wire \oc8051_golden_model_1.n1709 ;
  wire \oc8051_golden_model_1.n1711 ;
  wire \oc8051_golden_model_1.n1717 ;
  wire [7:0] \oc8051_golden_model_1.n1718 ;
  wire \oc8051_golden_model_1.n1722 ;
  wire \oc8051_golden_model_1.n1724 ;
  wire \oc8051_golden_model_1.n1730 ;
  wire [7:0] \oc8051_golden_model_1.n1731 ;
  wire \oc8051_golden_model_1.n1733 ;
  wire [7:0] \oc8051_golden_model_1.n1734 ;
  wire [7:0] \oc8051_golden_model_1.n1735 ;
  wire [15:0] \oc8051_golden_model_1.n1739 ;
  wire \oc8051_golden_model_1.n1745 ;
  wire [7:0] \oc8051_golden_model_1.n1746 ;
  wire \oc8051_golden_model_1.n1749 ;
  wire [7:0] \oc8051_golden_model_1.n1750 ;
  wire \oc8051_golden_model_1.n1765 ;
  wire [7:0] \oc8051_golden_model_1.n1766 ;
  wire \oc8051_golden_model_1.n1771 ;
  wire [7:0] \oc8051_golden_model_1.n1772 ;
  wire \oc8051_golden_model_1.n1777 ;
  wire [7:0] \oc8051_golden_model_1.n1778 ;
  wire \oc8051_golden_model_1.n1783 ;
  wire [7:0] \oc8051_golden_model_1.n1784 ;
  wire \oc8051_golden_model_1.n1789 ;
  wire [7:0] \oc8051_golden_model_1.n1790 ;
  wire [7:0] \oc8051_golden_model_1.n1791 ;
  wire [3:0] \oc8051_golden_model_1.n1792 ;
  wire [7:0] \oc8051_golden_model_1.n1793 ;
  wire [7:0] \oc8051_golden_model_1.n1828 ;
  wire \oc8051_golden_model_1.n1847 ;
  wire [7:0] \oc8051_golden_model_1.n1848 ;
  wire [7:0] \oc8051_golden_model_1.n1852 ;
  wire [3:0] \oc8051_golden_model_1.n1853 ;
  wire [7:0] \oc8051_golden_model_1.n1854 ;
  wire \oc8051_golden_model_1.rst ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire \oc8051_top_1.ea_int ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff0 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff1 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff2 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff3 ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dack_ir ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_o ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dadr_ot ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_ir ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ddat_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire \oc8051_top_1.oc8051_memory_interface1.dstb_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.dwe_o ;
  wire \oc8051_top_1.oc8051_memory_interface1.ea_int ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.ea_int ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.txd ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [7:0] \oc8051_top_1.psw ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.txd_o ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [15:0] \oc8051_top_1.wbd_adr_o ;
  wire \oc8051_top_1.wbd_cyc_o ;
  wire [7:0] \oc8051_top_1.wbd_dat_o ;
  wire \oc8051_top_1.wbd_stb_o ;
  wire \oc8051_top_1.wbd_we_o ;
  wire op0_cnst;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid_acc;
  output property_invalid_iram;
  output property_invalid_pc;
  wire [7:0] psw;
  wire [3:0] rd_iram_addr;
  wire [15:0] rd_rom_0_addr;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  wire txd_o;
  wire [15:0] wbd_adr_o;
  wire wbd_cyc_o;
  wire [7:0] wbd_dat_o;
  wire wbd_stb_o;
  wire wbd_we_o;
  input [127:0] word_in;
  not _43812_ (_42882_, rst);
  not _43813_ (_18188_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  not _43814_ (_18199_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _43815_ (_18210_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _18199_);
  and _43816_ (_18221_, _18210_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _43817_ (_18232_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _18199_);
  and _43818_ (_18243_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _18199_);
  nor _43819_ (_18254_, _18243_, _18232_);
  and _43820_ (_18265_, _18254_, _18221_);
  nor _43821_ (_18276_, _18265_, _18188_);
  and _43822_ (_18287_, _18188_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _43823_ (_18298_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  and _43824_ (_18309_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _18298_);
  nor _43825_ (_18320_, _18309_, _18287_);
  not _43826_ (_18331_, _18320_);
  and _43827_ (_18342_, _18331_, _18265_);
  or _43828_ (_18353_, _18342_, _18276_);
  and _43829_ (_22216_, _18353_, _42882_);
  nor _43830_ (_18374_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  not _43831_ (_18385_, _18374_);
  and _43832_ (_18396_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  and _43833_ (_18407_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _43834_ (_18418_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not _43835_ (_18429_, _18418_);
  not _43836_ (_18440_, _18309_);
  nor _43837_ (_18451_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  not _43838_ (_18462_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _43839_ (_18473_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _18462_);
  nor _43840_ (_18483_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  not _43841_ (_18494_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor _43842_ (_18505_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _18494_);
  nor _43843_ (_18516_, _18505_, _18483_);
  nor _43844_ (_18527_, _18516_, _18473_);
  not _43845_ (_18538_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _43846_ (_18549_, _18473_, _18538_);
  nor _43847_ (_18560_, _18549_, _18527_);
  and _43848_ (_18571_, _18560_, _18451_);
  not _43849_ (_18582_, _18571_);
  and _43850_ (_18593_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _43851_ (_18604_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  not _43852_ (_18615_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _43853_ (_18626_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0], _18615_);
  and _43854_ (_18637_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _43855_ (_18648_, _18637_, _18604_);
  and _43856_ (_18669_, _18648_, _18582_);
  nor _43857_ (_18670_, _18669_, _18440_);
  not _43858_ (_18681_, _18287_);
  nor _43859_ (_18702_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nor _43860_ (_18703_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _18494_);
  nor _43861_ (_18714_, _18703_, _18702_);
  nor _43862_ (_18735_, _18714_, _18473_);
  not _43863_ (_18736_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and _43864_ (_18747_, _18473_, _18736_);
  nor _43865_ (_18768_, _18747_, _18735_);
  and _43866_ (_18769_, _18768_, _18451_);
  not _43867_ (_18780_, _18769_);
  and _43868_ (_18801_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and _43869_ (_18802_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _43870_ (_18813_, _18802_, _18801_);
  and _43871_ (_18834_, _18813_, _18780_);
  nor _43872_ (_18835_, _18834_, _18681_);
  nor _43873_ (_18845_, _18835_, _18670_);
  nor _43874_ (_18866_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nor _43875_ (_18867_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _18494_);
  nor _43876_ (_18878_, _18867_, _18866_);
  nor _43877_ (_18889_, _18878_, _18473_);
  not _43878_ (_18900_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _43879_ (_18911_, _18473_, _18900_);
  nor _43880_ (_18922_, _18911_, _18889_);
  and _43881_ (_18933_, _18922_, _18451_);
  not _43882_ (_18944_, _18933_);
  and _43883_ (_18955_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  and _43884_ (_18966_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _43885_ (_18977_, _18966_, _18955_);
  and _43886_ (_18988_, _18977_, _18944_);
  nor _43887_ (_18999_, _18988_, _18331_);
  nor _43888_ (_19010_, _18999_, _18374_);
  and _43889_ (_19021_, _19010_, _18845_);
  nor _43890_ (_19032_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nor _43891_ (_19043_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _18494_);
  nor _43892_ (_19054_, _19043_, _19032_);
  nor _43893_ (_19065_, _19054_, _18473_);
  not _43894_ (_19076_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and _43895_ (_19087_, _18473_, _19076_);
  nor _43896_ (_19098_, _19087_, _19065_);
  and _43897_ (_19109_, _19098_, _18451_);
  not _43898_ (_19120_, _19109_);
  and _43899_ (_19131_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and _43900_ (_19142_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _43901_ (_19153_, _19142_, _19131_);
  and _43902_ (_19164_, _19153_, _19120_);
  and _43903_ (_19175_, _19164_, _18374_);
  nor _43904_ (_19185_, _19175_, _19021_);
  not _43905_ (_19196_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _43906_ (_19207_, _19196_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _43907_ (_19218_, _19207_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _43908_ (_19229_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _43909_ (_19240_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _43910_ (_19251_, _19240_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _43911_ (_19262_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _43912_ (_19272_, _19262_, _19229_);
  nor _43913_ (_19283_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _43914_ (_19294_, _19283_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and _43915_ (_19305_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not _43916_ (_19316_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _43917_ (_19327_, _19207_, _19316_);
  and _43918_ (_19338_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  nor _43919_ (_19349_, _19338_, _19305_);
  and _43920_ (_19359_, _19349_, _19272_);
  and _43921_ (_19370_, _19283_, _19196_);
  and _43922_ (_19381_, _19370_, _19098_);
  and _43923_ (_19392_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _43924_ (_19403_, _19392_, _19316_);
  and _43925_ (_19414_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _43926_ (_19425_, _19392_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _43927_ (_19436_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  nor _43928_ (_19446_, _19436_, _19414_);
  not _43929_ (_19457_, _19446_);
  nor _43930_ (_19468_, _19457_, _19381_);
  and _43931_ (_19479_, _19468_, _19359_);
  not _43932_ (_19490_, _19479_);
  and _43933_ (_19501_, _19490_, _19185_);
  not _43934_ (_19512_, _19501_);
  nor _43935_ (_19522_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nor _43936_ (_19533_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _18494_);
  nor _43937_ (_19544_, _19533_, _19522_);
  nor _43938_ (_19555_, _19544_, _18473_);
  not _43939_ (_19566_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _43940_ (_19577_, _18473_, _19566_);
  nor _43941_ (_19588_, _19577_, _19555_);
  and _43942_ (_19599_, _19588_, _18451_);
  not _43943_ (_19609_, _19599_);
  and _43944_ (_19620_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  and _43945_ (_19631_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _43946_ (_19642_, _19631_, _19620_);
  and _43947_ (_19653_, _19642_, _19609_);
  nor _43948_ (_19664_, _19653_, _18440_);
  nor _43949_ (_19675_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nor _43950_ (_19686_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _18494_);
  nor _43951_ (_19696_, _19686_, _19675_);
  nor _43952_ (_19707_, _19696_, _18473_);
  not _43953_ (_19718_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _43954_ (_19729_, _18473_, _19718_);
  nor _43955_ (_19740_, _19729_, _19707_);
  and _43956_ (_19751_, _19740_, _18451_);
  not _43957_ (_19762_, _19751_);
  and _43958_ (_19773_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and _43959_ (_19783_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _43960_ (_19794_, _19783_, _19773_);
  and _43961_ (_19805_, _19794_, _19762_);
  nor _43962_ (_19816_, _19805_, _18681_);
  nor _43963_ (_19827_, _19816_, _19664_);
  nor _43964_ (_19838_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nor _43965_ (_19859_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _18494_);
  nor _43966_ (_19871_, _19859_, _19838_);
  nor _43967_ (_19883_, _19871_, _18473_);
  not _43968_ (_19895_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _43969_ (_19907_, _18473_, _19895_);
  nor _43970_ (_19919_, _19907_, _19883_);
  and _43971_ (_19931_, _19919_, _18451_);
  not _43972_ (_19932_, _19931_);
  and _43973_ (_19943_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  and _43974_ (_19953_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _43975_ (_19964_, _19953_, _19943_);
  and _43976_ (_19975_, _19964_, _19932_);
  nor _43977_ (_19986_, _19975_, _18331_);
  nor _43978_ (_19997_, _19986_, _18374_);
  and _43979_ (_20008_, _19997_, _19827_);
  nor _43980_ (_20019_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor _43981_ (_20030_, _18494_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor _43982_ (_20040_, _20030_, _20019_);
  nor _43983_ (_20051_, _20040_, _18473_);
  not _43984_ (_20062_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and _43985_ (_20073_, _18473_, _20062_);
  nor _43986_ (_20084_, _20073_, _20051_);
  and _43987_ (_20095_, _20084_, _18451_);
  not _43988_ (_20106_, _20095_);
  and _43989_ (_20116_, _18593_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _43990_ (_20127_, _18626_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _43991_ (_20138_, _20127_, _20116_);
  and _43992_ (_20149_, _20138_, _20106_);
  and _43993_ (_20160_, _20149_, _18374_);
  nor _43994_ (_20171_, _20160_, _20008_);
  and _43995_ (_20182_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _43996_ (_20193_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _43997_ (_20203_, _20193_, _20182_);
  and _43998_ (_20214_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _43999_ (_20225_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor _44000_ (_20236_, _20225_, _20214_);
  and _44001_ (_20247_, _20236_, _20203_);
  and _44002_ (_20258_, _20084_, _19370_);
  and _44003_ (_20269_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _44004_ (_20280_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor _44005_ (_20290_, _20280_, _20269_);
  not _44006_ (_20301_, _20290_);
  nor _44007_ (_20312_, _20301_, _20258_);
  and _44008_ (_20323_, _20312_, _20247_);
  not _44009_ (_20334_, _20323_);
  and _44010_ (_20345_, _20334_, _20171_);
  and _44011_ (_20356_, _20345_, _19512_);
  not _44012_ (_20366_, _20356_);
  and _44013_ (_20377_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _44014_ (_20388_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _44015_ (_20399_, _20388_, _20377_);
  and _44016_ (_20410_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  and _44017_ (_20421_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor _44018_ (_20432_, _20421_, _20410_);
  and _44019_ (_20443_, _20432_, _20399_);
  and _44020_ (_20453_, _19740_, _19370_);
  and _44021_ (_20464_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and _44022_ (_20475_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor _44023_ (_20486_, _20475_, _20464_);
  not _44024_ (_20497_, _20486_);
  nor _44025_ (_20508_, _20497_, _20453_);
  and _44026_ (_20519_, _20508_, _20443_);
  not _44027_ (_20530_, _20519_);
  and _44028_ (_20541_, _20530_, _20171_);
  and _44029_ (_20551_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _44030_ (_20562_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _44031_ (_20573_, _20562_, _20551_);
  and _44032_ (_20584_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and _44033_ (_20595_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor _44034_ (_20606_, _20595_, _20584_);
  and _44035_ (_20617_, _20606_, _20573_);
  and _44036_ (_20628_, _19370_, _18768_);
  and _44037_ (_20639_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _44038_ (_20649_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor _44039_ (_20660_, _20649_, _20639_);
  not _44040_ (_20671_, _20660_);
  nor _44041_ (_20682_, _20671_, _20628_);
  and _44042_ (_20693_, _20682_, _20617_);
  not _44043_ (_20704_, _20693_);
  and _44044_ (_20715_, _20704_, _19185_);
  and _44045_ (_20726_, _20541_, _20715_);
  and _44046_ (_20736_, _19490_, _20726_);
  nor _44047_ (_20747_, _19501_, _20726_);
  nor _44048_ (_20768_, _20747_, _20736_);
  and _44049_ (_20779_, _20768_, _20541_);
  and _44050_ (_20780_, _20345_, _19501_);
  and _44051_ (_20791_, _19490_, _20171_);
  and _44052_ (_20812_, _20334_, _19185_);
  nor _44053_ (_20823_, _20812_, _20791_);
  nor _44054_ (_20824_, _20823_, _20780_);
  and _44055_ (_20844_, _20824_, _20779_);
  nor _44056_ (_20855_, _20824_, _20779_);
  nor _44057_ (_20856_, _20855_, _20844_);
  and _44058_ (_20867_, _20856_, _20736_);
  nor _44059_ (_20878_, _20867_, _20844_);
  nor _44060_ (_20889_, _20878_, _20366_);
  and _44061_ (_20910_, _20171_, _20704_);
  and _44062_ (_20911_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _44063_ (_20921_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _44064_ (_20932_, _20921_, _20911_);
  and _44065_ (_20943_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and _44066_ (_20954_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [3]);
  nor _44067_ (_20965_, _20954_, _20943_);
  and _44068_ (_20976_, _20965_, _20932_);
  and _44069_ (_20987_, _19588_, _19370_);
  and _44070_ (_20998_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _44071_ (_21009_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  nor _44072_ (_21019_, _21009_, _20998_);
  not _44073_ (_21040_, _21019_);
  nor _44074_ (_21041_, _21040_, _20987_);
  and _44075_ (_21052_, _21041_, _20976_);
  not _44076_ (_21063_, _21052_);
  and _44077_ (_21074_, _21063_, _19185_);
  and _44078_ (_21085_, _21074_, _20910_);
  and _44079_ (_21096_, _20530_, _19185_);
  nor _44080_ (_21106_, _21096_, _20910_);
  nor _44081_ (_21117_, _21106_, _20726_);
  and _44082_ (_21128_, _21117_, _21085_);
  nor _44083_ (_21139_, _19501_, _20541_);
  nor _44084_ (_21150_, _21139_, _20779_);
  and _44085_ (_21161_, _21150_, _21128_);
  nor _44086_ (_21172_, _20856_, _20736_);
  nor _44087_ (_21183_, _21172_, _20867_);
  and _44088_ (_21194_, _21183_, _21161_);
  nor _44089_ (_21214_, _21183_, _21161_);
  nor _44090_ (_21215_, _21214_, _21194_);
  not _44091_ (_21226_, _21215_);
  and _44092_ (_21237_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _44093_ (_21248_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _44094_ (_21259_, _21248_, _21237_);
  and _44095_ (_21270_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [1]);
  and _44096_ (_21281_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nor _44097_ (_21291_, _21281_, _21270_);
  and _44098_ (_21302_, _21291_, _21259_);
  and _44099_ (_21313_, _19919_, _19370_);
  and _44100_ (_21324_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  and _44101_ (_21335_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _44102_ (_21346_, _21335_, _21324_);
  not _44103_ (_21357_, _21346_);
  nor _44104_ (_21368_, _21357_, _21313_);
  and _44105_ (_21379_, _21368_, _21302_);
  not _44106_ (_21389_, _21379_);
  and _44107_ (_21410_, _21389_, _20171_);
  and _44108_ (_21411_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _44109_ (_21422_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _44110_ (_21433_, _21422_, _21411_);
  and _44111_ (_21444_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [2]);
  and _44112_ (_21455_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nor _44113_ (_21466_, _21455_, _21444_);
  and _44114_ (_21476_, _21466_, _21433_);
  and _44115_ (_21487_, _19370_, _18560_);
  and _44116_ (_21498_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _44117_ (_21509_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nor _44118_ (_21520_, _21509_, _21498_);
  not _44119_ (_21531_, _21520_);
  nor _44120_ (_21542_, _21531_, _21487_);
  and _44121_ (_21553_, _21542_, _21476_);
  not _44122_ (_21564_, _21553_);
  and _44123_ (_21574_, _21564_, _19185_);
  and _44124_ (_21585_, _21574_, _21410_);
  and _44125_ (_21596_, _21389_, _19185_);
  not _44126_ (_21607_, _21596_);
  and _44127_ (_21618_, _21564_, _20171_);
  and _44128_ (_21629_, _21618_, _21607_);
  and _44129_ (_21640_, _21629_, _21074_);
  nor _44130_ (_21651_, _21640_, _21585_);
  and _44131_ (_21661_, _21063_, _20171_);
  nor _44132_ (_21672_, _21661_, _20715_);
  nor _44133_ (_21683_, _21672_, _21085_);
  not _44134_ (_21694_, _21683_);
  nor _44135_ (_21705_, _21694_, _21651_);
  nor _44136_ (_21716_, _21117_, _21085_);
  nor _44137_ (_21727_, _21716_, _21128_);
  and _44138_ (_21737_, _21727_, _21705_);
  nor _44139_ (_21758_, _21150_, _21128_);
  nor _44140_ (_21759_, _21758_, _21161_);
  and _44141_ (_21770_, _21759_, _21737_);
  and _44142_ (_21781_, _19218_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _44143_ (_21792_, _19251_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _44144_ (_21803_, _21792_, _21781_);
  and _44145_ (_21814_, _19294_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _44146_ (_21824_, _19327_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nor _44147_ (_21835_, _21824_, _21814_);
  and _44148_ (_21846_, _21835_, _21803_);
  and _44149_ (_21867_, _19370_, _18922_);
  and _44150_ (_21868_, _19425_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and _44151_ (_21879_, _19403_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _44152_ (_21890_, _21879_, _21868_);
  not _44153_ (_21901_, _21890_);
  nor _44154_ (_21911_, _21901_, _21867_);
  and _44155_ (_21922_, _21911_, _21846_);
  not _44156_ (_21933_, _21922_);
  and _44157_ (_21944_, _21933_, _20171_);
  and _44158_ (_21955_, _21944_, _21596_);
  nor _44159_ (_21966_, _21574_, _21410_);
  nor _44160_ (_21977_, _21966_, _21585_);
  and _44161_ (_21988_, _21977_, _21955_);
  nor _44162_ (_21998_, _21629_, _21074_);
  nor _44163_ (_22009_, _21998_, _21640_);
  and _44164_ (_22020_, _22009_, _21988_);
  and _44165_ (_22031_, _21694_, _21651_);
  nor _44166_ (_22042_, _22031_, _21705_);
  and _44167_ (_22053_, _22042_, _22020_);
  nor _44168_ (_22064_, _21727_, _21705_);
  nor _44169_ (_22075_, _22064_, _21737_);
  and _44170_ (_22085_, _22075_, _22053_);
  nor _44171_ (_22096_, _21759_, _21737_);
  nor _44172_ (_22107_, _22096_, _21770_);
  and _44173_ (_22118_, _22107_, _22085_);
  nor _44174_ (_22129_, _22118_, _21770_);
  nor _44175_ (_22140_, _22129_, _21226_);
  nor _44176_ (_22151_, _22140_, _21194_);
  and _44177_ (_22161_, _20878_, _20366_);
  nor _44178_ (_22172_, _22161_, _20889_);
  not _44179_ (_22183_, _22172_);
  nor _44180_ (_22194_, _22183_, _22151_);
  or _44181_ (_22205_, _22194_, _20780_);
  nor _44182_ (_22217_, _22205_, _20889_);
  nor _44183_ (_22228_, _22217_, _18429_);
  and _44184_ (_22239_, _22217_, _18429_);
  nor _44185_ (_22249_, _22239_, _22228_);
  not _44186_ (_22260_, _22249_);
  and _44187_ (_22271_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and _44188_ (_22282_, _22183_, _22151_);
  nor _44189_ (_22293_, _22282_, _22194_);
  and _44190_ (_22314_, _22293_, _22271_);
  and _44191_ (_22315_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  and _44192_ (_22325_, _22129_, _21226_);
  nor _44193_ (_22336_, _22325_, _22140_);
  and _44194_ (_22347_, _22336_, _22315_);
  nor _44195_ (_22358_, _22336_, _22315_);
  nor _44196_ (_22369_, _22358_, _22347_);
  not _44197_ (_22380_, _22369_);
  and _44198_ (_22391_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  nor _44199_ (_22402_, _22107_, _22085_);
  nor _44200_ (_22412_, _22402_, _22118_);
  and _44201_ (_22423_, _22412_, _22391_);
  nor _44202_ (_22434_, _22412_, _22391_);
  nor _44203_ (_22445_, _22434_, _22423_);
  and _44204_ (_22456_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  nor _44205_ (_22467_, _22075_, _22053_);
  nor _44206_ (_22478_, _22467_, _22085_);
  and _44207_ (_22489_, _22478_, _22456_);
  nor _44208_ (_22499_, _22478_, _22456_);
  nor _44209_ (_22510_, _22499_, _22489_);
  not _44210_ (_22521_, _22510_);
  and _44211_ (_22532_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  nor _44212_ (_22543_, _22042_, _22020_);
  nor _44213_ (_22554_, _22543_, _22053_);
  and _44214_ (_22565_, _22554_, _22532_);
  and _44215_ (_22576_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  nor _44216_ (_22586_, _22009_, _21988_);
  nor _44217_ (_22607_, _22586_, _22020_);
  and _44218_ (_22608_, _22607_, _22576_);
  and _44219_ (_22619_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nor _44220_ (_22630_, _21977_, _21955_);
  nor _44221_ (_22641_, _22630_, _21988_);
  and _44222_ (_22652_, _22641_, _22619_);
  nor _44223_ (_22662_, _22607_, _22576_);
  nor _44224_ (_22673_, _22662_, _22608_);
  and _44225_ (_22684_, _22673_, _22652_);
  nor _44226_ (_22695_, _22684_, _22608_);
  not _44227_ (_22716_, _22695_);
  nor _44228_ (_22717_, _22554_, _22532_);
  nor _44229_ (_22728_, _22717_, _22565_);
  and _44230_ (_22739_, _22728_, _22716_);
  nor _44231_ (_22749_, _22739_, _22565_);
  nor _44232_ (_22760_, _22749_, _22521_);
  nor _44233_ (_22771_, _22760_, _22489_);
  not _44234_ (_22782_, _22771_);
  and _44235_ (_22793_, _22782_, _22445_);
  nor _44236_ (_22804_, _22793_, _22423_);
  nor _44237_ (_22815_, _22804_, _22380_);
  nor _44238_ (_22826_, _22815_, _22347_);
  nor _44239_ (_22836_, _22293_, _22271_);
  nor _44240_ (_22847_, _22836_, _22314_);
  not _44241_ (_22858_, _22847_);
  nor _44242_ (_22869_, _22858_, _22826_);
  nor _44243_ (_22880_, _22869_, _22314_);
  nor _44244_ (_22891_, _22880_, _22260_);
  nor _44245_ (_22902_, _22891_, _22228_);
  not _44246_ (_22913_, _22902_);
  and _44247_ (_22933_, _22913_, _18407_);
  and _44248_ (_22934_, _22933_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _44249_ (_22945_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _44250_ (_22956_, _22945_, _22934_);
  and _44251_ (_22967_, _22956_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _44252_ (_22978_, _22967_, _18396_);
  not _44253_ (_22989_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nor _44254_ (_23000_, _18374_, _22989_);
  or _44255_ (_23011_, _23000_, _22978_);
  nand _44256_ (_23022_, _22978_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  and _44257_ (_23033_, _23022_, _23011_);
  and _44258_ (_24374_, _23033_, _42882_);
  nor _44259_ (_23053_, _18265_, _18298_);
  and _44260_ (_23064_, _18265_, _18298_);
  or _44261_ (_23075_, _23064_, _23053_);
  and _44262_ (_02356_, _23075_, _42882_);
  and _44263_ (_23096_, _21933_, _19185_);
  and _44264_ (_02542_, _23096_, _42882_);
  nor _44265_ (_23117_, _21944_, _21596_);
  nor _44266_ (_23128_, _23117_, _21955_);
  and _44267_ (_02695_, _23128_, _42882_);
  nor _44268_ (_23149_, _22641_, _22619_);
  nor _44269_ (_23159_, _23149_, _22652_);
  and _44270_ (_02877_, _23159_, _42882_);
  nor _44271_ (_23190_, _22673_, _22652_);
  nor _44272_ (_23191_, _23190_, _22684_);
  and _44273_ (_03117_, _23191_, _42882_);
  nor _44274_ (_23212_, _22728_, _22716_);
  nor _44275_ (_23223_, _23212_, _22739_);
  and _44276_ (_03361_, _23223_, _42882_);
  and _44277_ (_23244_, _22749_, _22521_);
  nor _44278_ (_23255_, _23244_, _22760_);
  and _44279_ (_03562_, _23255_, _42882_);
  nor _44280_ (_23275_, _22782_, _22445_);
  nor _44281_ (_23286_, _23275_, _22793_);
  and _44282_ (_03757_, _23286_, _42882_);
  and _44283_ (_23307_, _22804_, _22380_);
  nor _44284_ (_23318_, _23307_, _22815_);
  and _44285_ (_03954_, _23318_, _42882_);
  and _44286_ (_23339_, _22858_, _22826_);
  nor _44287_ (_23350_, _23339_, _22869_);
  and _44288_ (_04054_, _23350_, _42882_);
  and _44289_ (_23370_, _22880_, _22260_);
  nor _44290_ (_23381_, _23370_, _22891_);
  and _44291_ (_04147_, _23381_, _42882_);
  nor _44292_ (_23402_, _22913_, _18407_);
  nor _44293_ (_23413_, _23402_, _22933_);
  and _44294_ (_04246_, _23413_, _42882_);
  and _44295_ (_23434_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  nor _44296_ (_23445_, _23434_, _22933_);
  nor _44297_ (_23466_, _23445_, _22934_);
  and _44298_ (_04345_, _23466_, _42882_);
  nor _44299_ (_23476_, _22945_, _22934_);
  nor _44300_ (_23487_, _23476_, _22956_);
  and _44301_ (_04444_, _23487_, _42882_);
  and _44302_ (_23508_, _18385_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  nor _44303_ (_23519_, _23508_, _22956_);
  nor _44304_ (_23530_, _23519_, _22967_);
  and _44305_ (_04542_, _23530_, _42882_);
  nor _44306_ (_23551_, _22967_, _18396_);
  nor _44307_ (_23562_, _23551_, _22978_);
  and _44308_ (_04641_, _23562_, _42882_);
  and _44309_ (_23582_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _18199_);
  nor _44310_ (_23593_, _23582_, _18210_);
  not _44311_ (_23604_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _44312_ (_23615_, _18232_, _23604_);
  and _44313_ (_23626_, _23615_, _23593_);
  and _44314_ (_23637_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _44315_ (_23648_, _23637_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _44316_ (_23658_, _23637_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44317_ (_23669_, _23658_, _23648_);
  and _44318_ (_00925_, _23669_, _42882_);
  and _44319_ (_00956_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _42882_);
  not _44320_ (_23700_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _44321_ (_23711_, _19975_, _23700_);
  and _44322_ (_23722_, _19653_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44323_ (_23733_, _23722_, _23711_);
  nor _44324_ (_23743_, _23733_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44325_ (_23754_, _19805_, _23700_);
  and _44326_ (_23765_, _20149_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _44327_ (_23776_, _23765_, _23754_);
  and _44328_ (_23787_, _23776_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _44329_ (_23798_, _23787_, _23743_);
  nor _44330_ (_23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44331_ (_23820_, _23809_, _20323_);
  nor _44332_ (_23830_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  nor _44333_ (_23841_, _23830_, _23820_);
  not _44334_ (_23852_, _23841_);
  and _44335_ (_23863_, _18988_, _23700_);
  and _44336_ (_23874_, _18669_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44337_ (_23895_, _23874_, _23863_);
  nor _44338_ (_23896_, _23895_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44339_ (_23907_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44340_ (_23917_, _18834_, _23700_);
  and _44341_ (_23928_, _19164_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44342_ (_23939_, _23928_, _23917_);
  nor _44343_ (_23950_, _23939_, _23907_);
  nor _44344_ (_23961_, _23950_, _23896_);
  nor _44345_ (_23972_, _23961_, _23852_);
  and _44346_ (_23983_, _23961_, _23852_);
  nor _44347_ (_23994_, _23983_, _23972_);
  and _44348_ (_24004_, _23809_, _19479_);
  nor _44349_ (_24015_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  nor _44350_ (_24026_, _24015_, _24004_);
  not _44351_ (_24037_, _24026_);
  nor _44352_ (_24048_, _19975_, _23700_);
  nor _44353_ (_24059_, _24048_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44354_ (_24079_, _19653_, _23700_);
  and _44355_ (_24080_, _19805_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44356_ (_24091_, _24080_, _24079_);
  nor _44357_ (_24102_, _24091_, _23907_);
  nor _44358_ (_24113_, _24102_, _24059_);
  nor _44359_ (_24124_, _24113_, _24037_);
  and _44360_ (_24135_, _24113_, _24037_);
  nor _44361_ (_24146_, _24135_, _24124_);
  not _44362_ (_24157_, _24146_);
  and _44363_ (_24167_, _23809_, _20519_);
  nor _44364_ (_24178_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  nor _44365_ (_24189_, _24178_, _24167_);
  not _44366_ (_24200_, _24189_);
  nor _44367_ (_24211_, _18988_, _23700_);
  nor _44368_ (_24222_, _24211_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44369_ (_24233_, _18669_, _23700_);
  and _44370_ (_24243_, _18834_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44371_ (_24254_, _24243_, _24233_);
  nor _44372_ (_24265_, _24254_, _23907_);
  nor _44373_ (_24276_, _24265_, _24222_);
  nor _44374_ (_24287_, _24276_, _24200_);
  and _44375_ (_24298_, _24276_, _24200_);
  and _44376_ (_24309_, _23733_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44377_ (_24320_, _24309_);
  nor _44378_ (_24330_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  and _44379_ (_24341_, _23809_, _20693_);
  nor _44380_ (_24352_, _24341_, _24330_);
  and _44381_ (_24363_, _24352_, _24320_);
  and _44382_ (_24375_, _23895_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44383_ (_24386_, _24375_);
  and _44384_ (_24397_, _23809_, _21052_);
  nor _44385_ (_24408_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  nor _44386_ (_24418_, _24408_, _24397_);
  and _44387_ (_24429_, _24418_, _24386_);
  nor _44388_ (_24440_, _24418_, _24386_);
  nor _44389_ (_24451_, _24440_, _24429_);
  not _44390_ (_24462_, _24451_);
  and _44391_ (_24473_, _24048_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44392_ (_24484_, _24473_);
  and _44393_ (_24495_, _23809_, _21553_);
  nor _44394_ (_24505_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  nor _44395_ (_24516_, _24505_, _24495_);
  and _44396_ (_24527_, _24516_, _24484_);
  and _44397_ (_24538_, _24211_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _44398_ (_24549_, _24538_);
  nor _44399_ (_24560_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  and _44400_ (_24571_, _23809_, _21379_);
  nor _44401_ (_24581_, _24571_, _24560_);
  nor _44402_ (_24592_, _24581_, _24549_);
  not _44403_ (_24613_, _24592_);
  nor _44404_ (_24614_, _24516_, _24484_);
  nor _44405_ (_24625_, _24614_, _24527_);
  and _44406_ (_24636_, _24625_, _24613_);
  nor _44407_ (_24647_, _24636_, _24527_);
  nor _44408_ (_24658_, _24647_, _24462_);
  nor _44409_ (_24668_, _24658_, _24429_);
  nor _44410_ (_24679_, _24352_, _24320_);
  nor _44411_ (_24690_, _24679_, _24363_);
  not _44412_ (_24701_, _24690_);
  nor _44413_ (_24712_, _24701_, _24668_);
  nor _44414_ (_24723_, _24712_, _24363_);
  nor _44415_ (_24734_, _24723_, _24298_);
  nor _44416_ (_24745_, _24734_, _24287_);
  nor _44417_ (_24755_, _24745_, _24157_);
  nor _44418_ (_24766_, _24755_, _24124_);
  not _44419_ (_24777_, _24766_);
  and _44420_ (_24788_, _24777_, _23994_);
  or _44421_ (_24799_, _24788_, _23972_);
  and _44422_ (_24810_, _20149_, _19164_);
  or _44423_ (_24821_, _24810_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _44424_ (_24832_, _23939_);
  and _44425_ (_24843_, _23776_, _24832_);
  nor _44426_ (_24854_, _24254_, _24091_);
  and _44427_ (_24865_, _24854_, _24843_);
  or _44428_ (_24876_, _24865_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _44429_ (_24887_, _24876_, _24821_);
  and _44430_ (_24898_, _24887_, _24799_);
  and _44431_ (_24909_, _24898_, _23798_);
  nor _44432_ (_24920_, _24777_, _23994_);
  or _44433_ (_24931_, _24920_, _24788_);
  and _44434_ (_24942_, _24931_, _24909_);
  nor _44435_ (_24953_, _24909_, _23841_);
  nor _44436_ (_24964_, _24953_, _24942_);
  not _44437_ (_24975_, _24964_);
  and _44438_ (_24986_, _24964_, _23798_);
  not _44439_ (_24997_, _23961_);
  nor _44440_ (_25008_, _24909_, _24037_);
  and _44441_ (_25018_, _24745_, _24157_);
  nor _44442_ (_25029_, _25018_, _24755_);
  and _44443_ (_25040_, _25029_, _24909_);
  or _44444_ (_25051_, _25040_, _25008_);
  and _44445_ (_25062_, _25051_, _24997_);
  nor _44446_ (_25073_, _25051_, _24997_);
  nor _44447_ (_25084_, _25073_, _25062_);
  not _44448_ (_25095_, _25084_);
  not _44449_ (_25106_, _24113_);
  nor _44450_ (_25117_, _24909_, _24200_);
  nor _44451_ (_25128_, _24298_, _24287_);
  nor _44452_ (_25139_, _25128_, _24723_);
  and _44453_ (_25160_, _25128_, _24723_);
  or _44454_ (_25161_, _25160_, _25139_);
  and _44455_ (_25172_, _25161_, _24909_);
  or _44456_ (_25183_, _25172_, _25117_);
  and _44457_ (_25194_, _25183_, _25106_);
  nor _44458_ (_25205_, _25183_, _25106_);
  not _44459_ (_25216_, _24276_);
  and _44460_ (_25227_, _24701_, _24668_);
  or _44461_ (_25238_, _25227_, _24712_);
  and _44462_ (_25249_, _25238_, _24909_);
  nor _44463_ (_25260_, _24909_, _24352_);
  nor _44464_ (_25271_, _25260_, _25249_);
  and _44465_ (_25282_, _25271_, _25216_);
  and _44466_ (_25293_, _24647_, _24462_);
  nor _44467_ (_25304_, _25293_, _24658_);
  not _44468_ (_25315_, _25304_);
  and _44469_ (_25326_, _25315_, _24909_);
  nor _44470_ (_25337_, _24909_, _24418_);
  nor _44471_ (_25348_, _25337_, _25326_);
  and _44472_ (_25359_, _25348_, _24320_);
  nor _44473_ (_25370_, _25348_, _24320_);
  nor _44474_ (_25381_, _25370_, _25359_);
  not _44475_ (_25391_, _25381_);
  nor _44476_ (_25402_, _24625_, _24613_);
  nor _44477_ (_25423_, _25402_, _24636_);
  not _44478_ (_25424_, _25423_);
  and _44479_ (_25435_, _25424_, _24909_);
  nor _44480_ (_25446_, _24909_, _24516_);
  nor _44481_ (_25457_, _25446_, _25435_);
  and _44482_ (_25468_, _25457_, _24386_);
  not _44483_ (_25479_, _24581_);
  and _44484_ (_25490_, _24909_, _24538_);
  or _44485_ (_25501_, _25490_, _25479_);
  nand _44486_ (_25512_, _24909_, _24538_);
  or _44487_ (_25523_, _25512_, _24581_);
  and _44488_ (_25534_, _25523_, _25501_);
  nor _44489_ (_25545_, _25534_, _24473_);
  and _44490_ (_25556_, _25534_, _24473_);
  nor _44491_ (_25567_, _25556_, _25545_);
  and _44492_ (_25578_, _23809_, _21922_);
  nor _44493_ (_25589_, _23809_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor _44494_ (_25600_, _25589_, _25578_);
  nor _44495_ (_25611_, _25600_, _24549_);
  not _44496_ (_25622_, _25611_);
  and _44497_ (_25633_, _25622_, _25567_);
  nor _44498_ (_25644_, _25633_, _25545_);
  nor _44499_ (_25655_, _25457_, _24386_);
  nor _44500_ (_25666_, _25655_, _25468_);
  not _44501_ (_25677_, _25666_);
  nor _44502_ (_25688_, _25677_, _25644_);
  nor _44503_ (_25699_, _25688_, _25468_);
  nor _44504_ (_25710_, _25699_, _25391_);
  nor _44505_ (_25731_, _25710_, _25359_);
  nor _44506_ (_25732_, _25271_, _25216_);
  nor _44507_ (_25742_, _25732_, _25282_);
  not _44508_ (_25753_, _25742_);
  nor _44509_ (_25764_, _25753_, _25731_);
  nor _44510_ (_25775_, _25764_, _25282_);
  nor _44511_ (_25786_, _25775_, _25205_);
  nor _44512_ (_25797_, _25786_, _25194_);
  nor _44513_ (_25808_, _25797_, _25095_);
  or _44514_ (_25819_, _25808_, _25062_);
  or _44515_ (_25830_, _25819_, _24986_);
  and _44516_ (_25841_, _25830_, _24887_);
  nor _44517_ (_25852_, _25841_, _24975_);
  and _44518_ (_25863_, _24986_, _24887_);
  and _44519_ (_25874_, _25863_, _25819_);
  or _44520_ (_25885_, _25874_, _25852_);
  and _44521_ (_00976_, _25885_, _42882_);
  or _44522_ (_25906_, _24964_, _23798_);
  and _44523_ (_25917_, _25906_, _25841_);
  and _44524_ (_02832_, _25917_, _42882_);
  and _44525_ (_02844_, _24909_, _42882_);
  and _44526_ (_02866_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _42882_);
  and _44527_ (_02890_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _42882_);
  and _44528_ (_02914_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _42882_);
  or _44529_ (_25978_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _44530_ (_25989_, _23637_, rst);
  and _44531_ (_02924_, _25989_, _25978_);
  not _44532_ (_26010_, _25600_);
  and _44533_ (_26021_, _25917_, _24538_);
  nor _44534_ (_26032_, _26021_, _26010_);
  and _44535_ (_26053_, _26021_, _26010_);
  or _44536_ (_26054_, _26053_, _26032_);
  and _44537_ (_02936_, _26054_, _42882_);
  nor _44538_ (_26074_, _25917_, _25534_);
  nor _44539_ (_26085_, _25622_, _25567_);
  nor _44540_ (_26096_, _26085_, _25633_);
  and _44541_ (_26107_, _26096_, _25917_);
  or _44542_ (_26118_, _26107_, _26074_);
  and _44543_ (_02948_, _26118_, _42882_);
  and _44544_ (_26139_, _25677_, _25644_);
  or _44545_ (_26150_, _26139_, _25688_);
  nand _44546_ (_26161_, _26150_, _25917_);
  or _44547_ (_26172_, _25917_, _25457_);
  and _44548_ (_26183_, _26172_, _26161_);
  and _44549_ (_02960_, _26183_, _42882_);
  and _44550_ (_26204_, _25699_, _25391_);
  or _44551_ (_26215_, _26204_, _25710_);
  nand _44552_ (_26226_, _26215_, _25917_);
  or _44553_ (_26237_, _25917_, _25348_);
  and _44554_ (_26248_, _26237_, _26226_);
  and _44555_ (_02971_, _26248_, _42882_);
  and _44556_ (_26269_, _25753_, _25731_);
  or _44557_ (_26280_, _26269_, _25764_);
  nand _44558_ (_26291_, _26280_, _25917_);
  or _44559_ (_26302_, _25917_, _25271_);
  and _44560_ (_26313_, _26302_, _26291_);
  and _44561_ (_02984_, _26313_, _42882_);
  or _44562_ (_26334_, _25205_, _25194_);
  and _44563_ (_26345_, _26334_, _25775_);
  nor _44564_ (_26356_, _26334_, _25775_);
  or _44565_ (_26367_, _26356_, _26345_);
  nand _44566_ (_26378_, _26367_, _25917_);
  or _44567_ (_26389_, _25917_, _25183_);
  and _44568_ (_26400_, _26389_, _26378_);
  and _44569_ (_02997_, _26400_, _42882_);
  and _44570_ (_26420_, _25797_, _25095_);
  or _44571_ (_26431_, _26420_, _25808_);
  nand _44572_ (_26442_, _26431_, _25917_);
  or _44573_ (_26453_, _25917_, _25051_);
  and _44574_ (_26464_, _26453_, _26442_);
  and _44575_ (_03011_, _26464_, _42882_);
  not _44576_ (_26485_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44577_ (_26496_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _18199_);
  and _44578_ (_26507_, _26496_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _44579_ (_26528_, _26507_, _26485_);
  and _44580_ (_26529_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _44581_ (_26540_, _26529_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _44582_ (_26551_, _26529_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _44583_ (_26562_, _26551_, _26540_);
  and _44584_ (_26573_, _26562_, _26528_);
  not _44585_ (_26584_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _44586_ (_26595_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _18199_);
  and _44587_ (_26606_, _26595_, _26485_);
  and _44588_ (_26617_, _26606_, _26584_);
  and _44589_ (_26628_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _44590_ (_26639_, _26628_, _26573_);
  not _44591_ (_26650_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and _44592_ (_26661_, _26496_, _26650_);
  and _44593_ (_26672_, _26661_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44594_ (_26683_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _44595_ (_26694_, _26661_, _26485_);
  and _44596_ (_26705_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  or _44597_ (_26716_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44598_ (_26727_, _26716_, _18199_);
  nor _44599_ (_26738_, _26727_, _26496_);
  and _44600_ (_26759_, _26738_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _44601_ (_26760_, _26759_, _26705_);
  nor _44602_ (_26771_, _26760_, _26683_);
  and _44603_ (_26781_, _26771_, _26639_);
  and _44604_ (_26792_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor _44605_ (_26803_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _44606_ (_26814_, _26803_, _26529_);
  and _44607_ (_26825_, _26814_, _26528_);
  nor _44608_ (_26836_, _26825_, _26792_);
  and _44609_ (_26847_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and _44610_ (_26858_, _26738_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and _44611_ (_26869_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or _44612_ (_26880_, _26869_, _26858_);
  nor _44613_ (_26891_, _26880_, _26847_);
  and _44614_ (_26902_, _26891_, _26836_);
  and _44615_ (_26913_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and _44616_ (_26924_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _44617_ (_26935_, _26924_, _26913_);
  and _44618_ (_26946_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not _44619_ (_26957_, _26946_);
  not _44620_ (_26968_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _44621_ (_26979_, _26528_, _26968_);
  and _44622_ (_26990_, _26738_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _44623_ (_27001_, _26990_, _26979_);
  and _44624_ (_27012_, _27001_, _26957_);
  and _44625_ (_27023_, _27012_, _26935_);
  and _44626_ (_27034_, _27023_, _26902_);
  and _44627_ (_27045_, _27034_, _26781_);
  and _44628_ (_27056_, _26540_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _44629_ (_27067_, _27056_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and _44630_ (_27078_, _27067_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _44631_ (_27089_, _27078_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _44632_ (_27100_, _27089_);
  not _44633_ (_27111_, _26528_);
  nor _44634_ (_27122_, _27078_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _44635_ (_27132_, _27122_, _27111_);
  and _44636_ (_27143_, _27132_, _27100_);
  not _44637_ (_27154_, _27143_);
  and _44638_ (_27165_, _26507_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _44639_ (_27176_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nor _44640_ (_27187_, _27176_, _27165_);
  and _44641_ (_27198_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _44642_ (_27209_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nor _44643_ (_27220_, _27209_, _27198_);
  and _44644_ (_27231_, _27220_, _27187_);
  and _44645_ (_27242_, _27231_, _27154_);
  nor _44646_ (_27253_, _27067_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not _44647_ (_27264_, _27253_);
  nor _44648_ (_27275_, _27078_, _27111_);
  and _44649_ (_27286_, _27275_, _27264_);
  not _44650_ (_27297_, _27286_);
  and _44651_ (_27308_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nor _44652_ (_27319_, _27308_, _27165_);
  and _44653_ (_27340_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and _44654_ (_27341_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor _44655_ (_27352_, _27341_, _27340_);
  and _44656_ (_27363_, _27352_, _27319_);
  and _44657_ (_27374_, _27363_, _27297_);
  nor _44658_ (_27385_, _27374_, _27242_);
  not _44659_ (_27396_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _44660_ (_27407_, _27089_, _27396_);
  and _44661_ (_27418_, _27089_, _27396_);
  nor _44662_ (_27429_, _27418_, _27407_);
  nor _44663_ (_27440_, _27429_, _27111_);
  not _44664_ (_27451_, _27440_);
  and _44665_ (_27462_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  not _44666_ (_27473_, _27462_);
  not _44667_ (_27483_, _27165_);
  and _44668_ (_27494_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  and _44669_ (_27505_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [7]);
  nor _44670_ (_27516_, _27505_, _27494_);
  and _44671_ (_27527_, _27516_, _27483_);
  and _44672_ (_27538_, _27527_, _27473_);
  and _44673_ (_27549_, _27538_, _27451_);
  not _44674_ (_27560_, _27549_);
  and _44675_ (_27571_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _44676_ (_27582_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor _44677_ (_27593_, _27582_, _27571_);
  not _44678_ (_27604_, _27056_);
  nor _44679_ (_27615_, _26540_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _44680_ (_27626_, _27615_, _27111_);
  and _44681_ (_27637_, _27626_, _27604_);
  and _44682_ (_27648_, _26738_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and _44683_ (_27659_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _44684_ (_27670_, _27659_, _27648_);
  not _44685_ (_27681_, _27670_);
  nor _44686_ (_27692_, _27681_, _27637_);
  and _44687_ (_27703_, _27692_, _27593_);
  not _44688_ (_27714_, _27703_);
  and _44689_ (_27725_, _26672_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nor _44690_ (_27736_, _27725_, _27165_);
  nor _44691_ (_27747_, _27056_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  or _44692_ (_27758_, _27747_, _27111_);
  nor _44693_ (_27769_, _27758_, _27067_);
  and _44694_ (_27780_, _26694_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor _44695_ (_27791_, _27780_, _27769_);
  and _44696_ (_27801_, _27791_, _27736_);
  and _44697_ (_27812_, _26738_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  and _44698_ (_27823_, _26617_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor _44699_ (_27834_, _27823_, _27812_);
  and _44700_ (_27845_, _27834_, _27801_);
  nor _44701_ (_27856_, _27845_, _27714_);
  and _44702_ (_27867_, _27856_, _27560_);
  and _44703_ (_27878_, _27867_, _27385_);
  nand _44704_ (_27889_, _27878_, _27045_);
  and _44705_ (_27900_, _25885_, _23626_);
  not _44706_ (_27911_, _27900_);
  and _44707_ (_27922_, _23033_, _18265_);
  not _44708_ (_27933_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _44709_ (_27944_, _18210_, _27933_);
  and _44710_ (_27955_, _27944_, _18254_);
  not _44711_ (_27976_, _27955_);
  nor _44712_ (_27977_, _20323_, _20149_);
  and _44713_ (_27988_, _20323_, _20149_);
  nor _44714_ (_27999_, _27988_, _27977_);
  not _44715_ (_28010_, _19164_);
  nor _44716_ (_28021_, _19479_, _28010_);
  nor _44717_ (_28032_, _19479_, _19164_);
  and _44718_ (_28043_, _19479_, _19164_);
  nor _44719_ (_28054_, _28043_, _28032_);
  not _44720_ (_28065_, _19805_);
  nor _44721_ (_28076_, _20519_, _28065_);
  nor _44722_ (_28087_, _20519_, _19805_);
  and _44723_ (_28098_, _20519_, _19805_);
  nor _44724_ (_28109_, _28098_, _28087_);
  not _44725_ (_28120_, _18834_);
  and _44726_ (_28130_, _20693_, _28120_);
  nor _44727_ (_28141_, _28130_, _28109_);
  nor _44728_ (_28152_, _28141_, _28076_);
  nor _44729_ (_28163_, _28152_, _28054_);
  nor _44730_ (_28174_, _28163_, _28021_);
  and _44731_ (_28185_, _28152_, _28054_);
  nor _44732_ (_28196_, _28185_, _28163_);
  not _44733_ (_28207_, _28196_);
  and _44734_ (_28218_, _28130_, _28109_);
  nor _44735_ (_28229_, _28218_, _28141_);
  not _44736_ (_28240_, _28229_);
  nor _44737_ (_28251_, _20693_, _18834_);
  and _44738_ (_28262_, _20693_, _18834_);
  nor _44739_ (_28283_, _28262_, _28251_);
  not _44740_ (_28284_, _28283_);
  and _44741_ (_28295_, _21052_, _19653_);
  nor _44742_ (_28306_, _21052_, _19653_);
  nor _44743_ (_28317_, _28306_, _28295_);
  not _44744_ (_28328_, _28317_);
  nor _44745_ (_28339_, _21553_, _18669_);
  and _44746_ (_28350_, _21553_, _18669_);
  nor _44747_ (_28361_, _28350_, _28339_);
  nor _44748_ (_28372_, _21379_, _19975_);
  and _44749_ (_28383_, _21379_, _19975_);
  nor _44750_ (_28394_, _28383_, _28372_);
  not _44751_ (_28405_, _18988_);
  and _44752_ (_28416_, _21922_, _28405_);
  nor _44753_ (_28427_, _28416_, _28394_);
  not _44754_ (_28437_, _19975_);
  nor _44755_ (_28448_, _21379_, _28437_);
  nor _44756_ (_28459_, _28448_, _28427_);
  nor _44757_ (_28470_, _28459_, _28361_);
  not _44758_ (_28481_, _18669_);
  nor _44759_ (_28492_, _21553_, _28481_);
  nor _44760_ (_28503_, _28492_, _28470_);
  nor _44761_ (_28514_, _28503_, _28328_);
  and _44762_ (_28525_, _28503_, _28328_);
  nor _44763_ (_28536_, _28525_, _28514_);
  and _44764_ (_28547_, _28459_, _28361_);
  nor _44765_ (_28558_, _28547_, _28470_);
  not _44766_ (_28569_, _28558_);
  nor _44767_ (_28580_, _21922_, _18988_);
  and _44768_ (_28591_, _21922_, _18988_);
  nor _44769_ (_28602_, _28591_, _28580_);
  not _44770_ (_28613_, \oc8051_top_1.oc8051_sfr1.bit_out );
  and _44771_ (_28634_, _18473_, _28613_);
  not _44772_ (_28635_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not _44773_ (_28646_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44774_ (_28657_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _28646_);
  and _44775_ (_28668_, _28657_, _19696_);
  nor _44776_ (_28679_, _28668_, _28635_);
  nor _44777_ (_28690_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44778_ (_28701_, _28690_, _18714_);
  not _44779_ (_28712_, _28701_);
  and _44780_ (_28723_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44781_ (_28733_, _28723_, _20040_);
  not _44782_ (_28744_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  and _44783_ (_28755_, _28744_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  and _44784_ (_28766_, _28755_, _19054_);
  nor _44785_ (_28777_, _28766_, _28733_);
  and _44786_ (_28788_, _28777_, _28712_);
  and _44787_ (_28799_, _28788_, _28679_);
  and _44788_ (_28810_, _28657_, _19871_);
  nor _44789_ (_28821_, _28810_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _44790_ (_28832_, _28755_, _18516_);
  not _44791_ (_28843_, _28832_);
  and _44792_ (_28854_, _28723_, _19544_);
  and _44793_ (_28865_, _28690_, _18878_);
  nor _44794_ (_28876_, _28865_, _28854_);
  and _44795_ (_28887_, _28876_, _28843_);
  and _44796_ (_28898_, _28887_, _28821_);
  nor _44797_ (_28909_, _28898_, _28799_);
  nor _44798_ (_28920_, _28909_, _18473_);
  nor _44799_ (_28931_, _28920_, _28634_);
  and _44800_ (_28942_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _44801_ (_28953_, _28942_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not _44802_ (_28964_, _28953_);
  and _44803_ (_28975_, _28964_, _28931_);
  and _44804_ (_28986_, _28964_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _44805_ (_29007_, _28986_, _28975_);
  nor _44806_ (_29008_, _29007_, _28602_);
  and _44807_ (_29019_, _28416_, _28394_);
  nor _44808_ (_29030_, _29019_, _28427_);
  not _44809_ (_29040_, _29030_);
  and _44810_ (_29051_, _29040_, _29008_);
  and _44811_ (_29062_, _29051_, _28569_);
  and _44812_ (_29073_, _29062_, _28536_);
  not _44813_ (_29084_, _19653_);
  or _44814_ (_29095_, _21052_, _29084_);
  and _44815_ (_29106_, _21052_, _29084_);
  or _44816_ (_29117_, _28503_, _29106_);
  and _44817_ (_29128_, _29117_, _29095_);
  or _44818_ (_29139_, _29128_, _29073_);
  and _44819_ (_29150_, _29139_, _28284_);
  and _44820_ (_29161_, _29150_, _28240_);
  and _44821_ (_29172_, _29161_, _28207_);
  nor _44822_ (_29183_, _29172_, _28174_);
  nor _44823_ (_29194_, _29183_, _27999_);
  and _44824_ (_29205_, _29183_, _27999_);
  nor _44825_ (_29216_, _29205_, _29194_);
  nor _44826_ (_29227_, _29216_, _27976_);
  not _44827_ (_29238_, _29227_);
  not _44828_ (_29249_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _44829_ (_29260_, _23582_, _29249_);
  and _44830_ (_29271_, _29260_, _18254_);
  not _44831_ (_29282_, _27999_);
  not _44832_ (_29293_, _28054_);
  and _44833_ (_29304_, _28251_, _28109_);
  nor _44834_ (_29315_, _29304_, _28087_);
  nor _44835_ (_29326_, _29315_, _29293_);
  not _44836_ (_29337_, _28361_);
  and _44837_ (_29347_, _28580_, _28394_);
  nor _44838_ (_29358_, _29347_, _28372_);
  nor _44839_ (_29369_, _29358_, _29337_);
  nor _44840_ (_29380_, _29369_, _28339_);
  nor _44841_ (_29391_, _29380_, _28317_);
  and _44842_ (_29402_, _29380_, _28317_);
  nor _44843_ (_29413_, _29402_, _29391_);
  not _44844_ (_29424_, _28602_);
  nor _44845_ (_29435_, _29007_, _29424_);
  and _44846_ (_29446_, _29435_, _28394_);
  and _44847_ (_29457_, _29358_, _29337_);
  nor _44848_ (_29468_, _29457_, _29369_);
  and _44849_ (_29479_, _29468_, _29446_);
  not _44850_ (_29490_, _29479_);
  nor _44851_ (_29501_, _29490_, _29413_);
  nor _44852_ (_29512_, _29380_, _28295_);
  or _44853_ (_29533_, _29512_, _28306_);
  or _44854_ (_29534_, _29533_, _29501_);
  and _44855_ (_29545_, _29534_, _28283_);
  nor _44856_ (_29556_, _28251_, _28109_);
  nor _44857_ (_29567_, _29556_, _29304_);
  and _44858_ (_29578_, _29567_, _29545_);
  and _44859_ (_29589_, _29315_, _29293_);
  nor _44860_ (_29600_, _29589_, _29326_);
  and _44861_ (_29611_, _29600_, _29578_);
  or _44862_ (_29622_, _29611_, _29326_);
  nor _44863_ (_29633_, _29622_, _28032_);
  nor _44864_ (_29644_, _29633_, _29282_);
  and _44865_ (_29654_, _29633_, _29282_);
  nor _44866_ (_29665_, _29654_, _29644_);
  and _44867_ (_29676_, _29665_, _29271_);
  and _44868_ (_29687_, _18243_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _44869_ (_29698_, _29687_, _27944_);
  nor _44870_ (_29709_, _21922_, _21379_);
  and _44871_ (_29720_, _29709_, _21564_);
  and _44872_ (_29731_, _29720_, _21063_);
  and _44873_ (_29742_, _29731_, _20704_);
  and _44874_ (_29753_, _29742_, _20530_);
  and _44875_ (_29763_, _29753_, _19490_);
  and _44876_ (_29774_, _29763_, _29007_);
  not _44877_ (_29785_, _29007_);
  and _44878_ (_29806_, _19479_, _20519_);
  and _44879_ (_29807_, _21553_, _21379_);
  and _44880_ (_29818_, _29807_, _21922_);
  and _44881_ (_29829_, _29818_, _21052_);
  and _44882_ (_29840_, _29829_, _20693_);
  and _44883_ (_29851_, _29840_, _29806_);
  and _44884_ (_29862_, _29851_, _29785_);
  nor _44885_ (_29872_, _29862_, _29774_);
  and _44886_ (_29883_, _29872_, _20323_);
  nor _44887_ (_29894_, _29872_, _20323_);
  nor _44888_ (_29905_, _29894_, _29883_);
  and _44889_ (_29916_, _29905_, _29698_);
  not _44890_ (_29927_, _20149_);
  nor _44891_ (_29938_, _29007_, _29927_);
  not _44892_ (_29949_, _29938_);
  and _44893_ (_29960_, _29007_, _20323_);
  and _44894_ (_29971_, _29687_, _18221_);
  not _44895_ (_29981_, _29971_);
  nor _44896_ (_29992_, _29981_, _29960_);
  and _44897_ (_30003_, _29992_, _29949_);
  nor _44898_ (_30014_, _30003_, _29916_);
  and _44899_ (_30025_, _29260_, _23615_);
  not _44900_ (_30036_, _30025_);
  nor _44901_ (_30047_, _29807_, _21052_);
  and _44902_ (_30058_, _30047_, _30025_);
  and _44903_ (_30069_, _30058_, _20704_);
  not _44904_ (_30080_, _30069_);
  and _44905_ (_30090_, _30080_, _29806_);
  nor _44906_ (_30101_, _29806_, _20323_);
  nor _44907_ (_30112_, _30101_, _30058_);
  and _44908_ (_30123_, _30112_, _29007_);
  nor _44909_ (_30134_, _30123_, _30090_);
  and _44910_ (_30145_, _30134_, _20323_);
  nor _44911_ (_30156_, _30134_, _20323_);
  nor _44912_ (_30167_, _30156_, _30145_);
  nor _44913_ (_30178_, _30167_, _30036_);
  and _44914_ (_30189_, _29687_, _29260_);
  not _44915_ (_30199_, _30189_);
  nor _44916_ (_30210_, _30199_, _29007_);
  not _44917_ (_30221_, _30210_);
  not _44918_ (_30232_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _44919_ (_30243_, _18243_, _30232_);
  and _44920_ (_30254_, _30243_, _29260_);
  not _44921_ (_30265_, _30254_);
  nor _44922_ (_30276_, _30265_, _27988_);
  and _44923_ (_30287_, _30243_, _23593_);
  and _44924_ (_30298_, _30287_, _27999_);
  nor _44925_ (_30308_, _30298_, _30276_);
  and _44926_ (_30319_, _23615_, _18221_);
  and _44927_ (_30330_, _30319_, _27977_);
  and _44928_ (_30341_, _27944_, _23615_);
  and _44929_ (_30352_, _30341_, _20323_);
  nor _44930_ (_30363_, _30352_, _30330_);
  and _44931_ (_30374_, _23593_, _18254_);
  not _44932_ (_30385_, _30374_);
  nor _44933_ (_30396_, _30385_, _20323_);
  and _44934_ (_30407_, _29687_, _23593_);
  and _44935_ (_30427_, _30407_, _21933_);
  and _44936_ (_30428_, _30243_, _18210_);
  not _44937_ (_30439_, _30428_);
  nor _44938_ (_30450_, _30439_, _19479_);
  or _44939_ (_30461_, _30450_, _30427_);
  nor _44940_ (_30472_, _30461_, _30396_);
  and _44941_ (_30483_, _30472_, _30363_);
  and _44942_ (_30494_, _30483_, _30308_);
  and _44943_ (_30505_, _30494_, _30221_);
  not _44944_ (_30516_, _30505_);
  nor _44945_ (_30526_, _30516_, _30178_);
  and _44946_ (_30537_, _30526_, _30014_);
  not _44947_ (_30548_, _30537_);
  nor _44948_ (_30559_, _30548_, _29676_);
  and _44949_ (_30570_, _30559_, _29238_);
  not _44950_ (_30581_, _30570_);
  nor _44951_ (_30592_, _30581_, _27922_);
  and _44952_ (_30603_, _30592_, _27911_);
  not _44953_ (_30614_, _30603_);
  or _44954_ (_30625_, _30614_, _27889_);
  not _44955_ (_30635_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _44956_ (_30646_, \oc8051_top_1.oc8051_decoder1.wr , _18199_);
  not _44957_ (_30657_, _30646_);
  nor _44958_ (_30668_, _30657_, _26606_);
  and _44959_ (_30679_, _30668_, _30635_);
  not _44960_ (_30690_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _44961_ (_30701_, _27889_, _30690_);
  and _44962_ (_30712_, _30701_, _30679_);
  and _44963_ (_30723_, _30712_, _30625_);
  nor _44964_ (_30734_, _30668_, _30690_);
  not _44965_ (_30744_, _29271_);
  nor _44966_ (_30755_, _29644_, _27977_);
  nor _44967_ (_30766_, _30755_, _30744_);
  not _44968_ (_30777_, _30766_);
  and _44969_ (_30788_, _20323_, _29927_);
  nor _44970_ (_30799_, _30788_, _29194_);
  nor _44971_ (_30810_, _30799_, _27976_);
  nor _44972_ (_30821_, _30069_, _20530_);
  and _44973_ (_30832_, _29007_, _19479_);
  and _44974_ (_30843_, _30832_, _30821_);
  nor _44975_ (_30853_, _30843_, _29960_);
  nor _44976_ (_30864_, _29007_, _20323_);
  not _44977_ (_30875_, _30864_);
  nor _44978_ (_30886_, _30875_, _30090_);
  nor _44979_ (_30897_, _30886_, _30036_);
  and _44980_ (_30908_, _30897_, _30853_);
  or _44981_ (_30919_, _30908_, _30058_);
  nor _44982_ (_30930_, _28986_, _28931_);
  not _44983_ (_30941_, _30287_);
  nor _44984_ (_30952_, _30941_, _28975_);
  nor _44985_ (_30962_, _30952_, _30254_);
  nor _44986_ (_30973_, _30962_, _30930_);
  not _44987_ (_30984_, _30973_);
  and _44988_ (_30995_, _28953_, _28931_);
  and _44989_ (_31006_, _30243_, _27944_);
  and _44990_ (_31017_, _30319_, _28931_);
  nor _44991_ (_31028_, _31017_, _31006_);
  nor _44992_ (_31039_, _31028_, _30995_);
  nand _44993_ (_31050_, _30407_, _28986_);
  nor _44994_ (_31061_, _31050_, _28931_);
  nor _44995_ (_31071_, _30199_, _21922_);
  and _44996_ (_31082_, _30243_, _18221_);
  not _44997_ (_31093_, _31082_);
  nor _44998_ (_31104_, _31093_, _20323_);
  nor _44999_ (_31115_, _31104_, _31071_);
  not _45000_ (_31137_, _31115_);
  nor _45001_ (_31138_, _31137_, _31061_);
  not _45002_ (_31160_, _31138_);
  nor _45003_ (_31161_, _31160_, _31039_);
  nor _45004_ (_31183_, _30385_, _29007_);
  and _45005_ (_31184_, _30341_, _29007_);
  nor _45006_ (_31205_, _31184_, _31183_);
  and _45007_ (_31206_, _31205_, _31161_);
  and _45008_ (_31217_, _31206_, _30984_);
  not _45009_ (_31228_, _31217_);
  nor _45010_ (_31239_, _31228_, _30919_);
  not _45011_ (_31260_, _31239_);
  nor _45012_ (_31261_, _31260_, _30810_);
  and _45013_ (_31282_, _31261_, _30777_);
  not _45014_ (_31283_, _26781_);
  nor _45015_ (_31303_, _27023_, _26902_);
  and _45016_ (_31304_, _31303_, _31283_);
  and _45017_ (_31325_, _31304_, _27878_);
  nand _45018_ (_31326_, _31325_, _31282_);
  or _45019_ (_31347_, _31325_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _45020_ (_31348_, _30668_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _45021_ (_31369_, _31348_, _31347_);
  and _45022_ (_31370_, _31369_, _31326_);
  or _45023_ (_31391_, _31370_, _30734_);
  or _45024_ (_31392_, _31391_, _30723_);
  and _45025_ (_06662_, _31392_, _42882_);
  and _45026_ (_31412_, _26054_, _23626_);
  not _45027_ (_31433_, _31412_);
  and _45028_ (_31434_, _29007_, _29424_);
  nor _45029_ (_31455_, _31434_, _29435_);
  nand _45030_ (_31456_, _29271_, _31455_);
  nor _45031_ (_31477_, _31093_, _29007_);
  and _45032_ (_31478_, _30319_, _28580_);
  and _45033_ (_31499_, _30341_, _21922_);
  nor _45034_ (_31500_, _31499_, _31478_);
  nor _45035_ (_31520_, _29981_, _18988_);
  and _45036_ (_31521_, _29698_, _21922_);
  nor _45037_ (_31542_, _31521_, _31520_);
  nor _45038_ (_31543_, _30374_, _30025_);
  nor _45039_ (_31564_, _31543_, _21922_);
  not _45040_ (_31565_, _31564_);
  and _45041_ (_31586_, _31565_, _31542_);
  nand _45042_ (_31587_, _31586_, _31500_);
  nor _45043_ (_31608_, _31587_, _31477_);
  and _45044_ (_31609_, _23350_, _18265_);
  and _45045_ (_31629_, _31455_, _27955_);
  nor _45046_ (_31630_, _30941_, _28580_);
  nor _45047_ (_31651_, _31630_, _30254_);
  or _45048_ (_31652_, _31651_, _28591_);
  and _45049_ (_31673_, _29687_, _29249_);
  not _45050_ (_31674_, _31673_);
  nor _45051_ (_31695_, _31674_, _21379_);
  and _45052_ (_31696_, _31006_, _20334_);
  nor _45053_ (_31717_, _31696_, _31695_);
  nand _45054_ (_31718_, _31717_, _31652_);
  or _45055_ (_31738_, _31718_, _31629_);
  nor _45056_ (_31739_, _31738_, _31609_);
  and _45057_ (_31760_, _31739_, _31608_);
  and _45058_ (_31761_, _31760_, _31456_);
  and _45059_ (_31782_, _31761_, _31433_);
  not _45060_ (_31783_, _31782_);
  or _45061_ (_31804_, _31783_, _27889_);
  not _45062_ (_31805_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _45063_ (_31826_, _27889_, _31805_);
  and _45064_ (_31827_, _31826_, _30679_);
  and _45065_ (_31847_, _31827_, _31804_);
  nor _45066_ (_31848_, _30668_, _31805_);
  not _45067_ (_31859_, _31282_);
  or _45068_ (_31870_, _31859_, _27889_);
  and _45069_ (_31881_, _31826_, _31348_);
  and _45070_ (_31892_, _31881_, _31870_);
  or _45071_ (_31903_, _31892_, _31848_);
  or _45072_ (_31914_, _31903_, _31847_);
  and _45073_ (_08903_, _31914_, _42882_);
  and _45074_ (_31935_, _23381_, _18265_);
  not _45075_ (_31946_, _31935_);
  and _45076_ (_31956_, _26118_, _23626_);
  nor _45077_ (_31967_, _29981_, _19975_);
  and _45078_ (_31978_, _21922_, _21379_);
  nor _45079_ (_31989_, _31978_, _29709_);
  not _45080_ (_32000_, _31989_);
  nor _45081_ (_32011_, _32000_, _29007_);
  and _45082_ (_32022_, _32000_, _29007_);
  nor _45083_ (_32033_, _32022_, _32011_);
  and _45084_ (_32044_, _32033_, _29698_);
  nor _45085_ (_32054_, _32044_, _31967_);
  nor _45086_ (_32065_, _30047_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _45087_ (_32076_, _32065_, _21389_);
  nor _45088_ (_32087_, _32065_, _21389_);
  nor _45089_ (_32098_, _32087_, _32076_);
  nor _45090_ (_32109_, _32098_, _30036_);
  not _45091_ (_32120_, _32109_);
  and _45092_ (_32131_, _30287_, _28394_);
  nor _45093_ (_32142_, _30265_, _28383_);
  not _45094_ (_32153_, _32142_);
  and _45095_ (_32164_, _30319_, _28372_);
  and _45096_ (_32174_, _30341_, _21379_);
  nor _45097_ (_32185_, _32174_, _32164_);
  nand _45098_ (_32196_, _32185_, _32153_);
  nor _45099_ (_32207_, _32196_, _32131_);
  nor _45100_ (_32218_, _30439_, _21922_);
  not _45101_ (_32229_, _32218_);
  nor _45102_ (_32240_, _30385_, _21379_);
  nor _45103_ (_32251_, _31674_, _21553_);
  nor _45104_ (_32262_, _32251_, _32240_);
  and _45105_ (_32273_, _32262_, _32229_);
  and _45106_ (_32283_, _32273_, _32207_);
  and _45107_ (_32294_, _32283_, _32120_);
  and _45108_ (_32305_, _32294_, _32054_);
  nor _45109_ (_32316_, _28580_, _28394_);
  or _45110_ (_32327_, _32316_, _29347_);
  and _45111_ (_32338_, _32327_, _29435_);
  nor _45112_ (_32349_, _32327_, _29435_);
  or _45113_ (_32360_, _32349_, _32338_);
  and _45114_ (_32371_, _32360_, _29271_);
  nor _45115_ (_32382_, _29040_, _29008_);
  nor _45116_ (_32392_, _32382_, _29051_);
  nor _45117_ (_32403_, _32392_, _27976_);
  nor _45118_ (_32414_, _32403_, _32371_);
  and _45119_ (_32425_, _32414_, _32305_);
  not _45120_ (_32436_, _32425_);
  nor _45121_ (_32447_, _32436_, _31956_);
  and _45122_ (_32458_, _32447_, _31946_);
  not _45123_ (_32469_, _32458_);
  or _45124_ (_32480_, _32469_, _27889_);
  not _45125_ (_32491_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _45126_ (_32501_, _27889_, _32491_);
  and _45127_ (_32512_, _32501_, _30679_);
  and _45128_ (_32523_, _32512_, _32480_);
  nor _45129_ (_32534_, _30668_, _32491_);
  not _45130_ (_32545_, _27023_);
  and _45131_ (_32556_, _32545_, _26902_);
  and _45132_ (_32567_, _32556_, _26781_);
  and _45133_ (_32578_, _32567_, _27878_);
  nand _45134_ (_32589_, _32578_, _31282_);
  or _45135_ (_32600_, _32578_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _45136_ (_32610_, _32600_, _31348_);
  and _45137_ (_32621_, _32610_, _32589_);
  or _45138_ (_32632_, _32621_, _32534_);
  or _45139_ (_32643_, _32632_, _32523_);
  and _45140_ (_08914_, _32643_, _42882_);
  and _45141_ (_32664_, _23413_, _18265_);
  not _45142_ (_32675_, _32664_);
  and _45143_ (_32686_, _26183_, _23626_);
  nor _45144_ (_32697_, _29981_, _18669_);
  nor _45145_ (_32708_, _31978_, _29007_);
  nor _45146_ (_32718_, _29709_, _29785_);
  nor _45147_ (_32729_, _32718_, _32708_);
  nor _45148_ (_32740_, _32729_, _21564_);
  and _45149_ (_32751_, _32729_, _21564_);
  nor _45150_ (_32762_, _32751_, _32740_);
  and _45151_ (_32773_, _32762_, _29698_);
  nor _45152_ (_32784_, _32773_, _32697_);
  nor _45153_ (_32795_, _29051_, _28569_);
  nor _45154_ (_32806_, _32795_, _29062_);
  nor _45155_ (_32817_, _32806_, _27976_);
  and _45156_ (_32827_, _30287_, _28361_);
  not _45157_ (_32838_, _32827_);
  nor _45158_ (_32849_, _30265_, _28350_);
  not _45159_ (_32860_, _32849_);
  and _45160_ (_32871_, _30319_, _28339_);
  and _45161_ (_32882_, _30341_, _21553_);
  nor _45162_ (_32893_, _32882_, _32871_);
  and _45163_ (_32904_, _32893_, _32860_);
  and _45164_ (_32915_, _32904_, _32838_);
  nor _45165_ (_32926_, _30439_, _21379_);
  not _45166_ (_32936_, _32926_);
  nor _45167_ (_32947_, _30385_, _21553_);
  nor _45168_ (_32958_, _31674_, _21052_);
  nor _45169_ (_32969_, _32958_, _32947_);
  and _45170_ (_32980_, _32969_, _32936_);
  and _45171_ (_32991_, _32980_, _32915_);
  not _45172_ (_33002_, _32991_);
  nor _45173_ (_33013_, _33002_, _32817_);
  nor _45174_ (_33024_, _29468_, _29446_);
  nor _45175_ (_33035_, _33024_, _30744_);
  and _45176_ (_33045_, _33035_, _29490_);
  nor _45177_ (_33056_, _32087_, _21553_);
  and _45178_ (_33067_, _29807_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _45179_ (_33078_, _33067_, _33056_);
  nor _45180_ (_33089_, _33078_, _30036_);
  nor _45181_ (_33100_, _33089_, _33045_);
  and _45182_ (_33111_, _33100_, _33013_);
  and _45183_ (_33122_, _33111_, _32784_);
  not _45184_ (_33133_, _33122_);
  nor _45185_ (_33144_, _33133_, _32686_);
  and _45186_ (_33154_, _33144_, _32675_);
  not _45187_ (_33165_, _33154_);
  or _45188_ (_33176_, _33165_, _27889_);
  not _45189_ (_33187_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _45190_ (_33198_, _27889_, _33187_);
  and _45191_ (_33209_, _33198_, _30679_);
  and _45192_ (_33220_, _33209_, _33176_);
  nor _45193_ (_33231_, _30668_, _33187_);
  nand _45194_ (_33242_, _27878_, _26781_);
  or _45195_ (_33253_, _31303_, _33242_);
  and _45196_ (_33263_, _33253_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not _45197_ (_33274_, _26902_);
  and _45198_ (_33285_, _26781_, _27023_);
  and _45199_ (_33296_, _33285_, _33274_);
  not _45200_ (_33307_, _33296_);
  nor _45201_ (_33318_, _33307_, _31282_);
  and _45202_ (_33329_, _26781_, _26902_);
  and _45203_ (_33340_, _33329_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _45204_ (_33351_, _33340_, _33318_);
  and _45205_ (_33362_, _33351_, _27878_);
  or _45206_ (_33372_, _33362_, _33263_);
  and _45207_ (_33383_, _33372_, _31348_);
  or _45208_ (_33394_, _33383_, _33231_);
  or _45209_ (_33405_, _33394_, _33220_);
  and _45210_ (_08925_, _33405_, _42882_);
  and _45211_ (_33426_, _26248_, _23626_);
  not _45212_ (_33437_, _33426_);
  and _45213_ (_33448_, _23466_, _18265_);
  and _45214_ (_33459_, _29490_, _29413_);
  or _45215_ (_33470_, _33459_, _30744_);
  nor _45216_ (_33480_, _33470_, _29501_);
  not _45217_ (_33491_, _33480_);
  nor _45218_ (_33502_, _29062_, _28536_);
  nor _45219_ (_33513_, _33502_, _29073_);
  nor _45220_ (_33524_, _33513_, _27976_);
  nor _45221_ (_33535_, _29981_, _19653_);
  and _45222_ (_33546_, _29720_, _29007_);
  and _45223_ (_33557_, _29818_, _29785_);
  nor _45224_ (_33568_, _33557_, _33546_);
  nor _45225_ (_33579_, _33568_, _21052_);
  not _45226_ (_33589_, _29698_);
  and _45227_ (_33600_, _33568_, _21052_);
  or _45228_ (_33611_, _33600_, _33589_);
  nor _45229_ (_33622_, _33611_, _33579_);
  nor _45230_ (_33633_, _33622_, _33535_);
  not _45231_ (_33644_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _45232_ (_33655_, _29807_, _33644_);
  nor _45233_ (_33666_, _33655_, _21063_);
  nor _45234_ (_33677_, _30385_, _21052_);
  nor _45235_ (_33688_, _30047_, _30036_);
  nor _45236_ (_33698_, _33688_, _33677_);
  or _45237_ (_33709_, _33698_, _33666_);
  nor _45238_ (_33720_, _30265_, _28295_);
  and _45239_ (_33731_, _30287_, _28317_);
  nor _45240_ (_33742_, _33731_, _33720_);
  and _45241_ (_33753_, _30319_, _28306_);
  and _45242_ (_33764_, _30341_, _21052_);
  nor _45243_ (_33775_, _33764_, _33753_);
  nor _45244_ (_33786_, _31674_, _20693_);
  nor _45245_ (_33797_, _30439_, _21553_);
  nor _45246_ (_33807_, _33797_, _33786_);
  and _45247_ (_33818_, _33807_, _33775_);
  and _45248_ (_33829_, _33818_, _33742_);
  and _45249_ (_33840_, _33829_, _33709_);
  nand _45250_ (_33851_, _33840_, _33633_);
  nor _45251_ (_33862_, _33851_, _33524_);
  and _45252_ (_33873_, _33862_, _33491_);
  not _45253_ (_33884_, _33873_);
  nor _45254_ (_33895_, _33884_, _33448_);
  and _45255_ (_33906_, _33895_, _33437_);
  not _45256_ (_33916_, _33906_);
  or _45257_ (_33927_, _33916_, _27889_);
  not _45258_ (_33938_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _45259_ (_33949_, _27889_, _33938_);
  and _45260_ (_33960_, _33949_, _30679_);
  and _45261_ (_33971_, _33960_, _33927_);
  nor _45262_ (_33982_, _30668_, _33938_);
  and _45263_ (_33993_, _33242_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _45264_ (_34004_, _31303_, _26781_);
  and _45265_ (_34015_, _34004_, _31859_);
  or _45266_ (_34026_, _31303_, _31283_);
  nor _45267_ (_34036_, _34026_, _33938_);
  or _45268_ (_34047_, _34036_, _34015_);
  and _45269_ (_34058_, _34047_, _27878_);
  or _45270_ (_34069_, _34058_, _33993_);
  and _45271_ (_34080_, _34069_, _31348_);
  or _45272_ (_34091_, _34080_, _33982_);
  or _45273_ (_34102_, _34091_, _33971_);
  and _45274_ (_08936_, _34102_, _42882_);
  and _45275_ (_34123_, _26313_, _23626_);
  not _45276_ (_34134_, _34123_);
  and _45277_ (_34144_, _23487_, _18265_);
  nor _45278_ (_34155_, _29534_, _28283_);
  not _45279_ (_34166_, _34155_);
  nor _45280_ (_34177_, _30744_, _29545_);
  and _45281_ (_34188_, _34177_, _34166_);
  not _45282_ (_34199_, _34188_);
  nor _45283_ (_34210_, _29139_, _28283_);
  and _45284_ (_34221_, _29139_, _28283_);
  nor _45285_ (_34232_, _34221_, _34210_);
  and _45286_ (_34243_, _34232_, _27955_);
  and _45287_ (_34253_, _29731_, _29007_);
  and _45288_ (_34264_, _29829_, _29785_);
  nor _45289_ (_34277_, _34264_, _34253_);
  and _45290_ (_34296_, _34277_, _20693_);
  nor _45291_ (_34307_, _34277_, _20693_);
  nor _45292_ (_34318_, _34307_, _34296_);
  and _45293_ (_34329_, _34318_, _29698_);
  nor _45294_ (_34340_, _29007_, _18834_);
  and _45295_ (_34351_, _29007_, _20704_);
  nor _45296_ (_34361_, _34351_, _34340_);
  nor _45297_ (_34372_, _34361_, _29981_);
  and _45298_ (_34383_, _30319_, _28251_);
  and _45299_ (_34394_, _30341_, _20693_);
  nor _45300_ (_34405_, _34394_, _34383_);
  and _45301_ (_34416_, _30287_, _28283_);
  nor _45302_ (_34427_, _30265_, _28262_);
  or _45303_ (_34438_, _34427_, _34416_);
  not _45304_ (_34449_, _34438_);
  and _45305_ (_34460_, _34449_, _34405_);
  not _45306_ (_34470_, _34460_);
  or _45307_ (_34481_, _34470_, _34372_);
  nor _45308_ (_34492_, _34481_, _34329_);
  nor _45309_ (_34503_, _30058_, _20704_);
  nor _45310_ (_34514_, _30385_, _20693_);
  nor _45311_ (_34525_, _30069_, _30036_);
  nor _45312_ (_34536_, _34525_, _34514_);
  or _45313_ (_34547_, _34536_, _34503_);
  nor _45314_ (_34558_, _31674_, _20519_);
  nor _45315_ (_34569_, _30439_, _21052_);
  nor _45316_ (_34580_, _34569_, _34558_);
  and _45317_ (_34590_, _34580_, _34547_);
  and _45318_ (_34601_, _34590_, _34492_);
  not _45319_ (_34612_, _34601_);
  nor _45320_ (_34623_, _34612_, _34243_);
  and _45321_ (_34634_, _34623_, _34199_);
  not _45322_ (_34645_, _34634_);
  nor _45323_ (_34656_, _34645_, _34144_);
  and _45324_ (_34667_, _34656_, _34134_);
  not _45325_ (_34678_, _34667_);
  or _45326_ (_34689_, _34678_, _27889_);
  not _45327_ (_34699_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _45328_ (_34710_, _27889_, _34699_);
  and _45329_ (_34721_, _34710_, _30679_);
  and _45330_ (_34732_, _34721_, _34689_);
  nor _45331_ (_34743_, _30668_, _34699_);
  not _45332_ (_34754_, _27878_);
  and _45333_ (_34765_, _27034_, _31283_);
  nor _45334_ (_34776_, _27034_, _31283_);
  nor _45335_ (_34787_, _34776_, _34765_);
  or _45336_ (_34798_, _34787_, _34754_);
  and _45337_ (_34808_, _34798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _45338_ (_34819_, _34765_, _31859_);
  and _45339_ (_34830_, _34776_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or _45340_ (_34841_, _34830_, _34819_);
  and _45341_ (_34852_, _34841_, _27878_);
  or _45342_ (_34863_, _34852_, _34808_);
  and _45343_ (_34874_, _34863_, _31348_);
  or _45344_ (_34885_, _34874_, _34743_);
  or _45345_ (_34896_, _34885_, _34732_);
  and _45346_ (_08947_, _34896_, _42882_);
  and _45347_ (_34916_, _23530_, _18265_);
  not _45348_ (_34927_, _34916_);
  and _45349_ (_34938_, _26400_, _23626_);
  nor _45350_ (_34949_, _29150_, _28240_);
  nor _45351_ (_34960_, _34949_, _29161_);
  nor _45352_ (_34971_, _34960_, _27976_);
  not _45353_ (_34982_, _34971_);
  nor _45354_ (_34993_, _30265_, _28098_);
  and _45355_ (_35004_, _30287_, _28109_);
  nor _45356_ (_35015_, _35004_, _34993_);
  and _45357_ (_35025_, _30319_, _28087_);
  and _45358_ (_35036_, _30341_, _20519_);
  nor _45359_ (_35047_, _35036_, _35025_);
  nor _45360_ (_35058_, _31674_, _19479_);
  not _45361_ (_35069_, _35058_);
  nor _45362_ (_35080_, _30385_, _20519_);
  nor _45363_ (_35091_, _30439_, _20693_);
  nor _45364_ (_35101_, _35091_, _35080_);
  and _45365_ (_35112_, _35101_, _35069_);
  and _45366_ (_35123_, _35112_, _35047_);
  and _45367_ (_35134_, _35123_, _35015_);
  nor _45368_ (_35145_, _29567_, _29545_);
  not _45369_ (_35156_, _35145_);
  nor _45370_ (_35167_, _30744_, _29578_);
  and _45371_ (_35178_, _35167_, _35156_);
  nor _45372_ (_35189_, _29007_, _19805_);
  and _45373_ (_35200_, _29007_, _20530_);
  nor _45374_ (_35211_, _35200_, _35189_);
  nor _45375_ (_35221_, _35211_, _29981_);
  and _45376_ (_35232_, _29742_, _29007_);
  and _45377_ (_35243_, _29840_, _29785_);
  nor _45378_ (_35254_, _35243_, _35232_);
  and _45379_ (_35265_, _35254_, _20519_);
  nor _45380_ (_35276_, _35254_, _20519_);
  or _45381_ (_35287_, _35276_, _33589_);
  nor _45382_ (_35298_, _35287_, _35265_);
  nor _45383_ (_35309_, _35298_, _35221_);
  not _45384_ (_35320_, _30123_);
  and _45385_ (_35331_, _35320_, _30821_);
  nor _45386_ (_35341_, _30123_, _30069_);
  nor _45387_ (_35352_, _35341_, _20519_);
  nor _45388_ (_35363_, _35352_, _35331_);
  nor _45389_ (_35374_, _35363_, _30036_);
  not _45390_ (_35385_, _35374_);
  nand _45391_ (_35396_, _35385_, _35309_);
  nor _45392_ (_35407_, _35396_, _35178_);
  and _45393_ (_35418_, _35407_, _35134_);
  and _45394_ (_35429_, _35418_, _34982_);
  not _45395_ (_35440_, _35429_);
  nor _45396_ (_35451_, _35440_, _34938_);
  and _45397_ (_35461_, _35451_, _34927_);
  not _45398_ (_35472_, _35461_);
  or _45399_ (_35483_, _35472_, _27889_);
  not _45400_ (_35494_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _45401_ (_35505_, _27889_, _35494_);
  and _45402_ (_35516_, _35505_, _30679_);
  and _45403_ (_35527_, _35516_, _35483_);
  nor _45404_ (_35538_, _30668_, _35494_);
  and _45405_ (_35549_, _32556_, _31283_);
  and _45406_ (_35560_, _35549_, _27878_);
  nand _45407_ (_35571_, _35560_, _31282_);
  or _45408_ (_35582_, _35560_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _45409_ (_35592_, _35582_, _31348_);
  and _45410_ (_35603_, _35592_, _35571_);
  or _45411_ (_35614_, _35603_, _35538_);
  or _45412_ (_35625_, _35614_, _35527_);
  and _45413_ (_08958_, _35625_, _42882_);
  and _45414_ (_35646_, _26464_, _23626_);
  not _45415_ (_35657_, _35646_);
  and _45416_ (_35668_, _23562_, _18265_);
  nor _45417_ (_35679_, _29600_, _29578_);
  not _45418_ (_35690_, _35679_);
  nor _45419_ (_35701_, _30744_, _29611_);
  and _45420_ (_35712_, _35701_, _35690_);
  not _45421_ (_35722_, _35712_);
  nor _45422_ (_35733_, _29161_, _28207_);
  nor _45423_ (_35744_, _35733_, _29172_);
  nor _45424_ (_35755_, _35744_, _27976_);
  nor _45425_ (_35766_, _29007_, _28010_);
  or _45426_ (_35777_, _35766_, _29981_);
  nor _45427_ (_35788_, _35777_, _30832_);
  or _45428_ (_35799_, _29007_, _20519_);
  or _45429_ (_35810_, _35243_, _29753_);
  and _45430_ (_35821_, _35810_, _35799_);
  and _45431_ (_35832_, _35821_, _19490_);
  nor _45432_ (_35842_, _35821_, _19490_);
  or _45433_ (_35853_, _35842_, _33589_);
  nor _45434_ (_35864_, _35853_, _35832_);
  nor _45435_ (_35875_, _35864_, _35788_);
  nor _45436_ (_35886_, _35331_, _19479_);
  and _45437_ (_35897_, _35331_, _19479_);
  nor _45438_ (_35908_, _35897_, _35886_);
  nor _45439_ (_35919_, _35908_, _30036_);
  and _45440_ (_35929_, _30287_, _28054_);
  nor _45441_ (_35940_, _30265_, _28043_);
  not _45442_ (_35951_, _35940_);
  and _45443_ (_35962_, _30319_, _28032_);
  and _45444_ (_35973_, _30341_, _19479_);
  nor _45445_ (_35984_, _35973_, _35962_);
  nand _45446_ (_35995_, _35984_, _35951_);
  nor _45447_ (_36006_, _35995_, _35929_);
  nor _45448_ (_36016_, _30439_, _20519_);
  not _45449_ (_36027_, _36016_);
  nor _45450_ (_36038_, _30385_, _19479_);
  nor _45451_ (_36049_, _31674_, _20323_);
  nor _45452_ (_36060_, _36049_, _36038_);
  and _45453_ (_36071_, _36060_, _36027_);
  and _45454_ (_36082_, _36071_, _36006_);
  not _45455_ (_36092_, _36082_);
  nor _45456_ (_36103_, _36092_, _35919_);
  and _45457_ (_36114_, _36103_, _35875_);
  not _45458_ (_36125_, _36114_);
  nor _45459_ (_36136_, _36125_, _35755_);
  and _45460_ (_36147_, _36136_, _35722_);
  not _45461_ (_36158_, _36147_);
  nor _45462_ (_36169_, _36158_, _35668_);
  and _45463_ (_36179_, _36169_, _35657_);
  not _45464_ (_36190_, _36179_);
  or _45465_ (_36201_, _36190_, _27889_);
  not _45466_ (_36212_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _45467_ (_36223_, _27889_, _36212_);
  and _45468_ (_36234_, _36223_, _30679_);
  and _45469_ (_36245_, _36234_, _36201_);
  nor _45470_ (_36256_, _30668_, _36212_);
  nor _45471_ (_36266_, _26781_, _26902_);
  and _45472_ (_36277_, _36266_, _27023_);
  and _45473_ (_36288_, _36277_, _27878_);
  nand _45474_ (_36299_, _36288_, _31282_);
  or _45475_ (_36310_, _36288_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _45476_ (_36321_, _36310_, _31348_);
  and _45477_ (_36332_, _36321_, _36299_);
  or _45478_ (_36343_, _36332_, _36256_);
  or _45479_ (_36353_, _36343_, _36245_);
  and _45480_ (_08969_, _36353_, _42882_);
  and _45481_ (_36374_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45482_ (_36385_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  or _45483_ (_36396_, _36385_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _45484_ (_36407_, _36396_);
  not _45485_ (_36418_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor _45486_ (_36428_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _45487_ (_36439_, _36428_, _36418_);
  and _45488_ (_36450_, _36385_, _18199_);
  and _45489_ (_36461_, _36450_, _36439_);
  not _45490_ (_36472_, _36461_);
  not _45491_ (_36483_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _45492_ (_36494_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _45493_ (_36505_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45494_ (_36516_, _36505_, _36494_);
  and _45495_ (_36527_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and _45496_ (_36537_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45497_ (_36548_, _36537_, _36494_);
  and _45498_ (_36559_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  not _45499_ (_36570_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45500_ (_36581_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _36570_);
  and _45501_ (_36592_, _36581_, _36494_);
  and _45502_ (_36603_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _45503_ (_36614_, _36603_, _36559_);
  or _45504_ (_36625_, _36614_, _36527_);
  and _45505_ (_36636_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _45506_ (_36646_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _45507_ (_36657_, _36646_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _45508_ (_36668_, _36657_, _36494_);
  and _45509_ (_36679_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _45510_ (_36690_, _36679_, _36636_);
  nor _45511_ (_36701_, _36505_, _36494_);
  and _45512_ (_36712_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _45513_ (_36723_, _36505_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _45514_ (_36734_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or _45515_ (_36745_, _36734_, _36712_);
  or _45516_ (_36756_, _36745_, _36690_);
  nor _45517_ (_36767_, _36756_, _36625_);
  and _45518_ (_36778_, _36767_, _36483_);
  nor _45519_ (_36789_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _36483_);
  nor _45520_ (_36800_, _36789_, _36778_);
  nor _45521_ (_36811_, _36800_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  not _45522_ (_36822_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45523_ (_36833_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _36822_);
  nor _45524_ (_36844_, _36833_, _36811_);
  nor _45525_ (_36855_, _36844_, _36472_);
  not _45526_ (_36866_, _36855_);
  not _45527_ (_36877_, _36439_);
  nor _45528_ (_36888_, _36450_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _45529_ (_36898_, _36888_, _36877_);
  and _45530_ (_36909_, _36898_, _36866_);
  not _45531_ (_36920_, _36909_);
  and _45532_ (_36931_, \oc8051_top_1.oc8051_memory_interface1.dack_ir , \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7]);
  and _45533_ (_36942_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _45534_ (_36953_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _45535_ (_36964_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _45536_ (_36975_, _36964_, _36953_);
  and _45537_ (_36986_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and _45538_ (_36997_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _45539_ (_37007_, _36997_, _36986_);
  and _45540_ (_37018_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  and _45541_ (_37029_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _45542_ (_37040_, _37029_, _37018_);
  and _45543_ (_37051_, _37040_, _37007_);
  and _45544_ (_37062_, _37051_, _36975_);
  or _45545_ (_37073_, _36636_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _45546_ (_37084_, _37073_, _37062_);
  nor _45547_ (_37095_, _37084_, _36942_);
  nor _45548_ (_37106_, _37095_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45549_ (_37117_, _37106_, _36931_);
  and _45550_ (_37127_, _37117_, _36461_);
  not _45551_ (_37138_, _37127_);
  nor _45552_ (_37149_, _36450_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _45553_ (_37160_, _37149_, _36877_);
  and _45554_ (_37171_, _37160_, _37138_);
  and _45555_ (_37182_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45556_ (_37193_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45557_ (_37204_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _45558_ (_37215_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor _45559_ (_37226_, _37215_, _37204_);
  and _45560_ (_37236_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _45561_ (_37247_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _45562_ (_37258_, _37247_, _37236_);
  and _45563_ (_37269_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and _45564_ (_37280_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _45565_ (_37291_, _37280_, _37269_);
  and _45566_ (_37302_, _37291_, _37258_);
  and _45567_ (_37313_, _37302_, _37226_);
  nor _45568_ (_37324_, _37313_, _37073_);
  or _45569_ (_37335_, _37324_, _37193_);
  and _45570_ (_37346_, _37335_, _36822_);
  nor _45571_ (_37357_, _37346_, _37182_);
  and _45572_ (_37368_, _37357_, _36461_);
  not _45573_ (_37379_, _37368_);
  nor _45574_ (_37390_, _36450_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _45575_ (_37401_, _37390_, _36877_);
  and _45576_ (_37410_, _37401_, _37379_);
  not _45577_ (_37421_, _37410_);
  and _45578_ (_37432_, _37421_, _37171_);
  and _45579_ (_37443_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45580_ (_37454_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45581_ (_37465_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and _45582_ (_37476_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _45583_ (_37487_, _37476_, _37465_);
  and _45584_ (_37498_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _45585_ (_37509_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _45586_ (_37520_, _37509_, _37498_);
  and _45587_ (_37531_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and _45588_ (_37542_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _45589_ (_37553_, _37542_, _37531_);
  and _45590_ (_37564_, _37553_, _37520_);
  and _45591_ (_37575_, _37564_, _37487_);
  nor _45592_ (_37586_, _37575_, _36636_);
  and _45593_ (_37597_, _37586_, _36483_);
  or _45594_ (_37608_, _37597_, _37454_);
  and _45595_ (_37619_, _37608_, _36822_);
  nor _45596_ (_37630_, _37619_, _37443_);
  and _45597_ (_37641_, _37630_, _36461_);
  not _45598_ (_37652_, _37641_);
  nor _45599_ (_37663_, _36450_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _45600_ (_37674_, _37663_, _36877_);
  and _45601_ (_37685_, _37674_, _37652_);
  and _45602_ (_37696_, _37685_, _37432_);
  and _45603_ (_37707_, _37696_, _36920_);
  and _45604_ (_37718_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45605_ (_37729_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45606_ (_37740_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and _45607_ (_37751_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _45608_ (_37762_, _37751_, _37740_);
  and _45609_ (_37773_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and _45610_ (_37784_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _45611_ (_37795_, _37784_, _37773_);
  and _45612_ (_37806_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _45613_ (_37817_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _45614_ (_37828_, _37817_, _37806_);
  and _45615_ (_37839_, _37828_, _37795_);
  and _45616_ (_37850_, _37839_, _37762_);
  nor _45617_ (_37861_, _37850_, _36636_);
  and _45618_ (_37872_, _37861_, _36483_);
  or _45619_ (_37883_, _37872_, _37729_);
  and _45620_ (_37894_, _37883_, _36822_);
  nor _45621_ (_37905_, _37894_, _37718_);
  and _45622_ (_37916_, _37905_, _36461_);
  not _45623_ (_37927_, _37916_);
  nor _45624_ (_37938_, _36450_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _45625_ (_37949_, _37938_, _36877_);
  and _45626_ (_37960_, _37949_, _37927_);
  and _45627_ (_37971_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45628_ (_37982_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45629_ (_37993_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and _45630_ (_38004_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _45631_ (_38015_, _38004_, _37993_);
  and _45632_ (_38026_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _45633_ (_38037_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _45634_ (_38048_, _38037_, _38026_);
  and _45635_ (_38059_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and _45636_ (_38069_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _45637_ (_38080_, _38069_, _38059_);
  and _45638_ (_38091_, _38080_, _38048_);
  and _45639_ (_38101_, _38091_, _38015_);
  nor _45640_ (_38112_, _38101_, _37073_);
  nor _45641_ (_38123_, _38112_, _37982_);
  nor _45642_ (_38134_, _38123_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45643_ (_38145_, _38134_, _37971_);
  nor _45644_ (_38156_, _38145_, _36472_);
  and _45645_ (_38165_, _36472_, \oc8051_top_1.oc8051_decoder1.op [2]);
  or _45646_ (_38166_, _38165_, _38156_);
  and _45647_ (_38167_, _38166_, _36439_);
  and _45648_ (_38168_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _45649_ (_38169_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and _45650_ (_38170_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _45651_ (_38171_, _38170_, _38169_);
  or _45652_ (_38172_, _38171_, _38168_);
  and _45653_ (_38173_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _45654_ (_38174_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _45655_ (_38175_, _38174_, _38173_);
  and _45656_ (_38176_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _45657_ (_38177_, _38176_, _36636_);
  nand _45658_ (_38178_, _38177_, _38175_);
  nor _45659_ (_38179_, _38178_, _38172_);
  and _45660_ (_38180_, _38179_, _36483_);
  nor _45661_ (_38181_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _36483_);
  nor _45662_ (_38182_, _38181_, _38180_);
  nor _45663_ (_38183_, _38182_, \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  nor _45664_ (_38184_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _36822_);
  nor _45665_ (_38185_, _38184_, _38183_);
  nor _45666_ (_38186_, _38185_, _36472_);
  not _45667_ (_38187_, _38186_);
  nor _45668_ (_38188_, _36450_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _45669_ (_38189_, _38188_, _36877_);
  and _45670_ (_38190_, _38189_, _38187_);
  not _45671_ (_38191_, _38190_);
  nor _45672_ (_38192_, _38191_, _38167_);
  and _45673_ (_38193_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], \oc8051_top_1.oc8051_memory_interface1.dack_ir );
  and _45674_ (_38194_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  and _45675_ (_38195_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and _45676_ (_38196_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _45677_ (_38197_, _38196_, _38195_);
  and _45678_ (_38198_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _45679_ (_38199_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _45680_ (_38200_, _38199_, _38198_);
  and _45681_ (_38201_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  and _45682_ (_38202_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _45683_ (_38203_, _38202_, _38201_);
  and _45684_ (_38204_, _38203_, _38200_);
  and _45685_ (_38205_, _38204_, _38197_);
  nor _45686_ (_38206_, _38205_, _36636_);
  and _45687_ (_38207_, _38206_, _36483_);
  or _45688_ (_38208_, _38207_, _38194_);
  and _45689_ (_38209_, _38208_, _36822_);
  nor _45690_ (_38210_, _38209_, _38193_);
  and _45691_ (_38211_, _38210_, _36461_);
  not _45692_ (_38212_, _38211_);
  nor _45693_ (_38213_, _36450_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _45694_ (_38214_, _38213_, _36877_);
  and _45695_ (_38215_, _38214_, _38212_);
  not _45696_ (_38216_, _38215_);
  and _45697_ (_38217_, _38216_, _38192_);
  and _45698_ (_38218_, _38217_, _37960_);
  and _45699_ (_38219_, _38218_, _37707_);
  not _45700_ (_38220_, _37171_);
  and _45701_ (_38221_, _37685_, _37410_);
  and _45702_ (_38222_, _38221_, _38220_);
  and _45703_ (_38223_, _38222_, _36909_);
  and _45704_ (_38224_, _38218_, _38223_);
  nor _45705_ (_38225_, _37685_, _37410_);
  and _45706_ (_38226_, _38225_, _37171_);
  and _45707_ (_38227_, _38226_, _36909_);
  and _45708_ (_38228_, _38218_, _38227_);
  nor _45709_ (_38229_, _38228_, _38224_);
  not _45710_ (_38230_, _38229_);
  nor _45711_ (_38231_, _38230_, _38219_);
  and _45712_ (_38232_, _38226_, _36920_);
  and _45713_ (_38233_, _38216_, _38167_);
  nor _45714_ (_38234_, _37960_, _38190_);
  and _45715_ (_38235_, _38234_, _38233_);
  and _45716_ (_38236_, _38235_, _38232_);
  and _45717_ (_38237_, _38235_, _37707_);
  nor _45718_ (_38238_, _38237_, _38236_);
  and _45719_ (_38239_, _38238_, _38231_);
  nor _45720_ (_38240_, _38239_, _36407_);
  not _45721_ (_38241_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _45722_ (_38242_, _18199_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _45723_ (_38243_, _38242_, _38241_);
  and _45724_ (_38244_, _37410_, _38220_);
  nor _45725_ (_38245_, _38215_, _38167_);
  and _45726_ (_38246_, _38234_, _38245_);
  and _45727_ (_38247_, _38246_, _38244_);
  and _45728_ (_38248_, _38247_, _38243_);
  and _45729_ (_38249_, _38237_, _18199_);
  and _45730_ (_38250_, _38236_, _18199_);
  nor _45731_ (_38251_, _38250_, _38249_);
  nor _45732_ (_38252_, _38251_, _36385_);
  nor _45733_ (_38253_, _38252_, _38248_);
  not _45734_ (_38254_, _38253_);
  nor _45735_ (_38255_, _38254_, _38240_);
  nor _45736_ (_38256_, _38255_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45737_ (_38257_, _38256_, _36374_);
  and _45738_ (_38258_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45739_ (_38259_, _37960_, _38215_);
  and _45740_ (_38260_, _38259_, _38192_);
  and _45741_ (_38261_, _38260_, _37707_);
  not _45742_ (_38262_, _37960_);
  nor _45743_ (_38263_, _37685_, _37421_);
  and _45744_ (_38264_, _38263_, _37171_);
  and _45745_ (_38265_, _38264_, _36909_);
  and _45746_ (_38266_, _38265_, _38217_);
  and _45747_ (_38267_, _38266_, _38262_);
  nor _45748_ (_38268_, _38267_, _38261_);
  and _45749_ (_38269_, _38190_, _38167_);
  nor _45750_ (_38270_, _38215_, _36909_);
  and _45751_ (_38271_, _38270_, _38269_);
  and _45752_ (_38272_, _38271_, _37696_);
  and _45753_ (_38273_, _38227_, _38260_);
  and _45754_ (_38274_, _37960_, _38191_);
  and _45755_ (_38275_, _38274_, _38233_);
  and _45756_ (_38276_, _38275_, _38232_);
  nor _45757_ (_38277_, _38276_, _38273_);
  not _45758_ (_38278_, _38277_);
  nor _45759_ (_38279_, _38278_, _38272_);
  and _45760_ (_38280_, _38221_, _37171_);
  and _45761_ (_38281_, _38280_, _36920_);
  and _45762_ (_38282_, _38281_, _38275_);
  and _45763_ (_38283_, _37432_, _36909_);
  and _45764_ (_38284_, _38283_, _38275_);
  nor _45765_ (_38285_, _38284_, _38282_);
  and _45766_ (_38286_, _38285_, _38279_);
  and _45767_ (_38287_, _38222_, _36920_);
  and _45768_ (_38288_, _38287_, _38275_);
  and _45769_ (_38289_, _38264_, _36920_);
  and _45770_ (_38290_, _38289_, _38275_);
  nor _45771_ (_38291_, _38290_, _38288_);
  and _45772_ (_38292_, _38215_, _37707_);
  not _45773_ (_38293_, _38292_);
  nor _45774_ (_38294_, _37410_, _37171_);
  and _45775_ (_38295_, _38294_, _37685_);
  and _45776_ (_38296_, _38295_, _38260_);
  not _45777_ (_38297_, _37685_);
  and _45778_ (_38298_, _38294_, _38297_);
  and _45779_ (_38299_, _38298_, _36920_);
  and _45780_ (_38300_, _38299_, _38275_);
  nor _45781_ (_38301_, _38300_, _38296_);
  and _45782_ (_38302_, _38301_, _38293_);
  and _45783_ (_38303_, _38302_, _38291_);
  and _45784_ (_38304_, _38303_, _38286_);
  and _45785_ (_38305_, _38304_, _38268_);
  and _45786_ (_38306_, _38275_, _38265_);
  and _45787_ (_38307_, _38298_, _36909_);
  and _45788_ (_38308_, _38307_, _38275_);
  nor _45789_ (_38309_, _38308_, _38306_);
  and _45790_ (_38310_, _38246_, _37696_);
  and _45791_ (_38311_, _38244_, _38297_);
  and _45792_ (_38312_, _38311_, _36920_);
  and _45793_ (_38313_, _38312_, _38275_);
  nor _45794_ (_38314_, _38313_, _38310_);
  and _45795_ (_38315_, _38314_, _38309_);
  and _45796_ (_38316_, _38289_, _38260_);
  and _45797_ (_38317_, _37696_, _36909_);
  and _45798_ (_38318_, _38317_, _38260_);
  nor _45799_ (_38319_, _38318_, _38316_);
  and _45800_ (_38320_, _38223_, _38260_);
  and _45801_ (_38321_, _38312_, _38217_);
  nor _45802_ (_38322_, _38321_, _38320_);
  and _45803_ (_38323_, _38322_, _38319_);
  and _45804_ (_38324_, _38323_, _38315_);
  and _45805_ (_38325_, _38232_, _38260_);
  and _45806_ (_38326_, _38311_, _36909_);
  and _45807_ (_38327_, _38326_, _38217_);
  nor _45808_ (_38328_, _38327_, _38325_);
  not _45809_ (_38329_, _38328_);
  nor _45810_ (_38330_, _38326_, _38295_);
  not _45811_ (_38331_, _38330_);
  and _45812_ (_38332_, _38331_, _38275_);
  nor _45813_ (_38333_, _38332_, _38329_);
  and _45814_ (_38334_, _38295_, _36909_);
  and _45815_ (_38335_, _38334_, _38246_);
  not _45816_ (_38336_, _38335_);
  and _45817_ (_38337_, _38295_, _36920_);
  and _45818_ (_38338_, _38337_, _38246_);
  and _45819_ (_38339_, _38246_, _38307_);
  nor _45820_ (_38340_, _38339_, _38338_);
  and _45821_ (_38341_, _38340_, _38336_);
  and _45822_ (_38342_, _38246_, _38264_);
  and _45823_ (_38343_, _38287_, _38217_);
  nor _45824_ (_38344_, _38343_, _38342_);
  and _45825_ (_38345_, _38344_, _38341_);
  and _45826_ (_38346_, _38345_, _38333_);
  and _45827_ (_38347_, _38346_, _38324_);
  and _45828_ (_38348_, _38347_, _38305_);
  nor _45829_ (_38349_, _38348_, _36407_);
  and _45830_ (_38350_, \oc8051_top_1.oc8051_decoder1.state [0], _18199_);
  and _45831_ (_38351_, _38350_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _45832_ (_38352_, _38351_, _38296_);
  nor _45833_ (_38353_, _38352_, _38248_);
  not _45834_ (_38354_, _38353_);
  nor _45835_ (_38355_, _38354_, _38349_);
  nor _45836_ (_38356_, _38355_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45837_ (_38357_, _38356_, _38258_);
  and _45838_ (_38358_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _45839_ (_38359_, _38269_, _38216_);
  and _45840_ (_38360_, _38359_, _38264_);
  nor _45841_ (_38361_, _38215_, _36920_);
  and _45842_ (_38362_, _38361_, _38269_);
  and _45843_ (_38363_, _38362_, _38226_);
  nor _45844_ (_38364_, _38363_, _38360_);
  and _45845_ (_38365_, _38362_, _37696_);
  and _45846_ (_38366_, _38298_, _38359_);
  nor _45847_ (_38367_, _38366_, _38365_);
  not _45848_ (_38368_, _38367_);
  and _45849_ (_38369_, _38362_, _38311_);
  and _45850_ (_38370_, _38295_, _38359_);
  or _45851_ (_38371_, _38370_, _38369_);
  nor _45852_ (_38372_, _38371_, _38368_);
  and _45853_ (_38373_, _38372_, _38364_);
  and _45854_ (_38374_, _37960_, _38216_);
  and _45855_ (_38375_, _38374_, _38192_);
  and _45856_ (_38376_, _38375_, _37707_);
  or _45857_ (_38377_, _38223_, _38227_);
  and _45858_ (_38378_, _38377_, _38375_);
  nor _45859_ (_38379_, _38378_, _38376_);
  and _45860_ (_38380_, _38246_, _38265_);
  and _45861_ (_38381_, _38226_, _38271_);
  nor _45862_ (_38382_, _38381_, _38380_);
  and _45863_ (_38383_, _38311_, _38271_);
  and _45864_ (_38384_, _38280_, _38271_);
  nor _45865_ (_38385_, _38384_, _38383_);
  and _45866_ (_38386_, _38222_, _38271_);
  nor _45867_ (_38387_, _38386_, _38296_);
  and _45868_ (_38388_, _38387_, _38385_);
  and _45869_ (_38389_, _38388_, _38382_);
  and _45870_ (_38390_, _38389_, _38379_);
  and _45871_ (_38391_, _38390_, _38373_);
  nor _45872_ (_38392_, _38391_, _36407_);
  and _45873_ (_38393_, _38243_, _38222_);
  and _45874_ (_38394_, _38393_, _38246_);
  or _45875_ (_38395_, _38394_, _38352_);
  nor _45876_ (_38396_, _38395_, _38392_);
  nor _45877_ (_38397_, _38396_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _45878_ (_38398_, _38397_, _38358_);
  nor _45879_ (_38399_, _38398_, _38357_);
  and _45880_ (_38400_, _38399_, _38257_);
  and _45881_ (_09519_, _38400_, _42882_);
  and _45882_ (_38401_, _30679_, _27703_);
  and _45883_ (_38402_, _38401_, _26781_);
  and _45884_ (_38403_, _27845_, _27374_);
  and _45885_ (_38404_, _27242_, _27560_);
  and _45886_ (_38405_, _38404_, _38403_);
  and _45887_ (_38406_, _38405_, _32556_);
  and _45888_ (_38407_, _38406_, _38402_);
  nor _45889_ (_38408_, _38407_, _27396_);
  not _45890_ (_38409_, _38407_);
  and _45891_ (_38410_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _45892_ (_38411_, _23626_, _18265_);
  and _45893_ (_38412_, _29260_, _23604_);
  nor _45894_ (_38413_, _30374_, _38412_);
  and _45895_ (_38414_, _38413_, _38411_);
  nor _45896_ (_38415_, _30428_, _31673_);
  and _45897_ (_38416_, _38415_, _38414_);
  nor _45898_ (_38417_, _38416_, _19479_);
  not _45899_ (_38418_, _38417_);
  and _45900_ (_38419_, _38418_, _36006_);
  and _45901_ (_38420_, _38419_, _35875_);
  nor _45902_ (_38421_, _38420_, _38409_);
  nor _45903_ (_38422_, _38421_, _38410_);
  and _45904_ (_38423_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _45905_ (_38424_, _38416_, _20519_);
  not _45906_ (_38425_, _38424_);
  and _45907_ (_38426_, _38425_, _35047_);
  and _45908_ (_38427_, _38426_, _35015_);
  and _45909_ (_38428_, _38427_, _35309_);
  nor _45910_ (_38429_, _38428_, _38409_);
  nor _45911_ (_38430_, _38429_, _38423_);
  and _45912_ (_38431_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _45913_ (_38432_, _38416_, _20693_);
  not _45914_ (_38433_, _38432_);
  and _45915_ (_38434_, _38433_, _34492_);
  nor _45916_ (_38435_, _38434_, _38409_);
  nor _45917_ (_38436_, _38435_, _38431_);
  and _45918_ (_38437_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _45919_ (_38438_, _38416_, _21052_);
  not _45920_ (_38439_, _38438_);
  and _45921_ (_38440_, _38439_, _33775_);
  and _45922_ (_38441_, _38440_, _33742_);
  and _45923_ (_38442_, _38441_, _33633_);
  nor _45924_ (_38443_, _38442_, _38409_);
  nor _45925_ (_38444_, _38443_, _38437_);
  and _45926_ (_38445_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _45927_ (_38446_, _38416_, _21553_);
  not _45928_ (_38447_, _38446_);
  and _45929_ (_38448_, _38447_, _32915_);
  and _45930_ (_38449_, _38448_, _32784_);
  nor _45931_ (_38450_, _38449_, _38409_);
  nor _45932_ (_38451_, _38450_, _38445_);
  and _45933_ (_38452_, _38409_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor _45934_ (_38453_, _38416_, _21379_);
  not _45935_ (_38454_, _38453_);
  and _45936_ (_38455_, _38454_, _32207_);
  and _45937_ (_38456_, _38455_, _32054_);
  nor _45938_ (_38457_, _38456_, _38409_);
  nor _45939_ (_38458_, _38457_, _38452_);
  nor _45940_ (_38459_, _38407_, _26968_);
  nor _45941_ (_38460_, _38416_, _21922_);
  not _45942_ (_38461_, _38460_);
  and _45943_ (_38462_, _38461_, _31542_);
  and _45944_ (_38463_, _38462_, _31500_);
  and _45945_ (_38464_, _38463_, _31652_);
  not _45946_ (_38465_, _38464_);
  and _45947_ (_38466_, _38465_, _38407_);
  nor _45948_ (_38467_, _38466_, _38459_);
  and _45949_ (_38468_, _38467_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _45950_ (_38469_, _38468_, _38458_);
  and _45951_ (_38470_, _38469_, _38451_);
  and _45952_ (_38471_, _38470_, _38444_);
  and _45953_ (_38472_, _38471_, _38436_);
  and _45954_ (_38473_, _38472_, _38430_);
  and _45955_ (_38474_, _38473_, _38422_);
  and _45956_ (_38475_, _38474_, _38408_);
  nor _45957_ (_38476_, _38474_, _38408_);
  nor _45958_ (_38477_, _38476_, _38475_);
  and _45959_ (_38478_, _38477_, _27111_);
  nor _45960_ (_38479_, _38407_, _27440_);
  not _45961_ (_38480_, _38479_);
  nor _45962_ (_38481_, _38480_, _38478_);
  or _45963_ (_38482_, _38416_, _20323_);
  and _45964_ (_38483_, _38482_, _30363_);
  and _45965_ (_38484_, _38483_, _30308_);
  and _45966_ (_38485_, _38484_, _30014_);
  and _45967_ (_38486_, _38485_, _38407_);
  or _45968_ (_38487_, _38486_, _38481_);
  nor _45969_ (_09540_, _38487_, rst);
  not _45970_ (_38488_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _45971_ (_38489_, _38467_, _38488_);
  nor _45972_ (_38490_, _38467_, _38488_);
  nor _45973_ (_38491_, _38490_, _38489_);
  and _45974_ (_38492_, _38491_, _27111_);
  nor _45975_ (_38493_, _38492_, _26979_);
  nor _45976_ (_38494_, _38493_, _38407_);
  nor _45977_ (_38495_, _38494_, _38466_);
  nand _45978_ (_10696_, _38495_, _42882_);
  nor _45979_ (_38496_, _38468_, _38458_);
  nor _45980_ (_38497_, _38496_, _38469_);
  nor _45981_ (_38498_, _38497_, _26528_);
  nor _45982_ (_38499_, _38498_, _26825_);
  nor _45983_ (_38500_, _38499_, _38407_);
  nor _45984_ (_38501_, _38500_, _38457_);
  nand _45985_ (_10707_, _38501_, _42882_);
  nor _45986_ (_38502_, _38469_, _38451_);
  nor _45987_ (_38503_, _38502_, _38470_);
  nor _45988_ (_38504_, _38503_, _26528_);
  nor _45989_ (_38505_, _38504_, _26573_);
  nor _45990_ (_38506_, _38505_, _38407_);
  nor _45991_ (_38507_, _38506_, _38450_);
  nand _45992_ (_10718_, _38507_, _42882_);
  nor _45993_ (_38508_, _38470_, _38444_);
  nor _45994_ (_38509_, _38508_, _38471_);
  nor _45995_ (_38510_, _38509_, _26528_);
  nor _45996_ (_38511_, _38510_, _27637_);
  nor _45997_ (_38512_, _38511_, _38407_);
  nor _45998_ (_38513_, _38512_, _38443_);
  nor _45999_ (_10729_, _38513_, rst);
  nor _46000_ (_38514_, _38471_, _38436_);
  nor _46001_ (_38515_, _38514_, _38472_);
  nor _46002_ (_38516_, _38515_, _26528_);
  nor _46003_ (_38517_, _38516_, _27769_);
  nor _46004_ (_38518_, _38517_, _38407_);
  nor _46005_ (_38519_, _38518_, _38435_);
  nor _46006_ (_10740_, _38519_, rst);
  nor _46007_ (_38520_, _38472_, _38430_);
  nor _46008_ (_38521_, _38520_, _38473_);
  nor _46009_ (_38522_, _38521_, _26528_);
  nor _46010_ (_38523_, _38522_, _27286_);
  nor _46011_ (_38524_, _38523_, _38407_);
  nor _46012_ (_38525_, _38524_, _38429_);
  nor _46013_ (_10751_, _38525_, rst);
  nor _46014_ (_38526_, _38473_, _38422_);
  nor _46015_ (_38527_, _38526_, _38474_);
  nor _46016_ (_38528_, _38527_, _26528_);
  nor _46017_ (_38529_, _38528_, _27143_);
  nor _46018_ (_38530_, _38529_, _38407_);
  nor _46019_ (_38531_, _38530_, _38421_);
  nor _46020_ (_10762_, _38531_, rst);
  and _46021_ (_38532_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _18199_);
  and _46022_ (_38533_, _38532_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not _46023_ (_38534_, _38533_);
  nor _46024_ (_38535_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not _46025_ (_38536_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _46026_ (_38537_, _38536_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46027_ (_38538_, _38537_, _38535_);
  nor _46028_ (_38539_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not _46029_ (_38540_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _46030_ (_38541_, _38540_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46031_ (_38542_, _38541_, _38539_);
  nor _46032_ (_38543_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not _46033_ (_38544_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _46034_ (_38545_, _38544_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46035_ (_38546_, _38545_, _38543_);
  nor _46036_ (_38547_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  not _46037_ (_38548_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _46038_ (_38549_, _38548_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46039_ (_38550_, _38549_, _38547_);
  nor _46040_ (_38551_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not _46041_ (_38552_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _46042_ (_38553_, _38552_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46043_ (_38554_, _38553_, _38551_);
  not _46044_ (_38555_, _38554_);
  nor _46045_ (_38556_, _38555_, _30755_);
  nor _46046_ (_38557_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  not _46047_ (_38558_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _46048_ (_38559_, _38558_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46049_ (_38560_, _38559_, _38557_);
  and _46050_ (_38561_, _38560_, _38556_);
  nor _46051_ (_38562_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  not _46052_ (_38563_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _46053_ (_38564_, _38563_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46054_ (_38565_, _38564_, _38562_);
  and _46055_ (_38566_, _38565_, _38561_);
  and _46056_ (_38567_, _38566_, _38550_);
  nor _46057_ (_38568_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  not _46058_ (_38569_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _46059_ (_38570_, _38569_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _46060_ (_38571_, _38570_, _38568_);
  and _46061_ (_38572_, _38571_, _38567_);
  and _46062_ (_38573_, _38572_, _38546_);
  and _46063_ (_38574_, _38573_, _38542_);
  nand _46064_ (_38575_, _38574_, _38538_);
  or _46065_ (_38576_, _38574_, _38538_);
  and _46066_ (_38577_, _38576_, _38575_);
  and _46067_ (_38578_, _38577_, _29271_);
  not _46068_ (_38579_, _38578_);
  and _46069_ (_38580_, _23318_, _18265_);
  and _46070_ (_38581_, _29763_, _20334_);
  and _46071_ (_38582_, _38581_, _28405_);
  and _46072_ (_38583_, _38582_, _28437_);
  and _46073_ (_38584_, _38583_, _28481_);
  and _46074_ (_38585_, _38584_, _29084_);
  nor _46075_ (_38586_, _38585_, _29785_);
  and _46076_ (_38587_, _29007_, _18834_);
  nor _46077_ (_38588_, _38587_, _38586_);
  and _46078_ (_38589_, _29851_, _20323_);
  and _46079_ (_38590_, _19653_, _18669_);
  and _46080_ (_38591_, _19975_, _18988_);
  and _46081_ (_38592_, _38591_, _38590_);
  and _46082_ (_38593_, _38592_, _38589_);
  and _46083_ (_38594_, _19805_, _18834_);
  and _46084_ (_38595_, _38594_, _38593_);
  nor _46085_ (_38596_, _38595_, _29007_);
  and _46086_ (_38597_, _29007_, _19805_);
  nor _46087_ (_38598_, _38597_, _38596_);
  and _46088_ (_38599_, _38598_, _38588_);
  nor _46089_ (_38600_, _29007_, _19164_);
  and _46090_ (_38601_, _29007_, _19164_);
  nor _46091_ (_38602_, _38601_, _38600_);
  and _46092_ (_38603_, _38602_, _38599_);
  and _46093_ (_38604_, _38603_, _29927_);
  nor _46094_ (_38605_, _38603_, _29927_);
  nor _46095_ (_38606_, _38605_, _38604_);
  and _46096_ (_38607_, _38606_, _29698_);
  and _46097_ (_38608_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  and _46098_ (_38609_, _29007_, _29927_);
  nor _46099_ (_38610_, _38609_, _30864_);
  nor _46100_ (_38611_, _38610_, _29981_);
  nor _46101_ (_38612_, _31093_, _21052_);
  nor _46102_ (_38613_, _30385_, _20149_);
  or _46103_ (_38614_, _38613_, _38612_);
  or _46104_ (_38615_, _38614_, _38611_);
  nor _46105_ (_38616_, _38615_, _38608_);
  not _46106_ (_38617_, _38616_);
  nor _46107_ (_38618_, _38617_, _38607_);
  not _46108_ (_38619_, _38618_);
  nor _46109_ (_38620_, _38619_, _38580_);
  and _46110_ (_38621_, _38620_, _38579_);
  nor _46111_ (_38622_, _38621_, _38534_);
  and _46112_ (_38623_, _38405_, _34004_);
  and _46113_ (_38624_, _38623_, _38401_);
  or _46114_ (_38625_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _46115_ (_38626_, _38625_, _38534_);
  nand _46116_ (_38627_, _38624_, _30603_);
  and _46117_ (_38628_, _38627_, _38626_);
  or _46118_ (_38629_, _38628_, _38622_);
  and _46119_ (_12713_, _38629_, _42882_);
  and _46120_ (_38630_, _38405_, _33296_);
  and _46121_ (_38631_, _38630_, _38401_);
  nor _46122_ (_38632_, _38631_, _38533_);
  not _46123_ (_38633_, _38632_);
  nand _46124_ (_38634_, _38633_, _30603_);
  or _46125_ (_38635_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _46126_ (_38636_, _38635_, _42882_);
  and _46127_ (_12734_, _38636_, _38634_);
  and _46128_ (_38637_, _25917_, _23626_);
  not _46129_ (_38638_, _38637_);
  and _46130_ (_38639_, _38555_, _30755_);
  nor _46131_ (_38640_, _38639_, _38556_);
  and _46132_ (_38641_, _38640_, _29271_);
  nor _46133_ (_38642_, _30864_, _29960_);
  not _46134_ (_38643_, _38642_);
  nor _46135_ (_38644_, _38643_, _29872_);
  nor _46136_ (_38645_, _38644_, _28405_);
  and _46137_ (_38646_, _38644_, _28405_);
  nor _46138_ (_38647_, _38646_, _38645_);
  and _46139_ (_38648_, _38647_, _29698_);
  nor _46140_ (_38649_, _30385_, _18988_);
  and _46141_ (_38650_, _23096_, _18265_);
  nor _46142_ (_38651_, _31093_, _20693_);
  nor _46143_ (_38652_, _29981_, _21922_);
  or _46144_ (_38653_, _38652_, _38651_);
  or _46145_ (_38654_, _38653_, _38650_);
  nor _46146_ (_38655_, _38654_, _38649_);
  not _46147_ (_38656_, _38655_);
  nor _46148_ (_38657_, _38656_, _38648_);
  not _46149_ (_38658_, _38657_);
  nor _46150_ (_38659_, _38658_, _38641_);
  and _46151_ (_38660_, _38659_, _38638_);
  nor _46152_ (_38661_, _38660_, _38534_);
  or _46153_ (_38662_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _46154_ (_38663_, _38662_, _38534_);
  nand _46155_ (_38664_, _38624_, _31782_);
  and _46156_ (_38665_, _38664_, _38663_);
  or _46157_ (_38666_, _38665_, _38661_);
  and _46158_ (_13647_, _38666_, _42882_);
  nor _46159_ (_38667_, _38560_, _38556_);
  nor _46160_ (_38668_, _38667_, _38561_);
  and _46161_ (_38669_, _38668_, _29271_);
  not _46162_ (_38670_, _38669_);
  and _46163_ (_38671_, _24909_, _23626_);
  nor _46164_ (_38672_, _20323_, _18988_);
  and _46165_ (_38673_, _38672_, _29763_);
  and _46166_ (_38674_, _38673_, _29007_);
  and _46167_ (_38675_, _38589_, _18988_);
  and _46168_ (_38676_, _38675_, _29785_);
  nor _46169_ (_38677_, _38676_, _38674_);
  nor _46170_ (_38678_, _38677_, _28437_);
  and _46171_ (_38679_, _38677_, _28437_);
  nor _46172_ (_38680_, _38679_, _38678_);
  nor _46173_ (_38681_, _38680_, _33589_);
  nor _46174_ (_38682_, _30385_, _19975_);
  and _46175_ (_38683_, _23128_, _18265_);
  nor _46176_ (_38684_, _31093_, _20519_);
  nor _46177_ (_38685_, _29981_, _21379_);
  or _46178_ (_38686_, _38685_, _38684_);
  or _46179_ (_38687_, _38686_, _38683_);
  nor _46180_ (_38688_, _38687_, _38682_);
  not _46181_ (_38689_, _38688_);
  nor _46182_ (_38690_, _38689_, _38681_);
  not _46183_ (_38691_, _38690_);
  nor _46184_ (_38692_, _38691_, _38671_);
  and _46185_ (_38693_, _38692_, _38670_);
  nor _46186_ (_38694_, _38693_, _38534_);
  or _46187_ (_38695_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _46188_ (_38696_, _38695_, _38534_);
  nand _46189_ (_38697_, _38624_, _32458_);
  and _46190_ (_38698_, _38697_, _38696_);
  or _46191_ (_38699_, _38698_, _38694_);
  and _46192_ (_13657_, _38699_, _42882_);
  nor _46193_ (_38700_, _38565_, _38561_);
  nor _46194_ (_38701_, _38700_, _38566_);
  and _46195_ (_38702_, _38701_, _29271_);
  not _46196_ (_38703_, _38702_);
  and _46197_ (_38704_, _38675_, _19975_);
  and _46198_ (_38705_, _38704_, _29785_);
  and _46199_ (_38706_, _38673_, _28437_);
  and _46200_ (_38707_, _38706_, _29007_);
  nor _46201_ (_38708_, _38707_, _38705_);
  and _46202_ (_38709_, _38708_, _18669_);
  nor _46203_ (_38710_, _38708_, _18669_);
  nor _46204_ (_38711_, _38710_, _38709_);
  and _46205_ (_38712_, _38711_, _29698_);
  not _46206_ (_38713_, _38712_);
  nor _46207_ (_38714_, _29981_, _21553_);
  and _46208_ (_38715_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor _46209_ (_38716_, _38715_, _38714_);
  and _46210_ (_38717_, _23159_, _18265_);
  nor _46211_ (_38718_, _31093_, _19479_);
  nor _46212_ (_38719_, _30385_, _18669_);
  or _46213_ (_38720_, _38719_, _38718_);
  nor _46214_ (_38721_, _38720_, _38717_);
  and _46215_ (_38722_, _38721_, _38716_);
  and _46216_ (_38723_, _38722_, _38713_);
  and _46217_ (_38724_, _38723_, _38703_);
  nor _46218_ (_38725_, _38724_, _38534_);
  or _46219_ (_38726_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _46220_ (_38727_, _38726_, _38534_);
  nand _46221_ (_38728_, _38624_, _33154_);
  and _46222_ (_38729_, _38728_, _38727_);
  or _46223_ (_38730_, _38729_, _38725_);
  and _46224_ (_13668_, _38730_, _42882_);
  nor _46225_ (_38731_, _38566_, _38550_);
  not _46226_ (_38732_, _38731_);
  nor _46227_ (_38733_, _38567_, _30744_);
  and _46228_ (_38734_, _38733_, _38732_);
  not _46229_ (_38735_, _38734_);
  and _46230_ (_38736_, _23191_, _18265_);
  not _46231_ (_38737_, _38736_);
  nor _46232_ (_38738_, _38584_, _29084_);
  not _46233_ (_38739_, _38738_);
  and _46234_ (_38740_, _38739_, _38586_);
  and _46235_ (_38741_, _38704_, _18669_);
  nor _46236_ (_38742_, _38741_, _19653_);
  nor _46237_ (_38743_, _38742_, _38593_);
  nor _46238_ (_38744_, _38743_, _29007_);
  nor _46239_ (_38745_, _38744_, _38740_);
  nor _46240_ (_38746_, _38745_, _33589_);
  nor _46241_ (_38747_, _30385_, _19653_);
  nor _46242_ (_38748_, _29981_, _21052_);
  and _46243_ (_38749_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or _46244_ (_38750_, _38749_, _38748_);
  or _46245_ (_38751_, _38750_, _31104_);
  nor _46246_ (_38752_, _38751_, _38747_);
  not _46247_ (_38753_, _38752_);
  nor _46248_ (_38754_, _38753_, _38746_);
  and _46249_ (_38755_, _38754_, _38737_);
  and _46250_ (_38756_, _38755_, _38735_);
  nor _46251_ (_38757_, _38756_, _38534_);
  or _46252_ (_38758_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _46253_ (_38759_, _38758_, _38534_);
  nand _46254_ (_38760_, _38624_, _33906_);
  and _46255_ (_38761_, _38760_, _38759_);
  or _46256_ (_38762_, _38761_, _38757_);
  and _46257_ (_13679_, _38762_, _42882_);
  nor _46258_ (_38763_, _38571_, _38567_);
  nor _46259_ (_38764_, _38763_, _38572_);
  and _46260_ (_38765_, _38764_, _29271_);
  not _46261_ (_38766_, _38765_);
  and _46262_ (_38767_, _23223_, _18265_);
  nor _46263_ (_38768_, _38593_, _29007_);
  nor _46264_ (_38769_, _38768_, _38586_);
  nor _46265_ (_38770_, _38769_, _28120_);
  and _46266_ (_38771_, _38769_, _28120_);
  nor _46267_ (_38772_, _38771_, _38770_);
  and _46268_ (_38773_, _38772_, _29698_);
  and _46269_ (_38774_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor _46270_ (_38775_, _29007_, _20704_);
  or _46271_ (_38776_, _38775_, _29981_);
  nor _46272_ (_38777_, _38776_, _38587_);
  nor _46273_ (_38778_, _31093_, _21922_);
  nor _46274_ (_38779_, _30385_, _18834_);
  or _46275_ (_38780_, _38779_, _38778_);
  or _46276_ (_38781_, _38780_, _38777_);
  nor _46277_ (_38782_, _38781_, _38774_);
  not _46278_ (_38783_, _38782_);
  nor _46279_ (_38784_, _38783_, _38773_);
  not _46280_ (_38785_, _38784_);
  nor _46281_ (_38786_, _38785_, _38767_);
  and _46282_ (_38787_, _38786_, _38766_);
  nor _46283_ (_38788_, _38787_, _38534_);
  or _46284_ (_38789_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _46285_ (_38790_, _38789_, _38534_);
  nand _46286_ (_38791_, _38624_, _34667_);
  and _46287_ (_38792_, _38791_, _38790_);
  or _46288_ (_38793_, _38792_, _38788_);
  and _46289_ (_13690_, _38793_, _42882_);
  nor _46290_ (_38794_, _38572_, _38546_);
  not _46291_ (_38795_, _38794_);
  nor _46292_ (_38796_, _38573_, _30744_);
  and _46293_ (_38797_, _38796_, _38795_);
  not _46294_ (_38798_, _38797_);
  and _46295_ (_38799_, _23255_, _18265_);
  and _46296_ (_38800_, _38593_, _18834_);
  nor _46297_ (_38801_, _38800_, _29007_);
  not _46298_ (_38802_, _38801_);
  and _46299_ (_38803_, _38802_, _38588_);
  and _46300_ (_38804_, _38803_, _19805_);
  nor _46301_ (_38805_, _38803_, _19805_);
  nor _46302_ (_38806_, _38805_, _38804_);
  nor _46303_ (_38807_, _38806_, _33589_);
  and _46304_ (_38808_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _46305_ (_38809_, _29007_, _20530_);
  or _46306_ (_38810_, _38809_, _29981_);
  nor _46307_ (_38811_, _38810_, _38597_);
  nor _46308_ (_38812_, _31093_, _21379_);
  nor _46309_ (_38813_, _30385_, _19805_);
  or _46310_ (_38814_, _38813_, _38812_);
  or _46311_ (_38815_, _38814_, _38811_);
  nor _46312_ (_38816_, _38815_, _38808_);
  not _46313_ (_38817_, _38816_);
  nor _46314_ (_38818_, _38817_, _38807_);
  not _46315_ (_38819_, _38818_);
  nor _46316_ (_38820_, _38819_, _38799_);
  and _46317_ (_38821_, _38820_, _38798_);
  nor _46318_ (_38822_, _38821_, _38534_);
  or _46319_ (_38823_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _46320_ (_38824_, _38823_, _38534_);
  nand _46321_ (_38825_, _38624_, _35461_);
  and _46322_ (_38826_, _38825_, _38824_);
  or _46323_ (_38827_, _38826_, _38822_);
  and _46324_ (_13701_, _38827_, _42882_);
  nor _46325_ (_38828_, _38573_, _38542_);
  nor _46326_ (_38829_, _38828_, _38574_);
  and _46327_ (_38830_, _38829_, _29271_);
  and _46328_ (_38831_, _23286_, _18265_);
  and _46329_ (_38832_, _38599_, _19164_);
  nor _46330_ (_38833_, _38599_, _19164_);
  or _46331_ (_38834_, _38833_, _38832_);
  and _46332_ (_38835_, _38834_, _29698_);
  or _46333_ (_38836_, _29007_, _19490_);
  nor _46334_ (_38837_, _38601_, _29981_);
  and _46335_ (_38838_, _38837_, _38836_);
  nor _46336_ (_38839_, _31093_, _21553_);
  nor _46337_ (_38840_, _30385_, _19164_);
  and _46338_ (_38841_, _23626_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  or _46339_ (_38842_, _38841_, _38840_);
  or _46340_ (_38843_, _38842_, _38839_);
  or _46341_ (_38844_, _38843_, _38838_);
  or _46342_ (_38845_, _38844_, _38835_);
  or _46343_ (_38846_, _38845_, _38831_);
  or _46344_ (_38847_, _38846_, _38830_);
  and _46345_ (_38848_, _38847_, _38533_);
  or _46346_ (_38849_, _38624_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and _46347_ (_38850_, _38849_, _38534_);
  nand _46348_ (_38851_, _38624_, _36179_);
  and _46349_ (_38852_, _38851_, _38850_);
  or _46350_ (_38853_, _38852_, _38848_);
  and _46351_ (_13712_, _38853_, _42882_);
  nand _46352_ (_38854_, _38633_, _31782_);
  or _46353_ (_38855_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _46354_ (_38856_, _38855_, _42882_);
  and _46355_ (_13723_, _38856_, _38854_);
  nand _46356_ (_38857_, _38633_, _32458_);
  or _46357_ (_38858_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _46358_ (_38859_, _38858_, _42882_);
  and _46359_ (_13733_, _38859_, _38857_);
  nand _46360_ (_38860_, _38633_, _33154_);
  or _46361_ (_38861_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _46362_ (_38862_, _38861_, _42882_);
  and _46363_ (_13744_, _38862_, _38860_);
  nand _46364_ (_38863_, _38633_, _33906_);
  or _46365_ (_38864_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _46366_ (_38865_, _38864_, _42882_);
  and _46367_ (_13755_, _38865_, _38863_);
  nand _46368_ (_38866_, _38633_, _34667_);
  or _46369_ (_38867_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _46370_ (_38868_, _38867_, _42882_);
  and _46371_ (_13766_, _38868_, _38866_);
  nand _46372_ (_38869_, _38633_, _35461_);
  or _46373_ (_38870_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _46374_ (_38871_, _38870_, _42882_);
  and _46375_ (_13777_, _38871_, _38869_);
  nand _46376_ (_38872_, _38633_, _36179_);
  or _46377_ (_38873_, _38633_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _46378_ (_38874_, _38873_, _42882_);
  and _46379_ (_13788_, _38874_, _38872_);
  nor _46380_ (_38875_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and _46381_ (_38876_, _38875_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _46382_ (_38877_, _38875_, _31282_);
  or _46383_ (_38878_, _38877_, _38876_);
  not _46384_ (_38879_, _27374_);
  nor _46385_ (_38880_, _38879_, _27242_);
  and _46386_ (_38881_, _38880_, _31348_);
  and _46387_ (_38882_, _38881_, _27867_);
  not _46388_ (_38883_, _38882_);
  and _46389_ (_38884_, _38883_, _38878_);
  and _46390_ (_38885_, _38880_, _27867_);
  and _46391_ (_38886_, _38885_, _31348_);
  not _46392_ (_38887_, _31304_);
  nor _46393_ (_38888_, _38887_, _31282_);
  not _46394_ (_38889_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _46395_ (_38890_, _31304_, _38889_);
  or _46396_ (_38891_, _38890_, _38888_);
  and _46397_ (_38892_, _38891_, _38886_);
  or _46398_ (_38893_, _38892_, _38884_);
  and _46399_ (_38894_, _38401_, _27045_);
  nor _46400_ (_38895_, _27242_, _27549_);
  nor _46401_ (_38896_, _27845_, _38879_);
  and _46402_ (_38897_, _38896_, _38895_);
  and _46403_ (_38898_, _38897_, _38894_);
  or _46404_ (_38899_, _38898_, _38893_);
  and _46405_ (_38900_, _38894_, _38895_);
  and _46406_ (_38901_, _38900_, _38896_);
  nand _46407_ (_38902_, _38901_, _38485_);
  and _46408_ (_38903_, _38902_, _42882_);
  and _46409_ (_15193_, _38903_, _38899_);
  not _46410_ (_38904_, _38901_);
  not _46411_ (_38905_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand _46412_ (_38906_, _38886_, _32567_);
  nand _46413_ (_38907_, _38906_, _38905_);
  and _46414_ (_38908_, _38907_, _38904_);
  or _46415_ (_38909_, _38906_, _31859_);
  and _46416_ (_38910_, _38909_, _38908_);
  nor _46417_ (_38911_, _38904_, _38456_);
  or _46418_ (_38912_, _38911_, _38910_);
  and _46419_ (_17374_, _38912_, _42882_);
  or _46420_ (_38913_, _30799_, _29183_);
  not _46421_ (_38914_, _30788_);
  nand _46422_ (_38915_, _38914_, _29183_);
  and _46423_ (_38916_, _38915_, _27955_);
  and _46424_ (_38917_, _38916_, _38913_);
  not _46425_ (_38918_, _27977_);
  nand _46426_ (_38919_, _29633_, _38918_);
  or _46427_ (_38920_, _29633_, _27988_);
  and _46428_ (_38921_, _29271_, _38920_);
  and _46429_ (_38922_, _38921_, _38919_);
  and _46430_ (_38923_, _38594_, _24810_);
  and _46431_ (_38924_, _38592_, _23626_);
  nand _46432_ (_38925_, _38924_, _38923_);
  nand _46433_ (_38926_, _38925_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _46434_ (_38927_, _38926_, _38922_);
  or _46435_ (_38928_, _38927_, _38917_);
  or _46436_ (_38929_, _23381_, _23350_);
  or _46437_ (_38930_, _38929_, _23413_);
  or _46438_ (_38931_, _38930_, _23466_);
  or _46439_ (_38932_, _38931_, _23487_);
  or _46440_ (_38933_, _38932_, _23530_);
  or _46441_ (_38934_, _38933_, _23562_);
  and _46442_ (_38935_, _38934_, _18265_);
  or _46443_ (_38936_, _38935_, _38928_);
  or _46444_ (_38937_, _38936_, _27922_);
  nor _46445_ (_38938_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _46446_ (_38939_, _38938_, _38882_);
  and _46447_ (_38940_, _38939_, _38937_);
  and _46448_ (_38941_, _33307_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _46449_ (_38942_, _38941_, _33318_);
  and _46450_ (_38943_, _38942_, _38886_);
  or _46451_ (_38944_, _38943_, _38898_);
  or _46452_ (_38945_, _38944_, _38940_);
  nand _46453_ (_38946_, _38901_, _38449_);
  and _46454_ (_38947_, _38946_, _42882_);
  and _46455_ (_17385_, _38947_, _38945_);
  not _46456_ (_38948_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nand _46457_ (_38949_, _38886_, _34004_);
  nand _46458_ (_38950_, _38949_, _38948_);
  and _46459_ (_38951_, _38950_, _38904_);
  or _46460_ (_38952_, _38949_, _31859_);
  and _46461_ (_38953_, _38952_, _38951_);
  nor _46462_ (_38954_, _38904_, _38442_);
  or _46463_ (_38957_, _38954_, _38953_);
  and _46464_ (_17396_, _38957_, _42882_);
  or _46465_ (_38959_, _38883_, _34787_);
  and _46466_ (_38960_, _38959_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _46467_ (_38961_, _34776_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _46468_ (_38962_, _38961_, _34819_);
  and _46469_ (_38963_, _38962_, _38886_);
  or _46470_ (_38964_, _38963_, _38960_);
  and _46471_ (_38965_, _38964_, _38904_);
  nor _46472_ (_38966_, _38904_, _38434_);
  or _46473_ (_38967_, _38966_, _38965_);
  and _46474_ (_17407_, _38967_, _42882_);
  not _46475_ (_38977_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand _46476_ (_38983_, _38886_, _35549_);
  nand _46477_ (_38989_, _38983_, _38977_);
  and _46478_ (_38992_, _38989_, _38904_);
  or _46479_ (_38993_, _38983_, _31859_);
  and _46480_ (_38994_, _38993_, _38992_);
  nor _46481_ (_38995_, _38904_, _38428_);
  or _46482_ (_38996_, _38995_, _38994_);
  and _46483_ (_17418_, _38996_, _42882_);
  nand _46484_ (_38997_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and _46485_ (_38998_, _29271_, _29534_);
  and _46486_ (_38999_, _29139_, _27955_);
  nor _46487_ (_39000_, _38999_, _38998_);
  nor _46488_ (_39001_, _39000_, _38997_);
  or _46489_ (_39002_, _38997_, _30374_);
  and _46490_ (_39003_, _39002_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _46491_ (_39004_, _39003_, _38882_);
  or _46492_ (_39005_, _39004_, _39001_);
  not _46493_ (_39006_, _36277_);
  nor _46494_ (_39007_, _39006_, _31282_);
  or _46495_ (_39008_, _36277_, _33644_);
  nand _46496_ (_39009_, _39008_, _38882_);
  or _46497_ (_39010_, _39009_, _39007_);
  and _46498_ (_39011_, _39010_, _39005_);
  or _46499_ (_39012_, _39011_, _38901_);
  nand _46500_ (_39013_, _38901_, _38420_);
  and _46501_ (_39014_, _39013_, _42882_);
  and _46502_ (_17429_, _39014_, _39012_);
  not _46503_ (_39017_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46504_ (_39018_, _38532_, _39017_);
  not _46505_ (_39019_, _39018_);
  nor _46506_ (_39020_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _46507_ (_39021_, _39020_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _46508_ (_39022_, _27045_, _27703_);
  and _46509_ (_39023_, _27845_, _38879_);
  and _46510_ (_39024_, _39023_, _38895_);
  and _46511_ (_39025_, _39024_, _39022_);
  and _46512_ (_39026_, _39025_, _30679_);
  nor _46513_ (_39027_, _39026_, _39021_);
  nor _46514_ (_39028_, _39027_, _30603_);
  and _46515_ (_39029_, _27845_, _27703_);
  not _46516_ (_39030_, _31348_);
  nor _46517_ (_39031_, _39030_, _27549_);
  and _46518_ (_39032_, _39031_, _27385_);
  and _46519_ (_39033_, _39032_, _39029_);
  and _46520_ (_39034_, _39033_, _31304_);
  and _46521_ (_39035_, _39034_, _31282_);
  nor _46522_ (_39036_, _39034_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _46523_ (_39037_, _39036_);
  and _46524_ (_39038_, _39027_, _39019_);
  and _46525_ (_39039_, _39038_, _39037_);
  not _46526_ (_39040_, _39039_);
  nor _46527_ (_39041_, _39040_, _39035_);
  or _46528_ (_39042_, _39041_, _39028_);
  and _46529_ (_39043_, _39042_, _39019_);
  nor _46530_ (_39044_, _39019_, _38621_);
  or _46531_ (_39045_, _39044_, _39043_);
  and _46532_ (_17998_, _39045_, _42882_);
  nor _46533_ (_39046_, _39019_, _38660_);
  nor _46534_ (_39047_, _39027_, _31783_);
  not _46535_ (_39048_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _46536_ (_39049_, _39029_, _27560_);
  and _46537_ (_39050_, _31348_, _27385_);
  and _46538_ (_39051_, _39050_, _39049_);
  nor _46539_ (_39052_, _39051_, _39048_);
  not _46540_ (_39053_, _39052_);
  and _46541_ (_39055_, _39053_, _39027_);
  not _46542_ (_39059_, _39055_);
  not _46543_ (_39065_, _27045_);
  nor _46544_ (_39070_, _31282_, _39065_);
  nor _46545_ (_39077_, _27045_, _39048_);
  nor _46546_ (_39085_, _39077_, _39070_);
  and _46547_ (_39093_, _39038_, _39051_);
  not _46548_ (_39094_, _39093_);
  nor _46549_ (_39095_, _39094_, _39085_);
  nor _46550_ (_39096_, _39095_, _39059_);
  nor _46551_ (_39097_, _39096_, _39018_);
  not _46552_ (_39098_, _39097_);
  nor _46553_ (_39099_, _39098_, _39047_);
  nor _46554_ (_39100_, _39099_, _39046_);
  nor _46555_ (_19849_, _39100_, rst);
  and _46556_ (_39101_, _39018_, _38693_);
  nor _46557_ (_39102_, _39027_, _32458_);
  and _46558_ (_39103_, _39033_, _32567_);
  and _46559_ (_39104_, _39103_, _31282_);
  nor _46560_ (_39105_, _39103_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  not _46561_ (_39106_, _39105_);
  and _46562_ (_39107_, _39106_, _39038_);
  not _46563_ (_39108_, _39107_);
  nor _46564_ (_39109_, _39108_, _39104_);
  nor _46565_ (_39110_, _39109_, _39018_);
  not _46566_ (_39111_, _39110_);
  nor _46567_ (_39112_, _39111_, _39102_);
  nor _46568_ (_39113_, _39112_, _39101_);
  and _46569_ (_19860_, _39113_, _42882_);
  nor _46570_ (_39114_, _39027_, _33154_);
  and _46571_ (_39115_, _39033_, _33296_);
  and _46572_ (_39116_, _39115_, _31282_);
  nor _46573_ (_39117_, _39115_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  not _46574_ (_39118_, _39117_);
  and _46575_ (_39119_, _39118_, _39038_);
  not _46576_ (_39120_, _39119_);
  nor _46577_ (_39121_, _39120_, _39116_);
  or _46578_ (_39122_, _39121_, _39114_);
  and _46579_ (_39123_, _39122_, _39019_);
  nor _46580_ (_39124_, _39019_, _38724_);
  or _46581_ (_39125_, _39124_, _39123_);
  and _46582_ (_19872_, _39125_, _42882_);
  nor _46583_ (_39126_, _39027_, _33906_);
  not _46584_ (_39127_, _39033_);
  and _46585_ (_39133_, _39038_, _39127_);
  and _46586_ (_39144_, _39133_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  not _46587_ (_39145_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor _46588_ (_39146_, _34004_, _39145_);
  nor _46589_ (_39147_, _39146_, _34015_);
  nor _46590_ (_39158_, _39147_, _39094_);
  nor _46591_ (_39164_, _39158_, _39144_);
  and _46592_ (_39165_, _39164_, _39019_);
  not _46593_ (_39166_, _39165_);
  nor _46594_ (_39167_, _39166_, _39126_);
  and _46595_ (_39168_, _39018_, _38756_);
  or _46596_ (_39169_, _39168_, _39167_);
  nor _46597_ (_19884_, _39169_, rst);
  nor _46598_ (_39170_, _39027_, _34667_);
  and _46599_ (_39171_, _39033_, _34765_);
  and _46600_ (_39172_, _39171_, _31282_);
  nor _46601_ (_39173_, _39171_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  not _46602_ (_39174_, _39173_);
  and _46603_ (_39175_, _39174_, _39038_);
  not _46604_ (_39176_, _39175_);
  nor _46605_ (_39177_, _39176_, _39172_);
  or _46606_ (_39178_, _39177_, _39170_);
  and _46607_ (_39179_, _39178_, _39019_);
  nor _46608_ (_39180_, _39019_, _38787_);
  or _46609_ (_39181_, _39180_, _39179_);
  and _46610_ (_19896_, _39181_, _42882_);
  nor _46611_ (_39182_, _39027_, _35461_);
  and _46612_ (_39183_, _39033_, _35549_);
  and _46613_ (_39184_, _39183_, _31282_);
  nor _46614_ (_39185_, _39183_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not _46615_ (_39186_, _39185_);
  and _46616_ (_39187_, _39186_, _39038_);
  not _46617_ (_39188_, _39187_);
  nor _46618_ (_39189_, _39188_, _39184_);
  or _46619_ (_39190_, _39189_, _39182_);
  and _46620_ (_39191_, _39190_, _39019_);
  nor _46621_ (_39192_, _39019_, _38821_);
  or _46622_ (_39193_, _39192_, _39191_);
  and _46623_ (_19908_, _39193_, _42882_);
  nor _46624_ (_39194_, _39027_, _36179_);
  and _46625_ (_39195_, _39133_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _46626_ (_39196_, _39006_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor _46627_ (_39197_, _39196_, _39007_);
  nor _46628_ (_39198_, _39197_, _39094_);
  nor _46629_ (_39199_, _39198_, _39195_);
  and _46630_ (_39200_, _39199_, _39019_);
  not _46631_ (_39201_, _39200_);
  nor _46632_ (_39202_, _39201_, _39194_);
  nor _46633_ (_39203_, _39019_, _38847_);
  or _46634_ (_39204_, _39203_, _39202_);
  nor _46635_ (_19920_, _39204_, rst);
  and _46636_ (_39205_, _27374_, _27242_);
  and _46637_ (_39206_, _39049_, _39205_);
  and _46638_ (_39207_, _39206_, _31304_);
  nand _46639_ (_39208_, _39207_, _31282_);
  or _46640_ (_39209_, _39207_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _46641_ (_39210_, _39209_, _31348_);
  and _46642_ (_39211_, _39210_, _39208_);
  and _46643_ (_39212_, _38405_, _39022_);
  nand _46644_ (_39213_, _39212_, _38485_);
  or _46645_ (_39214_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _46646_ (_39215_, _39214_, _30679_);
  and _46647_ (_39216_, _39215_, _39213_);
  not _46648_ (_39217_, _30668_);
  and _46649_ (_39218_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or _46650_ (_39219_, _39218_, rst);
  or _46651_ (_39220_, _39219_, _39216_);
  or _46652_ (_31126_, _39220_, _39211_);
  and _46653_ (_39221_, _39205_, _27867_);
  and _46654_ (_39222_, _39221_, _31304_);
  nand _46655_ (_39223_, _39222_, _31282_);
  or _46656_ (_39224_, _39222_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _46657_ (_39225_, _39224_, _31348_);
  and _46658_ (_39226_, _39225_, _39223_);
  and _46659_ (_39227_, _38896_, _38404_);
  and _46660_ (_39228_, _39227_, _39022_);
  nand _46661_ (_39229_, _39228_, _38485_);
  or _46662_ (_39230_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _46663_ (_39231_, _39230_, _30679_);
  and _46664_ (_39232_, _39231_, _39229_);
  and _46665_ (_39233_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or _46666_ (_39234_, _39233_, rst);
  or _46667_ (_39235_, _39234_, _39232_);
  or _46668_ (_31149_, _39235_, _39226_);
  and _46669_ (_39236_, _38879_, _27242_);
  and _46670_ (_39237_, _39236_, _39049_);
  and _46671_ (_39238_, _39237_, _31304_);
  nand _46672_ (_39239_, _39238_, _31282_);
  or _46673_ (_39240_, _39238_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _46674_ (_39241_, _39240_, _31348_);
  and _46675_ (_39242_, _39241_, _39239_);
  and _46676_ (_39243_, _39023_, _38404_);
  and _46677_ (_39244_, _39243_, _39022_);
  not _46678_ (_39245_, _39244_);
  nor _46679_ (_39246_, _39245_, _38485_);
  and _46680_ (_39247_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _46681_ (_39248_, _39247_, _39246_);
  and _46682_ (_39249_, _39248_, _30679_);
  and _46683_ (_39250_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or _46684_ (_39251_, _39250_, rst);
  or _46685_ (_39252_, _39251_, _39249_);
  or _46686_ (_31172_, _39252_, _39242_);
  and _46687_ (_39253_, _39236_, _27867_);
  and _46688_ (_39254_, _39253_, _31304_);
  nand _46689_ (_39255_, _39254_, _31282_);
  or _46690_ (_39256_, _39254_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _46691_ (_39257_, _39256_, _31348_);
  and _46692_ (_39258_, _39257_, _39255_);
  nor _46693_ (_39259_, _27845_, _27374_);
  and _46694_ (_39260_, _38404_, _39259_);
  and _46695_ (_39261_, _39260_, _39022_);
  not _46696_ (_39262_, _39261_);
  nor _46697_ (_39263_, _39262_, _38485_);
  and _46698_ (_39264_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _46699_ (_39265_, _39264_, _39263_);
  and _46700_ (_39266_, _39265_, _30679_);
  and _46701_ (_39267_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or _46702_ (_39268_, _39267_, rst);
  or _46703_ (_39269_, _39268_, _39266_);
  or _46704_ (_31194_, _39269_, _39258_);
  or _46705_ (_39270_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _46706_ (_39271_, _39270_, _31348_);
  nand _46707_ (_39272_, _39212_, _31282_);
  and _46708_ (_39273_, _39272_, _39271_);
  nand _46709_ (_39274_, _39212_, _38464_);
  and _46710_ (_39275_, _39274_, _30679_);
  and _46711_ (_39276_, _39275_, _39270_);
  and _46712_ (_39277_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or _46713_ (_39278_, _39277_, rst);
  or _46714_ (_39279_, _39278_, _39276_);
  or _46715_ (_40589_, _39279_, _39273_);
  and _46716_ (_39280_, _32567_, _27703_);
  and _46717_ (_39281_, _39280_, _38405_);
  nand _46718_ (_39282_, _39281_, _31282_);
  or _46719_ (_39283_, _39281_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _46720_ (_39284_, _39283_, _31348_);
  and _46721_ (_39285_, _39284_, _39282_);
  nand _46722_ (_39286_, _39212_, _38456_);
  or _46723_ (_39287_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _46724_ (_39288_, _39287_, _30679_);
  and _46725_ (_39289_, _39288_, _39286_);
  and _46726_ (_39290_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _46727_ (_39291_, _39290_, rst);
  or _46728_ (_39292_, _39291_, _39289_);
  or _46729_ (_40591_, _39292_, _39285_);
  not _46730_ (_39293_, _34026_);
  nand _46731_ (_39294_, _39206_, _39293_);
  and _46732_ (_39295_, _39294_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _46733_ (_39296_, _33329_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _46734_ (_39297_, _39296_, _33318_);
  and _46735_ (_39298_, _39297_, _39206_);
  or _46736_ (_39299_, _39298_, _39295_);
  and _46737_ (_39300_, _39299_, _31348_);
  nand _46738_ (_39301_, _39212_, _38449_);
  or _46739_ (_39302_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _46740_ (_39303_, _39302_, _30679_);
  and _46741_ (_39304_, _39303_, _39301_);
  and _46742_ (_39305_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _46743_ (_39306_, _39305_, rst);
  or _46744_ (_39307_, _39306_, _39304_);
  or _46745_ (_40593_, _39307_, _39300_);
  nand _46746_ (_39308_, _39206_, _26781_);
  and _46747_ (_39309_, _39308_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _46748_ (_39310_, _39293_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _46749_ (_39311_, _39310_, _34015_);
  and _46750_ (_39312_, _39311_, _39206_);
  or _46751_ (_39313_, _39312_, _39309_);
  and _46752_ (_39314_, _39313_, _31348_);
  nand _46753_ (_39315_, _39212_, _38442_);
  or _46754_ (_39316_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _46755_ (_39317_, _39316_, _30679_);
  and _46756_ (_39318_, _39317_, _39315_);
  and _46757_ (_39319_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _46758_ (_39320_, _39319_, rst);
  or _46759_ (_39321_, _39320_, _39318_);
  or _46760_ (_40595_, _39321_, _39314_);
  not _46761_ (_39322_, _39206_);
  or _46762_ (_39323_, _39322_, _34787_);
  and _46763_ (_39324_, _39323_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _46764_ (_39325_, _34776_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _46765_ (_39326_, _39325_, _34819_);
  and _46766_ (_39327_, _39326_, _39206_);
  or _46767_ (_39328_, _39327_, _39324_);
  and _46768_ (_39329_, _39328_, _31348_);
  nand _46769_ (_39330_, _39212_, _38434_);
  or _46770_ (_39331_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _46771_ (_39332_, _39331_, _30679_);
  and _46772_ (_39333_, _39332_, _39330_);
  and _46773_ (_39334_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or _46774_ (_39335_, _39334_, rst);
  or _46775_ (_39336_, _39335_, _39333_);
  or _46776_ (_40597_, _39336_, _39329_);
  and _46777_ (_39337_, _39206_, _35549_);
  nand _46778_ (_39338_, _39337_, _31282_);
  or _46779_ (_39347_, _39337_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _46780_ (_39358_, _39347_, _31348_);
  and _46781_ (_39369_, _39358_, _39338_);
  nand _46782_ (_39378_, _39212_, _38428_);
  or _46783_ (_39384_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _46784_ (_39395_, _39384_, _30679_);
  and _46785_ (_39406_, _39395_, _39378_);
  and _46786_ (_39417_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or _46787_ (_39428_, _39417_, rst);
  or _46788_ (_39439_, _39428_, _39406_);
  or _46789_ (_40599_, _39439_, _39369_);
  and _46790_ (_39460_, _39206_, _36277_);
  nand _46791_ (_39471_, _39460_, _31282_);
  or _46792_ (_39482_, _39460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _46793_ (_39493_, _39482_, _31348_);
  and _46794_ (_39504_, _39493_, _39471_);
  nand _46795_ (_39515_, _39212_, _38420_);
  or _46796_ (_39526_, _39212_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _46797_ (_39537_, _39526_, _30679_);
  and _46798_ (_39548_, _39537_, _39515_);
  and _46799_ (_39552_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _46800_ (_39553_, _39552_, rst);
  or _46801_ (_39554_, _39553_, _39548_);
  or _46802_ (_40601_, _39554_, _39504_);
  and _46803_ (_39555_, _39221_, _27045_);
  nand _46804_ (_39556_, _39555_, _31282_);
  or _46805_ (_39557_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _46806_ (_39558_, _39557_, _31348_);
  and _46807_ (_39559_, _39558_, _39556_);
  nand _46808_ (_39560_, _39228_, _38464_);
  and _46809_ (_39561_, _39560_, _30679_);
  and _46810_ (_39562_, _39561_, _39557_);
  and _46811_ (_39563_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or _46812_ (_39564_, _39563_, rst);
  or _46813_ (_39565_, _39564_, _39562_);
  or _46814_ (_40603_, _39565_, _39559_);
  and _46815_ (_39566_, _39221_, _32567_);
  nand _46816_ (_39567_, _39566_, _31282_);
  or _46817_ (_39568_, _39566_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _46818_ (_39569_, _39568_, _31348_);
  and _46819_ (_39570_, _39569_, _39567_);
  nand _46820_ (_39571_, _39228_, _38456_);
  or _46821_ (_39572_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _46822_ (_39573_, _39572_, _30679_);
  and _46823_ (_39574_, _39573_, _39571_);
  and _46824_ (_39575_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _46825_ (_39576_, _39575_, rst);
  or _46826_ (_39577_, _39576_, _39574_);
  or _46827_ (_40605_, _39577_, _39570_);
  and _46828_ (_39578_, _39221_, _33296_);
  nand _46829_ (_39579_, _39578_, _31282_);
  or _46830_ (_39580_, _39578_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _46831_ (_39581_, _39580_, _31348_);
  and _46832_ (_39582_, _39581_, _39579_);
  nand _46833_ (_39583_, _39228_, _38449_);
  or _46834_ (_39584_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _46835_ (_39585_, _39584_, _30679_);
  and _46836_ (_39586_, _39585_, _39583_);
  and _46837_ (_39587_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or _46838_ (_39588_, _39587_, rst);
  or _46839_ (_39589_, _39588_, _39586_);
  or _46840_ (_40607_, _39589_, _39582_);
  and _46841_ (_39590_, _39221_, _34004_);
  nand _46842_ (_39591_, _39590_, _31282_);
  or _46843_ (_39592_, _39590_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _46844_ (_39593_, _39592_, _31348_);
  and _46845_ (_39594_, _39593_, _39591_);
  nand _46846_ (_39595_, _39228_, _38442_);
  or _46847_ (_39596_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _46848_ (_39597_, _39596_, _30679_);
  and _46849_ (_39598_, _39597_, _39595_);
  and _46850_ (_39599_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _46851_ (_39600_, _39599_, rst);
  or _46852_ (_39601_, _39600_, _39598_);
  or _46853_ (_40609_, _39601_, _39594_);
  and _46854_ (_39602_, _39221_, _34765_);
  nand _46855_ (_39603_, _39602_, _31282_);
  or _46856_ (_39604_, _39602_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _46857_ (_39605_, _39604_, _31348_);
  and _46858_ (_39606_, _39605_, _39603_);
  nand _46859_ (_39607_, _39228_, _38434_);
  or _46860_ (_39608_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _46861_ (_39609_, _39608_, _30679_);
  and _46862_ (_39610_, _39609_, _39607_);
  and _46863_ (_39611_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or _46864_ (_39612_, _39611_, rst);
  or _46865_ (_39613_, _39612_, _39610_);
  or _46866_ (_40611_, _39613_, _39606_);
  and _46867_ (_39614_, _39221_, _35549_);
  nand _46868_ (_39615_, _39614_, _31282_);
  or _46869_ (_39616_, _39614_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _46870_ (_39617_, _39616_, _31348_);
  and _46871_ (_39618_, _39617_, _39615_);
  nand _46872_ (_39619_, _39228_, _38428_);
  or _46873_ (_39620_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _46874_ (_39621_, _39620_, _30679_);
  and _46875_ (_39622_, _39621_, _39619_);
  and _46876_ (_39623_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or _46877_ (_39624_, _39623_, rst);
  or _46878_ (_39625_, _39624_, _39622_);
  or _46879_ (_40612_, _39625_, _39618_);
  and _46880_ (_39626_, _39221_, _36277_);
  nand _46881_ (_39627_, _39626_, _31282_);
  or _46882_ (_39628_, _39626_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _46883_ (_39629_, _39628_, _31348_);
  and _46884_ (_39630_, _39629_, _39627_);
  nand _46885_ (_39631_, _39228_, _38420_);
  or _46886_ (_39632_, _39228_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _46887_ (_39633_, _39632_, _30679_);
  and _46888_ (_39634_, _39633_, _39631_);
  and _46889_ (_39635_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _46890_ (_39636_, _39635_, rst);
  or _46891_ (_39637_, _39636_, _39634_);
  or _46892_ (_40614_, _39637_, _39630_);
  nand _46893_ (_39638_, _39244_, _31282_);
  or _46894_ (_39639_, _39244_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _46895_ (_39640_, _39639_, _31348_);
  and _46896_ (_39641_, _39640_, _39638_);
  and _46897_ (_39642_, _39244_, _38465_);
  and _46898_ (_39643_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _46899_ (_39644_, _39643_, _39642_);
  and _46900_ (_39645_, _39644_, _30679_);
  and _46901_ (_39646_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or _46902_ (_39647_, _39646_, rst);
  or _46903_ (_39648_, _39647_, _39645_);
  or _46904_ (_40616_, _39648_, _39641_);
  and _46905_ (_39649_, _39237_, _32567_);
  nand _46906_ (_39650_, _39649_, _31282_);
  or _46907_ (_39651_, _39649_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _46908_ (_39652_, _39651_, _31348_);
  and _46909_ (_39653_, _39652_, _39650_);
  nor _46910_ (_39654_, _39245_, _38456_);
  and _46911_ (_39655_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _46912_ (_39656_, _39655_, _39654_);
  and _46913_ (_39657_, _39656_, _30679_);
  and _46914_ (_39658_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _46915_ (_39659_, _39658_, rst);
  or _46916_ (_39660_, _39659_, _39657_);
  or _46917_ (_40618_, _39660_, _39653_);
  and _46918_ (_39661_, _39237_, _33296_);
  nand _46919_ (_39662_, _39661_, _31282_);
  or _46920_ (_39663_, _39661_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _46921_ (_39664_, _39663_, _31348_);
  and _46922_ (_39665_, _39664_, _39662_);
  nor _46923_ (_39666_, _39245_, _38449_);
  and _46924_ (_39667_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _46925_ (_39668_, _39667_, _39666_);
  and _46926_ (_39669_, _39668_, _30679_);
  and _46927_ (_39670_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _46928_ (_39671_, _39670_, rst);
  or _46929_ (_39672_, _39671_, _39669_);
  or _46930_ (_40620_, _39672_, _39665_);
  and _46931_ (_39673_, _39237_, _34004_);
  nand _46932_ (_39674_, _39673_, _31282_);
  or _46933_ (_39675_, _39673_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _46934_ (_39676_, _39675_, _31348_);
  and _46935_ (_39677_, _39676_, _39674_);
  nor _46936_ (_39678_, _39245_, _38442_);
  and _46937_ (_39679_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _46938_ (_39680_, _39679_, _39678_);
  and _46939_ (_39681_, _39680_, _30679_);
  and _46940_ (_39682_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _46941_ (_39683_, _39682_, rst);
  or _46942_ (_39684_, _39683_, _39681_);
  or _46943_ (_40622_, _39684_, _39677_);
  and _46944_ (_39685_, _39237_, _34765_);
  nand _46945_ (_39686_, _39685_, _31282_);
  or _46946_ (_39687_, _39685_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _46947_ (_39688_, _39687_, _31348_);
  and _46948_ (_39689_, _39688_, _39686_);
  nor _46949_ (_39690_, _39245_, _38434_);
  and _46950_ (_39691_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _46951_ (_39692_, _39691_, _39690_);
  and _46952_ (_39693_, _39692_, _30679_);
  and _46953_ (_39694_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or _46954_ (_39695_, _39694_, rst);
  or _46955_ (_39696_, _39695_, _39693_);
  or _46956_ (_40624_, _39696_, _39689_);
  and _46957_ (_39697_, _39237_, _35549_);
  nand _46958_ (_39698_, _39697_, _31282_);
  or _46959_ (_39699_, _39697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _46960_ (_39700_, _39699_, _31348_);
  and _46961_ (_39701_, _39700_, _39698_);
  nor _46962_ (_39702_, _39245_, _38428_);
  and _46963_ (_39703_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _46964_ (_39704_, _39703_, _39702_);
  and _46965_ (_39705_, _39704_, _30679_);
  and _46966_ (_39706_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _46967_ (_39707_, _39706_, rst);
  or _46968_ (_39708_, _39707_, _39705_);
  or _46969_ (_40626_, _39708_, _39701_);
  and _46970_ (_39709_, _39237_, _36277_);
  nand _46971_ (_39710_, _39709_, _31282_);
  or _46972_ (_39711_, _39709_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _46973_ (_39712_, _39711_, _31348_);
  and _46974_ (_39713_, _39712_, _39710_);
  nor _46975_ (_39714_, _39245_, _38420_);
  and _46976_ (_39715_, _39245_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _46977_ (_39716_, _39715_, _39714_);
  and _46978_ (_39717_, _39716_, _30679_);
  and _46979_ (_39718_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _46980_ (_39719_, _39718_, rst);
  or _46981_ (_39720_, _39719_, _39717_);
  or _46982_ (_40628_, _39720_, _39713_);
  and _46983_ (_39721_, _39253_, _27045_);
  nand _46984_ (_39722_, _39721_, _31282_);
  or _46985_ (_39723_, _39721_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _46986_ (_39724_, _39723_, _31348_);
  and _46987_ (_39725_, _39724_, _39722_);
  and _46988_ (_39726_, _39261_, _38465_);
  and _46989_ (_39727_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _46990_ (_39728_, _39727_, _39726_);
  and _46991_ (_39729_, _39728_, _30679_);
  and _46992_ (_39730_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or _46993_ (_39731_, _39730_, rst);
  or _46994_ (_39732_, _39731_, _39729_);
  or _46995_ (_40630_, _39732_, _39725_);
  and _46996_ (_39733_, _39253_, _32567_);
  nand _46997_ (_39734_, _39733_, _31282_);
  or _46998_ (_39735_, _39733_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _46999_ (_39736_, _39735_, _31348_);
  and _47000_ (_39737_, _39736_, _39734_);
  nor _47001_ (_39738_, _39262_, _38456_);
  and _47002_ (_39739_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _47003_ (_39740_, _39739_, _39738_);
  and _47004_ (_39741_, _39740_, _30679_);
  and _47005_ (_39742_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _47006_ (_39743_, _39742_, rst);
  or _47007_ (_39744_, _39743_, _39741_);
  or _47008_ (_40632_, _39744_, _39737_);
  and _47009_ (_39745_, _39253_, _33296_);
  nand _47010_ (_39746_, _39745_, _31282_);
  or _47011_ (_39747_, _39745_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _47012_ (_39748_, _39747_, _31348_);
  and _47013_ (_39749_, _39748_, _39746_);
  nor _47014_ (_39750_, _39262_, _38449_);
  and _47015_ (_39751_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _47016_ (_39752_, _39751_, _39750_);
  and _47017_ (_39753_, _39752_, _30679_);
  and _47018_ (_39754_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or _47019_ (_39755_, _39754_, rst);
  or _47020_ (_39756_, _39755_, _39753_);
  or _47021_ (_40634_, _39756_, _39749_);
  and _47022_ (_39757_, _39253_, _34004_);
  nand _47023_ (_39758_, _39757_, _31282_);
  or _47024_ (_39759_, _39757_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _47025_ (_39761_, _39759_, _31348_);
  and _47026_ (_39766_, _39761_, _39758_);
  nor _47027_ (_39767_, _39262_, _38442_);
  and _47028_ (_39768_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _47029_ (_39769_, _39768_, _39767_);
  and _47030_ (_39770_, _39769_, _30679_);
  and _47031_ (_39771_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _47032_ (_39772_, _39771_, rst);
  or _47033_ (_39773_, _39772_, _39770_);
  or _47034_ (_40636_, _39773_, _39766_);
  and _47035_ (_39774_, _39253_, _34765_);
  nand _47036_ (_39775_, _39774_, _31282_);
  or _47037_ (_39776_, _39774_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _47038_ (_39777_, _39776_, _31348_);
  and _47039_ (_39778_, _39777_, _39775_);
  nor _47040_ (_39779_, _39262_, _38434_);
  and _47041_ (_39780_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _47042_ (_39781_, _39780_, _39779_);
  and _47043_ (_39782_, _39781_, _30679_);
  and _47044_ (_39783_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or _47045_ (_39784_, _39783_, rst);
  or _47046_ (_39785_, _39784_, _39782_);
  or _47047_ (_40638_, _39785_, _39778_);
  and _47048_ (_39786_, _39253_, _35549_);
  nand _47049_ (_39787_, _39786_, _31282_);
  or _47050_ (_39788_, _39786_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _47051_ (_39789_, _39788_, _31348_);
  and _47052_ (_39790_, _39789_, _39787_);
  nor _47053_ (_39791_, _39262_, _38428_);
  and _47054_ (_39802_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _47055_ (_39813_, _39802_, _39791_);
  and _47056_ (_39822_, _39813_, _30679_);
  and _47057_ (_39823_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or _47058_ (_39824_, _39823_, rst);
  or _47059_ (_39825_, _39824_, _39822_);
  or _47060_ (_40640_, _39825_, _39790_);
  and _47061_ (_39826_, _39253_, _36277_);
  nand _47062_ (_39827_, _39826_, _31282_);
  or _47063_ (_39828_, _39826_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _47064_ (_39829_, _39828_, _31348_);
  and _47065_ (_39830_, _39829_, _39827_);
  nor _47066_ (_39831_, _39262_, _38420_);
  and _47067_ (_39832_, _39262_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _47068_ (_39833_, _39832_, _39831_);
  and _47069_ (_39834_, _39833_, _30679_);
  and _47070_ (_39835_, _39217_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _47071_ (_39836_, _39835_, rst);
  or _47072_ (_39837_, _39836_, _39834_);
  or _47073_ (_40642_, _39837_, _39830_);
  and _47074_ (_41092_, t0_i, _42882_);
  and _47075_ (_41095_, t1_i, _42882_);
  not _47076_ (_39838_, _30679_);
  nor _47077_ (_39839_, _39838_, _27703_);
  and _47078_ (_39840_, _39839_, _34004_);
  and _47079_ (_39841_, _39840_, _38405_);
  nand _47080_ (_39842_, _39841_, _38485_);
  nor _47081_ (_39843_, _26781_, _27703_);
  and _47082_ (_39844_, _39843_, _38406_);
  and _47083_ (_39845_, _39844_, _30679_);
  not _47084_ (_39846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _47085_ (_39847_, _39846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _47086_ (_39848_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _47087_ (_39852_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _39848_);
  nor _47088_ (_39856_, _39852_, _39847_);
  nor _47089_ (_39857_, _39856_, _39845_);
  not _47090_ (_39858_, _39857_);
  and _47091_ (_39859_, _39858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not _47092_ (_39860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not _47093_ (_39861_, t1_i);
  and _47094_ (_39862_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _39861_);
  nor _47095_ (_39863_, _39862_, _39860_);
  not _47096_ (_39864_, _39863_);
  not _47097_ (_39865_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _47098_ (_39866_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _39865_);
  nor _47099_ (_39867_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _47100_ (_39868_, _39867_);
  and _47101_ (_39869_, _39868_, _39866_);
  and _47102_ (_39870_, _39869_, _39864_);
  not _47103_ (_39871_, _39870_);
  nand _47104_ (_39872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand _47105_ (_39873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or _47106_ (_39874_, _39873_, _39872_);
  nor _47107_ (_39875_, _39874_, _39871_);
  and _47108_ (_39876_, _39875_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _47109_ (_39877_, _39876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _47110_ (_39878_, _39877_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _47111_ (_39879_, _39878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not _47112_ (_39880_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _47113_ (_39881_, _39874_, _39880_);
  and _47114_ (_39882_, _39881_, _39870_);
  and _47115_ (_39883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _47116_ (_39884_, _39883_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _47117_ (_39885_, _39884_, _39882_);
  nor _47118_ (_39886_, _39885_, _39856_);
  and _47119_ (_39887_, _39886_, _39879_);
  and _47120_ (_39888_, _39885_, _39847_);
  and _47121_ (_39889_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47122_ (_39890_, _39889_, _39887_);
  nor _47123_ (_39891_, _39890_, _39845_);
  or _47124_ (_39892_, _39891_, _39859_);
  or _47125_ (_39893_, _39841_, _39892_);
  and _47126_ (_39894_, _39893_, _42882_);
  and _47127_ (_41098_, _39894_, _39842_);
  nand _47128_ (_39895_, _39845_, _38485_);
  and _47129_ (_39896_, _39839_, _38623_);
  not _47130_ (_39897_, _39896_);
  and _47131_ (_39898_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _47132_ (_39899_, _39898_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _47133_ (_39900_, _39884_, _39881_);
  and _47134_ (_39901_, _39900_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _47135_ (_39902_, _39901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _47136_ (_39903_, _39902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _47137_ (_39904_, _39903_, _39870_);
  and _47138_ (_39905_, _39904_, _39899_);
  and _47139_ (_39906_, _39905_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47140_ (_39907_, _39906_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47141_ (_39908_, _39906_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47142_ (_39909_, _39908_, _39907_);
  and _47143_ (_39910_, _39909_, _39852_);
  and _47144_ (_39911_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _47145_ (_39912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _47146_ (_39913_, _39912_, _39881_);
  and _47147_ (_39914_, _39913_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _47148_ (_39915_, _39914_, _39870_);
  and _47149_ (_39916_, _39915_, _39899_);
  and _47150_ (_39917_, _39916_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47151_ (_39918_, _39917_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor _47152_ (_39919_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _47153_ (_39920_, _39917_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _47154_ (_39921_, _39920_, _39919_);
  nor _47155_ (_39922_, _39921_, _39918_);
  or _47156_ (_39923_, _39922_, _39911_);
  or _47157_ (_39924_, _39923_, _39910_);
  or _47158_ (_39925_, _39924_, _39845_);
  and _47159_ (_39926_, _39925_, _39897_);
  and _47160_ (_39927_, _39926_, _39895_);
  and _47161_ (_39928_, _39896_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _47162_ (_39929_, _39928_, _39927_);
  and _47163_ (_41101_, _39929_, _42882_);
  not _47164_ (_39930_, _39845_);
  and _47165_ (_39931_, _39871_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  or _47166_ (_39932_, _39931_, _39907_);
  and _47167_ (_39933_, _39932_, _39852_);
  or _47168_ (_39934_, _39931_, _39918_);
  and _47169_ (_39942_, _39934_, _39919_);
  nand _47170_ (_39946_, _39870_, _39846_);
  and _47171_ (_39947_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  and _47172_ (_39948_, _39947_, _39946_);
  or _47173_ (_39949_, _39948_, _39888_);
  or _47174_ (_39950_, _39949_, _39942_);
  or _47175_ (_39951_, _39950_, _39933_);
  nor _47176_ (_39952_, _39896_, rst);
  and _47177_ (_39953_, _39952_, _39951_);
  and _47178_ (_41104_, _39953_, _39930_);
  and _47179_ (_39954_, _39839_, _34765_);
  and _47180_ (_39955_, _39954_, _38405_);
  nor _47181_ (_39956_, _39955_, rst);
  and _47182_ (_39957_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47183_ (_39958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _47184_ (_39959_, _39958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47185_ (_39960_, _39959_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47186_ (_39961_, _39960_, _39957_);
  and _47187_ (_39962_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _47188_ (_39963_, _39962_, _39961_);
  or _47189_ (_39964_, _39963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _47190_ (_39965_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _47191_ (_39966_, _39965_);
  and _47192_ (_39967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _47193_ (_39968_, _39967_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not _47194_ (_39969_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not _47195_ (_39970_, t0_i);
  and _47196_ (_39971_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _39970_);
  nor _47197_ (_39972_, _39971_, _39969_);
  not _47198_ (_39973_, _39972_);
  not _47199_ (_39974_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor _47200_ (_39975_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor _47201_ (_39976_, _39975_, _39974_);
  and _47202_ (_39977_, _39976_, _39973_);
  and _47203_ (_39978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _47204_ (_39979_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _47205_ (_39980_, _39979_, _39978_);
  and _47206_ (_39981_, _39980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _47207_ (_39982_, _39981_, _39977_);
  and _47208_ (_39983_, _39982_, _39968_);
  and _47209_ (_39984_, _39983_, _39966_);
  and _47210_ (_39985_, _39984_, _39964_);
  not _47211_ (_39986_, _39977_);
  and _47212_ (_39987_, _39986_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  and _47213_ (_39988_, _39982_, _39961_);
  and _47214_ (_39989_, _39988_, _39962_);
  and _47215_ (_39990_, _39989_, _39965_);
  or _47216_ (_39991_, _39990_, _39987_);
  nor _47217_ (_39992_, _39991_, _39985_);
  and _47218_ (_39993_, _39839_, _33296_);
  and _47219_ (_39994_, _39993_, _38405_);
  nor _47220_ (_39995_, _39994_, _39992_);
  and _47221_ (_41107_, _39995_, _39956_);
  and _47222_ (_39996_, _39839_, _38630_);
  nand _47223_ (_39997_, _39996_, _38485_);
  not _47224_ (_39998_, _39955_);
  or _47225_ (_39999_, _39998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _47226_ (_40000_, _39965_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _47227_ (_40001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _47228_ (_40002_, _40001_, _39982_);
  or _47229_ (_40003_, _40002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not _47230_ (_40004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _47231_ (_40005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _40004_);
  nand _47232_ (_40006_, _40005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _47233_ (_40007_, _40006_, _39983_);
  and _47234_ (_40008_, _40007_, _39966_);
  or _47235_ (_40009_, _40008_, _39955_);
  and _47236_ (_40010_, _40009_, _40003_);
  or _47237_ (_40011_, _40010_, _40000_);
  and _47238_ (_40012_, _40011_, _39999_);
  or _47239_ (_40013_, _40012_, _39996_);
  and _47240_ (_40014_, _40013_, _42882_);
  and _47241_ (_41110_, _40014_, _39997_);
  nand _47242_ (_40017_, _39955_, _38485_);
  not _47243_ (_40020_, _39994_);
  and _47244_ (_40021_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _40004_);
  or _47245_ (_40022_, _40005_, _40021_);
  not _47246_ (_40023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _47247_ (_40024_, _39981_, _39968_);
  and _47248_ (_40025_, _39977_, _40004_);
  and _47249_ (_40026_, _40025_, _40024_);
  and _47250_ (_40027_, _40026_, _39961_);
  and _47251_ (_40028_, _40027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _47252_ (_40029_, _40028_, _40023_);
  and _47253_ (_40030_, _40028_, _40023_);
  or _47254_ (_40031_, _40030_, _40029_);
  and _47255_ (_40032_, _40031_, _40022_);
  and _47256_ (_40033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47257_ (_40034_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _47258_ (_40035_, _40034_, _39960_);
  and _47259_ (_40038_, _40035_, _39957_);
  and _47260_ (_40046_, _40038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _47261_ (_40047_, _40046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _47262_ (_40048_, _40034_, _39963_);
  and _47263_ (_40049_, _40048_, _40047_);
  and _47264_ (_40050_, _40049_, _40033_);
  and _47265_ (_40051_, _39988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _47266_ (_40052_, _40051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _47267_ (_40053_, _39989_, _39966_);
  and _47268_ (_40054_, _40053_, _40052_);
  or _47269_ (_40055_, _40054_, _40050_);
  or _47270_ (_40056_, _40055_, _40032_);
  or _47271_ (_40057_, _40056_, _39955_);
  and _47272_ (_40058_, _40057_, _40020_);
  and _47273_ (_40059_, _40058_, _40017_);
  and _47274_ (_40060_, _39994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _47275_ (_40061_, _40060_, _40059_);
  and _47276_ (_41113_, _40061_, _42882_);
  and _47277_ (_40062_, _27023_, _33274_);
  nor _47278_ (_40063_, _31283_, _27703_);
  and _47279_ (_40064_, _40063_, _40062_);
  nand _47280_ (_40065_, _40064_, _38405_);
  or _47281_ (_40066_, _40065_, _39838_);
  not _47282_ (_40067_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  or _47283_ (_40068_, _40034_, _40067_);
  nand _47284_ (_40069_, _40068_, _40048_);
  nand _47285_ (_40070_, _40069_, _40033_);
  nor _47286_ (_40071_, _40070_, _39955_);
  and _47287_ (_40072_, _40071_, _40066_);
  and _47288_ (_41116_, _40072_, _42882_);
  and _47289_ (_40073_, _40063_, _38406_);
  and _47290_ (_40074_, _40073_, _30679_);
  or _47291_ (_40075_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _47292_ (_40076_, _40075_, _42882_);
  nand _47293_ (_40077_, _40074_, _38485_);
  and _47294_ (_41119_, _40077_, _40076_);
  not _47295_ (_40078_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _47296_ (_40079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _47297_ (_40080_, _40079_, _39845_);
  and _47298_ (_40081_, _40080_, _39870_);
  nor _47299_ (_40082_, _40081_, _40078_);
  and _47300_ (_40083_, _40081_, _40078_);
  or _47301_ (_40084_, _40083_, _40082_);
  nand _47302_ (_40085_, _39901_, _39847_);
  nor _47303_ (_40086_, _40085_, _39845_);
  or _47304_ (_40087_, _40086_, _39841_);
  or _47305_ (_40088_, _40087_, _40084_);
  nand _47306_ (_40089_, _39841_, _38464_);
  and _47307_ (_40090_, _40089_, _42882_);
  and _47308_ (_41601_, _40090_, _40088_);
  and _47309_ (_40091_, _39870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _47310_ (_40092_, _40091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _47311_ (_40093_, _40091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _47312_ (_40094_, _40093_, _40092_);
  nand _47313_ (_40095_, _40094_, _40080_);
  or _47314_ (_40096_, _40080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _47315_ (_40097_, _40096_, _40095_);
  nand _47316_ (_40098_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _47317_ (_40099_, _40098_, _39845_);
  or _47318_ (_40100_, _40099_, _39896_);
  or _47319_ (_40101_, _40100_, _40097_);
  nand _47320_ (_40102_, _39896_, _38456_);
  and _47321_ (_40103_, _40102_, _42882_);
  and _47322_ (_41603_, _40103_, _40101_);
  not _47323_ (_40104_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _47324_ (_40105_, _40080_, _40104_);
  nand _47325_ (_40106_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _47326_ (_40107_, _40106_, _39845_);
  or _47327_ (_40108_, _40107_, _40105_);
  nor _47328_ (_40109_, _40092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _47329_ (_40110_, _40092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _47330_ (_40111_, _40110_, _40109_);
  and _47331_ (_40112_, _40111_, _40080_);
  or _47332_ (_40113_, _40112_, _39841_);
  or _47333_ (_40114_, _40113_, _40108_);
  nand _47334_ (_40115_, _39841_, _38449_);
  and _47335_ (_40116_, _40115_, _42882_);
  and _47336_ (_41605_, _40116_, _40114_);
  not _47337_ (_40117_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _47338_ (_40118_, _40080_, _40117_);
  or _47339_ (_40119_, _40110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _47340_ (_40120_, _40079_, _39875_);
  and _47341_ (_40121_, _40120_, _40119_);
  and _47342_ (_40122_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _47343_ (_40123_, _40122_, _40121_);
  nor _47344_ (_40124_, _40123_, _39845_);
  or _47345_ (_40125_, _40124_, _40118_);
  and _47346_ (_40126_, _40125_, _39897_);
  nor _47347_ (_40127_, _39897_, _38442_);
  or _47348_ (_40128_, _40127_, _40126_);
  and _47349_ (_41606_, _40128_, _42882_);
  nor _47350_ (_40129_, _39875_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor _47351_ (_40130_, _40129_, _39882_);
  and _47352_ (_40131_, _40130_, _40080_);
  nor _47353_ (_40132_, _40080_, _39880_);
  nand _47354_ (_40133_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _47355_ (_40134_, _40133_, _39845_);
  or _47356_ (_40135_, _40134_, _40132_);
  or _47357_ (_40136_, _40135_, _40131_);
  or _47358_ (_40137_, _40136_, _39841_);
  nand _47359_ (_40138_, _39841_, _38434_);
  and _47360_ (_40139_, _40138_, _42882_);
  and _47361_ (_41608_, _40139_, _40137_);
  nand _47362_ (_40140_, _39841_, _38428_);
  and _47363_ (_40141_, _39882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _47364_ (_40142_, _39882_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor _47365_ (_40143_, _40142_, _40141_);
  and _47366_ (_40144_, _40143_, _39857_);
  and _47367_ (_40145_, _39858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nand _47368_ (_40146_, _39888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _47369_ (_40147_, _40146_, _39845_);
  or _47370_ (_40148_, _40147_, _40145_);
  or _47371_ (_40149_, _40148_, _40144_);
  or _47372_ (_40150_, _40149_, _39841_);
  and _47373_ (_40151_, _40150_, _42882_);
  and _47374_ (_41610_, _40151_, _40140_);
  nand _47375_ (_40152_, _39841_, _38420_);
  and _47376_ (_40153_, _39858_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _47377_ (_40154_, _39847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47378_ (_40155_, _40154_, _39870_);
  and _47379_ (_40156_, _40155_, _39900_);
  nor _47380_ (_40157_, _40141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _47381_ (_40158_, _40157_, _39856_);
  nor _47382_ (_40159_, _40158_, _39878_);
  nor _47383_ (_40160_, _40159_, _40156_);
  nor _47384_ (_40161_, _40160_, _39845_);
  or _47385_ (_40162_, _40161_, _40153_);
  or _47386_ (_40163_, _40162_, _39841_);
  and _47387_ (_40164_, _40163_, _42882_);
  and _47388_ (_41612_, _40164_, _40152_);
  nand _47389_ (_40165_, _39845_, _38464_);
  not _47390_ (_40166_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _47391_ (_40167_, _39882_, _39848_);
  nor _47392_ (_40168_, _39884_, _39846_);
  not _47393_ (_40169_, _40168_);
  and _47394_ (_40170_, _40169_, _40167_);
  nor _47395_ (_40171_, _40170_, _40166_);
  and _47396_ (_40172_, _40170_, _40166_);
  or _47397_ (_40173_, _40172_, _40171_);
  or _47398_ (_40174_, _40173_, _39845_);
  and _47399_ (_40175_, _40174_, _40165_);
  or _47400_ (_40176_, _40175_, _39896_);
  nand _47401_ (_40177_, _39896_, _40166_);
  and _47402_ (_40178_, _40177_, _42882_);
  and _47403_ (_41614_, _40178_, _40176_);
  not _47404_ (_40179_, _39852_);
  nor _47405_ (_40180_, _39885_, _40179_);
  not _47406_ (_40181_, _40180_);
  nor _47407_ (_40182_, _40167_, _39852_);
  nor _47408_ (_40183_, _40182_, _40166_);
  and _47409_ (_40184_, _40183_, _40181_);
  or _47410_ (_40185_, _40184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand _47411_ (_40186_, _40184_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _47412_ (_40187_, _40186_, _40185_);
  or _47413_ (_40188_, _40187_, _39845_);
  nand _47414_ (_40189_, _39845_, _38456_);
  and _47415_ (_40190_, _40189_, _40188_);
  or _47416_ (_40191_, _40190_, _39896_);
  or _47417_ (_40192_, _39897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _47418_ (_40193_, _40192_, _42882_);
  and _47419_ (_41616_, _40193_, _40191_);
  nand _47420_ (_40194_, _39845_, _38449_);
  and _47421_ (_40195_, _39912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _47422_ (_40196_, _40195_, _39882_);
  and _47423_ (_40197_, _40196_, _39848_);
  nand _47424_ (_40198_, _40197_, _40169_);
  and _47425_ (_40199_, _40198_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _47426_ (_40200_, _40168_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _47427_ (_40201_, _40200_);
  not _47428_ (_40202_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _47429_ (_40203_, _39912_, _40202_);
  and _47430_ (_40204_, _40203_, _39882_);
  and _47431_ (_40205_, _40204_, _40201_);
  or _47432_ (_40206_, _40205_, _40199_);
  or _47433_ (_40207_, _40206_, _39845_);
  and _47434_ (_40208_, _40207_, _40194_);
  or _47435_ (_40209_, _40208_, _39896_);
  nand _47436_ (_40210_, _39896_, _40202_);
  and _47437_ (_40211_, _40210_, _42882_);
  and _47438_ (_41618_, _40211_, _40209_);
  nand _47439_ (_40212_, _39845_, _38442_);
  nor _47440_ (_40213_, _39904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _47441_ (_40214_, _40196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _47442_ (_40215_, _40214_, _39884_);
  nor _47443_ (_40216_, _40215_, _40213_);
  or _47444_ (_40217_, _40216_, _40179_);
  not _47445_ (_40218_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _47446_ (_40219_, _40197_, _40218_);
  nor _47447_ (_40220_, _40197_, _40218_);
  or _47448_ (_40221_, _40220_, _39852_);
  or _47449_ (_40222_, _40221_, _40219_);
  and _47450_ (_40223_, _40222_, _40217_);
  or _47451_ (_40224_, _40223_, _39845_);
  and _47452_ (_40225_, _40224_, _40212_);
  or _47453_ (_40226_, _40225_, _39896_);
  nand _47454_ (_40227_, _39896_, _40218_);
  and _47455_ (_40228_, _40227_, _42882_);
  and _47456_ (_41620_, _40228_, _40226_);
  nand _47457_ (_40229_, _39845_, _38434_);
  and _47458_ (_40230_, _39904_, _39898_);
  or _47459_ (_40231_, _40215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _47460_ (_40232_, _40231_, _39852_);
  nor _47461_ (_40233_, _40232_, _40230_);
  and _47462_ (_40234_, _39915_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _47463_ (_40235_, _40234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _47464_ (_40236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  not _47465_ (_40237_, _39919_);
  and _47466_ (_40238_, _40214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor _47467_ (_40239_, _40238_, _40237_);
  or _47468_ (_40240_, _40239_, _40236_);
  and _47469_ (_40241_, _40240_, _40235_);
  or _47470_ (_40242_, _40241_, _40233_);
  nor _47471_ (_40243_, _40242_, _39845_);
  nor _47472_ (_40244_, _40243_, _39841_);
  and _47473_ (_40245_, _40244_, _40229_);
  and _47474_ (_40246_, _39896_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _47475_ (_40247_, _40246_, _40245_);
  and _47476_ (_41622_, _40247_, _42882_);
  nand _47477_ (_40248_, _39845_, _38428_);
  and _47478_ (_40249_, _40230_, _39848_);
  nor _47479_ (_40250_, _40249_, _39919_);
  nor _47480_ (_40251_, _40250_, _40239_);
  nand _47481_ (_40252_, _40251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _47482_ (_40253_, _40251_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _47483_ (_40254_, _40253_, _40252_);
  or _47484_ (_40255_, _40254_, _39845_);
  and _47485_ (_40256_, _40255_, _40248_);
  or _47486_ (_40257_, _40256_, _39896_);
  or _47487_ (_40258_, _39897_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _47488_ (_40259_, _40258_, _42882_);
  and _47489_ (_41623_, _40259_, _40257_);
  nand _47490_ (_40260_, _39845_, _38420_);
  and _47491_ (_40261_, _40238_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _47492_ (_40262_, _40201_, _40261_);
  or _47493_ (_40263_, _40262_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand _47494_ (_40264_, _40262_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _47495_ (_40265_, _40264_, _40263_);
  nor _47496_ (_40266_, _40265_, _39845_);
  nor _47497_ (_40267_, _40266_, _39841_);
  and _47498_ (_40268_, _40267_, _40260_);
  and _47499_ (_40269_, _39896_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _47500_ (_40270_, _40269_, _40268_);
  and _47501_ (_41625_, _40270_, _42882_);
  nor _47502_ (_40271_, _39986_, _39955_);
  or _47503_ (_40272_, _40271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _47504_ (_40273_, _39977_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _47505_ (_40274_, _40005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47506_ (_40275_, _40274_, _40024_);
  nand _47507_ (_40276_, _40275_, _40273_);
  or _47508_ (_40277_, _40276_, _39955_);
  and _47509_ (_40278_, _40277_, _40272_);
  or _47510_ (_40279_, _40278_, _39994_);
  nand _47511_ (_40280_, _39994_, _38464_);
  and _47512_ (_40281_, _40280_, _42882_);
  and _47513_ (_41627_, _40281_, _40279_);
  nand _47514_ (_40282_, _39994_, _38456_);
  and _47515_ (_40283_, _39955_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _47516_ (_40284_, _40273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _47517_ (_40285_, _40273_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _47518_ (_40286_, _40285_, _40284_);
  and _47519_ (_40287_, _40005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _47520_ (_40288_, _40287_, _39983_);
  nor _47521_ (_40289_, _40288_, _40286_);
  nor _47522_ (_40290_, _40289_, _39955_);
  or _47523_ (_40291_, _40290_, _40283_);
  or _47524_ (_40292_, _40291_, _39994_);
  and _47525_ (_40293_, _40292_, _42882_);
  and _47526_ (_41629_, _40293_, _40282_);
  not _47527_ (_40294_, _39996_);
  nor _47528_ (_40295_, _40285_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _47529_ (_40296_, _40273_, _39978_);
  nor _47530_ (_40297_, _40296_, _40295_);
  and _47531_ (_40298_, _40005_, _39983_);
  and _47532_ (_40299_, _40298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor _47533_ (_40300_, _40299_, _40297_);
  nor _47534_ (_40301_, _40300_, _39955_);
  and _47535_ (_40302_, _39955_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _47536_ (_40303_, _40302_, _40301_);
  and _47537_ (_40304_, _40303_, _40294_);
  nor _47538_ (_40305_, _40020_, _38449_);
  or _47539_ (_40306_, _40305_, _40304_);
  and _47540_ (_41631_, _40306_, _42882_);
  and _47541_ (_40307_, _39980_, _39977_);
  nor _47542_ (_40308_, _40296_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor _47543_ (_40309_, _40308_, _40307_);
  and _47544_ (_40310_, _40298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor _47545_ (_40311_, _40310_, _40309_);
  nor _47546_ (_40312_, _40311_, _39955_);
  and _47547_ (_40313_, _39955_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _47548_ (_40314_, _40313_, _40312_);
  and _47549_ (_40315_, _40314_, _40294_);
  nor _47550_ (_40316_, _40020_, _38442_);
  or _47551_ (_40317_, _40316_, _40315_);
  and _47552_ (_41633_, _40317_, _42882_);
  nand _47553_ (_40318_, _39994_, _38434_);
  or _47554_ (_40319_, _39998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _47555_ (_40320_, _40307_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor _47556_ (_40321_, _40320_, _39982_);
  and _47557_ (_40322_, _40298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _47558_ (_40323_, _40322_, _40321_);
  or _47559_ (_40324_, _40323_, _39955_);
  and _47560_ (_40325_, _40324_, _40319_);
  or _47561_ (_40326_, _40325_, _39994_);
  and _47562_ (_40327_, _40326_, _42882_);
  and _47563_ (_41635_, _40327_, _40318_);
  nand _47564_ (_40328_, _39994_, _38428_);
  not _47565_ (_40329_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _47566_ (_40330_, _39982_, _39966_);
  and _47567_ (_40331_, _40330_, _40329_);
  and _47568_ (_40332_, _40298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _47569_ (_40333_, _40332_, _40331_);
  nor _47570_ (_40334_, _40333_, _39955_);
  and _47571_ (_40335_, _40330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not _47572_ (_40336_, _40335_);
  or _47573_ (_40337_, _40336_, _39955_);
  and _47574_ (_40338_, _40337_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _47575_ (_40339_, _40338_, _40334_);
  or _47576_ (_40340_, _40339_, _39994_);
  and _47577_ (_40341_, _40340_, _42882_);
  and _47578_ (_41637_, _40341_, _40328_);
  and _47579_ (_40342_, _40005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _47580_ (_40343_, _40342_, _39977_);
  and _47581_ (_40344_, _40343_, _40024_);
  nor _47582_ (_40345_, _40336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor _47583_ (_40346_, _40345_, _40344_);
  nor _47584_ (_40347_, _40346_, _39955_);
  and _47585_ (_40348_, _40337_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _47586_ (_40349_, _40348_, _40347_);
  and _47587_ (_40350_, _40349_, _40294_);
  nor _47588_ (_40351_, _40020_, _38420_);
  or _47589_ (_40352_, _40351_, _40350_);
  and _47590_ (_41638_, _40352_, _42882_);
  or _47591_ (_40353_, _40026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47592_ (_40354_, _40353_, _40022_);
  and _47593_ (_40355_, _40026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _47594_ (_40356_, _40355_, _40354_);
  and _47595_ (_40357_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _47596_ (_40358_, _40034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47597_ (_40359_, _40358_, _40033_);
  nor _47598_ (_40360_, _40359_, _40357_);
  and _47599_ (_40361_, _39982_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _47600_ (_40362_, _39982_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _47601_ (_40363_, _40362_, _39965_);
  nor _47602_ (_40364_, _40363_, _40361_);
  or _47603_ (_40365_, _40364_, _40360_);
  or _47604_ (_40366_, _40365_, _40356_);
  or _47605_ (_40367_, _40366_, _39955_);
  nand _47606_ (_40368_, _39955_, _38464_);
  and _47607_ (_40369_, _40368_, _40367_);
  and _47608_ (_40370_, _40369_, _40066_);
  and _47609_ (_40371_, _39994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _47610_ (_40372_, _40371_, _40370_);
  and _47611_ (_41640_, _40372_, _42882_);
  nand _47612_ (_40373_, _39955_, _38456_);
  or _47613_ (_40374_, _40355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _47614_ (_40375_, _40024_, _39977_);
  and _47615_ (_40376_, _40375_, _39958_);
  not _47616_ (_40377_, _40376_);
  or _47617_ (_40378_, _40377_, _40005_);
  and _47618_ (_40379_, _40378_, _40022_);
  and _47619_ (_40380_, _40379_, _40374_);
  and _47620_ (_40381_, _40034_, _39958_);
  or _47621_ (_40382_, _40357_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _47622_ (_40383_, _40382_, _40033_);
  nor _47623_ (_40384_, _40383_, _40381_);
  and _47624_ (_40385_, _40361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _47625_ (_40386_, _40361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand _47626_ (_40387_, _40386_, _39965_);
  nor _47627_ (_40388_, _40387_, _40385_);
  or _47628_ (_40389_, _40388_, _40384_);
  or _47629_ (_40390_, _40389_, _40380_);
  or _47630_ (_40391_, _40390_, _39955_);
  and _47631_ (_40392_, _40391_, _40020_);
  and _47632_ (_40393_, _40392_, _40373_);
  and _47633_ (_40394_, _39994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or _47634_ (_40395_, _40394_, _40393_);
  and _47635_ (_41642_, _40395_, _42882_);
  nor _47636_ (_40396_, _39998_, _38449_);
  or _47637_ (_40397_, _40376_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47638_ (_40398_, _40375_, _39959_);
  not _47639_ (_40399_, _40398_);
  and _47640_ (_40400_, _40399_, _40021_);
  and _47641_ (_40401_, _40400_, _40397_);
  and _47642_ (_40402_, _39977_, _39958_);
  and _47643_ (_40403_, _40402_, _39981_);
  or _47644_ (_40404_, _40403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47645_ (_40405_, _39982_, _39959_);
  nor _47646_ (_40406_, _40405_, _39966_);
  and _47647_ (_40407_, _40406_, _40404_);
  and _47648_ (_40408_, _40381_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _47649_ (_40409_, _40408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47650_ (_40410_, _40034_, _39959_);
  nand _47651_ (_40411_, _40410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47652_ (_40412_, _40411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47653_ (_40413_, _40412_, _40409_);
  or _47654_ (_40414_, _40413_, _40407_);
  nor _47655_ (_40415_, _40414_, _40401_);
  nor _47656_ (_40416_, _40415_, _39955_);
  or _47657_ (_40417_, _40416_, _39996_);
  or _47658_ (_40418_, _40417_, _40396_);
  or _47659_ (_40419_, _40294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47660_ (_40420_, _40419_, _42882_);
  and _47661_ (_41644_, _40420_, _40418_);
  nor _47662_ (_40421_, _39998_, _38442_);
  not _47663_ (_40422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47664_ (_40423_, _40398_, _40004_);
  nor _47665_ (_40424_, _40423_, _40422_);
  and _47666_ (_40425_, _40423_, _40422_);
  or _47667_ (_40426_, _40425_, _40424_);
  and _47668_ (_40427_, _40426_, _40022_);
  or _47669_ (_40428_, _40410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _47670_ (_40429_, _40035_);
  and _47671_ (_40430_, _40429_, _40033_);
  and _47672_ (_40431_, _40430_, _40428_);
  or _47673_ (_40432_, _40405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47674_ (_40433_, _39982_, _39960_);
  nor _47675_ (_40434_, _40433_, _39966_);
  and _47676_ (_40435_, _40434_, _40432_);
  or _47677_ (_40436_, _40435_, _40431_);
  nor _47678_ (_40437_, _40436_, _40427_);
  nor _47679_ (_40438_, _40437_, _39955_);
  or _47680_ (_40439_, _40438_, _39996_);
  or _47681_ (_40440_, _40439_, _40421_);
  nand _47682_ (_40441_, _39996_, _40422_);
  and _47683_ (_40442_, _40441_, _42882_);
  and _47684_ (_41646_, _40442_, _40440_);
  nand _47685_ (_40443_, _39955_, _38434_);
  or _47686_ (_40444_, _40433_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47687_ (_40445_, _40403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _47688_ (_40446_, _40445_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _47689_ (_40447_, _40446_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor _47690_ (_40448_, _40447_, _39966_);
  and _47691_ (_40449_, _40448_, _40444_);
  and _47692_ (_40450_, _40375_, _39960_);
  nand _47693_ (_40451_, _40450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _47694_ (_40452_, _40450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47695_ (_40453_, _40452_, _40021_);
  and _47696_ (_40454_, _40453_, _40451_);
  and _47697_ (_40455_, _40035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _47698_ (_40456_, _40455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _47699_ (_40457_, _40456_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47700_ (_40458_, _40035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _47701_ (_40459_, _40458_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47702_ (_40460_, _40459_, _40457_);
  or _47703_ (_40461_, _40460_, _40454_);
  or _47704_ (_40462_, _40461_, _40449_);
  or _47705_ (_40463_, _40462_, _39955_);
  and _47706_ (_40464_, _40463_, _40020_);
  and _47707_ (_40465_, _40464_, _40443_);
  and _47708_ (_40466_, _39994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _47709_ (_40467_, _40466_, _40465_);
  and _47710_ (_41648_, _40467_, _42882_);
  nor _47711_ (_40468_, _39998_, _38428_);
  not _47712_ (_40469_, _40447_);
  nor _47713_ (_40470_, _40469_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47714_ (_40471_, _40469_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _47715_ (_40472_, _40471_, _40470_);
  and _47716_ (_40473_, _40472_, _39965_);
  nor _47717_ (_40474_, _40451_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _47718_ (_40475_, _40474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand _47719_ (_40476_, _40474_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47720_ (_40477_, _40476_, _40022_);
  and _47721_ (_40478_, _40477_, _40475_);
  not _47722_ (_40479_, _40038_);
  and _47723_ (_40480_, _40479_, _40033_);
  or _47724_ (_40481_, _40458_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47725_ (_40482_, _40481_, _40480_);
  or _47726_ (_40483_, _40482_, _40478_);
  nor _47727_ (_40484_, _40483_, _40473_);
  nor _47728_ (_40485_, _40484_, _39955_);
  or _47729_ (_40486_, _40485_, _39996_);
  or _47730_ (_40487_, _40486_, _40468_);
  or _47731_ (_40488_, _40294_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _47732_ (_40489_, _40488_, _42882_);
  and _47733_ (_41650_, _40489_, _40487_);
  nand _47734_ (_40490_, _39955_, _38420_);
  or _47735_ (_40491_, _40027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _47736_ (_40492_, _40491_, _40022_);
  nor _47737_ (_40493_, _40492_, _40028_);
  or _47738_ (_40494_, _40038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _47739_ (_40495_, _40046_);
  and _47740_ (_40496_, _40495_, _40033_);
  and _47741_ (_40497_, _40496_, _40494_);
  or _47742_ (_40498_, _39988_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor _47743_ (_40499_, _40051_, _39966_);
  and _47744_ (_40500_, _40499_, _40498_);
  or _47745_ (_40501_, _40500_, _40497_);
  or _47746_ (_40502_, _40501_, _40493_);
  or _47747_ (_40503_, _40502_, _39955_);
  and _47748_ (_40504_, _40503_, _40020_);
  and _47749_ (_40505_, _40504_, _40490_);
  and _47750_ (_40506_, _39994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _47751_ (_40507_, _40506_, _40505_);
  and _47752_ (_41652_, _40507_, _42882_);
  nand _47753_ (_40508_, _40074_, _38464_);
  or _47754_ (_40509_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _47755_ (_40510_, _40509_, _42882_);
  and _47756_ (_41653_, _40510_, _40508_);
  or _47757_ (_40511_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _47758_ (_40512_, _40511_, _42882_);
  nand _47759_ (_40513_, _40074_, _38456_);
  and _47760_ (_41655_, _40513_, _40512_);
  or _47761_ (_40514_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _47762_ (_40515_, _40514_, _42882_);
  nand _47763_ (_40516_, _40074_, _38449_);
  and _47764_ (_41657_, _40516_, _40515_);
  or _47765_ (_40517_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _47766_ (_40518_, _40517_, _42882_);
  nand _47767_ (_40519_, _40074_, _38442_);
  and _47768_ (_41659_, _40519_, _40518_);
  or _47769_ (_40520_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _47770_ (_40521_, _40520_, _42882_);
  nand _47771_ (_40522_, _40074_, _38434_);
  and _47772_ (_41660_, _40522_, _40521_);
  or _47773_ (_40523_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _47774_ (_40524_, _40523_, _42882_);
  nand _47775_ (_40525_, _40074_, _38428_);
  and _47776_ (_41662_, _40525_, _40524_);
  or _47777_ (_40526_, _40074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _47778_ (_40527_, _40526_, _42882_);
  nand _47779_ (_40528_, _40074_, _38420_);
  and _47780_ (_41664_, _40528_, _40527_);
  nor _47781_ (_40529_, _27845_, _27703_);
  and _47782_ (_40530_, _40529_, _39031_);
  and _47783_ (_40531_, _40530_, _39236_);
  and _47784_ (_40532_, _40531_, _31304_);
  nand _47785_ (_40533_, _40532_, _31282_);
  and _47786_ (_40534_, _38401_, _31304_);
  and _47787_ (_40535_, _40534_, _39260_);
  not _47788_ (_40536_, _40535_);
  or _47789_ (_40537_, _40532_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _47790_ (_40538_, _40537_, _40536_);
  and _47791_ (_40539_, _40538_, _40533_);
  nor _47792_ (_40540_, _40536_, _38485_);
  or _47793_ (_40541_, _40540_, _40539_);
  and _47794_ (_42827_, _40541_, _42882_);
  and _47795_ (_40542_, _39839_, _27045_);
  and _47796_ (_40543_, _40542_, _39243_);
  not _47797_ (_40544_, _40543_);
  and _47798_ (_40545_, _27845_, _27714_);
  and _47799_ (_40546_, _40545_, _39031_);
  and _47800_ (_40547_, _40546_, _39236_);
  and _47801_ (_40548_, _40547_, _31304_);
  or _47802_ (_40549_, _40548_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _47803_ (_40550_, _40549_, _40544_);
  nand _47804_ (_40551_, _40548_, _31282_);
  and _47805_ (_40552_, _40551_, _40550_);
  nor _47806_ (_40553_, _40544_, _38485_);
  or _47807_ (_40554_, _40553_, _40552_);
  and _47808_ (_42830_, _40554_, _42882_);
  and _47809_ (_40555_, _40542_, _38405_);
  nor _47810_ (_40556_, _39030_, _27703_);
  and _47811_ (_40557_, _40556_, _27845_);
  and _47812_ (_40558_, _40557_, _27560_);
  and _47813_ (_40559_, _40558_, _39205_);
  nand _47814_ (_40560_, _40559_, _27023_);
  and _47815_ (_40561_, _40560_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _47816_ (_40562_, _40561_, _40555_);
  or _47817_ (_40563_, _27034_, _33285_);
  and _47818_ (_40564_, _40563_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _47819_ (_40565_, _40564_, _39007_);
  and _47820_ (_40566_, _40565_, _40559_);
  or _47821_ (_40567_, _40566_, _40562_);
  nand _47822_ (_40568_, _40555_, _38420_);
  and _47823_ (_40569_, _40568_, _42882_);
  and _47824_ (_42832_, _40569_, _40567_);
  not _47825_ (_40570_, _40555_);
  nor _47826_ (_40571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _47827_ (_40572_, _40571_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff );
  not _47828_ (_40573_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not _47829_ (_40574_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _47830_ (_40575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _47831_ (_40576_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _40575_);
  and _47832_ (_40577_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47833_ (_40578_, _40577_, _40576_);
  nor _47834_ (_40579_, _40578_, _40574_);
  or _47835_ (_40580_, _40579_, _40573_);
  and _47836_ (_40581_, _40575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and _47837_ (_40582_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _47838_ (_40583_, _40582_, _40581_);
  nor _47839_ (_40584_, _40583_, _40574_);
  and _47840_ (_40585_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _40575_);
  and _47841_ (_40586_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _47842_ (_40587_, _40586_, _40585_);
  nand _47843_ (_40588_, _40587_, _40584_);
  or _47844_ (_40590_, _40588_, _40580_);
  and _47845_ (_40592_, _40590_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _47846_ (_40594_, _40592_, _40572_);
  and _47847_ (_40596_, _38405_, _31304_);
  and _47848_ (_40598_, _40596_, _40556_);
  or _47849_ (_40600_, _40598_, _40594_);
  and _47850_ (_40602_, _40600_, _40570_);
  nand _47851_ (_40604_, _40598_, _31282_);
  and _47852_ (_40606_, _40604_, _40602_);
  nor _47853_ (_40608_, _40570_, _38485_);
  or _47854_ (_40610_, _40608_, _40606_);
  and _47855_ (_42834_, _40610_, _42882_);
  and _47856_ (_40613_, _39844_, _31348_);
  nand _47857_ (_40615_, _40613_, _31282_);
  not _47858_ (_40617_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  and _47859_ (_40619_, _40617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _47860_ (_40621_, _40587_, _40574_);
  not _47861_ (_40623_, _40621_);
  or _47862_ (_40625_, _40623_, _40584_);
  or _47863_ (_40627_, _40625_, _40580_);
  and _47864_ (_40629_, _40627_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _47865_ (_40631_, _40629_, _40619_);
  or _47866_ (_40633_, _40631_, _40613_);
  and _47867_ (_40635_, _40633_, _40570_);
  and _47868_ (_40637_, _40635_, _40615_);
  nor _47869_ (_40639_, _40570_, _38428_);
  or _47870_ (_40641_, _40639_, _40637_);
  and _47871_ (_42836_, _40641_, _42882_);
  not _47872_ (_40643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _47873_ (_40644_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , _40643_);
  nand _47874_ (_40645_, _40579_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  or _47875_ (_40646_, _40621_, _40584_);
  or _47876_ (_40647_, _40646_, _40645_);
  and _47877_ (_40648_, _40647_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _47878_ (_40649_, _40648_, _40644_);
  and _47879_ (_40650_, _40073_, _31348_);
  or _47880_ (_40651_, _40650_, _40649_);
  and _47881_ (_40652_, _40651_, _40570_);
  nand _47882_ (_40653_, _40650_, _31282_);
  and _47883_ (_40654_, _40653_, _40652_);
  nor _47884_ (_40655_, _40570_, _38456_);
  or _47885_ (_40656_, _40655_, _40654_);
  and _47886_ (_42838_, _40656_, _42882_);
  and _47887_ (_40657_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or _47888_ (_40658_, _40645_, _40625_);
  and _47889_ (_40659_, _40658_, _40657_);
  and _47890_ (_40660_, _40556_, _38623_);
  or _47891_ (_40661_, _40660_, _40659_);
  and _47892_ (_40662_, _40661_, _40570_);
  nand _47893_ (_40663_, _40660_, _31282_);
  and _47894_ (_40664_, _40663_, _40662_);
  nor _47895_ (_40665_, _40570_, _38442_);
  or _47896_ (_40666_, _40665_, _40664_);
  and _47897_ (_42840_, _40666_, _42882_);
  and _47898_ (_40667_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _47899_ (_40668_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _40575_);
  nor _47900_ (_40669_, _40668_, _40667_);
  and _47901_ (_40670_, _40669_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor _47902_ (_40671_, _40670_, _40574_);
  and _47903_ (_40672_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _47904_ (_40673_, _40672_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _47905_ (_40674_, _40673_);
  and _47906_ (_40675_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _47907_ (_40676_, _40675_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _47908_ (_40677_, _40676_);
  and _47909_ (_40678_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _47910_ (_40679_, _40678_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _47911_ (_40680_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _47912_ (_40681_, _40680_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _47913_ (_40682_, _40681_, _40679_);
  and _47914_ (_40683_, _40682_, _40677_);
  and _47915_ (_40684_, _40683_, _40674_);
  not _47916_ (_40685_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _47917_ (_40686_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor _47918_ (_40687_, _40686_, _40685_);
  nand _47919_ (_40688_, _40687_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not _47920_ (_40689_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _47921_ (_40690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _47922_ (_40691_, _40690_, _40689_);
  and _47923_ (_40692_, _40691_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _47924_ (_40693_, _40692_);
  and _47925_ (_40694_, _40693_, _40688_);
  and _47926_ (_40695_, _40694_, _40684_);
  nor _47927_ (_40696_, _40695_, _40671_);
  and _47928_ (_40697_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor _47929_ (_40698_, _40697_, _40575_);
  and _47930_ (_40699_, _40698_, _40696_);
  not _47931_ (_40700_, _40699_);
  not _47932_ (_40701_, _40698_);
  and _47933_ (_40702_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _40574_);
  not _47934_ (_40703_, _40702_);
  not _47935_ (_40704_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _47936_ (_40705_, _40675_, _40704_);
  not _47937_ (_40706_, _40705_);
  not _47938_ (_40707_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _47939_ (_40708_, _40678_, _40707_);
  not _47940_ (_40709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _47941_ (_40710_, _40680_, _40709_);
  nor _47942_ (_40711_, _40710_, _40708_);
  and _47943_ (_40712_, _40711_, _40706_);
  nor _47944_ (_40713_, _40712_, _40703_);
  not _47945_ (_40714_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _47946_ (_40715_, _40687_, _40714_);
  not _47947_ (_40716_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _47948_ (_40717_, _40691_, _40716_);
  nor _47949_ (_40718_, _40717_, _40715_);
  not _47950_ (_40719_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _47951_ (_40720_, _40672_, _40719_);
  not _47952_ (_40721_, _40720_);
  and _47953_ (_40722_, _40721_, _40718_);
  nor _47954_ (_40723_, _40722_, _40703_);
  nor _47955_ (_40724_, _40723_, _40713_);
  or _47956_ (_40725_, _40724_, _40701_);
  and _47957_ (_40726_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42882_);
  and _47958_ (_40727_, _40726_, _40725_);
  and _47959_ (_42870_, _40727_, _40700_);
  nor _47960_ (_40728_, _40697_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not _47961_ (_40729_, _40728_);
  not _47962_ (_40730_, _40696_);
  and _47963_ (_40731_, _40724_, _40730_);
  nor _47964_ (_40732_, _40731_, _40729_);
  nand _47965_ (_40733_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42882_);
  nor _47966_ (_42872_, _40733_, _40732_);
  and _47967_ (_40734_, _40694_, _40674_);
  nand _47968_ (_40735_, _40734_, _40696_);
  or _47969_ (_40736_, _40723_, _40696_);
  and _47970_ (_40737_, _40736_, _40698_);
  and _47971_ (_40738_, _40737_, _40735_);
  or _47972_ (_40739_, _40738_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or _47973_ (_40740_, _40700_, _40683_);
  nor _47974_ (_40741_, _40701_, _40696_);
  nand _47975_ (_40742_, _40741_, _40713_);
  and _47976_ (_40743_, _40742_, _42882_);
  and _47977_ (_40744_, _40743_, _40740_);
  and _47978_ (_42873_, _40744_, _40739_);
  and _47979_ (_40745_, _40735_, _40728_);
  or _47980_ (_40746_, _40745_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and _47981_ (_40747_, _40728_, _40696_);
  not _47982_ (_40748_, _40747_);
  or _47983_ (_40749_, _40748_, _40683_);
  or _47984_ (_40750_, _40723_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nand _47985_ (_40754_, _40728_, _40713_);
  and _47986_ (_40755_, _40754_, _40750_);
  or _47987_ (_40761_, _40755_, _40696_);
  and _47988_ (_40767_, _40761_, _42882_);
  and _47989_ (_40773_, _40767_, _40749_);
  and _47990_ (_42875_, _40773_, _40746_);
  nand _47991_ (_40779_, _40731_, _40574_);
  nor _47992_ (_40780_, _40575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nand _47993_ (_40781_, _40780_, _40697_);
  and _47994_ (_40782_, _40781_, _42882_);
  and _47995_ (_42877_, _40782_, _40779_);
  and _47996_ (_40783_, _40731_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _47997_ (_40784_, _40575_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _47998_ (_40785_, _40784_, _40780_);
  nor _47999_ (_40786_, _40785_, _40730_);
  or _48000_ (_40787_, _40786_, _40697_);
  or _48001_ (_40788_, _40787_, _40783_);
  not _48002_ (_40789_, _40697_);
  or _48003_ (_40790_, _40785_, _40789_);
  and _48004_ (_40791_, _40790_, _42882_);
  and _48005_ (_42879_, _40791_, _40788_);
  and _48006_ (_40796_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42882_);
  and _48007_ (_42880_, _40796_, _40697_);
  nor _48008_ (_42885_, _40571_, rst);
  and _48009_ (_42886_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _42882_);
  nor _48010_ (_40804_, _40731_, _40697_);
  and _48011_ (_40810_, _40697_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _48012_ (_40811_, _40810_, _40804_);
  and _48013_ (_00130_, _40811_, _42882_);
  and _48014_ (_40812_, _40697_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _48015_ (_40817_, _40812_, _40804_);
  and _48016_ (_00132_, _40817_, _42882_);
  and _48017_ (_40822_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _42882_);
  and _48018_ (_00134_, _40822_, _40697_);
  not _48019_ (_40826_, _40710_);
  nor _48020_ (_40832_, _40717_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _48021_ (_40833_, _40832_, _40715_);
  or _48022_ (_40834_, _40833_, _40720_);
  and _48023_ (_40839_, _40834_, _40826_);
  or _48024_ (_40840_, _40839_, _40708_);
  nor _48025_ (_40845_, _40724_, _40696_);
  and _48026_ (_40846_, _40845_, _40706_);
  and _48027_ (_40847_, _40846_, _40840_);
  not _48028_ (_40852_, _40681_);
  or _48029_ (_40857_, _40692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _48030_ (_40858_, _40857_, _40688_);
  or _48031_ (_40859_, _40858_, _40673_);
  and _48032_ (_40868_, _40859_, _40852_);
  or _48033_ (_40869_, _40868_, _40679_);
  and _48034_ (_40870_, _40696_, _40677_);
  and _48035_ (_40871_, _40870_, _40869_);
  or _48036_ (_40875_, _40871_, _40697_);
  or _48037_ (_40881_, _40875_, _40847_);
  or _48038_ (_40882_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _48039_ (_40883_, _40882_, _42882_);
  and _48040_ (_00136_, _40883_, _40881_);
  not _48041_ (_40888_, _40679_);
  or _48042_ (_40893_, _40681_, _40673_);
  and _48043_ (_40894_, _40694_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _48044_ (_40895_, _40894_, _40893_);
  and _48045_ (_40900_, _40895_, _40888_);
  and _48046_ (_40905_, _40900_, _40870_);
  nor _48047_ (_40906_, _40708_, _40705_);
  or _48048_ (_40907_, _40720_, _40710_);
  and _48049_ (_40911_, _40718_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _48050_ (_40917_, _40911_, _40907_);
  and _48051_ (_40918_, _40917_, _40906_);
  and _48052_ (_40922_, _40918_, _40845_);
  or _48053_ (_40923_, _40922_, _40697_);
  or _48054_ (_40929_, _40923_, _40905_);
  or _48055_ (_40930_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _48056_ (_40931_, _40930_, _42882_);
  and _48057_ (_00138_, _40931_, _40929_);
  and _48058_ (_40938_, _40721_, _40702_);
  nand _48059_ (_40941_, _40938_, _40712_);
  nor _48060_ (_40942_, _40941_, _40718_);
  nor _48061_ (_40944_, _40694_, _40671_);
  or _48062_ (_40950_, _40944_, _40942_);
  or _48063_ (_40953_, _40684_, _40671_);
  and _48064_ (_40954_, _40953_, _40950_);
  or _48065_ (_40955_, _40954_, _40697_);
  or _48066_ (_40961_, _40789_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _48067_ (_40965_, _40961_, _42882_);
  and _48068_ (_00140_, _40965_, _40955_);
  and _48069_ (_40966_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _42882_);
  and _48070_ (_00141_, _40966_, _40697_);
  and _48071_ (_40974_, _40697_, _40575_);
  or _48072_ (_40975_, _40974_, _40732_);
  or _48073_ (_40976_, _40975_, _40741_);
  and _48074_ (_00143_, _40976_, _42882_);
  not _48075_ (_40977_, _40804_);
  and _48076_ (_40978_, _40977_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _48077_ (_40979_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _48078_ (_40980_, _40692_, _40575_);
  or _48079_ (_40981_, _40980_, _40979_);
  nor _48080_ (_40982_, _40688_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _48081_ (_40983_, _40982_, _40673_);
  nand _48082_ (_40984_, _40983_, _40981_);
  or _48083_ (_40985_, _40674_, _40577_);
  and _48084_ (_40986_, _40985_, _40984_);
  or _48085_ (_40987_, _40986_, _40681_);
  or _48086_ (_40988_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _40575_);
  or _48087_ (_40989_, _40988_, _40852_);
  and _48088_ (_40990_, _40989_, _40888_);
  and _48089_ (_40991_, _40990_, _40987_);
  and _48090_ (_40992_, _40679_, _40577_);
  or _48091_ (_40993_, _40992_, _40676_);
  or _48092_ (_40994_, _40993_, _40991_);
  or _48093_ (_40995_, _40988_, _40677_);
  and _48094_ (_40996_, _40995_, _40696_);
  and _48095_ (_40997_, _40996_, _40994_);
  and _48096_ (_40998_, _40717_, _40575_);
  or _48097_ (_40999_, _40998_, _40979_);
  and _48098_ (_41000_, _40715_, _40575_);
  nor _48099_ (_41001_, _41000_, _40720_);
  nand _48100_ (_41002_, _41001_, _40999_);
  or _48101_ (_41003_, _40721_, _40577_);
  and _48102_ (_41004_, _41003_, _41002_);
  or _48103_ (_41005_, _41004_, _40710_);
  not _48104_ (_41006_, _40708_);
  or _48105_ (_41007_, _40988_, _40826_);
  and _48106_ (_41008_, _41007_, _41006_);
  and _48107_ (_41009_, _41008_, _41005_);
  and _48108_ (_41010_, _40708_, _40577_);
  or _48109_ (_41011_, _41010_, _40705_);
  or _48110_ (_41012_, _41011_, _41009_);
  and _48111_ (_41013_, _40988_, _40845_);
  or _48112_ (_41014_, _41013_, _40846_);
  and _48113_ (_41015_, _41014_, _41012_);
  or _48114_ (_41016_, _41015_, _40997_);
  and _48115_ (_41017_, _41016_, _40789_);
  or _48116_ (_41018_, _41017_, _40978_);
  and _48117_ (_00145_, _41018_, _42882_);
  and _48118_ (_41019_, _40977_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  or _48119_ (_41020_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _40575_);
  and _48120_ (_41021_, _41020_, _40677_);
  or _48121_ (_41022_, _41021_, _40683_);
  or _48122_ (_41023_, _40980_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _48123_ (_41024_, _41023_, _40983_);
  nand _48124_ (_41025_, _40673_, _40586_);
  nand _48125_ (_41026_, _41025_, _40682_);
  or _48126_ (_41027_, _41026_, _41024_);
  and _48127_ (_41028_, _41027_, _41022_);
  and _48128_ (_41029_, _40676_, _40586_);
  or _48129_ (_41030_, _41029_, _41028_);
  and _48130_ (_41031_, _41030_, _40696_);
  and _48131_ (_41032_, _40705_, _40586_);
  and _48132_ (_41033_, _41020_, _40706_);
  or _48133_ (_41034_, _41033_, _40712_);
  and _48134_ (_41035_, _40720_, _40586_);
  not _48135_ (_41036_, _40711_);
  or _48136_ (_41037_, _40998_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _48137_ (_41038_, _41037_, _41001_);
  or _48138_ (_41039_, _41038_, _41036_);
  or _48139_ (_41040_, _41039_, _41035_);
  and _48140_ (_41041_, _41040_, _41034_);
  or _48141_ (_41042_, _41041_, _41032_);
  and _48142_ (_41043_, _41042_, _40845_);
  or _48143_ (_41044_, _41043_, _41031_);
  and _48144_ (_41045_, _41044_, _40789_);
  or _48145_ (_41046_, _41045_, _41019_);
  and _48146_ (_00147_, _41046_, _42882_);
  and _48147_ (_41047_, _40977_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _48148_ (_41048_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _48149_ (_41049_, _41048_, _40677_);
  and _48150_ (_41050_, _41049_, _40696_);
  not _48151_ (_41051_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _48152_ (_41052_, _40692_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _48153_ (_41053_, _41052_, _41051_);
  nor _48154_ (_41054_, _40688_, _40575_);
  nor _48155_ (_41055_, _41054_, _40673_);
  nand _48156_ (_41056_, _41055_, _41053_);
  or _48157_ (_41057_, _40674_, _40576_);
  and _48158_ (_41058_, _41057_, _41056_);
  or _48159_ (_41059_, _41058_, _40681_);
  or _48160_ (_41060_, _41048_, _40852_);
  and _48161_ (_41061_, _41060_, _40888_);
  and _48162_ (_41062_, _41061_, _41059_);
  and _48163_ (_41063_, _40679_, _40576_);
  or _48164_ (_41064_, _41063_, _40676_);
  or _48165_ (_41065_, _41064_, _41062_);
  and _48166_ (_41066_, _41065_, _41050_);
  or _48167_ (_41067_, _41048_, _40706_);
  and _48168_ (_41068_, _40717_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _48169_ (_41069_, _41068_, _41051_);
  and _48170_ (_41070_, _40715_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _48171_ (_41071_, _41070_, _40720_);
  nand _48172_ (_41072_, _41071_, _41069_);
  or _48173_ (_41073_, _40721_, _40576_);
  and _48174_ (_41074_, _41073_, _41072_);
  or _48175_ (_41075_, _41074_, _40710_);
  or _48176_ (_41076_, _41048_, _40826_);
  and _48177_ (_41077_, _41076_, _41006_);
  and _48178_ (_41078_, _41077_, _41075_);
  and _48179_ (_41079_, _40708_, _40576_);
  or _48180_ (_41080_, _41079_, _40705_);
  or _48181_ (_41081_, _41080_, _41078_);
  and _48182_ (_41082_, _41081_, _40845_);
  and _48183_ (_41083_, _41082_, _41067_);
  or _48184_ (_41084_, _41083_, _41066_);
  and _48185_ (_41085_, _41084_, _40789_);
  or _48186_ (_41086_, _41085_, _41047_);
  and _48187_ (_00149_, _41086_, _42882_);
  and _48188_ (_41087_, _40977_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  or _48189_ (_41088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _48190_ (_41089_, _41088_, _40677_);
  or _48191_ (_41090_, _41089_, _40683_);
  or _48192_ (_41091_, _41052_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _48193_ (_41093_, _41091_, _41055_);
  nand _48194_ (_41094_, _40673_, _40585_);
  nand _48195_ (_41096_, _41094_, _40682_);
  or _48196_ (_41097_, _41096_, _41093_);
  and _48197_ (_41099_, _41097_, _41090_);
  and _48198_ (_41100_, _40676_, _40585_);
  or _48199_ (_41102_, _41100_, _41099_);
  and _48200_ (_41103_, _41102_, _40696_);
  and _48201_ (_41105_, _40705_, _40585_);
  and _48202_ (_41106_, _41088_, _40706_);
  or _48203_ (_41108_, _41106_, _40712_);
  and _48204_ (_41109_, _40720_, _40585_);
  or _48205_ (_41111_, _41068_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _48206_ (_41112_, _41111_, _41071_);
  or _48207_ (_41114_, _41112_, _41036_);
  or _48208_ (_41115_, _41114_, _41109_);
  and _48209_ (_41117_, _41115_, _41108_);
  or _48210_ (_41118_, _41117_, _41105_);
  and _48211_ (_41120_, _41118_, _40845_);
  or _48212_ (_41121_, _41120_, _41103_);
  and _48213_ (_41122_, _41121_, _40789_);
  or _48214_ (_41123_, _41122_, _41087_);
  and _48215_ (_00151_, _41123_, _42882_);
  or _48216_ (_41124_, _40729_, _40724_);
  and _48217_ (_41125_, _41124_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  or _48218_ (_41126_, _41125_, _40747_);
  and _48219_ (_00152_, _41126_, _42882_);
  and _48220_ (_41127_, _40725_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  or _48221_ (_41128_, _41127_, _40699_);
  and _48222_ (_00154_, _41128_, _42882_);
  and _48223_ (_41129_, _40559_, _27045_);
  or _48224_ (_41130_, _41129_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _48225_ (_41131_, _41130_, _40570_);
  nand _48226_ (_41132_, _41129_, _31282_);
  and _48227_ (_41133_, _41132_, _41131_);
  and _48228_ (_41134_, _40555_, _38465_);
  or _48229_ (_41135_, _41134_, _41133_);
  and _48230_ (_00156_, _41135_, _42882_);
  and _48231_ (_41136_, _40559_, _33296_);
  or _48232_ (_41137_, _41136_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _48233_ (_41138_, _41137_, _40570_);
  nand _48234_ (_41139_, _41136_, _31282_);
  and _48235_ (_41140_, _41139_, _41138_);
  nor _48236_ (_41141_, _40570_, _38449_);
  or _48237_ (_41142_, _41141_, _41140_);
  and _48238_ (_00158_, _41142_, _42882_);
  and _48239_ (_41143_, _40559_, _34765_);
  or _48240_ (_41144_, _41143_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _48241_ (_41145_, _41144_, _40570_);
  nand _48242_ (_41146_, _41143_, _31282_);
  and _48243_ (_41147_, _41146_, _41145_);
  nor _48244_ (_41148_, _40570_, _38434_);
  or _48245_ (_41149_, _41148_, _41147_);
  and _48246_ (_00160_, _41149_, _42882_);
  and _48247_ (_41150_, _40547_, _27045_);
  or _48248_ (_41151_, _41150_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _48249_ (_41152_, _41151_, _40544_);
  nand _48250_ (_41153_, _41150_, _31282_);
  and _48251_ (_41154_, _41153_, _41152_);
  and _48252_ (_41155_, _40543_, _38465_);
  or _48253_ (_41156_, _41155_, _41154_);
  and _48254_ (_00162_, _41156_, _42882_);
  and _48255_ (_41157_, _40547_, _32567_);
  or _48256_ (_41158_, _41157_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _48257_ (_41159_, _41158_, _40544_);
  nand _48258_ (_41160_, _41157_, _31282_);
  and _48259_ (_41161_, _41160_, _41159_);
  nor _48260_ (_41162_, _40544_, _38456_);
  or _48261_ (_41163_, _41162_, _41161_);
  and _48262_ (_00163_, _41163_, _42882_);
  nand _48263_ (_41164_, _40547_, _39293_);
  and _48264_ (_41165_, _41164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _48265_ (_41166_, _41165_, _40543_);
  and _48266_ (_41167_, _33329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _48267_ (_41168_, _41167_, _33318_);
  and _48268_ (_41169_, _41168_, _40547_);
  or _48269_ (_41170_, _41169_, _41166_);
  nand _48270_ (_41171_, _40543_, _38449_);
  and _48271_ (_41172_, _41171_, _42882_);
  and _48272_ (_00165_, _41172_, _41170_);
  and _48273_ (_41173_, _40547_, _34004_);
  or _48274_ (_41174_, _41173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _48275_ (_41175_, _41174_, _40544_);
  nand _48276_ (_41176_, _41173_, _31282_);
  and _48277_ (_41177_, _41176_, _41175_);
  nor _48278_ (_41178_, _40544_, _38442_);
  or _48279_ (_41179_, _41178_, _41177_);
  and _48280_ (_00167_, _41179_, _42882_);
  and _48281_ (_41180_, _40547_, _34765_);
  or _48282_ (_41181_, _41180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _48283_ (_41182_, _41181_, _40544_);
  nand _48284_ (_41183_, _41180_, _31282_);
  and _48285_ (_41184_, _41183_, _41182_);
  nor _48286_ (_41185_, _40544_, _38434_);
  or _48287_ (_41186_, _41185_, _41184_);
  and _48288_ (_00169_, _41186_, _42882_);
  and _48289_ (_41187_, _40547_, _35549_);
  or _48290_ (_41188_, _41187_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _48291_ (_41189_, _41188_, _40544_);
  nand _48292_ (_41190_, _41187_, _31282_);
  and _48293_ (_41191_, _41190_, _41189_);
  nor _48294_ (_41192_, _40544_, _38428_);
  or _48295_ (_41193_, _41192_, _41191_);
  and _48296_ (_00171_, _41193_, _42882_);
  and _48297_ (_41194_, _40547_, _36277_);
  or _48298_ (_41195_, _41194_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _48299_ (_41196_, _41195_, _40544_);
  nand _48300_ (_41197_, _41194_, _31282_);
  and _48301_ (_41198_, _41197_, _41196_);
  nor _48302_ (_41199_, _40544_, _38420_);
  or _48303_ (_41200_, _41199_, _41198_);
  and _48304_ (_00173_, _41200_, _42882_);
  and _48305_ (_41201_, _40531_, _27045_);
  nand _48306_ (_41202_, _41201_, _31282_);
  or _48307_ (_41203_, _41201_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _48308_ (_41204_, _41203_, _40536_);
  and _48309_ (_41205_, _41204_, _41202_);
  and _48310_ (_41206_, _40535_, _38465_);
  or _48311_ (_41207_, _41206_, _41205_);
  and _48312_ (_00174_, _41207_, _42882_);
  and _48313_ (_41208_, _40531_, _32567_);
  nand _48314_ (_41209_, _41208_, _31282_);
  or _48315_ (_41210_, _41208_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _48316_ (_41211_, _41210_, _40536_);
  and _48317_ (_41212_, _41211_, _41209_);
  nor _48318_ (_41213_, _40536_, _38456_);
  or _48319_ (_41214_, _41213_, _41212_);
  and _48320_ (_00176_, _41214_, _42882_);
  and _48321_ (_41215_, _33329_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _48322_ (_41216_, _41215_, _33318_);
  and _48323_ (_41217_, _41216_, _40531_);
  nand _48324_ (_41218_, _40531_, _39293_);
  and _48325_ (_41219_, _41218_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _48326_ (_41220_, _41219_, _40535_);
  or _48327_ (_41221_, _41220_, _41217_);
  nand _48328_ (_41222_, _40535_, _38449_);
  and _48329_ (_41223_, _41222_, _42882_);
  and _48330_ (_00178_, _41223_, _41221_);
  and _48331_ (_41224_, _40531_, _34004_);
  nand _48332_ (_41225_, _41224_, _31282_);
  or _48333_ (_41226_, _41224_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _48334_ (_41227_, _41226_, _41225_);
  or _48335_ (_41228_, _41227_, _40535_);
  nand _48336_ (_41229_, _40535_, _38442_);
  and _48337_ (_41230_, _41229_, _42882_);
  and _48338_ (_00180_, _41230_, _41228_);
  and _48339_ (_41231_, _40531_, _34765_);
  nand _48340_ (_41232_, _41231_, _31282_);
  or _48341_ (_41233_, _41231_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _48342_ (_41234_, _41233_, _40536_);
  and _48343_ (_41235_, _41234_, _41232_);
  nor _48344_ (_41236_, _40536_, _38434_);
  or _48345_ (_41237_, _41236_, _41235_);
  and _48346_ (_00182_, _41237_, _42882_);
  and _48347_ (_41238_, _40531_, _35549_);
  nand _48348_ (_41239_, _41238_, _31282_);
  or _48349_ (_41240_, _41238_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _48350_ (_41241_, _41240_, _41239_);
  or _48351_ (_41242_, _41241_, _40535_);
  nand _48352_ (_41243_, _40535_, _38428_);
  and _48353_ (_41244_, _41243_, _42882_);
  and _48354_ (_00184_, _41244_, _41242_);
  and _48355_ (_41245_, _40531_, _36277_);
  nand _48356_ (_41246_, _41245_, _31282_);
  or _48357_ (_41247_, _41245_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _48358_ (_41248_, _41247_, _41246_);
  or _48359_ (_41249_, _41248_, _40535_);
  nand _48360_ (_41250_, _40535_, _38420_);
  and _48361_ (_41251_, _41250_, _42882_);
  and _48362_ (_00185_, _41251_, _41249_);
  and _48363_ (_41252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _48364_ (_41253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor _48365_ (_41254_, _40571_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  and _48366_ (_41255_, _41254_, _41253_);
  not _48367_ (_41256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _48368_ (_41257_, _41256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _48369_ (_41258_, _41257_, _41255_);
  nor _48370_ (_41259_, _41258_, _41252_);
  or _48371_ (_41260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _48372_ (_41261_, _41260_, _42882_);
  nor _48373_ (_00546_, _41261_, _41259_);
  nor _48374_ (_41262_, _41259_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _48375_ (_41263_, _41262_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _48376_ (_41264_, _41262_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _48377_ (_41265_, _41264_, _42882_);
  and _48378_ (_00548_, _41265_, _41263_);
  not _48379_ (_41266_, rxd_i);
  and _48380_ (_41267_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _41266_);
  nor _48381_ (_41268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _48382_ (_41269_, _41268_);
  and _48383_ (_41270_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  and _48384_ (_41271_, _41270_, _41269_);
  and _48385_ (_41272_, _41271_, _41267_);
  not _48386_ (_41273_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _48387_ (_41274_, _41273_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _48388_ (_41275_, _41274_, _41268_);
  or _48389_ (_41276_, _41275_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  or _48390_ (_41277_, _41276_, _41272_);
  and _48391_ (_41278_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _42882_);
  and _48392_ (_00551_, _41278_, _41277_);
  and _48393_ (_41279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _48394_ (_41280_, _41279_, _41269_);
  nor _48395_ (_41281_, _41268_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _48396_ (_41282_, _41281_, _41273_);
  nor _48397_ (_41283_, _41282_, _41280_);
  not _48398_ (_41284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _48399_ (_41285_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _41284_);
  not _48400_ (_41286_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _48401_ (_41287_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _41286_);
  and _48402_ (_41288_, _41287_, _41285_);
  not _48403_ (_41289_, _41288_);
  or _48404_ (_41290_, _41289_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  and _48405_ (_41291_, _41288_, _41280_);
  and _48406_ (_41292_, _41280_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48407_ (_41293_, _41292_, _41291_);
  and _48408_ (_41294_, _41293_, _41290_);
  or _48409_ (_41295_, _41294_, _41283_);
  not _48410_ (_41296_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nand _48411_ (_41297_, _41268_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor _48412_ (_41298_, _41297_, _41296_);
  not _48413_ (_41299_, _41298_);
  or _48414_ (_41300_, _41299_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand _48415_ (_41301_, _41300_, _41295_);
  nand _48416_ (_00554_, _41301_, _41278_);
  not _48417_ (_41302_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  not _48418_ (_41303_, _41280_);
  nor _48419_ (_41304_, _41273_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not _48420_ (_41305_, _41304_);
  not _48421_ (_41306_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _48422_ (_41307_, _41268_, _41306_);
  and _48423_ (_41308_, _41307_, _41305_);
  and _48424_ (_41309_, _41308_, _41303_);
  nor _48425_ (_41310_, _41309_, _41302_);
  and _48426_ (_41311_, _41309_, rxd_i);
  or _48427_ (_41312_, _41311_, rst);
  or _48428_ (_00556_, _41312_, _41310_);
  nor _48429_ (_41313_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _48430_ (_41314_, _41313_, _41285_);
  and _48431_ (_41315_, _41314_, _41292_);
  nand _48432_ (_41316_, _41315_, _41266_);
  or _48433_ (_41317_, _41315_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _48434_ (_41318_, _41317_, _42882_);
  and _48435_ (_00559_, _41318_, _41316_);
  and _48436_ (_41319_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _48437_ (_41320_, _41319_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _48438_ (_41321_, _41320_, _41284_);
  and _48439_ (_41322_, _41321_, _41292_);
  and _48440_ (_41323_, _41271_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _48441_ (_41324_, _41323_, _41292_);
  nor _48442_ (_41325_, _41320_, _41303_);
  or _48443_ (_41326_, _41325_, _41324_);
  and _48444_ (_41327_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _48445_ (_41328_, _41327_, _41322_);
  and _48446_ (_00562_, _41328_, _42882_);
  and _48447_ (_41329_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _42882_);
  nand _48448_ (_41330_, _41329_, _41306_);
  nand _48449_ (_41331_, _41278_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  nand _48450_ (_00564_, _41331_, _41330_);
  and _48451_ (_41332_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41306_);
  not _48452_ (_41333_, _41271_);
  nand _48453_ (_41334_, _41275_, _41296_);
  and _48454_ (_41335_, _41334_, _41333_);
  nand _48455_ (_41336_, _41335_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nand _48456_ (_41337_, _41336_, _41303_);
  or _48457_ (_41338_, _41288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor _48458_ (_41339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _48459_ (_41340_, _41339_, _41291_);
  and _48460_ (_41341_, _41340_, _41338_);
  and _48461_ (_41342_, _41341_, _41337_);
  or _48462_ (_41343_, _41342_, _41298_);
  nand _48463_ (_41344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nand _48464_ (_41345_, _41344_, _41280_);
  or _48465_ (_41346_, _41345_, _41289_);
  and _48466_ (_41347_, _41346_, _41299_);
  or _48467_ (_41348_, _41347_, rxd_i);
  and _48468_ (_41349_, _41348_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _48469_ (_41350_, _41349_, _41343_);
  or _48470_ (_41351_, _41350_, _41332_);
  and _48471_ (_00567_, _41351_, _42882_);
  and _48472_ (_41352_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _48473_ (_41353_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _48474_ (_41354_, _41254_, _41353_);
  or _48475_ (_41355_, _41354_, _41257_);
  nor _48476_ (_41356_, _41355_, _41352_);
  or _48477_ (_41357_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _48478_ (_41358_, _41357_, _42882_);
  nor _48479_ (_00570_, _41358_, _41356_);
  nor _48480_ (_41359_, _41356_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _48481_ (_41360_, _41359_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _48482_ (_41361_, _41359_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _48483_ (_41362_, _41361_, _42882_);
  and _48484_ (_00572_, _41362_, _41360_);
  not _48485_ (_41363_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _48486_ (_41364_, _41297_, _41363_);
  nor _48487_ (_41365_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not _48488_ (_41366_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _48489_ (_41367_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _48490_ (_41368_, _41367_, _41366_);
  and _48491_ (_41369_, _41368_, _41365_);
  not _48492_ (_41370_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _48493_ (_41371_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor _48494_ (_41372_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _48495_ (_41373_, _41372_, _41371_);
  and _48496_ (_41374_, _41373_, _41370_);
  and _48497_ (_41375_, _41374_, _41369_);
  or _48498_ (_41376_, _41375_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor _48499_ (_41377_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _48500_ (_41378_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _48501_ (_41379_, _41378_, _41377_);
  and _48502_ (_41380_, _41269_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _48503_ (_41381_, _41380_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _48504_ (_41382_, _41381_, _41379_);
  not _48505_ (_41383_, _41382_);
  or _48506_ (_41384_, _41383_, _41376_);
  and _48507_ (_41385_, _41379_, _41380_);
  or _48508_ (_41386_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _41363_);
  or _48509_ (_41387_, _41386_, _41385_);
  and _48510_ (_41388_, _41387_, _41384_);
  or _48511_ (_41389_, _41388_, _41364_);
  not _48512_ (_41390_, _41364_);
  not _48513_ (_41391_, _41375_);
  or _48514_ (_41392_, _41391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and _48515_ (_41393_, _41392_, _41376_);
  or _48516_ (_41394_, _41393_, _41390_);
  nand _48517_ (_41395_, _41394_, _41389_);
  and _48518_ (_41396_, _40063_, _32556_);
  and _48519_ (_41397_, _41396_, _30679_);
  and _48520_ (_41398_, _41397_, _39227_);
  nor _48521_ (_41399_, _41398_, rst);
  nand _48522_ (_41400_, _41399_, _41395_);
  not _48523_ (_41401_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  and _48524_ (_41402_, _41398_, _42882_);
  nand _48525_ (_41403_, _41402_, _41401_);
  and _48526_ (_00575_, _41403_, _41400_);
  nor _48527_ (_41404_, _41391_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand _48528_ (_41405_, _41385_, _41404_);
  and _48529_ (_41406_, _41375_, _41364_);
  or _48530_ (_41407_, _41363_, rst);
  nor _48531_ (_41408_, _41407_, _41406_);
  and _48532_ (_41409_, _41408_, _41405_);
  or _48533_ (_00578_, _41409_, _41402_);
  or _48534_ (_41410_, _41383_, _41404_);
  or _48535_ (_41411_, _41385_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _48536_ (_41412_, _41297_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _48537_ (_41413_, _41412_, _41411_);
  and _48538_ (_41414_, _41413_, _41410_);
  or _48539_ (_41415_, _41414_, _41406_);
  and _48540_ (_00580_, _41415_, _41399_);
  and _48541_ (_41416_, _41381_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _48542_ (_41417_, _41416_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _48543_ (_41418_, _41417_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or _48544_ (_41419_, _41418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand _48545_ (_41420_, _41418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _48546_ (_41421_, _41420_, _41419_);
  and _48547_ (_00583_, _41421_, _41399_);
  nor _48548_ (_41422_, _41382_, _41364_);
  and _48549_ (_41423_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _48550_ (_41424_, _41423_, _41399_);
  and _48551_ (_41425_, _41402_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _48552_ (_00586_, _41425_, _41424_);
  and _48553_ (_41426_, _40534_, _38405_);
  or _48554_ (_41427_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _48555_ (_41428_, _41427_, _42882_);
  nand _48556_ (_41429_, _41426_, _38485_);
  and _48557_ (_00588_, _41429_, _41428_);
  and _48558_ (_41430_, _40530_, _39205_);
  and _48559_ (_41431_, _41430_, _31304_);
  nand _48560_ (_41432_, _41431_, _31282_);
  and _48561_ (_41433_, _40542_, _39227_);
  not _48562_ (_41434_, _41433_);
  or _48563_ (_41435_, _41431_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _48564_ (_41436_, _41435_, _41434_);
  and _48565_ (_41437_, _41436_, _41432_);
  nor _48566_ (_41438_, _41434_, _38485_);
  or _48567_ (_41439_, _41438_, _41437_);
  and _48568_ (_00591_, _41439_, _42882_);
  nor _48569_ (_41440_, _41298_, _41291_);
  not _48570_ (_41441_, _41440_);
  nor _48571_ (_41442_, _41335_, _41280_);
  nor _48572_ (_41443_, _41442_, _41441_);
  nor _48573_ (_41444_, _41443_, _41306_);
  or _48574_ (_41445_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _48575_ (_41446_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _41306_);
  or _48576_ (_41447_, _41446_, _41440_);
  and _48577_ (_41448_, _41447_, _42882_);
  and _48578_ (_01210_, _41448_, _41445_);
  or _48579_ (_41449_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _48580_ (_41450_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _41306_);
  or _48581_ (_41451_, _41450_, _41440_);
  and _48582_ (_41452_, _41451_, _42882_);
  and _48583_ (_01212_, _41452_, _41449_);
  or _48584_ (_41453_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _48585_ (_41454_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41306_);
  or _48586_ (_41455_, _41454_, _41440_);
  and _48587_ (_41456_, _41455_, _42882_);
  and _48588_ (_01214_, _41456_, _41453_);
  or _48589_ (_41457_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _48590_ (_41458_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41306_);
  or _48591_ (_41459_, _41458_, _41440_);
  and _48592_ (_41460_, _41459_, _42882_);
  and _48593_ (_01216_, _41460_, _41457_);
  or _48594_ (_41461_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _48595_ (_41462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41306_);
  or _48596_ (_41463_, _41462_, _41440_);
  and _48597_ (_41464_, _41463_, _42882_);
  and _48598_ (_01218_, _41464_, _41461_);
  or _48599_ (_41465_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _48600_ (_41466_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41306_);
  or _48601_ (_41467_, _41466_, _41440_);
  and _48602_ (_41468_, _41467_, _42882_);
  and _48603_ (_01220_, _41468_, _41465_);
  or _48604_ (_41469_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _48605_ (_41470_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41306_);
  or _48606_ (_41471_, _41470_, _41440_);
  and _48607_ (_41472_, _41471_, _42882_);
  and _48608_ (_01222_, _41472_, _41469_);
  or _48609_ (_41473_, _41444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _48610_ (_41474_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _41306_);
  or _48611_ (_41475_, _41474_, _41440_);
  and _48612_ (_41476_, _41475_, _42882_);
  and _48613_ (_01224_, _41476_, _41473_);
  nor _48614_ (_41477_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and _48615_ (_41478_, _41477_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _48616_ (_41479_, _41289_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or _48617_ (_41480_, _41288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _48618_ (_41481_, _41480_, _41280_);
  and _48619_ (_41482_, _41481_, _41479_);
  or _48620_ (_41483_, _41271_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _48621_ (_41484_, _41483_, _41334_);
  and _48622_ (_41485_, _41484_, _41303_);
  or _48623_ (_41486_, _41485_, _41482_);
  or _48624_ (_41487_, _41486_, _41298_);
  or _48625_ (_41488_, _41299_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _48626_ (_41489_, _41488_, _41278_);
  and _48627_ (_41490_, _41489_, _41487_);
  or _48628_ (_01226_, _41490_, _41478_);
  and _48629_ (_41491_, _41288_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _48630_ (_41492_, _41491_, _41335_);
  or _48631_ (_41493_, _41492_, _41443_);
  and _48632_ (_41494_, _41493_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _48633_ (_41495_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _41306_);
  nand _48634_ (_41496_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _48635_ (_41497_, _41496_, _41440_);
  or _48636_ (_41498_, _41497_, _41495_);
  or _48637_ (_41499_, _41498_, _41494_);
  and _48638_ (_01228_, _41499_, _42882_);
  not _48639_ (_41500_, _41444_);
  and _48640_ (_41501_, _41500_, _41329_);
  or _48641_ (_41502_, _41492_, _41441_);
  and _48642_ (_41503_, _41278_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _48643_ (_41504_, _41503_, _41502_);
  or _48644_ (_01229_, _41504_, _41501_);
  or _48645_ (_41505_, _41322_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand _48646_ (_41506_, _41322_, _41266_);
  and _48647_ (_41507_, _41506_, _42882_);
  and _48648_ (_01231_, _41507_, _41505_);
  or _48649_ (_41508_, _41324_, _41286_);
  or _48650_ (_41509_, _41292_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _48651_ (_41510_, _41509_, _42882_);
  and _48652_ (_01233_, _41510_, _41508_);
  and _48653_ (_41511_, _41324_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _48654_ (_41512_, _41313_, _41319_);
  and _48655_ (_41513_, _41512_, _41292_);
  or _48656_ (_41514_, _41513_, _41511_);
  and _48657_ (_01235_, _41514_, _42882_);
  and _48658_ (_41515_, _41326_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _48659_ (_41516_, _41319_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _48660_ (_41517_, _41516_, _41325_);
  or _48661_ (_41518_, _41517_, _41515_);
  and _48662_ (_01237_, _41518_, _42882_);
  and _48663_ (_41519_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _41306_);
  and _48664_ (_41520_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48665_ (_41521_, _41520_, _41519_);
  and _48666_ (_01239_, _41521_, _42882_);
  and _48667_ (_41522_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _41306_);
  and _48668_ (_41523_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48669_ (_41524_, _41523_, _41522_);
  and _48670_ (_01241_, _41524_, _42882_);
  and _48671_ (_41525_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _41306_);
  and _48672_ (_41526_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48673_ (_41527_, _41526_, _41525_);
  and _48674_ (_01243_, _41527_, _42882_);
  and _48675_ (_41528_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _41306_);
  and _48676_ (_41529_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48677_ (_41530_, _41529_, _41528_);
  and _48678_ (_01245_, _41530_, _42882_);
  and _48679_ (_41531_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _41306_);
  and _48680_ (_41532_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48681_ (_41533_, _41532_, _41531_);
  and _48682_ (_01247_, _41533_, _42882_);
  and _48683_ (_41534_, _41278_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _48684_ (_01249_, _41534_, _41478_);
  and _48685_ (_41535_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _48686_ (_41536_, _41535_, _41495_);
  and _48687_ (_01251_, _41536_, _42882_);
  nor _48688_ (_41537_, _41381_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _48689_ (_41538_, _41537_, _41416_);
  and _48690_ (_01253_, _41538_, _41399_);
  nor _48691_ (_41539_, _41416_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _48692_ (_41540_, _41539_, _41417_);
  and _48693_ (_01255_, _41540_, _41399_);
  nor _48694_ (_41541_, _41417_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _48695_ (_41542_, _41541_, _41418_);
  and _48696_ (_01257_, _41542_, _41399_);
  or _48697_ (_41543_, _41382_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _48698_ (_41544_, _41383_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _48699_ (_41545_, _41544_, _41543_);
  and _48700_ (_41546_, _41545_, _41390_);
  and _48701_ (_41547_, _41375_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _48702_ (_41548_, _41547_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _48703_ (_41549_, _41548_, _41364_);
  or _48704_ (_41550_, _41549_, _41546_);
  and _48705_ (_41551_, _41550_, _41399_);
  nor _48706_ (_41552_, _41269_, _38464_);
  and _48707_ (_41553_, _41552_, _41402_);
  or _48708_ (_01259_, _41553_, _41551_);
  not _48709_ (_41554_, _41422_);
  and _48710_ (_41555_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _48711_ (_41556_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _48712_ (_41557_, _41556_, _41555_);
  and _48713_ (_41558_, _41557_, _41399_);
  nand _48714_ (_41559_, _41268_, _38456_);
  nand _48715_ (_41560_, _41269_, _38464_);
  and _48716_ (_41561_, _41560_, _41402_);
  and _48717_ (_41562_, _41561_, _41559_);
  or _48718_ (_01261_, _41562_, _41558_);
  nor _48719_ (_41563_, _41422_, _41370_);
  and _48720_ (_41564_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  or _48721_ (_41565_, _41564_, _41563_);
  and _48722_ (_41566_, _41565_, _41399_);
  nand _48723_ (_41567_, _41268_, _38449_);
  nand _48724_ (_41568_, _41269_, _38456_);
  and _48725_ (_41569_, _41568_, _41402_);
  and _48726_ (_41570_, _41569_, _41567_);
  or _48727_ (_01263_, _41570_, _41566_);
  nor _48728_ (_41571_, _41422_, _41366_);
  and _48729_ (_41572_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or _48730_ (_41573_, _41572_, _41571_);
  and _48731_ (_41574_, _41573_, _41399_);
  nand _48732_ (_41575_, _41269_, _38449_);
  nand _48733_ (_41576_, _41268_, _38442_);
  and _48734_ (_41577_, _41576_, _41402_);
  and _48735_ (_41578_, _41577_, _41575_);
  or _48736_ (_01264_, _41578_, _41574_);
  and _48737_ (_41579_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _48738_ (_41580_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  or _48739_ (_41581_, _41580_, _41579_);
  and _48740_ (_41582_, _41581_, _41399_);
  nand _48741_ (_41583_, _41268_, _38434_);
  nand _48742_ (_41584_, _41269_, _38442_);
  and _48743_ (_41585_, _41584_, _41402_);
  and _48744_ (_41586_, _41585_, _41583_);
  or _48745_ (_01266_, _41586_, _41582_);
  and _48746_ (_41587_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _48747_ (_41588_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or _48748_ (_41589_, _41588_, _41587_);
  and _48749_ (_41590_, _41589_, _41399_);
  nand _48750_ (_41591_, _41269_, _38434_);
  nand _48751_ (_41592_, _41268_, _38428_);
  and _48752_ (_41593_, _41592_, _41402_);
  and _48753_ (_41594_, _41593_, _41591_);
  or _48754_ (_01268_, _41594_, _41590_);
  and _48755_ (_41595_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _48756_ (_41596_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  or _48757_ (_41597_, _41596_, _41595_);
  and _48758_ (_41598_, _41597_, _41399_);
  nand _48759_ (_41599_, _41268_, _38420_);
  nand _48760_ (_41600_, _41269_, _38428_);
  and _48761_ (_41602_, _41600_, _41402_);
  and _48762_ (_41604_, _41602_, _41599_);
  or _48763_ (_01270_, _41604_, _41598_);
  and _48764_ (_41607_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _48765_ (_41609_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or _48766_ (_41611_, _41609_, _41607_);
  and _48767_ (_41613_, _41611_, _41399_);
  nand _48768_ (_41615_, _41268_, _38485_);
  nand _48769_ (_41617_, _41269_, _38420_);
  and _48770_ (_41619_, _41617_, _41402_);
  and _48771_ (_41621_, _41619_, _41615_);
  or _48772_ (_01272_, _41621_, _41613_);
  and _48773_ (_41624_, _41398_, _41269_);
  nand _48774_ (_41626_, _41624_, _38485_);
  and _48775_ (_41628_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _48776_ (_41630_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _48777_ (_41632_, _41630_, _41628_);
  or _48778_ (_41634_, _41632_, _41398_);
  and _48779_ (_41636_, _41634_, _42882_);
  and _48780_ (_01274_, _41636_, _41626_);
  and _48781_ (_41639_, _41554_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _48782_ (_41641_, _41422_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _48783_ (_41643_, _41641_, _41639_);
  and _48784_ (_41645_, _41643_, _41399_);
  or _48785_ (_41647_, _41256_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _48786_ (_41649_, _41647_, _41269_);
  and _48787_ (_41651_, _41649_, _41402_);
  or _48788_ (_01276_, _41651_, _41645_);
  nand _48789_ (_41654_, _41426_, _38464_);
  or _48790_ (_41656_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _48791_ (_41658_, _41656_, _42882_);
  and _48792_ (_01278_, _41658_, _41654_);
  or _48793_ (_41661_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _48794_ (_41663_, _41661_, _42882_);
  nand _48795_ (_41665_, _41426_, _38456_);
  and _48796_ (_01280_, _41665_, _41663_);
  or _48797_ (_41666_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _48798_ (_41667_, _41666_, _42882_);
  nand _48799_ (_41668_, _41426_, _38449_);
  and _48800_ (_01282_, _41668_, _41667_);
  or _48801_ (_41669_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _48802_ (_41670_, _41669_, _42882_);
  nand _48803_ (_41671_, _41426_, _38442_);
  and _48804_ (_01284_, _41671_, _41670_);
  or _48805_ (_41672_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _48806_ (_41673_, _41672_, _42882_);
  nand _48807_ (_41674_, _41426_, _38434_);
  and _48808_ (_01286_, _41674_, _41673_);
  or _48809_ (_41675_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _48810_ (_41676_, _41675_, _42882_);
  nand _48811_ (_41677_, _41426_, _38428_);
  and _48812_ (_01288_, _41677_, _41676_);
  or _48813_ (_41678_, _41426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _48814_ (_41679_, _41678_, _42882_);
  nand _48815_ (_41680_, _41426_, _38420_);
  and _48816_ (_01290_, _41680_, _41679_);
  not _48817_ (_41681_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _48818_ (_41682_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _41681_);
  or _48819_ (_41683_, _41682_, _41268_);
  nor _48820_ (_41684_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _48821_ (_41685_, _41684_, _41683_);
  or _48822_ (_41686_, _41685_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _48823_ (_41687_, _41686_, _41430_);
  nand _48824_ (_41688_, _39065_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand _48825_ (_41689_, _41688_, _41430_);
  or _48826_ (_41690_, _41689_, _39070_);
  and _48827_ (_41691_, _41690_, _41687_);
  or _48828_ (_41692_, _41691_, _41433_);
  nand _48829_ (_41693_, _41433_, _38464_);
  and _48830_ (_41694_, _41693_, _42882_);
  and _48831_ (_01292_, _41694_, _41692_);
  or _48832_ (_41695_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or _48833_ (_41696_, _41695_, _41430_);
  not _48834_ (_41697_, _32567_);
  nor _48835_ (_41698_, _41697_, _31282_);
  nand _48836_ (_41699_, _41697_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _48837_ (_41700_, _41699_, _41430_);
  or _48838_ (_41701_, _41700_, _41698_);
  and _48839_ (_41702_, _41701_, _41696_);
  or _48840_ (_41703_, _41702_, _41433_);
  nand _48841_ (_41704_, _41433_, _38456_);
  and _48842_ (_41705_, _41704_, _42882_);
  and _48843_ (_01294_, _41705_, _41703_);
  not _48844_ (_41706_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  not _48845_ (_41707_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and _48846_ (_41708_, _41281_, _41707_);
  nor _48847_ (_41709_, _41708_, _41706_);
  and _48848_ (_41710_, _41708_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or _48849_ (_41711_, _41710_, _41709_);
  or _48850_ (_41712_, _41711_, _41430_);
  or _48851_ (_41713_, _33296_, _41706_);
  nand _48852_ (_41714_, _41713_, _41430_);
  or _48853_ (_41715_, _41714_, _33318_);
  and _48854_ (_41716_, _41715_, _41712_);
  or _48855_ (_41717_, _41716_, _41433_);
  nand _48856_ (_41718_, _41433_, _38449_);
  and _48857_ (_41719_, _41718_, _42882_);
  and _48858_ (_01296_, _41719_, _41717_);
  and _48859_ (_41720_, _41430_, _34004_);
  nand _48860_ (_41721_, _41720_, _31282_);
  or _48861_ (_41722_, _41720_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _48862_ (_41723_, _41722_, _41434_);
  and _48863_ (_41724_, _41723_, _41721_);
  nor _48864_ (_41725_, _41434_, _38442_);
  or _48865_ (_41726_, _41725_, _41724_);
  and _48866_ (_01298_, _41726_, _42882_);
  and _48867_ (_41727_, _41430_, _34765_);
  nand _48868_ (_41728_, _41727_, _31282_);
  or _48869_ (_41729_, _41727_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _48870_ (_41730_, _41729_, _41434_);
  and _48871_ (_41731_, _41730_, _41728_);
  nor _48872_ (_41732_, _41434_, _38434_);
  or _48873_ (_41733_, _41732_, _41731_);
  and _48874_ (_01299_, _41733_, _42882_);
  and _48875_ (_41734_, _41430_, _35549_);
  nand _48876_ (_41735_, _41734_, _31282_);
  or _48877_ (_41736_, _41734_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _48878_ (_41737_, _41736_, _41434_);
  and _48879_ (_41738_, _41737_, _41735_);
  nor _48880_ (_41739_, _41434_, _38428_);
  or _48881_ (_41740_, _41739_, _41738_);
  and _48882_ (_01301_, _41740_, _42882_);
  and _48883_ (_41741_, _41430_, _36277_);
  nand _48884_ (_41742_, _41741_, _31282_);
  or _48885_ (_41743_, _41741_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _48886_ (_41744_, _41743_, _41434_);
  and _48887_ (_41745_, _41744_, _41742_);
  nor _48888_ (_41746_, _41434_, _38420_);
  or _48889_ (_41747_, _41746_, _41745_);
  and _48890_ (_01303_, _41747_, _42882_);
  and _48891_ (_01628_, t2_i, _42882_);
  nor _48892_ (_41748_, t2_i, rst);
  and _48893_ (_01631_, _41748_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  nand _48894_ (_41749_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _42882_);
  nor _48895_ (_01634_, _41749_, t2ex_i);
  and _48896_ (_01637_, t2ex_i, _42882_);
  and _48897_ (_41750_, _38403_, _38895_);
  and _48898_ (_41751_, _41750_, _39993_);
  nand _48899_ (_41752_, _41751_, _38485_);
  and _48900_ (_41753_, _41750_, _39840_);
  not _48901_ (_41754_, _41753_);
  and _48902_ (_41755_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _48903_ (_41756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _48904_ (_41757_, _41756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _48905_ (_41758_, _41757_, _41755_);
  not _48906_ (_41759_, _41758_);
  and _48907_ (_41760_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _48908_ (_41761_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _48909_ (_41762_, _41761_, _41760_);
  or _48910_ (_41763_, _41751_, _41762_);
  and _48911_ (_41764_, _41763_, _41754_);
  and _48912_ (_41765_, _41764_, _41752_);
  and _48913_ (_41766_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _48914_ (_41767_, _41766_, _41765_);
  and _48915_ (_01640_, _41767_, _42882_);
  nand _48916_ (_41768_, _41753_, _38485_);
  nor _48917_ (_41769_, _41751_, _41759_);
  or _48918_ (_41770_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not _48919_ (_41771_, _41769_);
  or _48920_ (_41772_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _48921_ (_41773_, _41772_, _41770_);
  or _48922_ (_41774_, _41773_, _41753_);
  and _48923_ (_41775_, _41774_, _42882_);
  and _48924_ (_01643_, _41775_, _41768_);
  not _48925_ (_41776_, _41756_);
  or _48926_ (_41777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _48927_ (_41778_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _48928_ (_41779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _41778_);
  and _48929_ (_41780_, _41779_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _48930_ (_41781_, _41780_, _41777_);
  and _48931_ (_41782_, _41781_, _41776_);
  and _48932_ (_41783_, _41750_, _39954_);
  and _48933_ (_41784_, _39839_, _35549_);
  and _48934_ (_41785_, _41784_, _41750_);
  nor _48935_ (_41786_, _41785_, _41783_);
  and _48936_ (_41787_, _41786_, _41782_);
  and _48937_ (_41788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _48938_ (_41789_, _41788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _48939_ (_41790_, _41789_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _48940_ (_41791_, _41790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _48941_ (_41792_, _41791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _48942_ (_41793_, _41792_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _48943_ (_41794_, _41793_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _48944_ (_41795_, _41794_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _48945_ (_41796_, _41795_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _48946_ (_41797_, _41796_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _48947_ (_41798_, _41797_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _48948_ (_41799_, _41798_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _48949_ (_41800_, _41799_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _48950_ (_41801_, _41800_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _48951_ (_41802_, _41801_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not _48952_ (_41803_, _41802_);
  nand _48953_ (_41804_, _41803_, _41787_);
  or _48954_ (_41805_, _41787_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _48955_ (_41806_, _41805_, _42882_);
  and _48956_ (_01646_, _41806_, _41804_);
  nand _48957_ (_41807_, _41783_, _38485_);
  and _48958_ (_41808_, _41750_, _35549_);
  and _48959_ (_41809_, _41808_, _39839_);
  not _48960_ (_41810_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _48961_ (_41811_, _41755_, _41810_);
  and _48962_ (_41812_, _41811_, _41756_);
  and _48963_ (_41813_, _41812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  not _48964_ (_41814_, _41812_);
  not _48965_ (_41815_, _41757_);
  and _48966_ (_41816_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _48967_ (_41817_, _41802_, _41781_);
  and _48968_ (_41818_, _41817_, _41816_);
  and _48969_ (_41819_, _41793_, _41781_);
  or _48970_ (_41820_, _41819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand _48971_ (_41821_, _41819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _48972_ (_41822_, _41821_, _41820_);
  or _48973_ (_41823_, _41822_, _41818_);
  and _48974_ (_41824_, _41823_, _41814_);
  or _48975_ (_41825_, _41824_, _41813_);
  nor _48976_ (_41826_, _41825_, _41783_);
  nor _48977_ (_41827_, _41826_, _41809_);
  and _48978_ (_41828_, _41827_, _41807_);
  and _48979_ (_41829_, _41809_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _48980_ (_41830_, _41829_, _41828_);
  and _48981_ (_01649_, _41830_, _42882_);
  and _48982_ (_41831_, _41801_, _41781_);
  or _48983_ (_41832_, _41831_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _48984_ (_41833_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nand _48985_ (_41834_, _41833_, _41817_);
  and _48986_ (_41835_, _41834_, _41832_);
  or _48987_ (_41836_, _41835_, _41812_);
  or _48988_ (_41837_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _48989_ (_41838_, _41837_, _41786_);
  and _48990_ (_41839_, _41838_, _41836_);
  and _48991_ (_41840_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not _48992_ (_41841_, _41785_);
  nor _48993_ (_41842_, _41841_, _38485_);
  or _48994_ (_41843_, _41842_, _41840_);
  or _48995_ (_41844_, _41843_, _41839_);
  and _48996_ (_01652_, _41844_, _42882_);
  and _48997_ (_41845_, _41814_, _41781_);
  and _48998_ (_41846_, _41845_, _41756_);
  nand _48999_ (_41847_, _41846_, _41802_);
  nand _49000_ (_41848_, _41847_, _41786_);
  or _49001_ (_41849_, _41786_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _49002_ (_41850_, _41849_, _42882_);
  and _49003_ (_01655_, _41850_, _41848_);
  or _49004_ (_41851_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _49005_ (_41852_, _40546_, _38880_);
  or _49006_ (_41853_, _41852_, _41851_);
  nand _49007_ (_41854_, _38887_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _49008_ (_41855_, _41854_, _41852_);
  or _49009_ (_41856_, _41855_, _38888_);
  and _49010_ (_41857_, _41856_, _41853_);
  and _49011_ (_41858_, _41750_, _40542_);
  or _49012_ (_41859_, _41858_, _41857_);
  nand _49013_ (_41860_, _41858_, _38485_);
  and _49014_ (_41861_, _41860_, _42882_);
  and _49015_ (_01658_, _41861_, _41859_);
  or _49016_ (_41862_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  not _49017_ (_41863_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand _49018_ (_41864_, _41758_, _41863_);
  and _49019_ (_41865_, _41864_, _41862_);
  or _49020_ (_41866_, _41865_, _41751_);
  nand _49021_ (_41867_, _41751_, _38464_);
  and _49022_ (_41868_, _41867_, _41866_);
  or _49023_ (_41869_, _41868_, _41753_);
  or _49024_ (_41870_, _41754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _49025_ (_41871_, _41870_, _42882_);
  and _49026_ (_02108_, _41871_, _41869_);
  nand _49027_ (_41872_, _41751_, _38456_);
  and _49028_ (_41873_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _49029_ (_41874_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _49030_ (_41875_, _41874_, _41873_);
  or _49031_ (_41876_, _41875_, _41751_);
  and _49032_ (_41877_, _41876_, _41754_);
  and _49033_ (_41878_, _41877_, _41872_);
  and _49034_ (_41879_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _49035_ (_41880_, _41879_, _41878_);
  and _49036_ (_02109_, _41880_, _42882_);
  nand _49037_ (_41881_, _41751_, _38449_);
  and _49038_ (_41882_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _49039_ (_41883_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _49040_ (_41884_, _41883_, _41882_);
  or _49041_ (_41885_, _41884_, _41751_);
  and _49042_ (_41886_, _41885_, _41754_);
  and _49043_ (_41887_, _41886_, _41881_);
  and _49044_ (_41888_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _49045_ (_41889_, _41888_, _41887_);
  and _49046_ (_02111_, _41889_, _42882_);
  or _49047_ (_41890_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _49048_ (_41891_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _49049_ (_41892_, _41891_, _41890_);
  or _49050_ (_41893_, _41892_, _41751_);
  nand _49051_ (_41894_, _41751_, _38442_);
  and _49052_ (_41895_, _41894_, _41893_);
  or _49053_ (_41896_, _41895_, _41753_);
  or _49054_ (_41897_, _41754_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _49055_ (_41898_, _41897_, _42882_);
  and _49056_ (_02113_, _41898_, _41896_);
  nand _49057_ (_41899_, _41751_, _38434_);
  and _49058_ (_41900_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _49059_ (_41901_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _49060_ (_41902_, _41901_, _41900_);
  or _49061_ (_41903_, _41902_, _41751_);
  and _49062_ (_41904_, _41903_, _41754_);
  and _49063_ (_41905_, _41904_, _41899_);
  and _49064_ (_41906_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _49065_ (_41907_, _41906_, _41905_);
  and _49066_ (_02115_, _41907_, _42882_);
  nand _49067_ (_41908_, _41751_, _38428_);
  and _49068_ (_41909_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _49069_ (_41910_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _49070_ (_41911_, _41910_, _41909_);
  or _49071_ (_41912_, _41911_, _41751_);
  and _49072_ (_41913_, _41912_, _41754_);
  and _49073_ (_41914_, _41913_, _41908_);
  and _49074_ (_41915_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _49075_ (_41916_, _41915_, _41914_);
  and _49076_ (_02116_, _41916_, _42882_);
  nand _49077_ (_41917_, _41751_, _38420_);
  and _49078_ (_41918_, _41759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _49079_ (_41919_, _41758_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _49080_ (_41920_, _41919_, _41918_);
  or _49081_ (_41921_, _41920_, _41751_);
  and _49082_ (_41922_, _41921_, _41754_);
  and _49083_ (_41923_, _41922_, _41917_);
  and _49084_ (_41924_, _41753_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or _49085_ (_41925_, _41924_, _41923_);
  and _49086_ (_02118_, _41925_, _42882_);
  or _49087_ (_41926_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not _49088_ (_41927_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _49089_ (_41928_, _41769_, _41927_);
  and _49090_ (_41929_, _41928_, _41926_);
  or _49091_ (_41930_, _41929_, _41753_);
  nand _49092_ (_41931_, _41753_, _38464_);
  and _49093_ (_41932_, _41931_, _42882_);
  and _49094_ (_02120_, _41932_, _41930_);
  nand _49095_ (_41933_, _41753_, _38456_);
  and _49096_ (_41934_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _49097_ (_41935_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _49098_ (_41936_, _41935_, _41934_);
  or _49099_ (_41937_, _41936_, _41753_);
  and _49100_ (_41938_, _41937_, _42882_);
  and _49101_ (_02122_, _41938_, _41933_);
  nand _49102_ (_41939_, _41753_, _38449_);
  and _49103_ (_41940_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _49104_ (_41941_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _49105_ (_41942_, _41941_, _41940_);
  or _49106_ (_41943_, _41942_, _41753_);
  and _49107_ (_41944_, _41943_, _42882_);
  and _49108_ (_02123_, _41944_, _41939_);
  nand _49109_ (_41945_, _41753_, _38442_);
  and _49110_ (_41946_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _49111_ (_41947_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _49112_ (_41948_, _41947_, _41946_);
  or _49113_ (_41949_, _41948_, _41753_);
  and _49114_ (_41950_, _41949_, _42882_);
  and _49115_ (_02125_, _41950_, _41945_);
  nand _49116_ (_41951_, _41753_, _38434_);
  and _49117_ (_41952_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _49118_ (_41953_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _49119_ (_41954_, _41953_, _41952_);
  or _49120_ (_41955_, _41954_, _41753_);
  and _49121_ (_41956_, _41955_, _42882_);
  and _49122_ (_02127_, _41956_, _41951_);
  nand _49123_ (_41957_, _41753_, _38428_);
  and _49124_ (_41958_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _49125_ (_41959_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _49126_ (_41960_, _41959_, _41958_);
  or _49127_ (_41961_, _41960_, _41753_);
  and _49128_ (_41962_, _41961_, _42882_);
  and _49129_ (_02129_, _41962_, _41957_);
  nand _49130_ (_41963_, _41753_, _38420_);
  and _49131_ (_41964_, _41771_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _49132_ (_41965_, _41769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _49133_ (_41966_, _41965_, _41964_);
  or _49134_ (_41967_, _41966_, _41753_);
  and _49135_ (_41968_, _41967_, _42882_);
  and _49136_ (_02130_, _41968_, _41963_);
  or _49137_ (_41969_, _41781_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _49138_ (_41970_, _41781_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _49139_ (_41971_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _49140_ (_41972_, _41971_, _41802_);
  nand _49141_ (_41973_, _41972_, _41970_);
  and _49142_ (_41974_, _41973_, _41969_);
  or _49143_ (_41975_, _41974_, _41812_);
  nor _49144_ (_41976_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor _49145_ (_41977_, _41976_, _41783_);
  and _49146_ (_41978_, _41977_, _41975_);
  and _49147_ (_41979_, _41783_, _38465_);
  or _49148_ (_41980_, _41979_, _41809_);
  or _49149_ (_41981_, _41980_, _41978_);
  nand _49150_ (_41982_, _41785_, _41863_);
  and _49151_ (_41983_, _41982_, _42882_);
  and _49152_ (_02132_, _41983_, _41981_);
  and _49153_ (_41984_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _49154_ (_41985_, _41984_, _41845_);
  and _49155_ (_41986_, _41985_, _41802_);
  and _49156_ (_41987_, _41812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _49157_ (_41988_, _41970_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand _49158_ (_41989_, _41788_, _41781_);
  and _49159_ (_41990_, _41989_, _41814_);
  and _49160_ (_41991_, _41990_, _41988_);
  nor _49161_ (_41992_, _41991_, _41987_);
  nand _49162_ (_41993_, _41992_, _41786_);
  or _49163_ (_41994_, _41993_, _41986_);
  nand _49164_ (_41995_, _41783_, _38456_);
  or _49165_ (_41996_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _49166_ (_41997_, _41996_, _42882_);
  and _49167_ (_41998_, _41997_, _41995_);
  and _49168_ (_02134_, _41998_, _41994_);
  not _49169_ (_41999_, _41783_);
  or _49170_ (_42000_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _49171_ (_42001_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _49172_ (_42002_, _42001_, _41817_);
  and _49173_ (_42003_, _41989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor _49174_ (_42004_, _41989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _49175_ (_42005_, _42004_, _41812_);
  or _49176_ (_42006_, _42005_, _42003_);
  or _49177_ (_42007_, _42006_, _42002_);
  nand _49178_ (_42008_, _42007_, _42000_);
  nand _49179_ (_42009_, _42008_, _41999_);
  nand _49180_ (_42010_, _41783_, _38449_);
  and _49181_ (_42011_, _42010_, _42009_);
  or _49182_ (_42012_, _42011_, _41785_);
  or _49183_ (_42013_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _49184_ (_42014_, _42013_, _42882_);
  and _49185_ (_02136_, _42014_, _42012_);
  or _49186_ (_42015_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _49187_ (_42016_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _49188_ (_42017_, _42016_, _41817_);
  nand _49189_ (_42018_, _41789_, _41781_);
  and _49190_ (_42019_, _42018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _49191_ (_42020_, _42018_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _49192_ (_42021_, _42020_, _41812_);
  or _49193_ (_42022_, _42021_, _42019_);
  or _49194_ (_42023_, _42022_, _42017_);
  nand _49195_ (_42024_, _42023_, _42015_);
  nand _49196_ (_42025_, _42024_, _41999_);
  nand _49197_ (_42026_, _41783_, _38442_);
  and _49198_ (_42027_, _42026_, _42025_);
  or _49199_ (_42028_, _42027_, _41785_);
  or _49200_ (_42029_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _49201_ (_42030_, _42029_, _42882_);
  and _49202_ (_02137_, _42030_, _42028_);
  and _49203_ (_42031_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _49204_ (_42032_, _42031_, _41817_);
  nand _49205_ (_42033_, _41790_, _41781_);
  and _49206_ (_42034_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nor _49207_ (_42035_, _42033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _49208_ (_42036_, _42035_, _41812_);
  or _49209_ (_42037_, _42036_, _42034_);
  or _49210_ (_42038_, _42037_, _42032_);
  nor _49211_ (_42039_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor _49212_ (_42040_, _42039_, _41783_);
  and _49213_ (_42041_, _42040_, _42038_);
  nor _49214_ (_42042_, _41999_, _38434_);
  or _49215_ (_42043_, _42042_, _42041_);
  or _49216_ (_42044_, _42043_, _41809_);
  or _49217_ (_42045_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _49218_ (_42046_, _42045_, _42882_);
  and _49219_ (_02139_, _42046_, _42044_);
  and _49220_ (_42047_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _49221_ (_42048_, _42047_, _41817_);
  nand _49222_ (_42049_, _41791_, _41781_);
  and _49223_ (_42050_, _42049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor _49224_ (_42051_, _42049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _49225_ (_42052_, _42051_, _41812_);
  or _49226_ (_42053_, _42052_, _42050_);
  or _49227_ (_42054_, _42053_, _42048_);
  nor _49228_ (_42055_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor _49229_ (_42056_, _42055_, _41783_);
  and _49230_ (_42057_, _42056_, _42054_);
  nor _49231_ (_42058_, _41999_, _38428_);
  or _49232_ (_42059_, _42058_, _42057_);
  or _49233_ (_42060_, _42059_, _41809_);
  or _49234_ (_42061_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _49235_ (_42062_, _42061_, _42882_);
  and _49236_ (_02141_, _42062_, _42060_);
  nor _49237_ (_42063_, _41999_, _38420_);
  and _49238_ (_42064_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _49239_ (_42065_, _42064_, _41817_);
  and _49240_ (_42066_, _41792_, _41781_);
  nor _49241_ (_42067_, _42066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor _49242_ (_42068_, _42067_, _41819_);
  or _49243_ (_42069_, _42068_, _41812_);
  or _49244_ (_42070_, _42069_, _42065_);
  nor _49245_ (_42071_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor _49246_ (_42072_, _42071_, _41783_);
  and _49247_ (_42073_, _42072_, _42070_);
  or _49248_ (_42074_, _42073_, _41809_);
  or _49249_ (_42075_, _42074_, _42063_);
  or _49250_ (_42076_, _41841_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _49251_ (_42077_, _42076_, _42882_);
  and _49252_ (_02143_, _42077_, _42075_);
  and _49253_ (_42078_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _49254_ (_42079_, _42078_, _41817_);
  nand _49255_ (_42080_, _41821_, _41927_);
  or _49256_ (_42081_, _41821_, _41927_);
  and _49257_ (_42082_, _42081_, _42080_);
  or _49258_ (_42083_, _42082_, _41812_);
  or _49259_ (_42084_, _42083_, _42079_);
  nor _49260_ (_42085_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor _49261_ (_42086_, _42085_, _41783_);
  and _49262_ (_42087_, _42086_, _42084_);
  and _49263_ (_42088_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _49264_ (_42089_, _42088_, _41809_);
  or _49265_ (_42090_, _42089_, _42087_);
  nand _49266_ (_42091_, _41785_, _38464_);
  and _49267_ (_42092_, _42091_, _42882_);
  and _49268_ (_02144_, _42092_, _42090_);
  and _49269_ (_42093_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _49270_ (_42094_, _42093_, _41817_);
  and _49271_ (_42095_, _41795_, _41781_);
  or _49272_ (_42096_, _42095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand _49273_ (_42097_, _42095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _49274_ (_42098_, _42097_, _42096_);
  or _49275_ (_42099_, _42098_, _41812_);
  or _49276_ (_42100_, _42099_, _42094_);
  nor _49277_ (_42101_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _49278_ (_42102_, _42101_, _41783_);
  and _49279_ (_42103_, _42102_, _42100_);
  and _49280_ (_42104_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _49281_ (_42105_, _42104_, _41809_);
  or _49282_ (_42106_, _42105_, _42103_);
  nand _49283_ (_42107_, _41809_, _38456_);
  and _49284_ (_42108_, _42107_, _42882_);
  and _49285_ (_02145_, _42108_, _42106_);
  and _49286_ (_42109_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _49287_ (_42110_, _42109_, _41817_);
  nand _49288_ (_42111_, _41796_, _41781_);
  and _49289_ (_42112_, _42111_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor _49290_ (_42113_, _42111_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _49291_ (_42114_, _42113_, _41812_);
  or _49292_ (_42115_, _42114_, _42112_);
  or _49293_ (_42116_, _42115_, _42110_);
  nor _49294_ (_42117_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _49295_ (_42118_, _42117_, _41783_);
  and _49296_ (_42119_, _42118_, _42116_);
  and _49297_ (_42120_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _49298_ (_42121_, _42120_, _41809_);
  or _49299_ (_42122_, _42121_, _42119_);
  nand _49300_ (_42123_, _41809_, _38449_);
  and _49301_ (_42124_, _42123_, _42882_);
  and _49302_ (_02146_, _42124_, _42122_);
  and _49303_ (_42125_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _49304_ (_42126_, _42125_, _41817_);
  nand _49305_ (_42127_, _41797_, _41781_);
  and _49306_ (_42128_, _42127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor _49307_ (_42129_, _42127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _49308_ (_42130_, _42129_, _41812_);
  or _49309_ (_42131_, _42130_, _42128_);
  or _49310_ (_42132_, _42131_, _42126_);
  nor _49311_ (_42133_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor _49312_ (_42134_, _42133_, _41783_);
  and _49313_ (_42135_, _42134_, _42132_);
  and _49314_ (_42136_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _49315_ (_42137_, _42136_, _41809_);
  or _49316_ (_42138_, _42137_, _42135_);
  nand _49317_ (_42139_, _41809_, _38442_);
  and _49318_ (_42140_, _42139_, _42882_);
  and _49319_ (_02147_, _42140_, _42138_);
  nand _49320_ (_42141_, _41785_, _38434_);
  and _49321_ (_42142_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _49322_ (_42143_, _42142_, _41817_);
  nand _49323_ (_42144_, _41798_, _41781_);
  and _49324_ (_42145_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _49325_ (_42146_, _42144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _49326_ (_42147_, _42146_, _41812_);
  or _49327_ (_42148_, _42147_, _42145_);
  or _49328_ (_42149_, _42148_, _42143_);
  nor _49329_ (_42150_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor _49330_ (_42151_, _42150_, _41783_);
  and _49331_ (_42152_, _42151_, _42149_);
  and _49332_ (_42153_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _49333_ (_42154_, _42153_, _41809_);
  or _49334_ (_42155_, _42154_, _42152_);
  and _49335_ (_42156_, _42155_, _42882_);
  and _49336_ (_02148_, _42156_, _42141_);
  and _49337_ (_42157_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _49338_ (_42158_, _42157_, _41817_);
  nand _49339_ (_42159_, _41799_, _41781_);
  and _49340_ (_42160_, _42159_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor _49341_ (_42161_, _42159_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _49342_ (_42162_, _42161_, _41812_);
  or _49343_ (_42163_, _42162_, _42160_);
  or _49344_ (_42164_, _42163_, _42158_);
  nor _49345_ (_42165_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor _49346_ (_42166_, _42165_, _41783_);
  and _49347_ (_42167_, _42166_, _42164_);
  and _49348_ (_42168_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _49349_ (_42169_, _42168_, _41809_);
  or _49350_ (_42170_, _42169_, _42167_);
  nand _49351_ (_42171_, _41809_, _38428_);
  and _49352_ (_42172_, _42171_, _42882_);
  and _49353_ (_02149_, _42172_, _42170_);
  and _49354_ (_42173_, _41815_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _49355_ (_42174_, _42173_, _41817_);
  and _49356_ (_42175_, _41800_, _41781_);
  nor _49357_ (_42176_, _42175_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _49358_ (_42177_, _42176_, _41831_);
  or _49359_ (_42178_, _42177_, _41812_);
  or _49360_ (_42179_, _42178_, _42174_);
  nor _49361_ (_42180_, _41814_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor _49362_ (_42181_, _42180_, _41783_);
  and _49363_ (_42182_, _42181_, _42179_);
  and _49364_ (_42183_, _41783_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _49365_ (_42184_, _42183_, _41809_);
  or _49366_ (_42185_, _42184_, _42182_);
  nand _49367_ (_42186_, _41809_, _38420_);
  and _49368_ (_42187_, _42186_, _42882_);
  and _49369_ (_02150_, _42187_, _42185_);
  and _49370_ (_42188_, _41852_, _27045_);
  nand _49371_ (_42189_, _42188_, _31282_);
  or _49372_ (_42190_, _42188_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _49373_ (_42191_, _42190_, _42189_);
  or _49374_ (_42192_, _42191_, _41858_);
  nand _49375_ (_42193_, _41858_, _38464_);
  and _49376_ (_42194_, _42193_, _42882_);
  and _49377_ (_02151_, _42194_, _42192_);
  not _49378_ (_42195_, _41858_);
  and _49379_ (_42196_, _41852_, _32567_);
  or _49380_ (_42197_, _42196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _49381_ (_42198_, _42197_, _42195_);
  nand _49382_ (_42199_, _42196_, _31282_);
  and _49383_ (_42200_, _42199_, _42198_);
  nor _49384_ (_42201_, _42195_, _38456_);
  or _49385_ (_42202_, _42201_, _42200_);
  and _49386_ (_02152_, _42202_, _42882_);
  nand _49387_ (_42203_, _41852_, _39293_);
  and _49388_ (_42204_, _42203_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _49389_ (_42205_, _42204_, _41858_);
  and _49390_ (_42206_, _33329_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _49391_ (_42207_, _42206_, _33318_);
  and _49392_ (_42208_, _42207_, _41852_);
  or _49393_ (_42209_, _42208_, _42205_);
  nand _49394_ (_42210_, _41858_, _38449_);
  and _49395_ (_42211_, _42210_, _42882_);
  and _49396_ (_02153_, _42211_, _42209_);
  and _49397_ (_42212_, _41852_, _34004_);
  or _49398_ (_42213_, _42212_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _49399_ (_42214_, _42213_, _42195_);
  nand _49400_ (_42215_, _42212_, _31282_);
  and _49401_ (_42216_, _42215_, _42214_);
  nor _49402_ (_42217_, _42195_, _38442_);
  or _49403_ (_42218_, _42217_, _42216_);
  and _49404_ (_02154_, _42218_, _42882_);
  and _49405_ (_42219_, _41852_, _34765_);
  or _49406_ (_42220_, _42219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _49407_ (_42221_, _42220_, _42195_);
  nand _49408_ (_42222_, _42219_, _31282_);
  and _49409_ (_42223_, _42222_, _42221_);
  nor _49410_ (_42224_, _42195_, _38434_);
  or _49411_ (_42225_, _42224_, _42223_);
  and _49412_ (_02155_, _42225_, _42882_);
  and _49413_ (_42226_, _41852_, _35549_);
  nand _49414_ (_42227_, _42226_, _31282_);
  or _49415_ (_42228_, _42226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _49416_ (_42229_, _42228_, _42227_);
  or _49417_ (_42230_, _42229_, _41858_);
  nand _49418_ (_42231_, _41858_, _38428_);
  and _49419_ (_42232_, _42231_, _42882_);
  and _49420_ (_02156_, _42232_, _42230_);
  not _49421_ (_42233_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _49422_ (_42234_, _41755_, _42233_);
  or _49423_ (_42235_, _42234_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _49424_ (_42236_, _42235_, _41852_);
  nand _49425_ (_42237_, _39006_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _49426_ (_42238_, _42237_, _41852_);
  or _49427_ (_42239_, _42238_, _39007_);
  and _49428_ (_42240_, _42239_, _42236_);
  or _49429_ (_42241_, _42240_, _41858_);
  nand _49430_ (_42242_, _41858_, _38420_);
  and _49431_ (_42243_, _42242_, _42882_);
  and _49432_ (_02157_, _42243_, _42241_);
  and _49433_ (_42244_, _30646_, _27527_);
  not _49434_ (_42245_, _38487_);
  and _49435_ (_42246_, _42245_, _38399_);
  not _49436_ (_42247_, _42246_);
  not _49437_ (_42248_, _38398_);
  nor _49438_ (_42249_, _42248_, _38357_);
  not _49439_ (_42250_, _36450_);
  and _49440_ (_42251_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [7]);
  and _49441_ (_42252_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _49442_ (_42253_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _49443_ (_42254_, _42253_, _42252_);
  and _49444_ (_42255_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _49445_ (_42256_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _49446_ (_42257_, _42256_, _42255_);
  and _49447_ (_42258_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _49448_ (_42259_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _49449_ (_42260_, _42259_, _42258_);
  and _49450_ (_42261_, _42260_, _42257_);
  and _49451_ (_42262_, _42261_, _42254_);
  nor _49452_ (_42263_, _36636_, _42250_);
  not _49453_ (_42264_, _42263_);
  nor _49454_ (_42265_, _42264_, _42262_);
  nor _49455_ (_42266_, _42265_, _42251_);
  not _49456_ (_42267_, _42266_);
  and _49457_ (_42268_, _42267_, _42249_);
  not _49458_ (_42269_, _42268_);
  not _49459_ (_42270_, _38257_);
  and _49460_ (_42271_, _42248_, _38357_);
  nor _49461_ (_42272_, _38901_, _38948_);
  nor _49462_ (_42273_, _42272_, _38954_);
  and _49463_ (_42274_, _42273_, _27714_);
  nor _49464_ (_42275_, _30657_, \oc8051_top_1.oc8051_indi_addr1.wr_bit_r );
  and _49465_ (_42276_, _42275_, _33329_);
  not _49466_ (_42277_, _42276_);
  nor _49467_ (_42278_, _42277_, _42274_);
  nor _49468_ (_42279_, _42273_, _27714_);
  and _49469_ (_42280_, _37960_, _27023_);
  nor _49470_ (_42281_, _37960_, _27023_);
  nor _49471_ (_42282_, _42281_, _42280_);
  not _49472_ (_42283_, _42282_);
  nor _49473_ (_42284_, _42283_, _42279_);
  and _49474_ (_42285_, _42284_, _42278_);
  not _49475_ (_42286_, _42285_);
  and _49476_ (_42287_, _42273_, _38262_);
  and _49477_ (_42288_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor _49478_ (_42289_, _42273_, _37960_);
  and _49479_ (_42290_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor _49480_ (_42291_, _42290_, _42288_);
  nor _49481_ (_42292_, _42273_, _38262_);
  and _49482_ (_42293_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _49483_ (_42294_, _42273_, _37960_);
  and _49484_ (_42295_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor _49485_ (_42296_, _42295_, _42293_);
  and _49486_ (_42297_, _42296_, _42291_);
  and _49487_ (_42298_, _42297_, _42286_);
  and _49488_ (_42299_, _42285_, _38485_);
  nor _49489_ (_42300_, _42299_, _42298_);
  and _49490_ (_42301_, _42300_, _42271_);
  nor _49491_ (_42302_, _42301_, _42270_);
  and _49492_ (_42303_, _42302_, _42269_);
  and _49493_ (_42304_, _42303_, _42247_);
  and _49494_ (_42305_, _38246_, _38317_);
  nor _49495_ (_42306_, _42305_, _38325_);
  not _49496_ (_42307_, _42306_);
  nor _49497_ (_42308_, _42307_, _38273_);
  and _49498_ (_42309_, _42308_, _38319_);
  and _49499_ (_42310_, _38246_, _37707_);
  nor _49500_ (_42311_, _42310_, _38320_);
  and _49501_ (_42312_, _42311_, _38341_);
  and _49502_ (_42313_, _42312_, _42309_);
  and _49503_ (_42314_, _42313_, _38268_);
  nor _49504_ (_42315_, _42314_, _36407_);
  nor _49505_ (_42316_, _38339_, _38335_);
  not _49506_ (_42317_, _38243_);
  nor _49507_ (_42318_, _42317_, _42316_);
  nor _49508_ (_42319_, _42318_, _42315_);
  not _49509_ (_42320_, _42319_);
  and _49510_ (_42321_, _42320_, _42304_);
  and _49511_ (_42322_, _42249_, _38257_);
  and _49512_ (_42323_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [4]);
  and _49513_ (_42324_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _49514_ (_42325_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _49515_ (_42326_, _42325_, _42324_);
  and _49516_ (_42327_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _49517_ (_42328_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _49518_ (_42329_, _42328_, _42327_);
  and _49519_ (_42330_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _49520_ (_42331_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _49521_ (_42332_, _42331_, _42330_);
  and _49522_ (_42333_, _42332_, _42329_);
  and _49523_ (_42334_, _42333_, _42326_);
  nor _49524_ (_42335_, _42334_, _42264_);
  nor _49525_ (_42336_, _42335_, _42323_);
  not _49526_ (_42337_, _42336_);
  and _49527_ (_42338_, _42337_, _42322_);
  and _49528_ (_42339_, _38398_, _38357_);
  and _49529_ (_42340_, _42339_, _38257_);
  and _49530_ (_42341_, _38904_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor _49531_ (_42342_, _42341_, _38966_);
  not _49532_ (_42343_, _42342_);
  and _49533_ (_42344_, _42343_, _42340_);
  nor _49534_ (_42345_, _42344_, _42338_);
  and _49535_ (_42346_, _42271_, _38257_);
  nor _49536_ (_42347_, _42286_, _38434_);
  and _49537_ (_42348_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _49538_ (_42349_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _49539_ (_42350_, _42349_, _42348_);
  and _49540_ (_42351_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _49541_ (_42352_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor _49542_ (_42353_, _42352_, _42351_);
  and _49543_ (_42354_, _42353_, _42350_);
  nor _49544_ (_42355_, _42354_, _42285_);
  nor _49545_ (_42356_, _42355_, _42347_);
  not _49546_ (_42357_, _42356_);
  and _49547_ (_42358_, _42357_, _42346_);
  not _49548_ (_42359_, _42358_);
  not _49549_ (_42360_, _38519_);
  and _49550_ (_42361_, _42360_, _38400_);
  and _49551_ (_42362_, _42270_, _38398_);
  nor _49552_ (_42363_, _42362_, _42361_);
  and _49553_ (_42364_, _42363_, _42359_);
  and _49554_ (_42365_, _42364_, _42345_);
  not _49555_ (_42366_, _42365_);
  and _49556_ (_42367_, _42366_, _42321_);
  and _49557_ (_42368_, _42271_, _42270_);
  and _49558_ (_42369_, _42340_, _38190_);
  or _49559_ (_42370_, _42369_, _42368_);
  and _49560_ (_42371_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [1]);
  and _49561_ (_42372_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _49562_ (_42373_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _49563_ (_42374_, _42373_, _42372_);
  and _49564_ (_42375_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _49565_ (_42376_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _49566_ (_42377_, _42376_, _42375_);
  and _49567_ (_42378_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _49568_ (_42379_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _49569_ (_42380_, _42379_, _42378_);
  and _49570_ (_42381_, _42380_, _42377_);
  and _49571_ (_42382_, _42381_, _42374_);
  nor _49572_ (_42383_, _42382_, _42264_);
  nor _49573_ (_42384_, _42383_, _42371_);
  not _49574_ (_42385_, _42384_);
  and _49575_ (_42386_, _42385_, _42322_);
  not _49576_ (_42387_, _38501_);
  and _49577_ (_42388_, _42387_, _38400_);
  and _49578_ (_42389_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _49579_ (_42390_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _49580_ (_42391_, _42390_, _42389_);
  and _49581_ (_42392_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _49582_ (_42393_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor _49583_ (_42394_, _42393_, _42392_);
  and _49584_ (_42395_, _42394_, _42391_);
  and _49585_ (_42396_, _42395_, _42286_);
  and _49586_ (_42397_, _42285_, _38456_);
  nor _49587_ (_42398_, _42397_, _42396_);
  and _49588_ (_42399_, _42398_, _42346_);
  or _49589_ (_42400_, _42399_, _42388_);
  or _49590_ (_42401_, _42400_, _42386_);
  nor _49591_ (_42402_, _42401_, _42370_);
  nor _49592_ (_42403_, _42402_, _42320_);
  nor _49593_ (_42404_, _42403_, _42367_);
  not _49594_ (_42405_, _27845_);
  and _49595_ (_42406_, _27549_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49596_ (_42407_, _42406_, _42405_);
  nor _49597_ (_42408_, _26902_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _49598_ (_42409_, _42408_, _42407_);
  nand _49599_ (_42410_, _42409_, _42404_);
  or _49600_ (_42411_, _42409_, _42404_);
  and _49601_ (_42412_, _42411_, _42410_);
  not _49602_ (_42413_, _42412_);
  not _49603_ (_42414_, _42273_);
  and _49604_ (_42415_, _42340_, _42414_);
  and _49605_ (_42416_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [3]);
  and _49606_ (_42417_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _49607_ (_42418_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _49608_ (_42419_, _42418_, _42417_);
  and _49609_ (_42420_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _49610_ (_42421_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _49611_ (_42422_, _42421_, _42420_);
  and _49612_ (_42423_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _49613_ (_42424_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _49614_ (_42425_, _42424_, _42423_);
  and _49615_ (_42426_, _42425_, _42422_);
  and _49616_ (_42427_, _42426_, _42419_);
  nor _49617_ (_42428_, _42427_, _42264_);
  nor _49618_ (_42429_, _42428_, _42416_);
  not _49619_ (_42430_, _42429_);
  and _49620_ (_42431_, _42430_, _42322_);
  nor _49621_ (_42432_, _42431_, _42415_);
  not _49622_ (_42433_, _38513_);
  and _49623_ (_42434_, _42433_, _38400_);
  and _49624_ (_42435_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _49625_ (_42436_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor _49626_ (_42437_, _42436_, _42435_);
  and _49627_ (_42438_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and _49628_ (_42439_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor _49629_ (_42440_, _42439_, _42438_);
  and _49630_ (_42441_, _42440_, _42437_);
  nor _49631_ (_42442_, _42441_, _42285_);
  nor _49632_ (_42443_, _42286_, _38442_);
  nor _49633_ (_42444_, _42443_, _42442_);
  not _49634_ (_42445_, _42444_);
  and _49635_ (_42446_, _42445_, _42346_);
  nor _49636_ (_42447_, _42446_, _42434_);
  and _49637_ (_42448_, _42447_, _42432_);
  not _49638_ (_42449_, _42448_);
  and _49639_ (_42450_, _42449_, _42321_);
  and _49640_ (_42451_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [0]);
  and _49641_ (_42452_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _49642_ (_42453_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor _49643_ (_42454_, _42453_, _42452_);
  and _49644_ (_42455_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _49645_ (_42456_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _49646_ (_42457_, _42456_, _42455_);
  and _49647_ (_42458_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _49648_ (_42459_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _49649_ (_42460_, _42459_, _42458_);
  and _49650_ (_42461_, _42460_, _42457_);
  and _49651_ (_42462_, _42461_, _42454_);
  nor _49652_ (_42463_, _42462_, _42264_);
  nor _49653_ (_42464_, _42463_, _42451_);
  not _49654_ (_42465_, _42464_);
  and _49655_ (_42466_, _42465_, _42322_);
  and _49656_ (_42467_, _42285_, _38465_);
  and _49657_ (_42468_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _49658_ (_42469_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _49659_ (_42470_, _42469_, _42468_);
  and _49660_ (_42471_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and _49661_ (_42472_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor _49662_ (_42473_, _42472_, _42471_);
  and _49663_ (_42474_, _42473_, _42470_);
  nor _49664_ (_42475_, _42474_, _42285_);
  nor _49665_ (_42476_, _42475_, _42467_);
  not _49666_ (_42477_, _42476_);
  and _49667_ (_42478_, _42477_, _42346_);
  nor _49668_ (_42479_, _42478_, _42466_);
  not _49669_ (_42480_, _38495_);
  and _49670_ (_42481_, _42480_, _38400_);
  and _49671_ (_42482_, _42340_, _37960_);
  nor _49672_ (_42483_, _42482_, _42481_);
  and _49673_ (_42484_, _42483_, _42479_);
  nor _49674_ (_42485_, _42484_, _42320_);
  nor _49675_ (_42486_, _42485_, _42450_);
  and _49676_ (_42487_, _42406_, _27714_);
  nor _49677_ (_42488_, _27023_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _49678_ (_42489_, _42488_, _42487_);
  not _49679_ (_42490_, _42489_);
  and _49680_ (_42491_, _42490_, _42486_);
  nor _49681_ (_42492_, _42490_, _42486_);
  nor _49682_ (_42493_, _42492_, _42491_);
  and _49683_ (_42494_, _42493_, _42413_);
  nor _49684_ (_42495_, _42271_, _38257_);
  and _49685_ (_42496_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _49686_ (_42497_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor _49687_ (_42498_, _42497_, _42496_);
  and _49688_ (_42499_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _49689_ (_42500_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor _49690_ (_42501_, _42500_, _42499_);
  and _49691_ (_42502_, _42501_, _42498_);
  and _49692_ (_42503_, _42502_, _42286_);
  and _49693_ (_42504_, _42285_, _38420_);
  nor _49694_ (_42505_, _42504_, _42503_);
  and _49695_ (_42506_, _42505_, _42346_);
  nor _49696_ (_42507_, _42506_, _42495_);
  not _49697_ (_42508_, _38531_);
  and _49698_ (_42509_, _42508_, _38400_);
  and _49699_ (_42510_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [6]);
  and _49700_ (_42511_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _49701_ (_42512_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _49702_ (_42513_, _42512_, _42511_);
  and _49703_ (_42514_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _49704_ (_42515_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _49705_ (_42516_, _42515_, _42514_);
  and _49706_ (_42517_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _49707_ (_42518_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _49708_ (_42519_, _42518_, _42517_);
  and _49709_ (_42520_, _42519_, _42516_);
  and _49710_ (_42521_, _42520_, _42513_);
  nor _49711_ (_42522_, _42521_, _42264_);
  nor _49712_ (_42523_, _42522_, _42510_);
  not _49713_ (_42524_, _42523_);
  and _49714_ (_42525_, _42524_, _42322_);
  nor _49715_ (_42526_, _42525_, _42509_);
  and _49716_ (_42527_, _42526_, _42507_);
  and _49717_ (_42528_, _42527_, _42321_);
  nor _49718_ (_42529_, _42449_, _42321_);
  nor _49719_ (_42530_, _42529_, _42528_);
  nor _49720_ (_42531_, _42406_, _27714_);
  and _49721_ (_42532_, _42406_, _27242_);
  nor _49722_ (_42533_, _42532_, _42531_);
  not _49723_ (_42534_, _42533_);
  and _49724_ (_42535_, _42534_, _42530_);
  nor _49725_ (_42536_, _42534_, _42530_);
  nor _49726_ (_42537_, _42536_, _42535_);
  and _49727_ (_42538_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [5]);
  and _49728_ (_42539_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _49729_ (_42540_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _49730_ (_42541_, _42540_, _42539_);
  and _49731_ (_42542_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _49732_ (_42543_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _49733_ (_42544_, _42543_, _42542_);
  and _49734_ (_42545_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _49735_ (_42546_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _49736_ (_42547_, _42546_, _42545_);
  and _49737_ (_42548_, _42547_, _42544_);
  and _49738_ (_42549_, _42548_, _42541_);
  nor _49739_ (_42550_, _42549_, _42264_);
  nor _49740_ (_42551_, _42550_, _42538_);
  not _49741_ (_42552_, _42551_);
  and _49742_ (_42553_, _42552_, _42322_);
  and _49743_ (_42554_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  not _49744_ (_42555_, _42554_);
  and _49745_ (_42556_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _49746_ (_42557_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor _49747_ (_42558_, _42557_, _42556_);
  and _49748_ (_42559_, _42558_, _42555_);
  and _49749_ (_42560_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor _49750_ (_42561_, _42560_, _42285_);
  and _49751_ (_42562_, _42561_, _42559_);
  and _49752_ (_42563_, _42285_, _38428_);
  or _49753_ (_42564_, _42563_, _42562_);
  not _49754_ (_42565_, _42564_);
  and _49755_ (_42566_, _42565_, _42346_);
  nor _49756_ (_42567_, _42566_, _42553_);
  nor _49757_ (_42568_, _38525_, _38398_);
  nor _49758_ (_42569_, _42568_, _42270_);
  or _49759_ (_42570_, _42249_, _42271_);
  nor _49760_ (_42571_, _42570_, _42569_);
  not _49761_ (_42572_, _42571_);
  and _49762_ (_42573_, _42572_, _42567_);
  not _49763_ (_42574_, _42573_);
  and _49764_ (_42575_, _42574_, _42321_);
  and _49765_ (_42576_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op2_buff [2]);
  and _49766_ (_42577_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _49767_ (_42578_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _49768_ (_42579_, _42578_, _42577_);
  and _49769_ (_42580_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _49770_ (_42581_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _49771_ (_42582_, _42581_, _42580_);
  and _49772_ (_42583_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _49773_ (_42584_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _49774_ (_42585_, _42584_, _42583_);
  and _49775_ (_42586_, _42585_, _42582_);
  and _49776_ (_42587_, _42586_, _42579_);
  nor _49777_ (_42588_, _42587_, _42264_);
  nor _49778_ (_42589_, _42588_, _42576_);
  not _49779_ (_42590_, _42589_);
  and _49780_ (_42591_, _42590_, _42322_);
  and _49781_ (_42592_, _42294_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _49782_ (_42593_, _42289_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _49783_ (_42594_, _42593_, _42592_);
  and _49784_ (_42595_, _42292_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _49785_ (_42596_, _42287_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor _49786_ (_42597_, _42596_, _42595_);
  and _49787_ (_42598_, _42597_, _42594_);
  nor _49788_ (_42599_, _42598_, _42285_);
  not _49789_ (_42600_, _38449_);
  and _49790_ (_42601_, _42285_, _42600_);
  nor _49791_ (_42602_, _42601_, _42599_);
  not _49792_ (_42603_, _42602_);
  and _49793_ (_42604_, _42603_, _42346_);
  nor _49794_ (_42605_, _42604_, _42591_);
  not _49795_ (_42606_, _38507_);
  and _49796_ (_42607_, _42606_, _38400_);
  and _49797_ (_42608_, _42340_, _38167_);
  nor _49798_ (_42609_, _42608_, _42607_);
  and _49799_ (_42610_, _42609_, _42605_);
  nor _49800_ (_42611_, _42610_, _42320_);
  nor _49801_ (_42612_, _42611_, _42575_);
  and _49802_ (_42613_, _42406_, _38879_);
  nor _49803_ (_42614_, _26781_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor _49804_ (_42615_, _42614_, _42613_);
  not _49805_ (_42616_, _42615_);
  nor _49806_ (_42617_, _42616_, _42612_);
  and _49807_ (_42618_, _42616_, _42612_);
  nor _49808_ (_42619_, _42618_, _42617_);
  and _49809_ (_42620_, _42619_, _42537_);
  and _49810_ (_42621_, _42620_, _42494_);
  and _49811_ (_42622_, _42621_, _42244_);
  nor _49812_ (_42623_, _42365_, _42321_);
  nor _49813_ (_42624_, _42406_, _27845_);
  not _49814_ (_42625_, _42624_);
  and _49815_ (_42626_, _42625_, _42623_);
  nor _49816_ (_42627_, _42625_, _42623_);
  nor _49817_ (_42628_, _42627_, _42626_);
  nor _49818_ (_42629_, _42574_, _42321_);
  nor _49819_ (_42630_, _42406_, _38879_);
  not _49820_ (_42631_, _42630_);
  and _49821_ (_42632_, _42631_, _42629_);
  nor _49822_ (_42633_, _42631_, _42629_);
  nor _49823_ (_42634_, _42633_, _42632_);
  and _49824_ (_42635_, _42634_, _42628_);
  nor _49825_ (_42636_, _42304_, _27549_);
  and _49826_ (_42637_, _42304_, _27549_);
  nor _49827_ (_42638_, _42637_, _42636_);
  not _49828_ (_42639_, _42638_);
  nor _49829_ (_42640_, _42527_, _42321_);
  nor _49830_ (_42641_, _42406_, _27242_);
  not _49831_ (_42642_, _42641_);
  nor _49832_ (_42643_, _42642_, _42640_);
  and _49833_ (_42644_, _42642_, _42640_);
  nor _49834_ (_42645_, _42644_, _42643_);
  and _49835_ (_42646_, _42645_, _42639_);
  and _49836_ (_42647_, _42646_, _42635_);
  and _49837_ (_42648_, _42647_, _42622_);
  not _49838_ (_42649_, _42612_);
  not _49839_ (_42650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor _49840_ (_42651_, _42486_, _42650_);
  and _49841_ (_42652_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  or _49842_ (_42653_, _42652_, _42404_);
  or _49843_ (_42654_, _42653_, _42651_);
  and _49844_ (_42655_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  not _49845_ (_42656_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  or _49846_ (_42657_, _42486_, _42656_);
  nand _49847_ (_42658_, _42657_, _42404_);
  or _49848_ (_42659_, _42658_, _42655_);
  and _49849_ (_42660_, _42659_, _42654_);
  or _49850_ (_42661_, _42660_, _42649_);
  not _49851_ (_42662_, _42530_);
  not _49852_ (_42663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor _49853_ (_42664_, _42486_, _42663_);
  and _49854_ (_42665_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  or _49855_ (_42666_, _42665_, _42404_);
  or _49856_ (_42667_, _42666_, _42664_);
  and _49857_ (_42668_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not _49858_ (_42669_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  or _49859_ (_42670_, _42486_, _42669_);
  nand _49860_ (_42671_, _42670_, _42404_);
  or _49861_ (_42672_, _42671_, _42668_);
  and _49862_ (_42673_, _42672_, _42667_);
  or _49863_ (_42674_, _42673_, _42612_);
  and _49864_ (_42675_, _42674_, _42662_);
  and _49865_ (_42676_, _42675_, _42661_);
  not _49866_ (_42677_, _42404_);
  not _49867_ (_42678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand _49868_ (_42679_, _42486_, _42678_);
  or _49869_ (_42680_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  and _49870_ (_42681_, _42680_, _42679_);
  or _49871_ (_42682_, _42681_, _42677_);
  or _49872_ (_42683_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  not _49873_ (_42684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nand _49874_ (_42685_, _42486_, _42684_);
  and _49875_ (_42686_, _42685_, _42683_);
  or _49876_ (_42687_, _42686_, _42404_);
  and _49877_ (_42688_, _42687_, _42682_);
  or _49878_ (_42689_, _42688_, _42649_);
  not _49879_ (_42690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand _49880_ (_42691_, _42486_, _42690_);
  or _49881_ (_42692_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  and _49882_ (_42693_, _42692_, _42691_);
  or _49883_ (_42694_, _42693_, _42677_);
  or _49884_ (_42695_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  not _49885_ (_42696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nand _49886_ (_42697_, _42486_, _42696_);
  and _49887_ (_42698_, _42697_, _42695_);
  or _49888_ (_42699_, _42698_, _42404_);
  and _49889_ (_42700_, _42699_, _42694_);
  or _49890_ (_42701_, _42700_, _42612_);
  and _49891_ (_42702_, _42701_, _42530_);
  and _49892_ (_42703_, _42702_, _42689_);
  nor _49893_ (_42704_, _42703_, _42676_);
  nor _49894_ (_42705_, _42704_, _42648_);
  not _49895_ (_42706_, _42622_);
  nor _49896_ (_42707_, _42648_, _42706_);
  and _49897_ (_42708_, _42648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  or _49898_ (_42709_, _42708_, _42707_);
  or _49899_ (_42710_, _42709_, _42705_);
  nor _49900_ (_42711_, _42707_, rst);
  and _49901_ (_42712_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nand _49902_ (_42713_, _42712_, _28723_);
  nor _49903_ (_42714_, _42713_, _31282_);
  nand _49904_ (_42715_, _28723_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _49905_ (_42716_, _20040_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49906_ (_42717_, _42716_, _42715_);
  nor _49907_ (_42718_, _38485_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or _49908_ (_42719_, _42718_, _42717_);
  or _49909_ (_42720_, _42719_, _42714_);
  and _49910_ (_40016_, _42720_, _42882_);
  or _49911_ (_42721_, _40016_, _42711_);
  and _49912_ (_02563_, _42721_, _42710_);
  not _49913_ (_42722_, _42244_);
  nor _49914_ (_42723_, _42489_, _42722_);
  nor _49915_ (_42724_, _42722_, _42409_);
  and _49916_ (_42725_, _42724_, _42723_);
  and _49917_ (_42726_, _42533_, _42244_);
  nor _49918_ (_42727_, _42722_, _42615_);
  and _49919_ (_42728_, _42727_, _42726_);
  and _49920_ (_42729_, _42728_, _42725_);
  and _49921_ (_42730_, _42720_, _42244_);
  and _49922_ (_42731_, _42730_, _42729_);
  not _49923_ (_42732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor _49924_ (_42733_, _42729_, _42732_);
  or _49925_ (_02573_, _42733_, _42731_);
  nor _49926_ (_42734_, _42727_, _42726_);
  nor _49927_ (_42735_, _42724_, _42723_);
  and _49928_ (_42736_, _42735_, _42244_);
  and _49929_ (_42737_, _42736_, _42734_);
  and _49930_ (_42738_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , _28635_);
  and _49931_ (_42739_, _42738_, _28690_);
  not _49932_ (_42740_, _42739_);
  nor _49933_ (_42741_, _42740_, _31282_);
  not _49934_ (_42742_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _49935_ (_42743_, _38464_, _42742_);
  or _49936_ (_42744_, _18878_, _42742_);
  and _49937_ (_42745_, _42744_, _42740_);
  and _49938_ (_42746_, _42745_, _42743_);
  or _49939_ (_42747_, _42746_, _42741_);
  and _49940_ (_42748_, _42747_, _42737_);
  not _49941_ (_42749_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor _49942_ (_42750_, _42737_, _42749_);
  or _49943_ (_02796_, _42750_, _42748_);
  nand _49944_ (_42751_, _42738_, _28657_);
  nor _49945_ (_42752_, _42751_, _31282_);
  nor _49946_ (_42753_, _38456_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49947_ (_42754_, _42738_, _28744_);
  and _49948_ (_42755_, _42738_, _28723_);
  or _49949_ (_42756_, _42755_, _42712_);
  or _49950_ (_42757_, _42756_, _42754_);
  and _49951_ (_42758_, _42757_, _19871_);
  or _49952_ (_42759_, _42758_, _42753_);
  or _49953_ (_42760_, _42759_, _42752_);
  and _49954_ (_42761_, _42760_, _42737_);
  not _49955_ (_42762_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _49956_ (_42763_, _42737_, _42762_);
  or _49957_ (_02801_, _42763_, _42761_);
  not _49958_ (_42764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _49959_ (_42765_, _42737_, _42764_);
  nand _49960_ (_42766_, _42738_, _28755_);
  nor _49961_ (_42767_, _42766_, _31282_);
  nor _49962_ (_42768_, _38449_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49963_ (_42769_, _42738_, _28646_);
  or _49964_ (_42770_, _42769_, _42756_);
  and _49965_ (_42771_, _42770_, _18516_);
  or _49966_ (_42772_, _42771_, _42768_);
  or _49967_ (_42773_, _42772_, _42767_);
  and _49968_ (_42774_, _42773_, _42737_);
  or _49969_ (_02806_, _42774_, _42765_);
  and _49970_ (_42775_, _42755_, _31859_);
  nor _49971_ (_42776_, _38442_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  or _49972_ (_42777_, _42754_, _42712_);
  or _49973_ (_42778_, _42777_, _42769_);
  and _49974_ (_42779_, _42778_, _19544_);
  or _49975_ (_42780_, _42779_, _42776_);
  or _49976_ (_42781_, _42780_, _42775_);
  and _49977_ (_42782_, _42781_, _42737_);
  not _49978_ (_42783_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _49979_ (_42784_, _42737_, _42783_);
  or _49980_ (_02811_, _42784_, _42782_);
  not _49981_ (_42785_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _49982_ (_42786_, _42737_, _42785_);
  nand _49983_ (_42787_, _42712_, _28690_);
  nor _49984_ (_42788_, _42787_, _31282_);
  nor _49985_ (_42789_, _38434_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _49986_ (_42790_, _28690_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _49987_ (_42791_, _18714_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49988_ (_42792_, _42791_, _42790_);
  or _49989_ (_42793_, _42792_, _42789_);
  or _49990_ (_42794_, _42793_, _42788_);
  and _49991_ (_42795_, _42794_, _42737_);
  or _49992_ (_02815_, _42795_, _42786_);
  nand _49993_ (_42796_, _42712_, _28657_);
  nor _49994_ (_42797_, _42796_, _31282_);
  nor _49995_ (_42798_, _38428_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _49996_ (_42799_, _28657_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _49997_ (_42800_, _19696_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _49998_ (_42801_, _42800_, _42799_);
  or _49999_ (_42802_, _42801_, _42798_);
  or _50000_ (_42803_, _42802_, _42797_);
  and _50001_ (_42804_, _42803_, _42737_);
  not _50002_ (_42805_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _50003_ (_42806_, _42737_, _42805_);
  or _50004_ (_02820_, _42806_, _42804_);
  nand _50005_ (_42807_, _42712_, _28755_);
  nor _50006_ (_42808_, _42807_, _31282_);
  nor _50007_ (_42809_, _38420_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nand _50008_ (_42810_, _28755_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  and _50009_ (_42811_, _19054_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  and _50010_ (_42812_, _42811_, _42810_);
  or _50011_ (_42813_, _42812_, _42809_);
  or _50012_ (_42814_, _42813_, _42808_);
  and _50013_ (_42815_, _42814_, _42737_);
  not _50014_ (_42816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _50015_ (_42817_, _42737_, _42816_);
  or _50016_ (_02825_, _42817_, _42815_);
  not _50017_ (_42818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor _50018_ (_42819_, _42737_, _42818_);
  and _50019_ (_42820_, _42737_, _42720_);
  or _50020_ (_02827_, _42820_, _42819_);
  and _50021_ (_42821_, _42747_, _42244_);
  and _50022_ (_42822_, _42723_, _42409_);
  and _50023_ (_42823_, _42822_, _42734_);
  and _50024_ (_42824_, _42823_, _42821_);
  not _50025_ (_42825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor _50026_ (_42826_, _42823_, _42825_);
  or _50027_ (_02835_, _42826_, _42824_);
  and _50028_ (_42828_, _42760_, _42244_);
  and _50029_ (_42829_, _42823_, _42828_);
  not _50030_ (_42831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor _50031_ (_42833_, _42823_, _42831_);
  or _50032_ (_02838_, _42833_, _42829_);
  and _50033_ (_42835_, _42773_, _42244_);
  and _50034_ (_42837_, _42823_, _42835_);
  not _50035_ (_42839_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor _50036_ (_42841_, _42823_, _42839_);
  or _50037_ (_02841_, _42841_, _42837_);
  and _50038_ (_42842_, _42781_, _42244_);
  and _50039_ (_42843_, _42823_, _42842_);
  not _50040_ (_42844_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor _50041_ (_42845_, _42823_, _42844_);
  or _50042_ (_02845_, _42845_, _42843_);
  and _50043_ (_42846_, _42794_, _42244_);
  and _50044_ (_42847_, _42823_, _42846_);
  not _50045_ (_42848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor _50046_ (_42849_, _42823_, _42848_);
  or _50047_ (_02849_, _42849_, _42847_);
  and _50048_ (_42850_, _42803_, _42244_);
  and _50049_ (_42851_, _42823_, _42850_);
  not _50050_ (_42852_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _50051_ (_42853_, _42823_, _42852_);
  or _50052_ (_02852_, _42853_, _42851_);
  and _50053_ (_42854_, _42814_, _42244_);
  and _50054_ (_42855_, _42823_, _42854_);
  not _50055_ (_42856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor _50056_ (_42857_, _42823_, _42856_);
  or _50057_ (_02855_, _42857_, _42855_);
  and _50058_ (_42858_, _42823_, _42730_);
  nor _50059_ (_42859_, _42823_, _42656_);
  or _50060_ (_02858_, _42859_, _42858_);
  and _50061_ (_42860_, _42724_, _42489_);
  and _50062_ (_42861_, _42860_, _42734_);
  and _50063_ (_42862_, _42861_, _42821_);
  not _50064_ (_42863_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor _50065_ (_42864_, _42861_, _42863_);
  or _50066_ (_02864_, _42864_, _42862_);
  and _50067_ (_42865_, _42861_, _42828_);
  not _50068_ (_42866_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor _50069_ (_42867_, _42861_, _42866_);
  or _50070_ (_02868_, _42867_, _42865_);
  and _50071_ (_42868_, _42861_, _42835_);
  not _50072_ (_42869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor _50073_ (_42871_, _42861_, _42869_);
  or _50074_ (_02871_, _42871_, _42868_);
  and _50075_ (_42874_, _42861_, _42842_);
  not _50076_ (_42876_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor _50077_ (_42878_, _42861_, _42876_);
  or _50078_ (_02875_, _42878_, _42874_);
  and _50079_ (_42881_, _42861_, _42846_);
  not _50080_ (_42883_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor _50081_ (_42884_, _42861_, _42883_);
  or _50082_ (_02878_, _42884_, _42881_);
  and _50083_ (_42887_, _42861_, _42850_);
  not _50084_ (_42888_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor _50085_ (_42889_, _42861_, _42888_);
  or _50086_ (_02882_, _42889_, _42887_);
  and _50087_ (_42890_, _42861_, _42854_);
  not _50088_ (_42891_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor _50089_ (_42892_, _42861_, _42891_);
  or _50090_ (_02885_, _42892_, _42890_);
  and _50091_ (_42893_, _42861_, _42730_);
  not _50092_ (_42894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor _50093_ (_42895_, _42861_, _42894_);
  or _50094_ (_02888_, _42895_, _42893_);
  and _50095_ (_42896_, _42734_, _42725_);
  and _50096_ (_42897_, _42896_, _42821_);
  not _50097_ (_42898_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor _50098_ (_42899_, _42896_, _42898_);
  or _50099_ (_02894_, _42899_, _42897_);
  and _50100_ (_42900_, _42896_, _42828_);
  not _50101_ (_42901_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor _50102_ (_42902_, _42896_, _42901_);
  or _50103_ (_02898_, _42902_, _42900_);
  and _50104_ (_42903_, _42896_, _42835_);
  not _50105_ (_42904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor _50106_ (_42905_, _42896_, _42904_);
  or _50107_ (_02902_, _42905_, _42903_);
  and _50108_ (_42906_, _42896_, _42842_);
  not _50109_ (_42907_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor _50110_ (_42908_, _42896_, _42907_);
  or _50111_ (_02905_, _42908_, _42906_);
  and _50112_ (_42909_, _42896_, _42846_);
  not _50113_ (_42910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor _50114_ (_42911_, _42896_, _42910_);
  or _50115_ (_02909_, _42911_, _42909_);
  and _50116_ (_42912_, _42896_, _42850_);
  not _50117_ (_42913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor _50118_ (_42914_, _42896_, _42913_);
  or _50119_ (_02912_, _42914_, _42912_);
  and _50120_ (_42915_, _42896_, _42854_);
  not _50121_ (_42916_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nor _50122_ (_42917_, _42896_, _42916_);
  or _50123_ (_02916_, _42917_, _42915_);
  and _50124_ (_42918_, _42896_, _42730_);
  nor _50125_ (_42919_, _42896_, _42650_);
  or _50126_ (_02919_, _42919_, _42918_);
  and _50127_ (_42920_, _42727_, _42534_);
  and _50128_ (_42921_, _42920_, _42735_);
  and _50129_ (_42922_, _42921_, _42821_);
  not _50130_ (_42923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor _50131_ (_42924_, _42921_, _42923_);
  or _50132_ (_02926_, _42924_, _42922_);
  and _50133_ (_42925_, _42921_, _42828_);
  not _50134_ (_42926_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _50135_ (_42927_, _42921_, _42926_);
  or _50136_ (_02929_, _42927_, _42925_);
  and _50137_ (_42928_, _42921_, _42835_);
  not _50138_ (_42929_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor _50139_ (_42930_, _42921_, _42929_);
  or _50140_ (_02933_, _42930_, _42928_);
  and _50141_ (_42931_, _42921_, _42842_);
  not _50142_ (_42932_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor _50143_ (_42933_, _42921_, _42932_);
  or _50144_ (_02937_, _42933_, _42931_);
  and _50145_ (_42934_, _42921_, _42846_);
  not _50146_ (_42935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor _50147_ (_42936_, _42921_, _42935_);
  or _50148_ (_02940_, _42936_, _42934_);
  and _50149_ (_42937_, _42921_, _42850_);
  not _50150_ (_42938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor _50151_ (_42939_, _42921_, _42938_);
  or _50152_ (_02943_, _42939_, _42937_);
  and _50153_ (_42940_, _42921_, _42854_);
  not _50154_ (_42941_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _50155_ (_42942_, _42921_, _42941_);
  or _50156_ (_02947_, _42942_, _42940_);
  and _50157_ (_42943_, _42921_, _42730_);
  not _50158_ (_42944_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor _50159_ (_42945_, _42921_, _42944_);
  or _50160_ (_02950_, _42945_, _42943_);
  and _50161_ (_42946_, _42920_, _42822_);
  and _50162_ (_42947_, _42946_, _42821_);
  not _50163_ (_42948_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor _50164_ (_42949_, _42946_, _42948_);
  or _50165_ (_02954_, _42949_, _42947_);
  and _50166_ (_42950_, _42946_, _42828_);
  not _50167_ (_42951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor _50168_ (_42952_, _42946_, _42951_);
  or _50169_ (_02957_, _42952_, _42950_);
  and _50170_ (_42953_, _42946_, _42835_);
  not _50171_ (_42954_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor _50172_ (_42955_, _42946_, _42954_);
  or _50173_ (_02962_, _42955_, _42953_);
  and _50174_ (_42956_, _42946_, _42842_);
  not _50175_ (_42957_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor _50176_ (_42958_, _42946_, _42957_);
  or _50177_ (_02965_, _42958_, _42956_);
  and _50178_ (_42959_, _42946_, _42846_);
  not _50179_ (_42960_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nor _50180_ (_42961_, _42946_, _42960_);
  or _50181_ (_02968_, _42961_, _42959_);
  and _50182_ (_42962_, _42946_, _42850_);
  not _50183_ (_42963_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor _50184_ (_42964_, _42946_, _42963_);
  or _50185_ (_02972_, _42964_, _42962_);
  and _50186_ (_42965_, _42946_, _42854_);
  not _50187_ (_42966_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor _50188_ (_42967_, _42946_, _42966_);
  or _50189_ (_02976_, _42967_, _42965_);
  and _50190_ (_42968_, _42946_, _42730_);
  nor _50191_ (_42969_, _42946_, _42669_);
  or _50192_ (_02978_, _42969_, _42968_);
  and _50193_ (_42970_, _42920_, _42860_);
  and _50194_ (_42971_, _42970_, _42821_);
  not _50195_ (_42972_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor _50196_ (_42973_, _42970_, _42972_);
  or _50197_ (_02983_, _42973_, _42971_);
  and _50198_ (_42974_, _42970_, _42828_);
  not _50199_ (_42975_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor _50200_ (_42976_, _42970_, _42975_);
  or _50201_ (_02987_, _42976_, _42974_);
  and _50202_ (_42977_, _42970_, _42835_);
  not _50203_ (_42978_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor _50204_ (_42979_, _42970_, _42978_);
  or _50205_ (_02991_, _42979_, _42977_);
  and _50206_ (_42980_, _42970_, _42842_);
  not _50207_ (_42981_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor _50208_ (_42982_, _42970_, _42981_);
  or _50209_ (_02994_, _42982_, _42980_);
  and _50210_ (_42983_, _42970_, _42846_);
  not _50211_ (_42984_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor _50212_ (_42985_, _42970_, _42984_);
  or _50213_ (_02999_, _42985_, _42983_);
  and _50214_ (_42986_, _42970_, _42850_);
  not _50215_ (_42987_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor _50216_ (_42988_, _42970_, _42987_);
  or _50217_ (_03002_, _42988_, _42986_);
  and _50218_ (_42989_, _42970_, _42854_);
  not _50219_ (_42990_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor _50220_ (_42991_, _42970_, _42990_);
  or _50221_ (_03006_, _42991_, _42989_);
  and _50222_ (_42992_, _42970_, _42730_);
  not _50223_ (_42993_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor _50224_ (_42994_, _42970_, _42993_);
  or _50225_ (_03009_, _42994_, _42992_);
  and _50226_ (_42995_, _42920_, _42725_);
  and _50227_ (_42996_, _42995_, _42821_);
  not _50228_ (_42997_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor _50229_ (_42998_, _42995_, _42997_);
  or _50230_ (_03014_, _42998_, _42996_);
  and _50231_ (_42999_, _42995_, _42828_);
  not _50232_ (_43000_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor _50233_ (_43001_, _42995_, _43000_);
  or _50234_ (_03018_, _43001_, _42999_);
  and _50235_ (_43002_, _42995_, _42835_);
  not _50236_ (_43003_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor _50237_ (_43004_, _42995_, _43003_);
  or _50238_ (_03021_, _43004_, _43002_);
  and _50239_ (_43005_, _42995_, _42842_);
  not _50240_ (_43006_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor _50241_ (_43007_, _42995_, _43006_);
  or _50242_ (_03025_, _43007_, _43005_);
  and _50243_ (_43008_, _42995_, _42846_);
  not _50244_ (_43009_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor _50245_ (_43010_, _42995_, _43009_);
  or _50246_ (_03028_, _43010_, _43008_);
  and _50247_ (_43011_, _42995_, _42850_);
  not _50248_ (_43012_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nor _50249_ (_43013_, _42995_, _43012_);
  or _50250_ (_03032_, _43013_, _43011_);
  and _50251_ (_43014_, _42995_, _42854_);
  not _50252_ (_43015_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor _50253_ (_43016_, _42995_, _43015_);
  or _50254_ (_03036_, _43016_, _43014_);
  and _50255_ (_43017_, _42995_, _42730_);
  nor _50256_ (_43018_, _42995_, _42663_);
  or _50257_ (_03038_, _43018_, _43017_);
  and _50258_ (_43019_, _42726_, _42615_);
  and _50259_ (_43020_, _43019_, _42735_);
  and _50260_ (_43021_, _43020_, _42821_);
  not _50261_ (_43022_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor _50262_ (_43023_, _43020_, _43022_);
  or _50263_ (_03045_, _43023_, _43021_);
  and _50264_ (_43024_, _43020_, _42828_);
  not _50265_ (_43025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor _50266_ (_43026_, _43020_, _43025_);
  or _50267_ (_03048_, _43026_, _43024_);
  and _50268_ (_43027_, _43020_, _42835_);
  not _50269_ (_43028_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor _50270_ (_43029_, _43020_, _43028_);
  or _50271_ (_03051_, _43029_, _43027_);
  and _50272_ (_43030_, _43020_, _42842_);
  not _50273_ (_43031_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor _50274_ (_43032_, _43020_, _43031_);
  or _50275_ (_03054_, _43032_, _43030_);
  and _50276_ (_43033_, _43020_, _42846_);
  not _50277_ (_43034_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor _50278_ (_43035_, _43020_, _43034_);
  or _50279_ (_03058_, _43035_, _43033_);
  and _50280_ (_43036_, _43020_, _42850_);
  not _50281_ (_43037_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor _50282_ (_43038_, _43020_, _43037_);
  or _50283_ (_03061_, _43038_, _43036_);
  and _50284_ (_43039_, _43020_, _42854_);
  not _50285_ (_43040_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor _50286_ (_43041_, _43020_, _43040_);
  or _50287_ (_03064_, _43041_, _43039_);
  and _50288_ (_43042_, _43020_, _42730_);
  nor _50289_ (_43043_, _43020_, _42678_);
  or _50290_ (_03067_, _43043_, _43042_);
  and _50291_ (_43044_, _43019_, _42822_);
  and _50292_ (_43045_, _43044_, _42821_);
  not _50293_ (_43046_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor _50294_ (_43047_, _43044_, _43046_);
  or _50295_ (_03071_, _43047_, _43045_);
  and _50296_ (_43048_, _43044_, _42828_);
  not _50297_ (_43049_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor _50298_ (_43050_, _43044_, _43049_);
  or _50299_ (_03074_, _43050_, _43048_);
  and _50300_ (_43051_, _43044_, _42835_);
  not _50301_ (_43052_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor _50302_ (_43053_, _43044_, _43052_);
  or _50303_ (_03078_, _43053_, _43051_);
  and _50304_ (_43054_, _43044_, _42842_);
  not _50305_ (_43055_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor _50306_ (_43056_, _43044_, _43055_);
  or _50307_ (_03081_, _43056_, _43054_);
  and _50308_ (_43057_, _43044_, _42846_);
  not _50309_ (_43058_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor _50310_ (_43059_, _43044_, _43058_);
  or _50311_ (_03085_, _43059_, _43057_);
  and _50312_ (_43060_, _43044_, _42850_);
  not _50313_ (_43061_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor _50314_ (_43062_, _43044_, _43061_);
  or _50315_ (_03089_, _43062_, _43060_);
  and _50316_ (_43063_, _43044_, _42854_);
  not _50317_ (_43064_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor _50318_ (_43065_, _43044_, _43064_);
  or _50319_ (_03093_, _43065_, _43063_);
  and _50320_ (_43066_, _43044_, _42730_);
  not _50321_ (_43067_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor _50322_ (_43068_, _43044_, _43067_);
  or _50323_ (_03096_, _43068_, _43066_);
  and _50324_ (_43069_, _43019_, _42860_);
  and _50325_ (_43070_, _43069_, _42821_);
  not _50326_ (_43071_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor _50327_ (_43072_, _43069_, _43071_);
  or _50328_ (_03101_, _43072_, _43070_);
  and _50329_ (_43073_, _43069_, _42828_);
  not _50330_ (_43074_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor _50331_ (_43075_, _43069_, _43074_);
  or _50332_ (_03105_, _43075_, _43073_);
  and _50333_ (_43076_, _43069_, _42835_);
  not _50334_ (_43077_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor _50335_ (_43078_, _43069_, _43077_);
  or _50336_ (_03109_, _43078_, _43076_);
  and _50337_ (_43079_, _43069_, _42842_);
  not _50338_ (_43080_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor _50339_ (_43081_, _43069_, _43080_);
  or _50340_ (_03113_, _43081_, _43079_);
  and _50341_ (_43082_, _43069_, _42846_);
  not _50342_ (_43083_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor _50343_ (_43084_, _43069_, _43083_);
  or _50344_ (_03118_, _43084_, _43082_);
  and _50345_ (_43085_, _43069_, _42850_);
  not _50346_ (_43086_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor _50347_ (_43087_, _43069_, _43086_);
  or _50348_ (_03122_, _43087_, _43085_);
  and _50349_ (_43088_, _43069_, _42854_);
  not _50350_ (_43089_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor _50351_ (_43090_, _43069_, _43089_);
  or _50352_ (_03126_, _43090_, _43088_);
  and _50353_ (_43091_, _43069_, _42730_);
  nor _50354_ (_43092_, _43069_, _42684_);
  or _50355_ (_03129_, _43092_, _43091_);
  and _50356_ (_43093_, _43019_, _42725_);
  and _50357_ (_43094_, _43093_, _42821_);
  not _50358_ (_43095_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor _50359_ (_43096_, _43093_, _43095_);
  or _50360_ (_03134_, _43096_, _43094_);
  and _50361_ (_43097_, _43093_, _42828_);
  not _50362_ (_43098_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor _50363_ (_43099_, _43093_, _43098_);
  or _50364_ (_03138_, _43099_, _43097_);
  and _50365_ (_43100_, _43093_, _42835_);
  not _50366_ (_43101_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor _50367_ (_43102_, _43093_, _43101_);
  or _50368_ (_03142_, _43102_, _43100_);
  and _50369_ (_43103_, _43093_, _42842_);
  not _50370_ (_43104_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor _50371_ (_43105_, _43093_, _43104_);
  or _50372_ (_03146_, _43105_, _43103_);
  and _50373_ (_43106_, _43093_, _42846_);
  not _50374_ (_43107_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor _50375_ (_43108_, _43093_, _43107_);
  or _50376_ (_03150_, _43108_, _43106_);
  and _50377_ (_43109_, _43093_, _42850_);
  not _50378_ (_43110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor _50379_ (_43111_, _43093_, _43110_);
  or _50380_ (_03154_, _43111_, _43109_);
  and _50381_ (_43112_, _43093_, _42854_);
  not _50382_ (_43113_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor _50383_ (_43114_, _43093_, _43113_);
  or _50384_ (_03158_, _43114_, _43112_);
  and _50385_ (_43115_, _43093_, _42730_);
  not _50386_ (_43116_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor _50387_ (_43117_, _43093_, _43116_);
  or _50388_ (_03161_, _43117_, _43115_);
  and _50389_ (_43118_, _42735_, _42728_);
  and _50390_ (_43119_, _43118_, _42821_);
  not _50391_ (_43120_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor _50392_ (_43121_, _43118_, _43120_);
  or _50393_ (_03167_, _43121_, _43119_);
  and _50394_ (_43122_, _43118_, _42828_);
  not _50395_ (_43123_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor _50396_ (_43124_, _43118_, _43123_);
  or _50397_ (_03171_, _43124_, _43122_);
  and _50398_ (_43125_, _43118_, _42835_);
  not _50399_ (_43126_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nor _50400_ (_43127_, _43118_, _43126_);
  or _50401_ (_03175_, _43127_, _43125_);
  and _50402_ (_43128_, _43118_, _42842_);
  not _50403_ (_43129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor _50404_ (_43130_, _43118_, _43129_);
  or _50405_ (_03179_, _43130_, _43128_);
  and _50406_ (_43131_, _43118_, _42846_);
  not _50407_ (_43132_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor _50408_ (_43133_, _43118_, _43132_);
  or _50409_ (_03183_, _43133_, _43131_);
  and _50410_ (_43134_, _43118_, _42850_);
  not _50411_ (_43135_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor _50412_ (_43136_, _43118_, _43135_);
  or _50413_ (_03187_, _43136_, _43134_);
  and _50414_ (_43137_, _43118_, _42854_);
  not _50415_ (_43138_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor _50416_ (_43139_, _43118_, _43138_);
  or _50417_ (_03191_, _43139_, _43137_);
  and _50418_ (_43140_, _43118_, _42730_);
  nor _50419_ (_43141_, _43118_, _42690_);
  or _50420_ (_03194_, _43141_, _43140_);
  and _50421_ (_43142_, _42822_, _42728_);
  and _50422_ (_43143_, _43142_, _42821_);
  not _50423_ (_43144_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor _50424_ (_43145_, _43142_, _43144_);
  or _50425_ (_03199_, _43145_, _43143_);
  and _50426_ (_43146_, _43142_, _42828_);
  not _50427_ (_43147_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor _50428_ (_43148_, _43142_, _43147_);
  or _50429_ (_03203_, _43148_, _43146_);
  and _50430_ (_43149_, _43142_, _42835_);
  not _50431_ (_43150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor _50432_ (_43151_, _43142_, _43150_);
  or _50433_ (_03207_, _43151_, _43149_);
  and _50434_ (_43152_, _43142_, _42842_);
  not _50435_ (_43153_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor _50436_ (_43154_, _43142_, _43153_);
  or _50437_ (_03211_, _43154_, _43152_);
  and _50438_ (_43155_, _43142_, _42846_);
  not _50439_ (_43156_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor _50440_ (_43157_, _43142_, _43156_);
  or _50441_ (_03215_, _43157_, _43155_);
  and _50442_ (_43158_, _43142_, _42850_);
  not _50443_ (_43159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor _50444_ (_43160_, _43142_, _43159_);
  or _50445_ (_03219_, _43160_, _43158_);
  and _50446_ (_43161_, _43142_, _42854_);
  not _50447_ (_43162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor _50448_ (_43163_, _43142_, _43162_);
  or _50449_ (_03223_, _43163_, _43161_);
  and _50450_ (_43164_, _43142_, _42730_);
  not _50451_ (_43165_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor _50452_ (_43166_, _43142_, _43165_);
  or _50453_ (_03226_, _43166_, _43164_);
  and _50454_ (_43167_, _42860_, _42728_);
  and _50455_ (_43168_, _43167_, _42821_);
  not _50456_ (_43169_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor _50457_ (_43170_, _43167_, _43169_);
  or _50458_ (_03231_, _43170_, _43168_);
  and _50459_ (_43171_, _43167_, _42828_);
  not _50460_ (_43172_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor _50461_ (_43173_, _43167_, _43172_);
  or _50462_ (_03235_, _43173_, _43171_);
  and _50463_ (_43174_, _43167_, _42835_);
  not _50464_ (_43175_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor _50465_ (_43176_, _43167_, _43175_);
  or _50466_ (_03239_, _43176_, _43174_);
  and _50467_ (_43177_, _43167_, _42842_);
  not _50468_ (_43178_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor _50469_ (_43179_, _43167_, _43178_);
  or _50470_ (_03243_, _43179_, _43177_);
  and _50471_ (_43180_, _43167_, _42846_);
  not _50472_ (_43181_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor _50473_ (_43182_, _43167_, _43181_);
  or _50474_ (_03247_, _43182_, _43180_);
  and _50475_ (_43183_, _43167_, _42850_);
  not _50476_ (_43184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor _50477_ (_43185_, _43167_, _43184_);
  or _50478_ (_03251_, _43185_, _43183_);
  and _50479_ (_43186_, _43167_, _42854_);
  not _50480_ (_43187_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor _50481_ (_43188_, _43167_, _43187_);
  or _50482_ (_03255_, _43188_, _43186_);
  and _50483_ (_43189_, _43167_, _42730_);
  nor _50484_ (_43190_, _43167_, _42696_);
  or _50485_ (_03258_, _43190_, _43189_);
  and _50486_ (_43191_, _42821_, _42729_);
  not _50487_ (_43192_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor _50488_ (_43193_, _42729_, _43192_);
  or _50489_ (_03263_, _43193_, _43191_);
  and _50490_ (_43194_, _42828_, _42729_);
  not _50491_ (_43195_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor _50492_ (_43196_, _42729_, _43195_);
  or _50493_ (_03267_, _43196_, _43194_);
  and _50494_ (_43197_, _42835_, _42729_);
  not _50495_ (_43198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor _50496_ (_43199_, _42729_, _43198_);
  or _50497_ (_03271_, _43199_, _43197_);
  and _50498_ (_43200_, _42842_, _42729_);
  not _50499_ (_43201_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor _50500_ (_43202_, _42729_, _43201_);
  or _50501_ (_03275_, _43202_, _43200_);
  and _50502_ (_43203_, _42846_, _42729_);
  not _50503_ (_43204_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor _50504_ (_43205_, _42729_, _43204_);
  or _50505_ (_03279_, _43205_, _43203_);
  and _50506_ (_43206_, _42850_, _42729_);
  not _50507_ (_43207_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor _50508_ (_43208_, _42729_, _43207_);
  or _50509_ (_03283_, _43208_, _43206_);
  and _50510_ (_43209_, _42854_, _42729_);
  not _50511_ (_43210_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor _50512_ (_43211_, _42729_, _43210_);
  or _50513_ (_03287_, _43211_, _43209_);
  nor _50514_ (_43212_, _42486_, _42898_);
  and _50515_ (_43213_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  or _50516_ (_43214_, _43213_, _42404_);
  or _50517_ (_43215_, _43214_, _43212_);
  and _50518_ (_43216_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  or _50519_ (_43217_, _42486_, _42825_);
  nand _50520_ (_43218_, _43217_, _42404_);
  or _50521_ (_43219_, _43218_, _43216_);
  and _50522_ (_43220_, _43219_, _43215_);
  or _50523_ (_43221_, _43220_, _42649_);
  nor _50524_ (_43222_, _42486_, _42997_);
  and _50525_ (_43223_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  or _50526_ (_43224_, _43223_, _42404_);
  or _50527_ (_43225_, _43224_, _43222_);
  and _50528_ (_43226_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  or _50529_ (_43227_, _42486_, _42948_);
  nand _50530_ (_43228_, _43227_, _42404_);
  or _50531_ (_43229_, _43228_, _43226_);
  and _50532_ (_43230_, _43229_, _43225_);
  or _50533_ (_43231_, _43230_, _42612_);
  and _50534_ (_43232_, _43231_, _42662_);
  and _50535_ (_43233_, _43232_, _43221_);
  nand _50536_ (_43234_, _42486_, _43022_);
  or _50537_ (_43235_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  and _50538_ (_43236_, _43235_, _43234_);
  or _50539_ (_43237_, _43236_, _42677_);
  or _50540_ (_43238_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nand _50541_ (_43239_, _42486_, _43071_);
  and _50542_ (_43240_, _43239_, _43238_);
  or _50543_ (_43241_, _43240_, _42404_);
  and _50544_ (_43242_, _43241_, _43237_);
  or _50545_ (_43243_, _43242_, _42649_);
  nand _50546_ (_43244_, _42486_, _43120_);
  or _50547_ (_43245_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _50548_ (_43246_, _43245_, _43244_);
  or _50549_ (_43247_, _43246_, _42677_);
  or _50550_ (_43248_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nand _50551_ (_43249_, _42486_, _43169_);
  and _50552_ (_43250_, _43249_, _43248_);
  or _50553_ (_43251_, _43250_, _42404_);
  and _50554_ (_43252_, _43251_, _43247_);
  or _50555_ (_43253_, _43252_, _42612_);
  and _50556_ (_43254_, _43253_, _42530_);
  and _50557_ (_43255_, _43254_, _43243_);
  or _50558_ (_43256_, _43255_, _43233_);
  or _50559_ (_43257_, _43256_, _42648_);
  not _50560_ (_43258_, _42648_);
  or _50561_ (_43259_, _43258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  and _50562_ (_43260_, _43259_, _42711_);
  and _50563_ (_43261_, _43260_, _43257_);
  and _50564_ (_40036_, _42747_, _42882_);
  and _50565_ (_43262_, _40036_, _42707_);
  or _50566_ (_05081_, _43262_, _43261_);
  nor _50567_ (_43263_, _42486_, _42901_);
  and _50568_ (_43264_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  or _50569_ (_43265_, _43264_, _42404_);
  or _50570_ (_43266_, _43265_, _43263_);
  and _50571_ (_43267_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  or _50572_ (_43268_, _42486_, _42831_);
  nand _50573_ (_43269_, _43268_, _42404_);
  or _50574_ (_43270_, _43269_, _43267_);
  and _50575_ (_43271_, _43270_, _43266_);
  or _50576_ (_43272_, _43271_, _42649_);
  nor _50577_ (_43273_, _42486_, _43000_);
  and _50578_ (_43274_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  or _50579_ (_43275_, _43274_, _42404_);
  or _50580_ (_43276_, _43275_, _43273_);
  and _50581_ (_43277_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  or _50582_ (_43278_, _42486_, _42951_);
  nand _50583_ (_43279_, _43278_, _42404_);
  or _50584_ (_43280_, _43279_, _43277_);
  and _50585_ (_43281_, _43280_, _43276_);
  or _50586_ (_43282_, _43281_, _42612_);
  and _50587_ (_43283_, _43282_, _42662_);
  and _50588_ (_43284_, _43283_, _43272_);
  nand _50589_ (_43285_, _42486_, _43025_);
  or _50590_ (_43286_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _50591_ (_43287_, _43286_, _43285_);
  or _50592_ (_43288_, _43287_, _42677_);
  or _50593_ (_43289_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nand _50594_ (_43290_, _42486_, _43074_);
  and _50595_ (_43291_, _43290_, _43289_);
  or _50596_ (_43292_, _43291_, _42404_);
  and _50597_ (_43293_, _43292_, _43288_);
  or _50598_ (_43294_, _43293_, _42649_);
  nand _50599_ (_43295_, _42486_, _43123_);
  or _50600_ (_43296_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _50601_ (_43297_, _43296_, _43295_);
  or _50602_ (_43298_, _43297_, _42677_);
  or _50603_ (_43299_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nand _50604_ (_43300_, _42486_, _43172_);
  and _50605_ (_43301_, _43300_, _43299_);
  or _50606_ (_43302_, _43301_, _42404_);
  and _50607_ (_43303_, _43302_, _43298_);
  or _50608_ (_43304_, _43303_, _42612_);
  and _50609_ (_43305_, _43304_, _42530_);
  and _50610_ (_43306_, _43305_, _43294_);
  nor _50611_ (_43307_, _43306_, _43284_);
  nor _50612_ (_43308_, _43307_, _42648_);
  and _50613_ (_43309_, _42648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  or _50614_ (_43310_, _43309_, _42707_);
  or _50615_ (_43311_, _43310_, _43308_);
  and _50616_ (_40037_, _42760_, _42882_);
  or _50617_ (_43312_, _40037_, _42711_);
  and _50618_ (_05083_, _43312_, _43311_);
  or _50619_ (_43313_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nand _50620_ (_43314_, _42486_, _43175_);
  and _50621_ (_43315_, _43314_, _43313_);
  or _50622_ (_43316_, _43315_, _42404_);
  nand _50623_ (_43317_, _42486_, _43126_);
  or _50624_ (_43318_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and _50625_ (_43319_, _43318_, _43317_);
  or _50626_ (_43320_, _43319_, _42677_);
  and _50627_ (_43321_, _43320_, _42530_);
  and _50628_ (_43322_, _43321_, _43316_);
  and _50629_ (_43323_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor _50630_ (_43331_, _42486_, _42954_);
  or _50631_ (_43337_, _43331_, _42677_);
  or _50632_ (_43341_, _43337_, _43323_);
  nor _50633_ (_43348_, _42486_, _43003_);
  and _50634_ (_43356_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  or _50635_ (_43360_, _43356_, _42404_);
  or _50636_ (_43365_, _43360_, _43348_);
  and _50637_ (_43373_, _43365_, _42662_);
  and _50638_ (_43379_, _43373_, _43341_);
  or _50639_ (_43383_, _43379_, _43322_);
  and _50640_ (_43390_, _43383_, _42649_);
  or _50641_ (_43398_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nand _50642_ (_43402_, _42486_, _43077_);
  and _50643_ (_43407_, _43402_, _43398_);
  or _50644_ (_43415_, _43407_, _42404_);
  nand _50645_ (_43416_, _42486_, _43028_);
  or _50646_ (_43424_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _50647_ (_43433_, _43424_, _43416_);
  or _50648_ (_43439_, _43433_, _42677_);
  and _50649_ (_43443_, _43439_, _42530_);
  and _50650_ (_43450_, _43443_, _43415_);
  and _50651_ (_43458_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _50652_ (_43462_, _42486_, _42839_);
  or _50653_ (_43467_, _43462_, _42677_);
  or _50654_ (_43475_, _43467_, _43458_);
  nor _50655_ (_43481_, _42486_, _42904_);
  and _50656_ (_43485_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  or _50657_ (_43492_, _43485_, _42404_);
  or _50658_ (_43500_, _43492_, _43481_);
  and _50659_ (_43504_, _43500_, _42662_);
  and _50660_ (_43509_, _43504_, _43475_);
  or _50661_ (_43517_, _43509_, _43450_);
  and _50662_ (_43518_, _43517_, _42612_);
  or _50663_ (_43519_, _43518_, _42622_);
  or _50664_ (_43520_, _43519_, _43390_);
  or _50665_ (_43521_, _43258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  and _50666_ (_40039_, _42773_, _42882_);
  or _50667_ (_43522_, _40039_, _42711_);
  and _50668_ (_43523_, _43522_, _43521_);
  and _50669_ (_05084_, _43523_, _43520_);
  nor _50670_ (_43524_, _42486_, _42907_);
  and _50671_ (_43525_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  or _50672_ (_43526_, _43525_, _42404_);
  or _50673_ (_43527_, _43526_, _43524_);
  and _50674_ (_43528_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  or _50675_ (_43529_, _42486_, _42844_);
  nand _50676_ (_43530_, _43529_, _42404_);
  or _50677_ (_43531_, _43530_, _43528_);
  and _50678_ (_43532_, _43531_, _43527_);
  or _50679_ (_43533_, _43532_, _42649_);
  nor _50680_ (_43534_, _42486_, _43006_);
  and _50681_ (_43535_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  or _50682_ (_43536_, _43535_, _42404_);
  or _50683_ (_43537_, _43536_, _43534_);
  and _50684_ (_43538_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  or _50685_ (_43539_, _42486_, _42957_);
  nand _50686_ (_43540_, _43539_, _42404_);
  or _50687_ (_43541_, _43540_, _43538_);
  and _50688_ (_43542_, _43541_, _43537_);
  or _50689_ (_43543_, _43542_, _42612_);
  and _50690_ (_43544_, _43543_, _42662_);
  and _50691_ (_43545_, _43544_, _43533_);
  nand _50692_ (_43546_, _42486_, _43031_);
  or _50693_ (_43547_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  and _50694_ (_43548_, _43547_, _43546_);
  or _50695_ (_43549_, _43548_, _42677_);
  or _50696_ (_43550_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nand _50697_ (_43551_, _42486_, _43080_);
  and _50698_ (_43552_, _43551_, _43550_);
  or _50699_ (_43553_, _43552_, _42404_);
  and _50700_ (_43554_, _43553_, _43549_);
  or _50701_ (_43555_, _43554_, _42649_);
  nand _50702_ (_43556_, _42486_, _43129_);
  or _50703_ (_43557_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  and _50704_ (_43558_, _43557_, _43556_);
  or _50705_ (_43559_, _43558_, _42677_);
  or _50706_ (_43560_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nand _50707_ (_43561_, _42486_, _43178_);
  and _50708_ (_43562_, _43561_, _43560_);
  or _50709_ (_43563_, _43562_, _42404_);
  and _50710_ (_43564_, _43563_, _43559_);
  or _50711_ (_43565_, _43564_, _42612_);
  and _50712_ (_43566_, _43565_, _42530_);
  and _50713_ (_43567_, _43566_, _43555_);
  nor _50714_ (_43568_, _43567_, _43545_);
  nor _50715_ (_43569_, _43568_, _42648_);
  and _50716_ (_43570_, _42648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  or _50717_ (_43571_, _43570_, _42707_);
  or _50718_ (_43572_, _43571_, _43569_);
  and _50719_ (_40040_, _42781_, _42882_);
  or _50720_ (_43573_, _40040_, _42711_);
  and _50721_ (_05086_, _43573_, _43572_);
  and _50722_ (_43574_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  or _50723_ (_43575_, _42486_, _42848_);
  nand _50724_ (_43576_, _43575_, _42404_);
  or _50725_ (_43577_, _43576_, _43574_);
  nor _50726_ (_43578_, _42486_, _42910_);
  and _50727_ (_43579_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  or _50728_ (_43580_, _43579_, _42404_);
  or _50729_ (_43581_, _43580_, _43578_);
  and _50730_ (_43582_, _43581_, _43577_);
  or _50731_ (_43583_, _43582_, _42649_);
  nor _50732_ (_43584_, _42486_, _43009_);
  and _50733_ (_43585_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  or _50734_ (_43586_, _43585_, _42404_);
  or _50735_ (_43587_, _43586_, _43584_);
  and _50736_ (_43588_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  or _50737_ (_43589_, _42486_, _42960_);
  nand _50738_ (_43590_, _43589_, _42404_);
  or _50739_ (_43591_, _43590_, _43588_);
  and _50740_ (_43592_, _43591_, _43587_);
  or _50741_ (_43593_, _43592_, _42612_);
  and _50742_ (_43594_, _43593_, _42662_);
  and _50743_ (_43595_, _43594_, _43583_);
  nor _50744_ (_43596_, _42486_, _43107_);
  and _50745_ (_43597_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  or _50746_ (_43598_, _43597_, _42404_);
  or _50747_ (_43599_, _43598_, _43596_);
  and _50748_ (_43600_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  or _50749_ (_43601_, _42486_, _43058_);
  nand _50750_ (_43602_, _43601_, _42404_);
  or _50751_ (_43603_, _43602_, _43600_);
  and _50752_ (_43604_, _43603_, _43599_);
  or _50753_ (_43605_, _43604_, _42649_);
  nor _50754_ (_43606_, _42486_, _43204_);
  and _50755_ (_43607_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  or _50756_ (_43608_, _43607_, _42404_);
  or _50757_ (_43609_, _43608_, _43606_);
  and _50758_ (_43610_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  or _50759_ (_43611_, _42486_, _43156_);
  nand _50760_ (_43612_, _43611_, _42404_);
  or _50761_ (_43613_, _43612_, _43610_);
  and _50762_ (_43614_, _43613_, _43609_);
  or _50763_ (_43615_, _43614_, _42612_);
  and _50764_ (_43616_, _43615_, _42530_);
  and _50765_ (_43617_, _43616_, _43605_);
  or _50766_ (_43618_, _43617_, _43595_);
  and _50767_ (_43619_, _43618_, _42706_);
  and _50768_ (_43620_, _42794_, _42707_);
  and _50769_ (_43621_, _42648_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  or _50770_ (_43622_, _43621_, _43620_);
  or _50771_ (_43623_, _43622_, _43619_);
  and _50772_ (_05088_, _43623_, _42882_);
  nor _50773_ (_43624_, _42486_, _42913_);
  and _50774_ (_43625_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  or _50775_ (_43626_, _43625_, _42404_);
  or _50776_ (_43627_, _43626_, _43624_);
  and _50777_ (_43628_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  or _50778_ (_43629_, _42486_, _42852_);
  nand _50779_ (_43630_, _43629_, _42404_);
  or _50780_ (_43631_, _43630_, _43628_);
  and _50781_ (_43632_, _43631_, _43627_);
  or _50782_ (_43633_, _43632_, _42649_);
  nor _50783_ (_43634_, _42486_, _43012_);
  and _50784_ (_43635_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  or _50785_ (_43636_, _43635_, _42404_);
  or _50786_ (_43637_, _43636_, _43634_);
  and _50787_ (_43638_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  or _50788_ (_43639_, _42486_, _42963_);
  nand _50789_ (_43640_, _43639_, _42404_);
  or _50790_ (_43641_, _43640_, _43638_);
  and _50791_ (_43642_, _43641_, _43637_);
  or _50792_ (_43643_, _43642_, _42612_);
  and _50793_ (_43644_, _43643_, _42662_);
  and _50794_ (_43645_, _43644_, _43633_);
  nand _50795_ (_43646_, _42486_, _43037_);
  or _50796_ (_43647_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  and _50797_ (_43648_, _43647_, _43646_);
  or _50798_ (_43649_, _43648_, _42677_);
  or _50799_ (_43650_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nand _50800_ (_43651_, _42486_, _43086_);
  and _50801_ (_43652_, _43651_, _43650_);
  or _50802_ (_43653_, _43652_, _42404_);
  and _50803_ (_43654_, _43653_, _43649_);
  or _50804_ (_43655_, _43654_, _42649_);
  nand _50805_ (_43656_, _42486_, _43135_);
  or _50806_ (_43657_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and _50807_ (_43658_, _43657_, _43656_);
  or _50808_ (_43659_, _43658_, _42677_);
  or _50809_ (_43660_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nand _50810_ (_43661_, _42486_, _43184_);
  and _50811_ (_43662_, _43661_, _43660_);
  or _50812_ (_43663_, _43662_, _42404_);
  and _50813_ (_43664_, _43663_, _43659_);
  or _50814_ (_43665_, _43664_, _42612_);
  and _50815_ (_43666_, _43665_, _42530_);
  and _50816_ (_43667_, _43666_, _43655_);
  or _50817_ (_43668_, _43667_, _43645_);
  or _50818_ (_43669_, _43668_, _42648_);
  or _50819_ (_43670_, _43258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  and _50820_ (_43671_, _43670_, _42711_);
  and _50821_ (_43672_, _43671_, _43669_);
  and _50822_ (_40042_, _42803_, _42882_);
  and _50823_ (_43673_, _40042_, _42707_);
  or _50824_ (_05090_, _43673_, _43672_);
  nor _50825_ (_43674_, _42486_, _42916_);
  and _50826_ (_43675_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  or _50827_ (_43676_, _43675_, _42404_);
  or _50828_ (_43677_, _43676_, _43674_);
  and _50829_ (_43678_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  or _50830_ (_43679_, _42486_, _42856_);
  nand _50831_ (_43680_, _43679_, _42404_);
  or _50832_ (_43681_, _43680_, _43678_);
  and _50833_ (_43682_, _43681_, _43677_);
  or _50834_ (_43683_, _43682_, _42649_);
  nor _50835_ (_43684_, _42486_, _43015_);
  and _50836_ (_43685_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  or _50837_ (_43686_, _43685_, _42404_);
  or _50838_ (_43687_, _43686_, _43684_);
  and _50839_ (_43688_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  or _50840_ (_43689_, _42486_, _42966_);
  nand _50841_ (_43690_, _43689_, _42404_);
  or _50842_ (_43691_, _43690_, _43688_);
  and _50843_ (_43692_, _43691_, _43687_);
  or _50844_ (_43693_, _43692_, _42612_);
  and _50845_ (_43694_, _43693_, _42662_);
  and _50846_ (_43695_, _43694_, _43683_);
  nand _50847_ (_43696_, _42486_, _43040_);
  or _50848_ (_43697_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  and _50849_ (_43698_, _43697_, _43696_);
  or _50850_ (_43699_, _43698_, _42677_);
  or _50851_ (_43700_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nand _50852_ (_43701_, _42486_, _43089_);
  and _50853_ (_43702_, _43701_, _43700_);
  or _50854_ (_43703_, _43702_, _42404_);
  and _50855_ (_43704_, _43703_, _43699_);
  or _50856_ (_43705_, _43704_, _42649_);
  nand _50857_ (_43706_, _42486_, _43138_);
  or _50858_ (_43707_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _50859_ (_43708_, _43707_, _43706_);
  or _50860_ (_43709_, _43708_, _42677_);
  or _50861_ (_43710_, _42486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nand _50862_ (_43711_, _42486_, _43187_);
  and _50863_ (_43712_, _43711_, _43710_);
  or _50864_ (_43713_, _43712_, _42404_);
  and _50865_ (_43714_, _43713_, _43709_);
  or _50866_ (_43715_, _43714_, _42612_);
  and _50867_ (_43716_, _43715_, _42530_);
  and _50868_ (_43717_, _43716_, _43705_);
  or _50869_ (_43718_, _43717_, _43695_);
  or _50870_ (_43719_, _43718_, _42648_);
  or _50871_ (_43720_, _43258_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  and _50872_ (_43721_, _43720_, _42711_);
  and _50873_ (_43722_, _43721_, _43719_);
  and _50874_ (_40043_, _42814_, _42882_);
  and _50875_ (_43723_, _40043_, _42707_);
  or _50876_ (_05092_, _43723_, _43722_);
  or _50877_ (_43724_, \oc8051_gm_cxrom_1.cell0.valid , word_in[7]);
  not _50878_ (_43725_, \oc8051_gm_cxrom_1.cell0.valid );
  or _50879_ (_43726_, _43725_, \oc8051_gm_cxrom_1.cell0.data [7]);
  nand _50880_ (_43727_, _43726_, _43724_);
  nand _50881_ (_43728_, _43727_, _42882_);
  or _50882_ (_43729_, \oc8051_gm_cxrom_1.cell0.data [7], _42882_);
  and _50883_ (_05100_, _43729_, _43728_);
  or _50884_ (_43730_, word_in[0], \oc8051_gm_cxrom_1.cell0.valid );
  or _50885_ (_43731_, \oc8051_gm_cxrom_1.cell0.data [0], _43725_);
  nand _50886_ (_43732_, _43731_, _43730_);
  nand _50887_ (_43733_, _43732_, _42882_);
  or _50888_ (_43734_, \oc8051_gm_cxrom_1.cell0.data [0], _42882_);
  and _50889_ (_05107_, _43734_, _43733_);
  or _50890_ (_43735_, word_in[1], \oc8051_gm_cxrom_1.cell0.valid );
  or _50891_ (_43736_, \oc8051_gm_cxrom_1.cell0.data [1], _43725_);
  nand _50892_ (_43737_, _43736_, _43735_);
  nand _50893_ (_43738_, _43737_, _42882_);
  or _50894_ (_43739_, \oc8051_gm_cxrom_1.cell0.data [1], _42882_);
  and _50895_ (_05111_, _43739_, _43738_);
  or _50896_ (_43740_, word_in[2], \oc8051_gm_cxrom_1.cell0.valid );
  or _50897_ (_43741_, \oc8051_gm_cxrom_1.cell0.data [2], _43725_);
  nand _50898_ (_43742_, _43741_, _43740_);
  nand _50899_ (_43743_, _43742_, _42882_);
  or _50900_ (_43744_, \oc8051_gm_cxrom_1.cell0.data [2], _42882_);
  and _50901_ (_05115_, _43744_, _43743_);
  or _50902_ (_43745_, word_in[3], \oc8051_gm_cxrom_1.cell0.valid );
  or _50903_ (_43746_, \oc8051_gm_cxrom_1.cell0.data [3], _43725_);
  nand _50904_ (_43747_, _43746_, _43745_);
  nand _50905_ (_43748_, _43747_, _42882_);
  or _50906_ (_43749_, \oc8051_gm_cxrom_1.cell0.data [3], _42882_);
  and _50907_ (_05119_, _43749_, _43748_);
  or _50908_ (_43750_, word_in[4], \oc8051_gm_cxrom_1.cell0.valid );
  or _50909_ (_43751_, \oc8051_gm_cxrom_1.cell0.data [4], _43725_);
  nand _50910_ (_43752_, _43751_, _43750_);
  nand _50911_ (_43753_, _43752_, _42882_);
  or _50912_ (_43754_, \oc8051_gm_cxrom_1.cell0.data [4], _42882_);
  and _50913_ (_05123_, _43754_, _43753_);
  nor _50914_ (_43755_, word_in[5], \oc8051_gm_cxrom_1.cell0.valid );
  nor _50915_ (_43756_, \oc8051_gm_cxrom_1.cell0.data [5], _43725_);
  or _50916_ (_43757_, _43756_, _43755_);
  nand _50917_ (_43758_, _43757_, _42882_);
  or _50918_ (_43759_, \oc8051_gm_cxrom_1.cell0.data [5], _42882_);
  and _50919_ (_05126_, _43759_, _43758_);
  or _50920_ (_43760_, word_in[6], \oc8051_gm_cxrom_1.cell0.valid );
  or _50921_ (_43761_, \oc8051_gm_cxrom_1.cell0.data [6], _43725_);
  nand _50922_ (_43762_, _43761_, _43760_);
  nand _50923_ (_43763_, _43762_, _42882_);
  or _50924_ (_43764_, \oc8051_gm_cxrom_1.cell0.data [6], _42882_);
  and _50925_ (_05130_, _43764_, _43763_);
  or _50926_ (_43765_, \oc8051_gm_cxrom_1.cell1.valid , word_in[15]);
  not _50927_ (_43766_, \oc8051_gm_cxrom_1.cell1.valid );
  or _50928_ (_43767_, _43766_, \oc8051_gm_cxrom_1.cell1.data [7]);
  nand _50929_ (_43768_, _43767_, _43765_);
  nand _50930_ (_43769_, _43768_, _42882_);
  or _50931_ (_43770_, \oc8051_gm_cxrom_1.cell1.data [7], _42882_);
  and _50932_ (_05152_, _43770_, _43769_);
  or _50933_ (_43771_, word_in[8], \oc8051_gm_cxrom_1.cell1.valid );
  or _50934_ (_43772_, \oc8051_gm_cxrom_1.cell1.data [0], _43766_);
  nand _50935_ (_43773_, _43772_, _43771_);
  nand _50936_ (_43774_, _43773_, _42882_);
  or _50937_ (_43775_, \oc8051_gm_cxrom_1.cell1.data [0], _42882_);
  and _50938_ (_05159_, _43775_, _43774_);
  or _50939_ (_43776_, word_in[9], \oc8051_gm_cxrom_1.cell1.valid );
  or _50940_ (_43777_, \oc8051_gm_cxrom_1.cell1.data [1], _43766_);
  nand _50941_ (_43778_, _43777_, _43776_);
  nand _50942_ (_43779_, _43778_, _42882_);
  or _50943_ (_43780_, \oc8051_gm_cxrom_1.cell1.data [1], _42882_);
  and _50944_ (_05162_, _43780_, _43779_);
  or _50945_ (_43781_, word_in[10], \oc8051_gm_cxrom_1.cell1.valid );
  or _50946_ (_43782_, \oc8051_gm_cxrom_1.cell1.data [2], _43766_);
  nand _50947_ (_43783_, _43782_, _43781_);
  nand _50948_ (_43784_, _43783_, _42882_);
  or _50949_ (_43785_, \oc8051_gm_cxrom_1.cell1.data [2], _42882_);
  and _50950_ (_05166_, _43785_, _43784_);
  or _50951_ (_43786_, word_in[11], \oc8051_gm_cxrom_1.cell1.valid );
  or _50952_ (_43787_, \oc8051_gm_cxrom_1.cell1.data [3], _43766_);
  nand _50953_ (_43788_, _43787_, _43786_);
  nand _50954_ (_43789_, _43788_, _42882_);
  or _50955_ (_43790_, \oc8051_gm_cxrom_1.cell1.data [3], _42882_);
  and _50956_ (_05170_, _43790_, _43789_);
  or _50957_ (_43791_, word_in[12], \oc8051_gm_cxrom_1.cell1.valid );
  or _50958_ (_43792_, \oc8051_gm_cxrom_1.cell1.data [4], _43766_);
  nand _50959_ (_43793_, _43792_, _43791_);
  nand _50960_ (_43794_, _43793_, _42882_);
  or _50961_ (_43795_, \oc8051_gm_cxrom_1.cell1.data [4], _42882_);
  and _50962_ (_05174_, _43795_, _43794_);
  nor _50963_ (_43796_, word_in[13], \oc8051_gm_cxrom_1.cell1.valid );
  nor _50964_ (_43797_, \oc8051_gm_cxrom_1.cell1.data [5], _43766_);
  or _50965_ (_43798_, _43797_, _43796_);
  nand _50966_ (_43799_, _43798_, _42882_);
  or _50967_ (_43800_, \oc8051_gm_cxrom_1.cell1.data [5], _42882_);
  and _50968_ (_05178_, _43800_, _43799_);
  or _50969_ (_43801_, word_in[14], \oc8051_gm_cxrom_1.cell1.valid );
  or _50970_ (_43802_, \oc8051_gm_cxrom_1.cell1.data [6], _43766_);
  nand _50971_ (_43803_, _43802_, _43801_);
  nand _50972_ (_43804_, _43803_, _42882_);
  or _50973_ (_43805_, \oc8051_gm_cxrom_1.cell1.data [6], _42882_);
  and _50974_ (_05182_, _43805_, _43804_);
  or _50975_ (_43806_, \oc8051_gm_cxrom_1.cell2.valid , word_in[23]);
  not _50976_ (_43807_, \oc8051_gm_cxrom_1.cell2.valid );
  or _50977_ (_43808_, _43807_, \oc8051_gm_cxrom_1.cell2.data [7]);
  nand _50978_ (_43809_, _43808_, _43806_);
  nand _50979_ (_43810_, _43809_, _42882_);
  or _50980_ (_43811_, \oc8051_gm_cxrom_1.cell2.data [7], _42882_);
  and _50981_ (_05203_, _43811_, _43810_);
  or _50982_ (_00002_, word_in[16], \oc8051_gm_cxrom_1.cell2.valid );
  or _50983_ (_00003_, \oc8051_gm_cxrom_1.cell2.data [0], _43807_);
  nand _50984_ (_00004_, _00003_, _00002_);
  nand _50985_ (_00005_, _00004_, _42882_);
  or _50986_ (_00006_, \oc8051_gm_cxrom_1.cell2.data [0], _42882_);
  and _50987_ (_05210_, _00006_, _00005_);
  or _50988_ (_00007_, word_in[17], \oc8051_gm_cxrom_1.cell2.valid );
  or _50989_ (_00008_, \oc8051_gm_cxrom_1.cell2.data [1], _43807_);
  nand _50990_ (_00009_, _00008_, _00007_);
  nand _50991_ (_00010_, _00009_, _42882_);
  or _50992_ (_00011_, \oc8051_gm_cxrom_1.cell2.data [1], _42882_);
  and _50993_ (_05214_, _00011_, _00010_);
  or _50994_ (_00012_, word_in[18], \oc8051_gm_cxrom_1.cell2.valid );
  or _50995_ (_00013_, \oc8051_gm_cxrom_1.cell2.data [2], _43807_);
  nand _50996_ (_00014_, _00013_, _00012_);
  nand _50997_ (_00015_, _00014_, _42882_);
  or _50998_ (_00016_, \oc8051_gm_cxrom_1.cell2.data [2], _42882_);
  and _50999_ (_05218_, _00016_, _00015_);
  or _51000_ (_00017_, word_in[19], \oc8051_gm_cxrom_1.cell2.valid );
  or _51001_ (_00018_, \oc8051_gm_cxrom_1.cell2.data [3], _43807_);
  nand _51002_ (_00019_, _00018_, _00017_);
  nand _51003_ (_00020_, _00019_, _42882_);
  or _51004_ (_00021_, \oc8051_gm_cxrom_1.cell2.data [3], _42882_);
  and _51005_ (_05222_, _00021_, _00020_);
  or _51006_ (_00022_, word_in[20], \oc8051_gm_cxrom_1.cell2.valid );
  or _51007_ (_00023_, \oc8051_gm_cxrom_1.cell2.data [4], _43807_);
  nand _51008_ (_00024_, _00023_, _00022_);
  nand _51009_ (_00025_, _00024_, _42882_);
  or _51010_ (_00026_, \oc8051_gm_cxrom_1.cell2.data [4], _42882_);
  and _51011_ (_05226_, _00026_, _00025_);
  nor _51012_ (_00027_, word_in[21], \oc8051_gm_cxrom_1.cell2.valid );
  nor _51013_ (_00028_, \oc8051_gm_cxrom_1.cell2.data [5], _43807_);
  or _51014_ (_00029_, _00028_, _00027_);
  nand _51015_ (_00030_, _00029_, _42882_);
  or _51016_ (_00031_, \oc8051_gm_cxrom_1.cell2.data [5], _42882_);
  and _51017_ (_05230_, _00031_, _00030_);
  or _51018_ (_00032_, word_in[22], \oc8051_gm_cxrom_1.cell2.valid );
  or _51019_ (_00033_, \oc8051_gm_cxrom_1.cell2.data [6], _43807_);
  nand _51020_ (_00034_, _00033_, _00032_);
  nand _51021_ (_00035_, _00034_, _42882_);
  or _51022_ (_00036_, \oc8051_gm_cxrom_1.cell2.data [6], _42882_);
  and _51023_ (_05234_, _00036_, _00035_);
  or _51024_ (_00037_, \oc8051_gm_cxrom_1.cell3.valid , word_in[31]);
  not _51025_ (_00038_, \oc8051_gm_cxrom_1.cell3.valid );
  or _51026_ (_00039_, _00038_, \oc8051_gm_cxrom_1.cell3.data [7]);
  nand _51027_ (_00040_, _00039_, _00037_);
  nand _51028_ (_00041_, _00040_, _42882_);
  or _51029_ (_00042_, \oc8051_gm_cxrom_1.cell3.data [7], _42882_);
  and _51030_ (_05255_, _00042_, _00041_);
  or _51031_ (_00043_, word_in[24], \oc8051_gm_cxrom_1.cell3.valid );
  or _51032_ (_00044_, \oc8051_gm_cxrom_1.cell3.data [0], _00038_);
  nand _51033_ (_00045_, _00044_, _00043_);
  nand _51034_ (_00046_, _00045_, _42882_);
  or _51035_ (_00047_, \oc8051_gm_cxrom_1.cell3.data [0], _42882_);
  and _51036_ (_05262_, _00047_, _00046_);
  or _51037_ (_00048_, word_in[25], \oc8051_gm_cxrom_1.cell3.valid );
  or _51038_ (_00049_, \oc8051_gm_cxrom_1.cell3.data [1], _00038_);
  nand _51039_ (_00050_, _00049_, _00048_);
  nand _51040_ (_00051_, _00050_, _42882_);
  or _51041_ (_00052_, \oc8051_gm_cxrom_1.cell3.data [1], _42882_);
  and _51042_ (_05266_, _00052_, _00051_);
  or _51043_ (_00053_, word_in[26], \oc8051_gm_cxrom_1.cell3.valid );
  or _51044_ (_00054_, \oc8051_gm_cxrom_1.cell3.data [2], _00038_);
  nand _51045_ (_00055_, _00054_, _00053_);
  nand _51046_ (_00056_, _00055_, _42882_);
  or _51047_ (_00057_, \oc8051_gm_cxrom_1.cell3.data [2], _42882_);
  and _51048_ (_05270_, _00057_, _00056_);
  or _51049_ (_00058_, word_in[27], \oc8051_gm_cxrom_1.cell3.valid );
  or _51050_ (_00059_, \oc8051_gm_cxrom_1.cell3.data [3], _00038_);
  nand _51051_ (_00060_, _00059_, _00058_);
  nand _51052_ (_00061_, _00060_, _42882_);
  or _51053_ (_00062_, \oc8051_gm_cxrom_1.cell3.data [3], _42882_);
  and _51054_ (_05273_, _00062_, _00061_);
  or _51055_ (_00063_, word_in[28], \oc8051_gm_cxrom_1.cell3.valid );
  or _51056_ (_00064_, \oc8051_gm_cxrom_1.cell3.data [4], _00038_);
  nand _51057_ (_00065_, _00064_, _00063_);
  nand _51058_ (_00066_, _00065_, _42882_);
  or _51059_ (_00067_, \oc8051_gm_cxrom_1.cell3.data [4], _42882_);
  and _51060_ (_05277_, _00067_, _00066_);
  nor _51061_ (_00068_, word_in[29], \oc8051_gm_cxrom_1.cell3.valid );
  nor _51062_ (_00069_, \oc8051_gm_cxrom_1.cell3.data [5], _00038_);
  or _51063_ (_00070_, _00069_, _00068_);
  nand _51064_ (_00071_, _00070_, _42882_);
  or _51065_ (_00072_, \oc8051_gm_cxrom_1.cell3.data [5], _42882_);
  and _51066_ (_05281_, _00072_, _00071_);
  or _51067_ (_00073_, word_in[30], \oc8051_gm_cxrom_1.cell3.valid );
  or _51068_ (_00074_, \oc8051_gm_cxrom_1.cell3.data [6], _00038_);
  nand _51069_ (_00075_, _00074_, _00073_);
  nand _51070_ (_00076_, _00075_, _42882_);
  or _51071_ (_00077_, \oc8051_gm_cxrom_1.cell3.data [6], _42882_);
  and _51072_ (_05285_, _00077_, _00076_);
  or _51073_ (_00078_, \oc8051_gm_cxrom_1.cell4.valid , word_in[39]);
  not _51074_ (_00079_, \oc8051_gm_cxrom_1.cell4.valid );
  or _51075_ (_00080_, _00079_, \oc8051_gm_cxrom_1.cell4.data [7]);
  nand _51076_ (_00081_, _00080_, _00078_);
  nand _51077_ (_00082_, _00081_, _42882_);
  or _51078_ (_00083_, \oc8051_gm_cxrom_1.cell4.data [7], _42882_);
  and _51079_ (_05306_, _00083_, _00082_);
  or _51080_ (_00084_, word_in[32], \oc8051_gm_cxrom_1.cell4.valid );
  or _51081_ (_00085_, \oc8051_gm_cxrom_1.cell4.data [0], _00079_);
  nand _51082_ (_00086_, _00085_, _00084_);
  nand _51083_ (_00087_, _00086_, _42882_);
  or _51084_ (_00088_, \oc8051_gm_cxrom_1.cell4.data [0], _42882_);
  and _51085_ (_05313_, _00088_, _00087_);
  or _51086_ (_00089_, word_in[33], \oc8051_gm_cxrom_1.cell4.valid );
  or _51087_ (_00090_, \oc8051_gm_cxrom_1.cell4.data [1], _00079_);
  nand _51088_ (_00091_, _00090_, _00089_);
  nand _51089_ (_00092_, _00091_, _42882_);
  or _51090_ (_00093_, \oc8051_gm_cxrom_1.cell4.data [1], _42882_);
  and _51091_ (_05317_, _00093_, _00092_);
  or _51092_ (_00094_, word_in[34], \oc8051_gm_cxrom_1.cell4.valid );
  or _51093_ (_00095_, \oc8051_gm_cxrom_1.cell4.data [2], _00079_);
  nand _51094_ (_00096_, _00095_, _00094_);
  nand _51095_ (_00097_, _00096_, _42882_);
  or _51096_ (_00098_, \oc8051_gm_cxrom_1.cell4.data [2], _42882_);
  and _51097_ (_05321_, _00098_, _00097_);
  or _51098_ (_00099_, word_in[35], \oc8051_gm_cxrom_1.cell4.valid );
  or _51099_ (_00100_, \oc8051_gm_cxrom_1.cell4.data [3], _00079_);
  nand _51100_ (_00101_, _00100_, _00099_);
  nand _51101_ (_00102_, _00101_, _42882_);
  or _51102_ (_00103_, \oc8051_gm_cxrom_1.cell4.data [3], _42882_);
  and _51103_ (_05325_, _00103_, _00102_);
  or _51104_ (_00104_, word_in[36], \oc8051_gm_cxrom_1.cell4.valid );
  or _51105_ (_00105_, \oc8051_gm_cxrom_1.cell4.data [4], _00079_);
  nand _51106_ (_00106_, _00105_, _00104_);
  nand _51107_ (_00107_, _00106_, _42882_);
  or _51108_ (_00108_, \oc8051_gm_cxrom_1.cell4.data [4], _42882_);
  and _51109_ (_05329_, _00108_, _00107_);
  nor _51110_ (_00109_, word_in[37], \oc8051_gm_cxrom_1.cell4.valid );
  nor _51111_ (_00110_, \oc8051_gm_cxrom_1.cell4.data [5], _00079_);
  or _51112_ (_00111_, _00110_, _00109_);
  nand _51113_ (_00112_, _00111_, _42882_);
  or _51114_ (_00113_, \oc8051_gm_cxrom_1.cell4.data [5], _42882_);
  and _51115_ (_05333_, _00113_, _00112_);
  or _51116_ (_00114_, word_in[38], \oc8051_gm_cxrom_1.cell4.valid );
  or _51117_ (_00115_, \oc8051_gm_cxrom_1.cell4.data [6], _00079_);
  nand _51118_ (_00116_, _00115_, _00114_);
  nand _51119_ (_00117_, _00116_, _42882_);
  or _51120_ (_00118_, \oc8051_gm_cxrom_1.cell4.data [6], _42882_);
  and _51121_ (_05337_, _00118_, _00117_);
  or _51122_ (_00119_, \oc8051_gm_cxrom_1.cell5.valid , word_in[47]);
  not _51123_ (_00120_, \oc8051_gm_cxrom_1.cell5.valid );
  or _51124_ (_00121_, _00120_, \oc8051_gm_cxrom_1.cell5.data [7]);
  nand _51125_ (_00122_, _00121_, _00119_);
  nand _51126_ (_00123_, _00122_, _42882_);
  or _51127_ (_00124_, \oc8051_gm_cxrom_1.cell5.data [7], _42882_);
  and _51128_ (_05359_, _00124_, _00123_);
  or _51129_ (_00125_, word_in[40], \oc8051_gm_cxrom_1.cell5.valid );
  or _51130_ (_00126_, \oc8051_gm_cxrom_1.cell5.data [0], _00120_);
  nand _51131_ (_00127_, _00126_, _00125_);
  nand _51132_ (_00128_, _00127_, _42882_);
  or _51133_ (_00129_, \oc8051_gm_cxrom_1.cell5.data [0], _42882_);
  and _51134_ (_05366_, _00129_, _00128_);
  or _51135_ (_00131_, word_in[41], \oc8051_gm_cxrom_1.cell5.valid );
  or _51136_ (_00133_, \oc8051_gm_cxrom_1.cell5.data [1], _00120_);
  nand _51137_ (_00135_, _00133_, _00131_);
  nand _51138_ (_00137_, _00135_, _42882_);
  or _51139_ (_00139_, \oc8051_gm_cxrom_1.cell5.data [1], _42882_);
  and _51140_ (_05370_, _00139_, _00137_);
  or _51141_ (_00142_, word_in[42], \oc8051_gm_cxrom_1.cell5.valid );
  or _51142_ (_00144_, \oc8051_gm_cxrom_1.cell5.data [2], _00120_);
  nand _51143_ (_00146_, _00144_, _00142_);
  nand _51144_ (_00148_, _00146_, _42882_);
  or _51145_ (_00150_, \oc8051_gm_cxrom_1.cell5.data [2], _42882_);
  and _51146_ (_05374_, _00150_, _00148_);
  or _51147_ (_00153_, word_in[43], \oc8051_gm_cxrom_1.cell5.valid );
  or _51148_ (_00155_, \oc8051_gm_cxrom_1.cell5.data [3], _00120_);
  nand _51149_ (_00157_, _00155_, _00153_);
  nand _51150_ (_00159_, _00157_, _42882_);
  or _51151_ (_00161_, \oc8051_gm_cxrom_1.cell5.data [3], _42882_);
  and _51152_ (_05378_, _00161_, _00159_);
  or _51153_ (_00164_, word_in[44], \oc8051_gm_cxrom_1.cell5.valid );
  or _51154_ (_00166_, \oc8051_gm_cxrom_1.cell5.data [4], _00120_);
  nand _51155_ (_00168_, _00166_, _00164_);
  nand _51156_ (_00170_, _00168_, _42882_);
  or _51157_ (_00172_, \oc8051_gm_cxrom_1.cell5.data [4], _42882_);
  and _51158_ (_05382_, _00172_, _00170_);
  nor _51159_ (_00175_, word_in[45], \oc8051_gm_cxrom_1.cell5.valid );
  nor _51160_ (_00177_, \oc8051_gm_cxrom_1.cell5.data [5], _00120_);
  or _51161_ (_00179_, _00177_, _00175_);
  nand _51162_ (_00181_, _00179_, _42882_);
  or _51163_ (_00183_, \oc8051_gm_cxrom_1.cell5.data [5], _42882_);
  and _51164_ (_05386_, _00183_, _00181_);
  or _51165_ (_00186_, word_in[46], \oc8051_gm_cxrom_1.cell5.valid );
  or _51166_ (_00187_, \oc8051_gm_cxrom_1.cell5.data [6], _00120_);
  nand _51167_ (_00188_, _00187_, _00186_);
  nand _51168_ (_00189_, _00188_, _42882_);
  or _51169_ (_00190_, \oc8051_gm_cxrom_1.cell5.data [6], _42882_);
  and _51170_ (_05390_, _00190_, _00189_);
  or _51171_ (_00191_, \oc8051_gm_cxrom_1.cell6.valid , word_in[55]);
  not _51172_ (_00192_, \oc8051_gm_cxrom_1.cell6.valid );
  or _51173_ (_00193_, _00192_, \oc8051_gm_cxrom_1.cell6.data [7]);
  nand _51174_ (_00194_, _00193_, _00191_);
  nand _51175_ (_00195_, _00194_, _42882_);
  or _51176_ (_00196_, \oc8051_gm_cxrom_1.cell6.data [7], _42882_);
  and _51177_ (_05412_, _00196_, _00195_);
  or _51178_ (_00197_, word_in[48], \oc8051_gm_cxrom_1.cell6.valid );
  or _51179_ (_00198_, \oc8051_gm_cxrom_1.cell6.data [0], _00192_);
  nand _51180_ (_00199_, _00198_, _00197_);
  nand _51181_ (_00200_, _00199_, _42882_);
  or _51182_ (_00201_, \oc8051_gm_cxrom_1.cell6.data [0], _42882_);
  and _51183_ (_05419_, _00201_, _00200_);
  or _51184_ (_00202_, word_in[49], \oc8051_gm_cxrom_1.cell6.valid );
  or _51185_ (_00203_, \oc8051_gm_cxrom_1.cell6.data [1], _00192_);
  nand _51186_ (_00204_, _00203_, _00202_);
  nand _51187_ (_00205_, _00204_, _42882_);
  or _51188_ (_00206_, \oc8051_gm_cxrom_1.cell6.data [1], _42882_);
  and _51189_ (_05423_, _00206_, _00205_);
  or _51190_ (_00207_, word_in[50], \oc8051_gm_cxrom_1.cell6.valid );
  or _51191_ (_00208_, \oc8051_gm_cxrom_1.cell6.data [2], _00192_);
  nand _51192_ (_00209_, _00208_, _00207_);
  nand _51193_ (_00210_, _00209_, _42882_);
  or _51194_ (_00211_, \oc8051_gm_cxrom_1.cell6.data [2], _42882_);
  and _51195_ (_05427_, _00211_, _00210_);
  or _51196_ (_00212_, word_in[51], \oc8051_gm_cxrom_1.cell6.valid );
  or _51197_ (_00213_, \oc8051_gm_cxrom_1.cell6.data [3], _00192_);
  nand _51198_ (_00214_, _00213_, _00212_);
  nand _51199_ (_00215_, _00214_, _42882_);
  or _51200_ (_00216_, \oc8051_gm_cxrom_1.cell6.data [3], _42882_);
  and _51201_ (_05431_, _00216_, _00215_);
  or _51202_ (_00217_, word_in[52], \oc8051_gm_cxrom_1.cell6.valid );
  or _51203_ (_00218_, \oc8051_gm_cxrom_1.cell6.data [4], _00192_);
  nand _51204_ (_00219_, _00218_, _00217_);
  nand _51205_ (_00220_, _00219_, _42882_);
  or _51206_ (_00221_, \oc8051_gm_cxrom_1.cell6.data [4], _42882_);
  and _51207_ (_05435_, _00221_, _00220_);
  nor _51208_ (_00222_, word_in[53], \oc8051_gm_cxrom_1.cell6.valid );
  nor _51209_ (_00223_, \oc8051_gm_cxrom_1.cell6.data [5], _00192_);
  or _51210_ (_00224_, _00223_, _00222_);
  nand _51211_ (_00225_, _00224_, _42882_);
  or _51212_ (_00226_, \oc8051_gm_cxrom_1.cell6.data [5], _42882_);
  and _51213_ (_05439_, _00226_, _00225_);
  or _51214_ (_00227_, word_in[54], \oc8051_gm_cxrom_1.cell6.valid );
  or _51215_ (_00228_, \oc8051_gm_cxrom_1.cell6.data [6], _00192_);
  nand _51216_ (_00229_, _00228_, _00227_);
  nand _51217_ (_00230_, _00229_, _42882_);
  or _51218_ (_00231_, \oc8051_gm_cxrom_1.cell6.data [6], _42882_);
  and _51219_ (_05443_, _00231_, _00230_);
  or _51220_ (_00232_, \oc8051_gm_cxrom_1.cell7.valid , word_in[63]);
  not _51221_ (_00233_, \oc8051_gm_cxrom_1.cell7.valid );
  or _51222_ (_00234_, _00233_, \oc8051_gm_cxrom_1.cell7.data [7]);
  nand _51223_ (_00235_, _00234_, _00232_);
  nand _51224_ (_00236_, _00235_, _42882_);
  or _51225_ (_00237_, \oc8051_gm_cxrom_1.cell7.data [7], _42882_);
  and _51226_ (_05465_, _00237_, _00236_);
  or _51227_ (_00238_, word_in[56], \oc8051_gm_cxrom_1.cell7.valid );
  or _51228_ (_00239_, \oc8051_gm_cxrom_1.cell7.data [0], _00233_);
  nand _51229_ (_00240_, _00239_, _00238_);
  nand _51230_ (_00241_, _00240_, _42882_);
  or _51231_ (_00242_, \oc8051_gm_cxrom_1.cell7.data [0], _42882_);
  and _51232_ (_05472_, _00242_, _00241_);
  or _51233_ (_00243_, word_in[57], \oc8051_gm_cxrom_1.cell7.valid );
  or _51234_ (_00244_, \oc8051_gm_cxrom_1.cell7.data [1], _00233_);
  nand _51235_ (_00245_, _00244_, _00243_);
  nand _51236_ (_00246_, _00245_, _42882_);
  or _51237_ (_00247_, \oc8051_gm_cxrom_1.cell7.data [1], _42882_);
  and _51238_ (_05476_, _00247_, _00246_);
  or _51239_ (_00248_, word_in[58], \oc8051_gm_cxrom_1.cell7.valid );
  or _51240_ (_00249_, \oc8051_gm_cxrom_1.cell7.data [2], _00233_);
  nand _51241_ (_00250_, _00249_, _00248_);
  nand _51242_ (_00251_, _00250_, _42882_);
  or _51243_ (_00252_, \oc8051_gm_cxrom_1.cell7.data [2], _42882_);
  and _51244_ (_05480_, _00252_, _00251_);
  or _51245_ (_00253_, word_in[59], \oc8051_gm_cxrom_1.cell7.valid );
  or _51246_ (_00254_, \oc8051_gm_cxrom_1.cell7.data [3], _00233_);
  nand _51247_ (_00255_, _00254_, _00253_);
  nand _51248_ (_00256_, _00255_, _42882_);
  or _51249_ (_00257_, \oc8051_gm_cxrom_1.cell7.data [3], _42882_);
  and _51250_ (_05484_, _00257_, _00256_);
  or _51251_ (_00258_, word_in[60], \oc8051_gm_cxrom_1.cell7.valid );
  or _51252_ (_00259_, \oc8051_gm_cxrom_1.cell7.data [4], _00233_);
  nand _51253_ (_00260_, _00259_, _00258_);
  nand _51254_ (_00261_, _00260_, _42882_);
  or _51255_ (_00262_, \oc8051_gm_cxrom_1.cell7.data [4], _42882_);
  and _51256_ (_05488_, _00262_, _00261_);
  nor _51257_ (_00263_, word_in[61], \oc8051_gm_cxrom_1.cell7.valid );
  nor _51258_ (_00264_, \oc8051_gm_cxrom_1.cell7.data [5], _00233_);
  or _51259_ (_00265_, _00264_, _00263_);
  nand _51260_ (_00266_, _00265_, _42882_);
  or _51261_ (_00267_, \oc8051_gm_cxrom_1.cell7.data [5], _42882_);
  and _51262_ (_05492_, _00267_, _00266_);
  or _51263_ (_00268_, word_in[62], \oc8051_gm_cxrom_1.cell7.valid );
  or _51264_ (_00269_, \oc8051_gm_cxrom_1.cell7.data [6], _00233_);
  nand _51265_ (_00270_, _00269_, _00268_);
  nand _51266_ (_00271_, _00270_, _42882_);
  or _51267_ (_00272_, \oc8051_gm_cxrom_1.cell7.data [6], _42882_);
  and _51268_ (_05496_, _00272_, _00271_);
  or _51269_ (_00273_, \oc8051_gm_cxrom_1.cell8.valid , word_in[71]);
  not _51270_ (_00274_, \oc8051_gm_cxrom_1.cell8.valid );
  or _51271_ (_00275_, _00274_, \oc8051_gm_cxrom_1.cell8.data [7]);
  nand _51272_ (_00276_, _00275_, _00273_);
  nand _51273_ (_00277_, _00276_, _42882_);
  or _51274_ (_00278_, \oc8051_gm_cxrom_1.cell8.data [7], _42882_);
  and _51275_ (_05518_, _00278_, _00277_);
  or _51276_ (_00279_, word_in[64], \oc8051_gm_cxrom_1.cell8.valid );
  or _51277_ (_00280_, \oc8051_gm_cxrom_1.cell8.data [0], _00274_);
  nand _51278_ (_00281_, _00280_, _00279_);
  nand _51279_ (_00282_, _00281_, _42882_);
  or _51280_ (_00283_, \oc8051_gm_cxrom_1.cell8.data [0], _42882_);
  and _51281_ (_05525_, _00283_, _00282_);
  or _51282_ (_00284_, word_in[65], \oc8051_gm_cxrom_1.cell8.valid );
  or _51283_ (_00285_, \oc8051_gm_cxrom_1.cell8.data [1], _00274_);
  nand _51284_ (_00286_, _00285_, _00284_);
  nand _51285_ (_00287_, _00286_, _42882_);
  or _51286_ (_00288_, \oc8051_gm_cxrom_1.cell8.data [1], _42882_);
  and _51287_ (_05529_, _00288_, _00287_);
  or _51288_ (_00289_, word_in[66], \oc8051_gm_cxrom_1.cell8.valid );
  or _51289_ (_00290_, \oc8051_gm_cxrom_1.cell8.data [2], _00274_);
  nand _51290_ (_00291_, _00290_, _00289_);
  nand _51291_ (_00292_, _00291_, _42882_);
  or _51292_ (_00293_, \oc8051_gm_cxrom_1.cell8.data [2], _42882_);
  and _51293_ (_05533_, _00293_, _00292_);
  or _51294_ (_00294_, word_in[67], \oc8051_gm_cxrom_1.cell8.valid );
  or _51295_ (_00295_, \oc8051_gm_cxrom_1.cell8.data [3], _00274_);
  nand _51296_ (_00296_, _00295_, _00294_);
  nand _51297_ (_00297_, _00296_, _42882_);
  or _51298_ (_00298_, \oc8051_gm_cxrom_1.cell8.data [3], _42882_);
  and _51299_ (_05537_, _00298_, _00297_);
  or _51300_ (_00299_, word_in[68], \oc8051_gm_cxrom_1.cell8.valid );
  or _51301_ (_00300_, \oc8051_gm_cxrom_1.cell8.data [4], _00274_);
  nand _51302_ (_00301_, _00300_, _00299_);
  nand _51303_ (_00302_, _00301_, _42882_);
  or _51304_ (_00303_, \oc8051_gm_cxrom_1.cell8.data [4], _42882_);
  and _51305_ (_05541_, _00303_, _00302_);
  nor _51306_ (_00304_, word_in[69], \oc8051_gm_cxrom_1.cell8.valid );
  nor _51307_ (_00305_, \oc8051_gm_cxrom_1.cell8.data [5], _00274_);
  or _51308_ (_00306_, _00305_, _00304_);
  nand _51309_ (_00307_, _00306_, _42882_);
  or _51310_ (_00308_, \oc8051_gm_cxrom_1.cell8.data [5], _42882_);
  and _51311_ (_05545_, _00308_, _00307_);
  or _51312_ (_00309_, word_in[70], \oc8051_gm_cxrom_1.cell8.valid );
  or _51313_ (_00310_, \oc8051_gm_cxrom_1.cell8.data [6], _00274_);
  nand _51314_ (_00311_, _00310_, _00309_);
  nand _51315_ (_00312_, _00311_, _42882_);
  or _51316_ (_00313_, \oc8051_gm_cxrom_1.cell8.data [6], _42882_);
  and _51317_ (_05549_, _00313_, _00312_);
  or _51318_ (_00314_, \oc8051_gm_cxrom_1.cell9.valid , word_in[79]);
  not _51319_ (_00315_, \oc8051_gm_cxrom_1.cell9.valid );
  or _51320_ (_00316_, _00315_, \oc8051_gm_cxrom_1.cell9.data [7]);
  nand _51321_ (_00317_, _00316_, _00314_);
  nand _51322_ (_00318_, _00317_, _42882_);
  or _51323_ (_00319_, \oc8051_gm_cxrom_1.cell9.data [7], _42882_);
  and _51324_ (_05571_, _00319_, _00318_);
  or _51325_ (_00320_, word_in[72], \oc8051_gm_cxrom_1.cell9.valid );
  or _51326_ (_00321_, \oc8051_gm_cxrom_1.cell9.data [0], _00315_);
  nand _51327_ (_00322_, _00321_, _00320_);
  nand _51328_ (_00323_, _00322_, _42882_);
  or _51329_ (_00324_, \oc8051_gm_cxrom_1.cell9.data [0], _42882_);
  and _51330_ (_05578_, _00324_, _00323_);
  or _51331_ (_00325_, word_in[73], \oc8051_gm_cxrom_1.cell9.valid );
  or _51332_ (_00326_, \oc8051_gm_cxrom_1.cell9.data [1], _00315_);
  nand _51333_ (_00327_, _00326_, _00325_);
  nand _51334_ (_00328_, _00327_, _42882_);
  or _51335_ (_00329_, \oc8051_gm_cxrom_1.cell9.data [1], _42882_);
  and _51336_ (_05582_, _00329_, _00328_);
  or _51337_ (_00330_, word_in[74], \oc8051_gm_cxrom_1.cell9.valid );
  or _51338_ (_00331_, \oc8051_gm_cxrom_1.cell9.data [2], _00315_);
  nand _51339_ (_00332_, _00331_, _00330_);
  nand _51340_ (_00333_, _00332_, _42882_);
  or _51341_ (_00334_, \oc8051_gm_cxrom_1.cell9.data [2], _42882_);
  and _51342_ (_05586_, _00334_, _00333_);
  or _51343_ (_00335_, word_in[75], \oc8051_gm_cxrom_1.cell9.valid );
  or _51344_ (_00336_, \oc8051_gm_cxrom_1.cell9.data [3], _00315_);
  nand _51345_ (_00337_, _00336_, _00335_);
  nand _51346_ (_00338_, _00337_, _42882_);
  or _51347_ (_00339_, \oc8051_gm_cxrom_1.cell9.data [3], _42882_);
  and _51348_ (_05590_, _00339_, _00338_);
  or _51349_ (_00340_, word_in[76], \oc8051_gm_cxrom_1.cell9.valid );
  or _51350_ (_00341_, \oc8051_gm_cxrom_1.cell9.data [4], _00315_);
  nand _51351_ (_00342_, _00341_, _00340_);
  nand _51352_ (_00343_, _00342_, _42882_);
  or _51353_ (_00344_, \oc8051_gm_cxrom_1.cell9.data [4], _42882_);
  and _51354_ (_05594_, _00344_, _00343_);
  nor _51355_ (_00345_, word_in[77], \oc8051_gm_cxrom_1.cell9.valid );
  nor _51356_ (_00346_, \oc8051_gm_cxrom_1.cell9.data [5], _00315_);
  or _51357_ (_00347_, _00346_, _00345_);
  nand _51358_ (_00348_, _00347_, _42882_);
  or _51359_ (_00349_, \oc8051_gm_cxrom_1.cell9.data [5], _42882_);
  and _51360_ (_05598_, _00349_, _00348_);
  or _51361_ (_00350_, word_in[78], \oc8051_gm_cxrom_1.cell9.valid );
  or _51362_ (_00351_, \oc8051_gm_cxrom_1.cell9.data [6], _00315_);
  nand _51363_ (_00352_, _00351_, _00350_);
  nand _51364_ (_00353_, _00352_, _42882_);
  or _51365_ (_00354_, \oc8051_gm_cxrom_1.cell9.data [6], _42882_);
  and _51366_ (_05602_, _00354_, _00353_);
  or _51367_ (_00355_, \oc8051_gm_cxrom_1.cell10.valid , word_in[87]);
  not _51368_ (_00356_, \oc8051_gm_cxrom_1.cell10.valid );
  or _51369_ (_00357_, _00356_, \oc8051_gm_cxrom_1.cell10.data [7]);
  nand _51370_ (_00358_, _00357_, _00355_);
  nand _51371_ (_00359_, _00358_, _42882_);
  or _51372_ (_00360_, \oc8051_gm_cxrom_1.cell10.data [7], _42882_);
  and _51373_ (_05624_, _00360_, _00359_);
  or _51374_ (_00361_, word_in[80], \oc8051_gm_cxrom_1.cell10.valid );
  or _51375_ (_00362_, \oc8051_gm_cxrom_1.cell10.data [0], _00356_);
  nand _51376_ (_00363_, _00362_, _00361_);
  nand _51377_ (_00364_, _00363_, _42882_);
  or _51378_ (_00365_, \oc8051_gm_cxrom_1.cell10.data [0], _42882_);
  and _51379_ (_05631_, _00365_, _00364_);
  or _51380_ (_00366_, word_in[81], \oc8051_gm_cxrom_1.cell10.valid );
  or _51381_ (_00367_, \oc8051_gm_cxrom_1.cell10.data [1], _00356_);
  nand _51382_ (_00368_, _00367_, _00366_);
  nand _51383_ (_00369_, _00368_, _42882_);
  or _51384_ (_00370_, \oc8051_gm_cxrom_1.cell10.data [1], _42882_);
  and _51385_ (_05635_, _00370_, _00369_);
  or _51386_ (_00371_, word_in[82], \oc8051_gm_cxrom_1.cell10.valid );
  or _51387_ (_00372_, \oc8051_gm_cxrom_1.cell10.data [2], _00356_);
  nand _51388_ (_00373_, _00372_, _00371_);
  nand _51389_ (_00374_, _00373_, _42882_);
  or _51390_ (_00375_, \oc8051_gm_cxrom_1.cell10.data [2], _42882_);
  and _51391_ (_05639_, _00375_, _00374_);
  or _51392_ (_00376_, word_in[83], \oc8051_gm_cxrom_1.cell10.valid );
  or _51393_ (_00377_, \oc8051_gm_cxrom_1.cell10.data [3], _00356_);
  nand _51394_ (_00378_, _00377_, _00376_);
  nand _51395_ (_00379_, _00378_, _42882_);
  or _51396_ (_00380_, \oc8051_gm_cxrom_1.cell10.data [3], _42882_);
  and _51397_ (_05643_, _00380_, _00379_);
  or _51398_ (_00381_, word_in[84], \oc8051_gm_cxrom_1.cell10.valid );
  or _51399_ (_00382_, \oc8051_gm_cxrom_1.cell10.data [4], _00356_);
  nand _51400_ (_00383_, _00382_, _00381_);
  nand _51401_ (_00384_, _00383_, _42882_);
  or _51402_ (_00385_, \oc8051_gm_cxrom_1.cell10.data [4], _42882_);
  and _51403_ (_05647_, _00385_, _00384_);
  nor _51404_ (_00386_, word_in[85], \oc8051_gm_cxrom_1.cell10.valid );
  nor _51405_ (_00387_, \oc8051_gm_cxrom_1.cell10.data [5], _00356_);
  or _51406_ (_00388_, _00387_, _00386_);
  nand _51407_ (_00389_, _00388_, _42882_);
  or _51408_ (_00390_, \oc8051_gm_cxrom_1.cell10.data [5], _42882_);
  and _51409_ (_05651_, _00390_, _00389_);
  or _51410_ (_00391_, word_in[86], \oc8051_gm_cxrom_1.cell10.valid );
  or _51411_ (_00392_, \oc8051_gm_cxrom_1.cell10.data [6], _00356_);
  nand _51412_ (_00393_, _00392_, _00391_);
  nand _51413_ (_00394_, _00393_, _42882_);
  or _51414_ (_00395_, \oc8051_gm_cxrom_1.cell10.data [6], _42882_);
  and _51415_ (_05655_, _00395_, _00394_);
  or _51416_ (_00396_, \oc8051_gm_cxrom_1.cell11.valid , word_in[95]);
  not _51417_ (_00397_, \oc8051_gm_cxrom_1.cell11.valid );
  or _51418_ (_00398_, _00397_, \oc8051_gm_cxrom_1.cell11.data [7]);
  nand _51419_ (_00399_, _00398_, _00396_);
  nand _51420_ (_00400_, _00399_, _42882_);
  or _51421_ (_00401_, \oc8051_gm_cxrom_1.cell11.data [7], _42882_);
  and _51422_ (_05677_, _00401_, _00400_);
  or _51423_ (_00402_, word_in[88], \oc8051_gm_cxrom_1.cell11.valid );
  or _51424_ (_00403_, \oc8051_gm_cxrom_1.cell11.data [0], _00397_);
  nand _51425_ (_00404_, _00403_, _00402_);
  nand _51426_ (_00405_, _00404_, _42882_);
  or _51427_ (_00406_, \oc8051_gm_cxrom_1.cell11.data [0], _42882_);
  and _51428_ (_05684_, _00406_, _00405_);
  or _51429_ (_00407_, word_in[89], \oc8051_gm_cxrom_1.cell11.valid );
  or _51430_ (_00408_, \oc8051_gm_cxrom_1.cell11.data [1], _00397_);
  nand _51431_ (_00409_, _00408_, _00407_);
  nand _51432_ (_00410_, _00409_, _42882_);
  or _51433_ (_00411_, \oc8051_gm_cxrom_1.cell11.data [1], _42882_);
  and _51434_ (_05688_, _00411_, _00410_);
  or _51435_ (_00412_, word_in[90], \oc8051_gm_cxrom_1.cell11.valid );
  or _51436_ (_00413_, \oc8051_gm_cxrom_1.cell11.data [2], _00397_);
  nand _51437_ (_00414_, _00413_, _00412_);
  nand _51438_ (_00415_, _00414_, _42882_);
  or _51439_ (_00416_, \oc8051_gm_cxrom_1.cell11.data [2], _42882_);
  and _51440_ (_05692_, _00416_, _00415_);
  or _51441_ (_00417_, word_in[91], \oc8051_gm_cxrom_1.cell11.valid );
  or _51442_ (_00418_, \oc8051_gm_cxrom_1.cell11.data [3], _00397_);
  nand _51443_ (_00419_, _00418_, _00417_);
  nand _51444_ (_00420_, _00419_, _42882_);
  or _51445_ (_00421_, \oc8051_gm_cxrom_1.cell11.data [3], _42882_);
  and _51446_ (_05696_, _00421_, _00420_);
  or _51447_ (_00422_, word_in[92], \oc8051_gm_cxrom_1.cell11.valid );
  or _51448_ (_00423_, \oc8051_gm_cxrom_1.cell11.data [4], _00397_);
  nand _51449_ (_00424_, _00423_, _00422_);
  nand _51450_ (_00425_, _00424_, _42882_);
  or _51451_ (_00426_, \oc8051_gm_cxrom_1.cell11.data [4], _42882_);
  and _51452_ (_05700_, _00426_, _00425_);
  nor _51453_ (_00427_, word_in[93], \oc8051_gm_cxrom_1.cell11.valid );
  nor _51454_ (_00428_, \oc8051_gm_cxrom_1.cell11.data [5], _00397_);
  or _51455_ (_00429_, _00428_, _00427_);
  nand _51456_ (_00430_, _00429_, _42882_);
  or _51457_ (_00431_, \oc8051_gm_cxrom_1.cell11.data [5], _42882_);
  and _51458_ (_05704_, _00431_, _00430_);
  or _51459_ (_00432_, word_in[94], \oc8051_gm_cxrom_1.cell11.valid );
  or _51460_ (_00433_, \oc8051_gm_cxrom_1.cell11.data [6], _00397_);
  nand _51461_ (_00434_, _00433_, _00432_);
  nand _51462_ (_00435_, _00434_, _42882_);
  or _51463_ (_00436_, \oc8051_gm_cxrom_1.cell11.data [6], _42882_);
  and _51464_ (_05708_, _00436_, _00435_);
  or _51465_ (_00437_, \oc8051_gm_cxrom_1.cell12.valid , word_in[103]);
  not _51466_ (_00438_, \oc8051_gm_cxrom_1.cell12.valid );
  or _51467_ (_00439_, _00438_, \oc8051_gm_cxrom_1.cell12.data [7]);
  nand _51468_ (_00440_, _00439_, _00437_);
  nand _51469_ (_00441_, _00440_, _42882_);
  or _51470_ (_00442_, \oc8051_gm_cxrom_1.cell12.data [7], _42882_);
  and _51471_ (_05730_, _00442_, _00441_);
  or _51472_ (_00443_, word_in[96], \oc8051_gm_cxrom_1.cell12.valid );
  or _51473_ (_00444_, \oc8051_gm_cxrom_1.cell12.data [0], _00438_);
  nand _51474_ (_00445_, _00444_, _00443_);
  nand _51475_ (_00446_, _00445_, _42882_);
  or _51476_ (_00447_, \oc8051_gm_cxrom_1.cell12.data [0], _42882_);
  and _51477_ (_05737_, _00447_, _00446_);
  or _51478_ (_00448_, word_in[97], \oc8051_gm_cxrom_1.cell12.valid );
  or _51479_ (_00449_, \oc8051_gm_cxrom_1.cell12.data [1], _00438_);
  nand _51480_ (_00450_, _00449_, _00448_);
  nand _51481_ (_00451_, _00450_, _42882_);
  or _51482_ (_00452_, \oc8051_gm_cxrom_1.cell12.data [1], _42882_);
  and _51483_ (_05741_, _00452_, _00451_);
  or _51484_ (_00453_, word_in[98], \oc8051_gm_cxrom_1.cell12.valid );
  or _51485_ (_00454_, \oc8051_gm_cxrom_1.cell12.data [2], _00438_);
  nand _51486_ (_00455_, _00454_, _00453_);
  nand _51487_ (_00456_, _00455_, _42882_);
  or _51488_ (_00457_, \oc8051_gm_cxrom_1.cell12.data [2], _42882_);
  and _51489_ (_05745_, _00457_, _00456_);
  or _51490_ (_00458_, word_in[99], \oc8051_gm_cxrom_1.cell12.valid );
  or _51491_ (_00459_, \oc8051_gm_cxrom_1.cell12.data [3], _00438_);
  nand _51492_ (_00460_, _00459_, _00458_);
  nand _51493_ (_00461_, _00460_, _42882_);
  or _51494_ (_00462_, \oc8051_gm_cxrom_1.cell12.data [3], _42882_);
  and _51495_ (_05749_, _00462_, _00461_);
  or _51496_ (_00463_, word_in[100], \oc8051_gm_cxrom_1.cell12.valid );
  or _51497_ (_00464_, \oc8051_gm_cxrom_1.cell12.data [4], _00438_);
  nand _51498_ (_00465_, _00464_, _00463_);
  nand _51499_ (_00466_, _00465_, _42882_);
  or _51500_ (_00467_, \oc8051_gm_cxrom_1.cell12.data [4], _42882_);
  and _51501_ (_05753_, _00467_, _00466_);
  nor _51502_ (_00468_, word_in[101], \oc8051_gm_cxrom_1.cell12.valid );
  nor _51503_ (_00469_, \oc8051_gm_cxrom_1.cell12.data [5], _00438_);
  or _51504_ (_00470_, _00469_, _00468_);
  nand _51505_ (_00471_, _00470_, _42882_);
  or _51506_ (_00472_, \oc8051_gm_cxrom_1.cell12.data [5], _42882_);
  and _51507_ (_05757_, _00472_, _00471_);
  or _51508_ (_00473_, word_in[102], \oc8051_gm_cxrom_1.cell12.valid );
  or _51509_ (_00474_, \oc8051_gm_cxrom_1.cell12.data [6], _00438_);
  nand _51510_ (_00475_, _00474_, _00473_);
  nand _51511_ (_00476_, _00475_, _42882_);
  or _51512_ (_00477_, \oc8051_gm_cxrom_1.cell12.data [6], _42882_);
  and _51513_ (_05761_, _00477_, _00476_);
  or _51514_ (_00478_, \oc8051_gm_cxrom_1.cell13.valid , word_in[111]);
  not _51515_ (_00479_, \oc8051_gm_cxrom_1.cell13.valid );
  or _51516_ (_00480_, _00479_, \oc8051_gm_cxrom_1.cell13.data [7]);
  nand _51517_ (_00481_, _00480_, _00478_);
  nand _51518_ (_00482_, _00481_, _42882_);
  or _51519_ (_00483_, \oc8051_gm_cxrom_1.cell13.data [7], _42882_);
  and _51520_ (_05783_, _00483_, _00482_);
  or _51521_ (_00484_, word_in[104], \oc8051_gm_cxrom_1.cell13.valid );
  or _51522_ (_00485_, \oc8051_gm_cxrom_1.cell13.data [0], _00479_);
  nand _51523_ (_00486_, _00485_, _00484_);
  nand _51524_ (_00487_, _00486_, _42882_);
  or _51525_ (_00488_, \oc8051_gm_cxrom_1.cell13.data [0], _42882_);
  and _51526_ (_05790_, _00488_, _00487_);
  or _51527_ (_00489_, word_in[105], \oc8051_gm_cxrom_1.cell13.valid );
  or _51528_ (_00490_, \oc8051_gm_cxrom_1.cell13.data [1], _00479_);
  nand _51529_ (_00491_, _00490_, _00489_);
  nand _51530_ (_00492_, _00491_, _42882_);
  or _51531_ (_00493_, \oc8051_gm_cxrom_1.cell13.data [1], _42882_);
  and _51532_ (_05794_, _00493_, _00492_);
  or _51533_ (_00494_, word_in[106], \oc8051_gm_cxrom_1.cell13.valid );
  or _51534_ (_00495_, \oc8051_gm_cxrom_1.cell13.data [2], _00479_);
  nand _51535_ (_00496_, _00495_, _00494_);
  nand _51536_ (_00497_, _00496_, _42882_);
  or _51537_ (_00498_, \oc8051_gm_cxrom_1.cell13.data [2], _42882_);
  and _51538_ (_05798_, _00498_, _00497_);
  or _51539_ (_00499_, word_in[107], \oc8051_gm_cxrom_1.cell13.valid );
  or _51540_ (_00500_, \oc8051_gm_cxrom_1.cell13.data [3], _00479_);
  nand _51541_ (_00501_, _00500_, _00499_);
  nand _51542_ (_00502_, _00501_, _42882_);
  or _51543_ (_00503_, \oc8051_gm_cxrom_1.cell13.data [3], _42882_);
  and _51544_ (_05802_, _00503_, _00502_);
  or _51545_ (_00504_, word_in[108], \oc8051_gm_cxrom_1.cell13.valid );
  or _51546_ (_00505_, \oc8051_gm_cxrom_1.cell13.data [4], _00479_);
  nand _51547_ (_00506_, _00505_, _00504_);
  nand _51548_ (_00507_, _00506_, _42882_);
  or _51549_ (_00508_, \oc8051_gm_cxrom_1.cell13.data [4], _42882_);
  and _51550_ (_05806_, _00508_, _00507_);
  nor _51551_ (_00509_, word_in[109], \oc8051_gm_cxrom_1.cell13.valid );
  nor _51552_ (_00510_, \oc8051_gm_cxrom_1.cell13.data [5], _00479_);
  or _51553_ (_00511_, _00510_, _00509_);
  nand _51554_ (_00512_, _00511_, _42882_);
  or _51555_ (_00513_, \oc8051_gm_cxrom_1.cell13.data [5], _42882_);
  and _51556_ (_05810_, _00513_, _00512_);
  or _51557_ (_00514_, word_in[110], \oc8051_gm_cxrom_1.cell13.valid );
  or _51558_ (_00515_, \oc8051_gm_cxrom_1.cell13.data [6], _00479_);
  nand _51559_ (_00516_, _00515_, _00514_);
  nand _51560_ (_00517_, _00516_, _42882_);
  or _51561_ (_00518_, \oc8051_gm_cxrom_1.cell13.data [6], _42882_);
  and _51562_ (_05814_, _00518_, _00517_);
  or _51563_ (_00519_, \oc8051_gm_cxrom_1.cell14.valid , word_in[119]);
  not _51564_ (_00520_, \oc8051_gm_cxrom_1.cell14.valid );
  or _51565_ (_00521_, _00520_, \oc8051_gm_cxrom_1.cell14.data [7]);
  nand _51566_ (_00522_, _00521_, _00519_);
  nand _51567_ (_00523_, _00522_, _42882_);
  or _51568_ (_00524_, \oc8051_gm_cxrom_1.cell14.data [7], _42882_);
  and _51569_ (_05836_, _00524_, _00523_);
  or _51570_ (_00525_, word_in[112], \oc8051_gm_cxrom_1.cell14.valid );
  or _51571_ (_00526_, \oc8051_gm_cxrom_1.cell14.data [0], _00520_);
  nand _51572_ (_00527_, _00526_, _00525_);
  nand _51573_ (_00528_, _00527_, _42882_);
  or _51574_ (_00529_, \oc8051_gm_cxrom_1.cell14.data [0], _42882_);
  and _51575_ (_05843_, _00529_, _00528_);
  or _51576_ (_00530_, word_in[113], \oc8051_gm_cxrom_1.cell14.valid );
  or _51577_ (_00531_, \oc8051_gm_cxrom_1.cell14.data [1], _00520_);
  nand _51578_ (_00532_, _00531_, _00530_);
  nand _51579_ (_00533_, _00532_, _42882_);
  or _51580_ (_00534_, \oc8051_gm_cxrom_1.cell14.data [1], _42882_);
  and _51581_ (_05847_, _00534_, _00533_);
  or _51582_ (_00535_, word_in[114], \oc8051_gm_cxrom_1.cell14.valid );
  or _51583_ (_00536_, \oc8051_gm_cxrom_1.cell14.data [2], _00520_);
  nand _51584_ (_00537_, _00536_, _00535_);
  nand _51585_ (_00538_, _00537_, _42882_);
  or _51586_ (_00539_, \oc8051_gm_cxrom_1.cell14.data [2], _42882_);
  and _51587_ (_05851_, _00539_, _00538_);
  or _51588_ (_00540_, word_in[115], \oc8051_gm_cxrom_1.cell14.valid );
  or _51589_ (_00541_, \oc8051_gm_cxrom_1.cell14.data [3], _00520_);
  nand _51590_ (_00542_, _00541_, _00540_);
  nand _51591_ (_00544_, _00542_, _42882_);
  or _51592_ (_00545_, \oc8051_gm_cxrom_1.cell14.data [3], _42882_);
  and _51593_ (_05855_, _00545_, _00544_);
  or _51594_ (_00547_, word_in[116], \oc8051_gm_cxrom_1.cell14.valid );
  or _51595_ (_00549_, \oc8051_gm_cxrom_1.cell14.data [4], _00520_);
  nand _51596_ (_00550_, _00549_, _00547_);
  nand _51597_ (_00552_, _00550_, _42882_);
  or _51598_ (_00553_, \oc8051_gm_cxrom_1.cell14.data [4], _42882_);
  and _51599_ (_05859_, _00553_, _00552_);
  nor _51600_ (_00555_, word_in[117], \oc8051_gm_cxrom_1.cell14.valid );
  nor _51601_ (_00557_, \oc8051_gm_cxrom_1.cell14.data [5], _00520_);
  or _51602_ (_00558_, _00557_, _00555_);
  nand _51603_ (_00560_, _00558_, _42882_);
  or _51604_ (_00561_, \oc8051_gm_cxrom_1.cell14.data [5], _42882_);
  and _51605_ (_05863_, _00561_, _00560_);
  or _51606_ (_00563_, word_in[118], \oc8051_gm_cxrom_1.cell14.valid );
  or _51607_ (_00565_, \oc8051_gm_cxrom_1.cell14.data [6], _00520_);
  nand _51608_ (_00566_, _00565_, _00563_);
  nand _51609_ (_00568_, _00566_, _42882_);
  or _51610_ (_00569_, \oc8051_gm_cxrom_1.cell14.data [6], _42882_);
  and _51611_ (_05867_, _00569_, _00568_);
  or _51612_ (_00571_, \oc8051_gm_cxrom_1.cell15.valid , word_in[127]);
  not _51613_ (_00573_, \oc8051_gm_cxrom_1.cell15.valid );
  or _51614_ (_00574_, _00573_, \oc8051_gm_cxrom_1.cell15.data [7]);
  nand _51615_ (_00576_, _00574_, _00571_);
  nand _51616_ (_00577_, _00576_, _42882_);
  or _51617_ (_00579_, \oc8051_gm_cxrom_1.cell15.data [7], _42882_);
  and _51618_ (_05889_, _00579_, _00577_);
  or _51619_ (_00581_, word_in[120], \oc8051_gm_cxrom_1.cell15.valid );
  or _51620_ (_00582_, \oc8051_gm_cxrom_1.cell15.data [0], _00573_);
  nand _51621_ (_00584_, _00582_, _00581_);
  nand _51622_ (_00585_, _00584_, _42882_);
  or _51623_ (_00587_, \oc8051_gm_cxrom_1.cell15.data [0], _42882_);
  and _51624_ (_05896_, _00587_, _00585_);
  or _51625_ (_00589_, word_in[121], \oc8051_gm_cxrom_1.cell15.valid );
  or _51626_ (_00590_, \oc8051_gm_cxrom_1.cell15.data [1], _00573_);
  nand _51627_ (_00592_, _00590_, _00589_);
  nand _51628_ (_00593_, _00592_, _42882_);
  or _51629_ (_00594_, \oc8051_gm_cxrom_1.cell15.data [1], _42882_);
  and _51630_ (_05900_, _00594_, _00593_);
  or _51631_ (_00595_, word_in[122], \oc8051_gm_cxrom_1.cell15.valid );
  or _51632_ (_00596_, \oc8051_gm_cxrom_1.cell15.data [2], _00573_);
  nand _51633_ (_00597_, _00596_, _00595_);
  nand _51634_ (_00598_, _00597_, _42882_);
  or _51635_ (_00599_, \oc8051_gm_cxrom_1.cell15.data [2], _42882_);
  and _51636_ (_05904_, _00599_, _00598_);
  or _51637_ (_00600_, word_in[123], \oc8051_gm_cxrom_1.cell15.valid );
  or _51638_ (_00601_, \oc8051_gm_cxrom_1.cell15.data [3], _00573_);
  nand _51639_ (_00602_, _00601_, _00600_);
  nand _51640_ (_00603_, _00602_, _42882_);
  or _51641_ (_00604_, \oc8051_gm_cxrom_1.cell15.data [3], _42882_);
  and _51642_ (_05908_, _00604_, _00603_);
  or _51643_ (_00605_, word_in[124], \oc8051_gm_cxrom_1.cell15.valid );
  or _51644_ (_00606_, \oc8051_gm_cxrom_1.cell15.data [4], _00573_);
  nand _51645_ (_00607_, _00606_, _00605_);
  nand _51646_ (_00608_, _00607_, _42882_);
  or _51647_ (_00609_, \oc8051_gm_cxrom_1.cell15.data [4], _42882_);
  and _51648_ (_05912_, _00609_, _00608_);
  nor _51649_ (_00610_, word_in[125], \oc8051_gm_cxrom_1.cell15.valid );
  nor _51650_ (_00611_, \oc8051_gm_cxrom_1.cell15.data [5], _00573_);
  or _51651_ (_00612_, _00611_, _00610_);
  nand _51652_ (_00613_, _00612_, _42882_);
  or _51653_ (_00614_, \oc8051_gm_cxrom_1.cell15.data [5], _42882_);
  and _51654_ (_05916_, _00614_, _00613_);
  or _51655_ (_00615_, word_in[126], \oc8051_gm_cxrom_1.cell15.valid );
  or _51656_ (_00616_, \oc8051_gm_cxrom_1.cell15.data [6], _00573_);
  nand _51657_ (_00617_, _00616_, _00615_);
  nand _51658_ (_00618_, _00617_, _42882_);
  or _51659_ (_00619_, \oc8051_gm_cxrom_1.cell15.data [6], _42882_);
  and _51660_ (_05920_, _00619_, _00618_);
  nor _51661_ (_09695_, _38255_, rst);
  and _51662_ (_00620_, _38246_, _38280_);
  and _51663_ (_00621_, _00620_, _36920_);
  not _51664_ (_00622_, _00621_);
  and _51665_ (_00623_, _38218_, _38226_);
  and _51666_ (_00624_, _38281_, _38217_);
  nor _51667_ (_00625_, _00624_, _00623_);
  and _51668_ (_00626_, _00625_, _00622_);
  and _51669_ (_00627_, _38280_, _36909_);
  or _51670_ (_00628_, _38246_, _38217_);
  nand _51671_ (_00629_, _00628_, _00627_);
  and _51672_ (_00630_, _00629_, _00626_);
  and _51673_ (_00631_, _36450_, _42882_);
  not _51674_ (_00632_, _00631_);
  or _51675_ (_00633_, _00632_, _00623_);
  or _51676_ (_09698_, _00633_, _00630_);
  not _51677_ (_00634_, _37117_);
  and _51678_ (_00635_, _37357_, _00634_);
  and _51679_ (_00636_, _00635_, _37630_);
  not _51680_ (_00637_, _37905_);
  and _51681_ (_00638_, _38210_, _38145_);
  and _51682_ (_00639_, _00638_, _38185_);
  and _51683_ (_00640_, _00639_, _00637_);
  and _51684_ (_00641_, _00640_, _00636_);
  not _51685_ (_00642_, _36844_);
  nor _51686_ (_00643_, _38210_, _00642_);
  nor _51687_ (_00644_, _37357_, _37117_);
  and _51688_ (_00645_, _00644_, _37630_);
  and _51689_ (_00646_, _00645_, _00643_);
  not _51690_ (_00647_, _38185_);
  not _51691_ (_00648_, _38145_);
  and _51692_ (_00649_, _38210_, _00648_);
  and _51693_ (_00650_, _00649_, _00647_);
  nor _51694_ (_00651_, _37630_, _00642_);
  and _51695_ (_00652_, _00651_, _00635_);
  and _51696_ (_00653_, _00652_, _00650_);
  or _51697_ (_00654_, _00653_, _00646_);
  or _51698_ (_00655_, _00654_, _00641_);
  not _51699_ (_00656_, _37357_);
  and _51700_ (_00657_, _00656_, _37117_);
  and _51701_ (_00658_, _00657_, _00651_);
  and _51702_ (_00659_, _00658_, _00640_);
  and _51703_ (_00660_, _00639_, _37905_);
  and _51704_ (_00661_, _37357_, _37117_);
  and _51705_ (_00662_, _00661_, _37630_);
  and _51706_ (_00663_, _00662_, _00660_);
  or _51707_ (_00664_, _00663_, _00659_);
  or _51708_ (_00665_, _00664_, _00655_);
  and _51709_ (_00666_, _37905_, _00647_);
  and _51710_ (_00667_, _00666_, _00638_);
  and _51711_ (_00668_, _00667_, _00661_);
  and _51712_ (_00669_, _37630_, _00642_);
  nor _51713_ (_00670_, _00669_, _00651_);
  and _51714_ (_00671_, _00670_, _00668_);
  and _51715_ (_00672_, _00667_, _36844_);
  and _51716_ (_00673_, _00672_, _00657_);
  or _51717_ (_00674_, _00673_, _00671_);
  or _51718_ (_00675_, _00674_, _00665_);
  and _51719_ (_00676_, _00638_, _00647_);
  not _51720_ (_00677_, _00676_);
  nor _51721_ (_00678_, _37630_, _36844_);
  and _51722_ (_00679_, _00678_, _00657_);
  nor _51723_ (_00680_, _00679_, _00637_);
  nor _51724_ (_00681_, _00680_, _00677_);
  not _51725_ (_00682_, _00681_);
  and _51726_ (_00683_, _00669_, _00657_);
  and _51727_ (_00684_, _00683_, _00667_);
  and _51728_ (_00685_, _00661_, _00651_);
  and _51729_ (_00686_, _00685_, _00667_);
  nor _51730_ (_00687_, _00686_, _00684_);
  and _51731_ (_00688_, _00687_, _00682_);
  not _51732_ (_00689_, _37630_);
  and _51733_ (_00690_, _00644_, _00689_);
  and _51734_ (_00691_, _00690_, _00639_);
  and _51735_ (_00692_, _00635_, _00689_);
  and _51736_ (_00693_, _38185_, _36844_);
  and _51737_ (_00694_, _00693_, _00649_);
  and _51738_ (_00695_, _00694_, _00692_);
  nor _51739_ (_00696_, _37630_, _00656_);
  and _51740_ (_00697_, _00696_, _00643_);
  and _51741_ (_00698_, _00697_, _00634_);
  or _51742_ (_00699_, _00698_, _00695_);
  and _51743_ (_00700_, _00690_, _00667_);
  or _51744_ (_00701_, _00700_, _00699_);
  or _51745_ (_00702_, _00701_, _00691_);
  and _51746_ (_00703_, _00666_, _00649_);
  and _51747_ (_00704_, _00703_, _00642_);
  and _51748_ (_00705_, _00704_, _00635_);
  and _51749_ (_00706_, _37630_, _36844_);
  and _51750_ (_00707_, _00706_, _00644_);
  and _51751_ (_00708_, _00650_, _00637_);
  and _51752_ (_00709_, _00708_, _00707_);
  or _51753_ (_00710_, _00709_, _00705_);
  and _51754_ (_00711_, _00669_, _00635_);
  and _51755_ (_00712_, _00711_, _00667_);
  and _51756_ (_00713_, _00661_, _00689_);
  and _51757_ (_00714_, _00713_, _00660_);
  or _51758_ (_00715_, _00714_, _00712_);
  or _51759_ (_00716_, _00715_, _00710_);
  nor _51760_ (_00717_, _00716_, _00702_);
  nand _51761_ (_00718_, _00717_, _00688_);
  or _51762_ (_00719_, _00718_, _00675_);
  and _51763_ (_00720_, _00719_, _36461_);
  not _51764_ (_00721_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _51765_ (_00722_, _36439_, _18199_);
  and _51766_ (_00723_, _00722_, _38241_);
  nor _51767_ (_00724_, _00723_, _00721_);
  or _51768_ (_00725_, _00724_, rst);
  or _51769_ (_09701_, _00725_, _00720_);
  nand _51770_ (_00726_, _37117_, _36385_);
  or _51771_ (_00727_, _36385_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _51772_ (_00728_, _00727_, _42882_);
  and _51773_ (_09704_, _00728_, _00726_);
  and _51774_ (_00729_, \oc8051_top_1.oc8051_sfr1.wait_data , _42882_);
  and _51775_ (_00730_, _00729_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _51776_ (_00731_, _38246_, _38232_);
  or _51777_ (_00732_, _00731_, _38247_);
  or _51778_ (_00733_, _00732_, _38316_);
  and _51779_ (_00734_, _38218_, _38289_);
  or _51780_ (_00735_, _00734_, _38266_);
  or _51781_ (_00736_, _00735_, _00733_);
  and _51782_ (_00737_, _38235_, _38281_);
  and _51783_ (_00738_, _00623_, _36920_);
  nor _51784_ (_00739_, _00738_, _00737_);
  nand _51785_ (_00740_, _00739_, _38341_);
  or _51786_ (_00741_, _00740_, _00736_);
  and _51787_ (_00742_, _00741_, _00631_);
  or _51788_ (_09707_, _00742_, _00730_);
  and _51789_ (_00743_, _38233_, _38191_);
  and _51790_ (_00744_, _00743_, _38289_);
  and _51791_ (_00745_, _38215_, _36920_);
  and _51792_ (_00746_, _00745_, _38264_);
  or _51793_ (_00747_, _00746_, _38360_);
  and _51794_ (_00748_, _38246_, _38227_);
  or _51795_ (_00749_, _00748_, _38219_);
  or _51796_ (_00750_, _00749_, _00747_);
  or _51797_ (_00751_, _00750_, _00744_);
  and _51798_ (_00752_, _00751_, _36450_);
  and _51799_ (_00753_, _38350_, _00721_);
  not _51800_ (_00754_, _38238_);
  and _51801_ (_00755_, _00754_, _00753_);
  and _51802_ (_00756_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _51803_ (_00757_, _00756_, _00755_);
  or _51804_ (_00758_, _00757_, _00752_);
  and _51805_ (_09710_, _00758_, _42882_);
  and _51806_ (_00759_, _00729_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _51807_ (_00760_, _38235_, _38299_);
  or _51808_ (_00761_, _38299_, _38265_);
  and _51809_ (_00762_, _00761_, _38275_);
  or _51810_ (_00763_, _00762_, _00760_);
  and _51811_ (_00764_, _00743_, _38307_);
  or _51812_ (_00765_, _00764_, _00763_);
  and _51813_ (_00766_, _00761_, _38215_);
  and _51814_ (_00767_, _38215_, _36909_);
  and _51815_ (_00768_, _00767_, _38298_);
  or _51816_ (_00769_, _00768_, _00766_);
  or _51817_ (_00770_, _00769_, _38368_);
  and _51818_ (_00771_, _38235_, _38283_);
  and _51819_ (_00772_, _38317_, _38215_);
  or _51820_ (_00773_, _00772_, _00771_);
  or _51821_ (_00774_, _00773_, _00749_);
  or _51822_ (_00775_, _00774_, _00770_);
  or _51823_ (_00776_, _00775_, _00765_);
  and _51824_ (_00777_, _00776_, _00631_);
  or _51825_ (_09713_, _00777_, _00759_);
  and _51826_ (_00778_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _51827_ (_00779_, _38276_, _36450_);
  or _51828_ (_00780_, _00779_, _00778_);
  or _51829_ (_00781_, _00780_, _00755_);
  and _51830_ (_09716_, _00781_, _42882_);
  and _51831_ (_00782_, _38307_, _38260_);
  and _51832_ (_00783_, _38274_, _38245_);
  and _51833_ (_00784_, _00783_, _36909_);
  or _51834_ (_00785_, _00784_, _00782_);
  and _51835_ (_00786_, _00785_, _38243_);
  or _51836_ (_00787_, _00786_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _51837_ (_00788_, _00785_, _00738_);
  and _51838_ (_00789_, _00788_, _36396_);
  and _51839_ (_00790_, _38280_, _38192_);
  and _51840_ (_00791_, _00790_, _38270_);
  and _51841_ (_00792_, _38226_, _38375_);
  and _51842_ (_00793_, _38246_, _38281_);
  or _51843_ (_00794_, _00793_, _00792_);
  or _51844_ (_00795_, _00794_, _00791_);
  and _51845_ (_00796_, _00795_, _00753_);
  or _51846_ (_00797_, _00796_, _00789_);
  or _51847_ (_00798_, _00797_, _00787_);
  or _51848_ (_00799_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _18199_);
  and _51849_ (_00800_, _00799_, _42882_);
  and _51850_ (_09719_, _00800_, _00798_);
  and _51851_ (_00801_, _00729_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or _51852_ (_00802_, _00746_, _38290_);
  or _51853_ (_00803_, _38307_, _38289_);
  and _51854_ (_00804_, _00803_, _38359_);
  or _51855_ (_00805_, _00804_, _38266_);
  or _51856_ (_00806_, _00805_, _00802_);
  and _51857_ (_00807_, _38235_, _38307_);
  or _51858_ (_00808_, _00807_, _38308_);
  and _51859_ (_00809_, _00767_, _38264_);
  or _51860_ (_00810_, _00768_, _00809_);
  or _51861_ (_00811_, _38376_, _38306_);
  or _51862_ (_00812_, _00811_, _00810_);
  or _51863_ (_00813_, _00812_, _00808_);
  or _51864_ (_00814_, _38318_, _38261_);
  or _51865_ (_00815_, _00814_, _00813_);
  or _51866_ (_00816_, _00815_, _00806_);
  and _51867_ (_00817_, _00816_, _00631_);
  or _51868_ (_09722_, _00817_, _00801_);
  and _51869_ (_00818_, _00729_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _51870_ (_00819_, _00743_, _38287_);
  and _51871_ (_00820_, _38218_, _38294_);
  or _51872_ (_00821_, _00820_, _00744_);
  or _51873_ (_00822_, _00821_, _00819_);
  or _51874_ (_00823_, _00822_, _00769_);
  not _51875_ (_00824_, _38322_);
  and _51876_ (_00825_, _38235_, _38312_);
  or _51877_ (_00826_, _00825_, _00824_);
  and _51878_ (_00827_, _38271_, _38263_);
  or _51879_ (_00828_, _00827_, _38386_);
  and _51880_ (_00829_, _38359_, _38265_);
  or _51881_ (_00830_, _00829_, _00828_);
  or _51882_ (_00831_, _00830_, _00826_);
  or _51883_ (_00832_, _00831_, _00823_);
  and _51884_ (_00833_, _00745_, _38263_);
  and _51885_ (_00834_, _00745_, _38222_);
  or _51886_ (_00835_, _00834_, _00833_);
  nor _51887_ (_00836_, _38366_, _38343_);
  nand _51888_ (_00837_, _00836_, _38314_);
  or _51889_ (_00838_, _00837_, _00835_);
  or _51890_ (_00839_, _00838_, _00765_);
  or _51891_ (_00840_, _00839_, _00832_);
  and _51892_ (_00841_, _00840_, _00631_);
  or _51893_ (_09725_, _00841_, _00818_);
  and _51894_ (_00842_, _00743_, _38295_);
  or _51895_ (_00843_, _00842_, _38363_);
  and _51896_ (_00844_, _00767_, _38225_);
  and _51897_ (_00845_, _00844_, _37171_);
  or _51898_ (_00846_, _00845_, _38370_);
  and _51899_ (_00847_, _38295_, _38215_);
  or _51900_ (_00848_, _00847_, _00846_);
  or _51901_ (_00849_, _00848_, _00843_);
  and _51902_ (_00850_, _00743_, _38227_);
  or _51903_ (_00851_, _00850_, _00849_);
  and _51904_ (_00852_, _00851_, _36450_);
  nand _51905_ (_00853_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand _51906_ (_00854_, _00853_, _38251_);
  or _51907_ (_00855_, _00854_, _00852_);
  and _51908_ (_09728_, _00855_, _42882_);
  nand _51909_ (_00856_, _38344_, _38319_);
  or _51910_ (_00857_, _00856_, _00762_);
  or _51911_ (_00858_, _38290_, _38267_);
  and _51912_ (_00859_, _38221_, _36909_);
  and _51913_ (_00860_, _00859_, _38275_);
  or _51914_ (_00861_, _00860_, _38308_);
  or _51915_ (_00862_, _00861_, _00782_);
  or _51916_ (_00863_, _38321_, _38278_);
  or _51917_ (_00864_, _00863_, _00862_);
  or _51918_ (_00865_, _00864_, _00858_);
  or _51919_ (_00866_, _00865_, _00857_);
  and _51920_ (_00867_, _00745_, _38226_);
  or _51921_ (_00868_, _00867_, _38292_);
  or _51922_ (_00869_, _00868_, _00784_);
  and _51923_ (_00870_, _00767_, _38221_);
  or _51924_ (_00871_, _00870_, _38381_);
  or _51925_ (_00872_, _00871_, _38327_);
  or _51926_ (_00873_, _00872_, _00869_);
  and _51927_ (_00874_, _38359_, _37707_);
  and _51928_ (_00875_, _38362_, _38221_);
  or _51929_ (_00876_, _00875_, _38366_);
  or _51930_ (_00877_, _00876_, _00874_);
  or _51931_ (_00878_, _00877_, _00747_);
  or _51932_ (_00879_, _00878_, _00873_);
  or _51933_ (_00880_, _00879_, _00769_);
  or _51934_ (_00881_, _00880_, _00866_);
  and _51935_ (_00882_, _00881_, _36450_);
  and _51936_ (_00883_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or _51937_ (_00884_, _00786_, _00755_);
  and _51938_ (_00885_, _38243_, _38339_);
  or _51939_ (_00886_, _00885_, _00884_);
  or _51940_ (_00887_, _00886_, _00883_);
  or _51941_ (_00888_, _00887_, _00882_);
  and _51942_ (_09731_, _00888_, _42882_);
  nor _51943_ (_09790_, _38396_, rst);
  nor _51944_ (_09792_, _38355_, rst);
  or _51945_ (_09795_, _00632_, _00626_);
  nor _51946_ (_00889_, _00623_, _00620_);
  or _51947_ (_09798_, _00889_, _00632_);
  or _51948_ (_00890_, _00714_, _00705_);
  or _51949_ (_00891_, _00641_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _51950_ (_00892_, _00891_, _00890_);
  and _51951_ (_00893_, _00892_, _00723_);
  nor _51952_ (_00894_, _00722_, _38241_);
  or _51953_ (_00895_, _00894_, rst);
  or _51954_ (_09801_, _00895_, _00893_);
  nand _51955_ (_00896_, _37905_, _36385_);
  or _51956_ (_00897_, _36385_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _51957_ (_00898_, _00897_, _42882_);
  and _51958_ (_09804_, _00898_, _00896_);
  not _51959_ (_00899_, _36385_);
  or _51960_ (_00900_, _38185_, _00899_);
  or _51961_ (_00901_, _36385_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _51962_ (_00902_, _00901_, _42882_);
  and _51963_ (_09807_, _00902_, _00900_);
  nand _51964_ (_00903_, _38145_, _36385_);
  or _51965_ (_00904_, _36385_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _51966_ (_00905_, _00904_, _42882_);
  and _51967_ (_09810_, _00905_, _00903_);
  nand _51968_ (_00906_, _38210_, _36385_);
  or _51969_ (_00907_, _36385_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _51970_ (_00908_, _00907_, _42882_);
  and _51971_ (_09813_, _00908_, _00906_);
  or _51972_ (_00909_, _36844_, _00899_);
  or _51973_ (_00910_, _36385_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _51974_ (_00911_, _00910_, _42882_);
  and _51975_ (_09816_, _00911_, _00909_);
  nand _51976_ (_00912_, _37630_, _36385_);
  or _51977_ (_00913_, _36385_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _51978_ (_00914_, _00913_, _42882_);
  and _51979_ (_09819_, _00914_, _00912_);
  nand _51980_ (_00915_, _37357_, _36385_);
  or _51981_ (_00916_, _36385_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _51982_ (_00917_, _00916_, _42882_);
  and _51983_ (_09822_, _00917_, _00915_);
  and _51984_ (_00918_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _51985_ (_00919_, _00918_, _00796_);
  and _51986_ (_00920_, _00919_, _42882_);
  and _51987_ (_00921_, _38311_, _38215_);
  and _51988_ (_00922_, _00921_, _36909_);
  or _51989_ (_00923_, _00922_, _00847_);
  and _51990_ (_00924_, _00743_, _38312_);
  or _51991_ (_00926_, _00924_, _00748_);
  or _51992_ (_00927_, _00926_, _00923_);
  or _51993_ (_00928_, _38295_, _38281_);
  and _51994_ (_00929_, _00928_, _00743_);
  or _51995_ (_00930_, _38298_, _38265_);
  and _51996_ (_00931_, _00930_, _38235_);
  or _51997_ (_00932_, _00931_, _00929_);
  or _51998_ (_00933_, _00932_, _00927_);
  and _51999_ (_00934_, _00743_, _38326_);
  or _52000_ (_00935_, _38311_, _38280_);
  and _52001_ (_00936_, _00935_, _00745_);
  or _52002_ (_00937_, _00936_, _00934_);
  and _52003_ (_00938_, _38235_, _38223_);
  and _52004_ (_00939_, _00627_, _38235_);
  or _52005_ (_00940_, _00939_, _00938_);
  or _52006_ (_00941_, _00940_, _00937_);
  or _52007_ (_00942_, _00834_, _00819_);
  or _52008_ (_00943_, _00846_, _38369_);
  or _52009_ (_00944_, _00943_, _00942_);
  and _52010_ (_00945_, _38227_, _38359_);
  or _52011_ (_00946_, _00945_, _38219_);
  or _52012_ (_00947_, _00850_, _00820_);
  or _52013_ (_00948_, _00947_, _00946_);
  and _52014_ (_00949_, _00935_, _38271_);
  and _52015_ (_00950_, _38287_, _38359_);
  or _52016_ (_00951_, _00950_, _00949_);
  or _52017_ (_00952_, _00951_, _00948_);
  or _52018_ (_00953_, _00952_, _00944_);
  or _52019_ (_00954_, _00953_, _00941_);
  or _52020_ (_00955_, _00954_, _00933_);
  and _52021_ (_00957_, _00955_, _00631_);
  or _52022_ (_09825_, _00957_, _00920_);
  and _52023_ (_00958_, _00729_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _52024_ (_00959_, _00926_, _00835_);
  or _52025_ (_00960_, _38312_, _38287_);
  and _52026_ (_00961_, _00960_, _38260_);
  and _52027_ (_00962_, _38235_, _38331_);
  or _52028_ (_00963_, _00962_, _00961_);
  or _52029_ (_00964_, _00963_, _00959_);
  and _52030_ (_00965_, _38235_, _38287_);
  and _52031_ (_00966_, _37685_, _37421_);
  and _52032_ (_00967_, _00767_, _00966_);
  and _52033_ (_00968_, _00967_, _37171_);
  nor _52034_ (_00969_, _00968_, _38365_);
  not _52035_ (_00970_, _00969_);
  or _52036_ (_00971_, _00970_, _00771_);
  or _52037_ (_00972_, _00971_, _00965_);
  nand _52038_ (_00973_, _00739_, _38291_);
  or _52039_ (_00974_, _00973_, _00972_);
  or _52040_ (_00975_, _00974_, _00830_);
  or _52041_ (_00977_, _00975_, _00964_);
  and _52042_ (_00978_, _00977_, _00631_);
  or _52043_ (_34273_, _00978_, _00958_);
  or _52044_ (_00979_, _00784_, _38327_);
  or _52045_ (_00980_, _00867_, _38381_);
  or _52046_ (_00981_, _00980_, _00866_);
  or _52047_ (_00982_, _00981_, _00979_);
  and _52048_ (_00983_, _00982_, _36450_);
  and _52049_ (_00984_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52050_ (_00985_, _00984_, _00886_);
  or _52051_ (_00986_, _00985_, _00983_);
  and _52052_ (_34275_, _00986_, _42882_);
  and _52053_ (_00987_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52054_ (_00988_, _00987_, _00884_);
  and _52055_ (_00989_, _00988_, _42882_);
  and _52056_ (_00990_, _38342_, _36920_);
  or _52057_ (_00991_, _00990_, _00785_);
  or _52058_ (_00992_, _00991_, _00877_);
  or _52059_ (_00993_, _00992_, _38360_);
  and _52060_ (_00994_, _00993_, _00631_);
  or _52061_ (_34278_, _00994_, _00989_);
  and _52062_ (_00995_, _00842_, _36909_);
  or _52063_ (_00996_, _00623_, _38237_);
  or _52064_ (_00997_, _00996_, _00934_);
  or _52065_ (_00998_, _00997_, _00995_);
  or _52066_ (_00999_, _00938_, _00825_);
  and _52067_ (_01000_, _00627_, _38275_);
  or _52068_ (_01001_, _01000_, _00965_);
  or _52069_ (_01002_, _01001_, _00999_);
  or _52070_ (_01003_, _01002_, _00998_);
  or _52071_ (_01004_, _00923_, _00820_);
  or _52072_ (_01005_, _01004_, _00943_);
  or _52073_ (_01006_, _01005_, _01003_);
  and _52074_ (_01007_, _00743_, _38317_);
  or _52075_ (_01008_, _01007_, _00850_);
  or _52076_ (_01009_, _01008_, _00737_);
  or _52077_ (_01010_, _01009_, _00939_);
  and _52078_ (_01011_, _38235_, _38289_);
  or _52079_ (_01012_, _01011_, _38236_);
  or _52080_ (_01013_, _01012_, _00931_);
  or _52081_ (_01014_, _01013_, _01010_);
  and _52082_ (_01015_, _00859_, _38359_);
  or _52083_ (_01016_, _00870_, _00945_);
  or _52084_ (_01017_, _01016_, _01015_);
  or _52085_ (_01018_, _01017_, _00785_);
  and _52086_ (_01019_, _38327_, _38262_);
  and _52087_ (_01020_, _00842_, _36920_);
  or _52088_ (_01021_, _01020_, _38224_);
  or _52089_ (_01022_, _01021_, _01019_);
  or _52090_ (_01023_, _01022_, _01018_);
  or _52091_ (_01024_, _01023_, _01014_);
  or _52092_ (_01025_, _01024_, _01006_);
  and _52093_ (_01026_, _01025_, _36450_);
  and _52094_ (_01027_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _52095_ (_01028_, _38238_, _36396_);
  or _52096_ (_01029_, _00796_, _01028_);
  or _52097_ (_01030_, _01029_, _01027_);
  or _52098_ (_01031_, _01030_, _01026_);
  and _52099_ (_34280_, _01031_, _42882_);
  and _52100_ (_01032_, _00627_, _38359_);
  or _52101_ (_01033_, _38237_, _00945_);
  or _52102_ (_01034_, _01033_, _38327_);
  or _52103_ (_01035_, _01034_, _01032_);
  or _52104_ (_01036_, _01035_, _01004_);
  or _52105_ (_01037_, _01036_, _00943_);
  and _52106_ (_01038_, _00767_, _38280_);
  or _52107_ (_01039_, _00860_, _00748_);
  or _52108_ (_01040_, _01039_, _01038_);
  or _52109_ (_01041_, _01040_, _38230_);
  and _52110_ (_01042_, _00960_, _38218_);
  or _52111_ (_01043_, _01042_, _38332_);
  or _52112_ (_01044_, _01043_, _01041_);
  or _52113_ (_01045_, _01044_, _01014_);
  or _52114_ (_01046_, _01045_, _01037_);
  and _52115_ (_01047_, _01046_, _36450_);
  and _52116_ (_01048_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52117_ (_01049_, _01048_, _01029_);
  or _52118_ (_01050_, _01049_, _01047_);
  and _52119_ (_34282_, _01050_, _42882_);
  and _52120_ (_01051_, _00729_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _52121_ (_01052_, _00850_, _42307_);
  or _52122_ (_01053_, _01052_, _00804_);
  or _52123_ (_01054_, _38307_, _38265_);
  and _52124_ (_01055_, _01054_, _38218_);
  and _52125_ (_01056_, _38235_, _38265_);
  or _52126_ (_01057_, _01056_, _00764_);
  or _52127_ (_01058_, _01057_, _01055_);
  or _52128_ (_01059_, _01058_, _01053_);
  or _52129_ (_01060_, _00945_, _38273_);
  or _52130_ (_01061_, _01060_, _00995_);
  or _52131_ (_01062_, _00845_, _00746_);
  and _52132_ (_01063_, _38317_, _38217_);
  and _52133_ (_01064_, _01063_, _37960_);
  or _52134_ (_01065_, _01064_, _01062_);
  or _52135_ (_01066_, _01065_, _01061_);
  and _52136_ (_01067_, _38218_, _38334_);
  and _52137_ (_01068_, _38362_, _38295_);
  and _52138_ (_01069_, _38334_, _38215_);
  or _52139_ (_01070_, _01069_, _01068_);
  nor _52140_ (_01071_, _01070_, _01067_);
  nand _52141_ (_01072_, _01071_, _42311_);
  or _52142_ (_01073_, _01072_, _01066_);
  or _52143_ (_01074_, _00858_, _00812_);
  or _52144_ (_01075_, _01074_, _01073_);
  or _52145_ (_01076_, _01075_, _01059_);
  and _52146_ (_01077_, _01076_, _00631_);
  or _52147_ (_34284_, _01077_, _01051_);
  or _52148_ (_01078_, _00923_, _38329_);
  or _52149_ (_01079_, _01067_, _01056_);
  or _52150_ (_01080_, _01079_, _01021_);
  or _52151_ (_01081_, _01080_, _01078_);
  or _52152_ (_01082_, _00744_, _38313_);
  or _52153_ (_01083_, _00829_, _00827_);
  or _52154_ (_01084_, _01083_, _01082_);
  and _52155_ (_01085_, _38218_, _38307_);
  or _52156_ (_01086_, _00833_, _38219_);
  or _52157_ (_01087_, _01086_, _01085_);
  or _52158_ (_01088_, _01087_, _38371_);
  or _52159_ (_01089_, _01088_, _01084_);
  or _52160_ (_01090_, _00998_, _00826_);
  or _52161_ (_01091_, _01090_, _01089_);
  or _52162_ (_01092_, _01091_, _01081_);
  and _52163_ (_01093_, _01092_, _00631_);
  and _52164_ (_01094_, \oc8051_top_1.oc8051_decoder1.alu_op [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _52165_ (_01095_, _38237_, _36407_);
  or _52166_ (_01096_, _01095_, _01094_);
  and _52167_ (_01097_, _01096_, _42882_);
  or _52168_ (_34286_, _01097_, _01093_);
  and _52169_ (_01098_, _38326_, _38359_);
  or _52170_ (_01099_, _01098_, _00744_);
  or _52171_ (_01100_, _01062_, _00922_);
  or _52172_ (_01101_, _01100_, _01099_);
  and _52173_ (_01102_, _38218_, _38295_);
  or _52174_ (_01103_, _00772_, _01063_);
  or _52175_ (_01104_, _01103_, _01102_);
  not _52176_ (_01105_, _38364_);
  or _52177_ (_01106_, _01105_, _42310_);
  or _52178_ (_01107_, _01106_, _01104_);
  or _52179_ (_01108_, _01107_, _01101_);
  not _52180_ (_01109_, _00934_);
  and _52181_ (_01110_, _01109_, _38328_);
  not _52182_ (_01111_, _01110_);
  or _52183_ (_01112_, _01111_, _01010_);
  or _52184_ (_01113_, _01112_, _01108_);
  or _52185_ (_01114_, _00770_, _00765_);
  or _52186_ (_01115_, _01114_, _01113_);
  and _52187_ (_01116_, _01115_, _36450_);
  and _52188_ (_01117_, \oc8051_top_1.oc8051_decoder1.alu_op [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52189_ (_01118_, _01117_, _38249_);
  or _52190_ (_01119_, _01118_, _01116_);
  and _52191_ (_34288_, _01119_, _42882_);
  and _52192_ (_01120_, _38218_, _38298_);
  or _52193_ (_01121_, _01120_, _01063_);
  or _52194_ (_01122_, _01121_, _38327_);
  or _52195_ (_01123_, _01098_, _42307_);
  or _52196_ (_01124_, _01123_, _01122_);
  or _52197_ (_01125_, _01057_, _00802_);
  or _52198_ (_01126_, _01125_, _01124_);
  or _52199_ (_01127_, _00939_, _00934_);
  or _52200_ (_01128_, _38360_, _38366_);
  or _52201_ (_01129_, _01128_, _00922_);
  or _52202_ (_01130_, _01129_, _01127_);
  or _52203_ (_01131_, _01130_, _00769_);
  or _52204_ (_01132_, _01131_, _00763_);
  or _52205_ (_01133_, _01132_, _01126_);
  and _52206_ (_01134_, _01133_, _36450_);
  and _52207_ (_01135_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _52208_ (_01136_, _01135_, _38250_);
  or _52209_ (_01137_, _01136_, _01134_);
  and _52210_ (_34290_, _01137_, _42882_);
  and _52211_ (_01138_, _00729_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not _52212_ (_01139_, _42311_);
  or _52213_ (_01140_, _01052_, _01139_);
  or _52214_ (_01141_, _01079_, _01055_);
  or _52215_ (_01142_, _01141_, _01140_);
  not _52216_ (_01143_, _38245_);
  or _52217_ (_01144_, _38218_, _01143_);
  and _52218_ (_01145_, _01144_, _38317_);
  or _52219_ (_01146_, _00734_, _38261_);
  or _52220_ (_01147_, _01146_, _01145_);
  or _52221_ (_01148_, _01147_, _00849_);
  or _52222_ (_01149_, _01148_, _01142_);
  and _52223_ (_01150_, _01149_, _00631_);
  or _52224_ (_34292_, _01150_, _01138_);
  nor _52225_ (_38955_, _37117_, rst);
  nor _52226_ (_38956_, _42266_, rst);
  and _52227_ (_01151_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  and _52228_ (_01152_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  and _52229_ (_01153_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _52230_ (_01154_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _52231_ (_01155_, _01154_, _01153_);
  and _52232_ (_01156_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _52233_ (_01157_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _52234_ (_01158_, _01157_, _01156_);
  and _52235_ (_01159_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and _52236_ (_01160_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _52237_ (_01161_, _01160_, _01159_);
  and _52238_ (_01162_, _01161_, _01158_);
  and _52239_ (_01163_, _01162_, _01155_);
  nor _52240_ (_01164_, _01163_, _36636_);
  nor _52241_ (_01165_, _01164_, _01152_);
  nor _52242_ (_01166_, _01165_, _42250_);
  nor _52243_ (_01167_, _01166_, _01151_);
  nor _52244_ (_38958_, _01167_, rst);
  nor _52245_ (_38968_, _37905_, rst);
  and _52246_ (_38969_, _38185_, _42882_);
  nor _52247_ (_38970_, _38145_, rst);
  nor _52248_ (_38971_, _38210_, rst);
  and _52249_ (_38972_, _36844_, _42882_);
  nor _52250_ (_38973_, _37630_, rst);
  nor _52251_ (_38974_, _37357_, rst);
  nor _52252_ (_38975_, _42464_, rst);
  nor _52253_ (_38976_, _42384_, rst);
  nor _52254_ (_38978_, _42589_, rst);
  nor _52255_ (_38979_, _42429_, rst);
  nor _52256_ (_38980_, _42336_, rst);
  nor _52257_ (_38981_, _42551_, rst);
  nor _52258_ (_38982_, _42523_, rst);
  and _52259_ (_01168_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [0]);
  and _52260_ (_01169_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  and _52261_ (_01170_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _52262_ (_01171_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _52263_ (_01172_, _01171_, _01170_);
  and _52264_ (_01173_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _52265_ (_01174_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _52266_ (_01175_, _01174_, _01173_);
  and _52267_ (_01176_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _52268_ (_01177_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _52269_ (_01178_, _01177_, _01176_);
  and _52270_ (_01179_, _01178_, _01175_);
  and _52271_ (_01180_, _01179_, _01172_);
  nor _52272_ (_01181_, _01180_, _36636_);
  nor _52273_ (_01182_, _01181_, _01169_);
  nor _52274_ (_01183_, _01182_, _42250_);
  nor _52275_ (_01184_, _01183_, _01168_);
  nor _52276_ (_38984_, _01184_, rst);
  and _52277_ (_01185_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  and _52278_ (_01186_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  and _52279_ (_01187_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _52280_ (_01188_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _52281_ (_01189_, _01188_, _01187_);
  and _52282_ (_01190_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _52283_ (_01191_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _52284_ (_01192_, _01191_, _01190_);
  and _52285_ (_01193_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and _52286_ (_01194_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _52287_ (_01195_, _01194_, _01193_);
  and _52288_ (_01196_, _01195_, _01192_);
  and _52289_ (_01197_, _01196_, _01189_);
  nor _52290_ (_01198_, _01197_, _36636_);
  nor _52291_ (_01199_, _01198_, _01186_);
  nor _52292_ (_01200_, _01199_, _42250_);
  nor _52293_ (_01201_, _01200_, _01185_);
  nor _52294_ (_38985_, _01201_, rst);
  and _52295_ (_01202_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  and _52296_ (_01203_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  and _52297_ (_01204_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _52298_ (_01205_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _52299_ (_01206_, _01205_, _01204_);
  and _52300_ (_01207_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _52301_ (_01208_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _52302_ (_01209_, _01208_, _01207_);
  and _52303_ (_01211_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and _52304_ (_01213_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor _52305_ (_01215_, _01213_, _01211_);
  and _52306_ (_01217_, _01215_, _01209_);
  and _52307_ (_01219_, _01217_, _01206_);
  nor _52308_ (_01221_, _01219_, _36636_);
  nor _52309_ (_01223_, _01221_, _01203_);
  nor _52310_ (_01225_, _01223_, _42250_);
  nor _52311_ (_01227_, _01225_, _01202_);
  nor _52312_ (_38986_, _01227_, rst);
  and _52313_ (_01230_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [3]);
  and _52314_ (_01232_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  and _52315_ (_01234_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _52316_ (_01236_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _52317_ (_01238_, _01236_, _01234_);
  and _52318_ (_01240_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _52319_ (_01242_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _52320_ (_01244_, _01242_, _01240_);
  and _52321_ (_01246_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _52322_ (_01248_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _52323_ (_01250_, _01248_, _01246_);
  and _52324_ (_01252_, _01250_, _01244_);
  and _52325_ (_01254_, _01252_, _01238_);
  nor _52326_ (_01256_, _01254_, _36636_);
  nor _52327_ (_01258_, _01256_, _01232_);
  nor _52328_ (_01260_, _01258_, _42250_);
  nor _52329_ (_01262_, _01260_, _01230_);
  nor _52330_ (_38987_, _01262_, rst);
  and _52331_ (_01265_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [4]);
  and _52332_ (_01267_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  and _52333_ (_01269_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _52334_ (_01271_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _52335_ (_01273_, _01271_, _01269_);
  and _52336_ (_01275_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _52337_ (_01277_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _52338_ (_01279_, _01277_, _01275_);
  and _52339_ (_01281_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _52340_ (_01283_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _52341_ (_01285_, _01283_, _01281_);
  and _52342_ (_01287_, _01285_, _01279_);
  and _52343_ (_01289_, _01287_, _01273_);
  nor _52344_ (_01291_, _01289_, _36636_);
  nor _52345_ (_01293_, _01291_, _01267_);
  nor _52346_ (_01295_, _01293_, _42250_);
  nor _52347_ (_01297_, _01295_, _01265_);
  nor _52348_ (_38988_, _01297_, rst);
  and _52349_ (_01300_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [5]);
  and _52350_ (_01302_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  and _52351_ (_01304_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _52352_ (_01305_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _52353_ (_01306_, _01305_, _01304_);
  and _52354_ (_01307_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _52355_ (_01308_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _52356_ (_01309_, _01308_, _01307_);
  and _52357_ (_01310_, _01309_, _01306_);
  and _52358_ (_01311_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _52359_ (_01312_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _52360_ (_01313_, _01312_, _01311_);
  and _52361_ (_01314_, _01313_, _01310_);
  nor _52362_ (_01315_, _01314_, _36636_);
  nor _52363_ (_01316_, _01315_, _01302_);
  nor _52364_ (_01317_, _01316_, _42250_);
  nor _52365_ (_01318_, _01317_, _01300_);
  nor _52366_ (_38990_, _01318_, rst);
  and _52367_ (_01319_, _42250_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [6]);
  and _52368_ (_01320_, _36636_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  and _52369_ (_01321_, _36701_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _52370_ (_01322_, _36668_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _52371_ (_01323_, _01322_, _01321_);
  and _52372_ (_01324_, _36548_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _52373_ (_01325_, _36516_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _52374_ (_01326_, _01325_, _01324_);
  and _52375_ (_01327_, _36723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _52376_ (_01328_, _36592_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _52377_ (_01329_, _01328_, _01327_);
  and _52378_ (_01330_, _01329_, _01326_);
  and _52379_ (_01331_, _01330_, _01323_);
  nor _52380_ (_01332_, _01331_, _36636_);
  nor _52381_ (_01333_, _01332_, _01320_);
  nor _52382_ (_01334_, _01333_, _42250_);
  nor _52383_ (_01335_, _01334_, _01319_);
  nor _52384_ (_38991_, _01335_, rst);
  and _52385_ (_01336_, _36461_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  or _52386_ (_01337_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand _52387_ (_01338_, _01336_, _38536_);
  and _52388_ (_01339_, _01338_, _42882_);
  and _52389_ (_39015_, _01339_, _01337_);
  not _52390_ (_01340_, _01336_);
  or _52391_ (_01341_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _52392_ (_01342_, _36461_, _42882_);
  and _52393_ (_00000_, _01342_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and _52394_ (_01343_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _42882_);
  or _52395_ (_01344_, _01343_, _00000_);
  and _52396_ (_39016_, _01344_, _01341_);
  nor _52397_ (_39054_, _42304_, rst);
  nor _52398_ (_39056_, _42342_, rst);
  and _52399_ (_39057_, _42300_, _42882_);
  not _52400_ (_01345_, _38352_);
  nor _52401_ (_01346_, _38341_, _38350_);
  nor _52402_ (_01347_, _42448_, _27703_);
  and _52403_ (_01348_, _42448_, _27703_);
  nor _52404_ (_01349_, _01348_, _01347_);
  nor _52405_ (_01350_, _42365_, _27845_);
  and _52406_ (_01351_, _42365_, _27845_);
  nor _52407_ (_01352_, _01351_, _01350_);
  nor _52408_ (_01353_, _01352_, _01349_);
  nor _52409_ (_01354_, _42573_, _27374_);
  and _52410_ (_01355_, _42573_, _27374_);
  nor _52411_ (_01356_, _01355_, _01354_);
  nor _52412_ (_01357_, _42527_, _27242_);
  and _52413_ (_01358_, _42527_, _27242_);
  nor _52414_ (_01359_, _01358_, _01357_);
  nor _52415_ (_01360_, _01359_, _01356_);
  and _52416_ (_01361_, _01360_, _01353_);
  and _52417_ (_01362_, _01361_, _42639_);
  nor _52418_ (_01363_, _31304_, _39838_);
  and _52419_ (_01364_, _01363_, _01362_);
  and _52420_ (_01365_, _01364_, _01346_);
  not _52421_ (_01366_, _01365_);
  nor _52422_ (_01367_, _42402_, _26902_);
  and _52423_ (_01368_, _42402_, _26902_);
  nor _52424_ (_01369_, _01368_, _01367_);
  and _52425_ (_01370_, _42484_, _32545_);
  nor _52426_ (_01371_, _01370_, _01369_);
  nor _52427_ (_01372_, _42610_, _26781_);
  and _52428_ (_01373_, _42610_, _26781_);
  nor _52429_ (_01374_, _01373_, _01372_);
  nor _52430_ (_01375_, _42484_, _32545_);
  or _52431_ (_01376_, _01375_, _39217_);
  nor _52432_ (_01377_, _01376_, _01374_);
  and _52433_ (_01378_, _01377_, _01362_);
  and _52434_ (_01379_, _01378_, _01371_);
  nor _52435_ (_01380_, _27549_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _52436_ (_01381_, _01380_, _01379_);
  not _52437_ (_01382_, _01381_);
  and _52438_ (_01383_, _38298_, _38260_);
  nor _52439_ (_01384_, _01383_, _00783_);
  nor _52440_ (_01385_, _01384_, _36407_);
  not _52441_ (_01386_, _38296_);
  and _52442_ (_01387_, _38223_, _38375_);
  nor _52443_ (_01388_, _01387_, _00731_);
  nor _52444_ (_01389_, _01346_, _38248_);
  not _52445_ (_01390_, _31455_);
  nand _52446_ (_01391_, _33513_, _01390_);
  or _52447_ (_01392_, _01391_, _29030_);
  nor _52448_ (_01393_, _01392_, _34232_);
  and _52449_ (_01394_, _01393_, _34960_);
  and _52450_ (_01395_, _01394_, _28569_);
  and _52451_ (_01396_, _01395_, _01389_);
  and _52452_ (_01397_, _01396_, _35744_);
  and _52453_ (_01398_, _01397_, _29216_);
  not _52454_ (_01399_, _01398_);
  and _52455_ (_01400_, _01346_, _28931_);
  not _52456_ (_01401_, _01400_);
  not _52457_ (_01402_, _38248_);
  nor _52458_ (_01403_, _01346_, _38297_);
  nor _52459_ (_01404_, _01403_, _01402_);
  and _52460_ (_01405_, _01404_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _52461_ (_01406_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _52462_ (_01407_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _52463_ (_01408_, _01407_, _01406_);
  nor _52464_ (_01409_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _52465_ (_01410_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _52466_ (_01411_, _01410_, _01409_);
  and _52467_ (_01412_, _01411_, _01408_);
  and _52468_ (_01413_, _01412_, _38394_);
  nor _52469_ (_01414_, _01413_, _01405_);
  and _52470_ (_01415_, _01414_, _01401_);
  and _52471_ (_01416_, _01415_, _01399_);
  or _52472_ (_01417_, _38334_, _38223_);
  or _52473_ (_01418_, _01417_, _38326_);
  and _52474_ (_01419_, _01418_, _38246_);
  not _52475_ (_01420_, _01419_);
  not _52476_ (_01421_, _00809_);
  nor _52477_ (_01422_, _01007_, _38306_);
  and _52478_ (_01423_, _01422_, _01421_);
  and _52479_ (_01424_, _01423_, _00969_);
  and _52480_ (_01425_, _01424_, _01420_);
  not _52481_ (_01426_, _01425_);
  and _52482_ (_01427_, _01426_, _01416_);
  and _52483_ (_01428_, _38247_, _36920_);
  not _52484_ (_01429_, _01428_);
  and _52485_ (_01430_, _01429_, _38340_);
  nor _52486_ (_01431_, _01430_, _01416_);
  nor _52487_ (_01432_, _01431_, _01427_);
  and _52488_ (_01433_, _01432_, _01388_);
  and _52489_ (_01434_, _01433_, _01386_);
  nor _52490_ (_01435_, _38352_, _38243_);
  nor _52491_ (_01436_, _01435_, _01434_);
  nor _52492_ (_01437_, _01436_, _01385_);
  not _52493_ (_01438_, _38875_);
  nor _52494_ (_01439_, _38901_, _01438_);
  and _52495_ (_01440_, _01439_, _38883_);
  not _52496_ (_01441_, _01440_);
  and _52497_ (_01442_, _01441_, _01404_);
  not _52498_ (_01443_, _39133_);
  and _52499_ (_01444_, _01443_, _38394_);
  nor _52500_ (_01445_, _01444_, _01442_);
  not _52501_ (_01446_, _01445_);
  nor _52502_ (_01447_, _01446_, _01437_);
  and _52503_ (_01448_, _01447_, _01382_);
  and _52504_ (_01449_, _01448_, _01366_);
  and _52505_ (_01450_, _01449_, _01345_);
  and _52506_ (_39061_, _01450_, _42882_);
  and _52507_ (_39062_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _42882_);
  and _52508_ (_39063_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _42882_);
  and _52509_ (_01451_, _00969_, _38341_);
  and _52510_ (_01452_, _01451_, _01422_);
  nor _52511_ (_01453_, _01452_, _42317_);
  and _52512_ (_01454_, _01383_, _36396_);
  not _52513_ (_01455_, _01454_);
  and _52514_ (_01456_, _38246_, _38295_);
  and _52515_ (_01457_, _01456_, _36396_);
  nor _52516_ (_01458_, _01457_, _38352_);
  and _52517_ (_01459_, _01458_, _01455_);
  not _52518_ (_01460_, _01459_);
  nor _52519_ (_01461_, _01460_, _01453_);
  and _52520_ (_01462_, _01461_, _42266_);
  not _52521_ (_01463_, _01167_);
  nor _52522_ (_01464_, _01461_, _01463_);
  nor _52523_ (_01465_, _01464_, _01462_);
  and _52524_ (_01466_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _52525_ (_01467_, _01466_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _52526_ (_01468_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _52527_ (_01469_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _52528_ (_01470_, _01461_, _42523_);
  not _52529_ (_01471_, _01335_);
  nor _52530_ (_01472_, _01461_, _01471_);
  nor _52531_ (_01473_, _01472_, _01470_);
  and _52532_ (_01474_, _01473_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _52533_ (_01475_, _01473_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _52534_ (_01476_, _01475_, _01474_);
  and _52535_ (_01477_, _01461_, _42551_);
  not _52536_ (_01478_, _01318_);
  nor _52537_ (_01479_, _01461_, _01478_);
  nor _52538_ (_01480_, _01479_, _01477_);
  and _52539_ (_01481_, _01480_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _52540_ (_01482_, _01480_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _52541_ (_01483_, _01461_, _42336_);
  not _52542_ (_01484_, _01297_);
  nor _52543_ (_01485_, _01461_, _01484_);
  nor _52544_ (_01486_, _01485_, _01483_);
  nand _52545_ (_01487_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _52546_ (_01488_, _01461_, _42429_);
  not _52547_ (_01489_, _01262_);
  nor _52548_ (_01490_, _01461_, _01489_);
  nor _52549_ (_01491_, _01490_, _01488_);
  and _52550_ (_01492_, _01491_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _52551_ (_01493_, _01491_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _52552_ (_01494_, _01461_, _42589_);
  not _52553_ (_01495_, _01227_);
  nor _52554_ (_01496_, _01461_, _01495_);
  nor _52555_ (_01497_, _01496_, _01494_);
  and _52556_ (_01498_, _01497_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _52557_ (_01499_, _01461_, _42384_);
  not _52558_ (_01500_, _01201_);
  nor _52559_ (_01501_, _01461_, _01500_);
  nor _52560_ (_01502_, _01501_, _01499_);
  and _52561_ (_01503_, _01502_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _52562_ (_01504_, _01461_, _42464_);
  not _52563_ (_01505_, _01184_);
  nor _52564_ (_01506_, _01461_, _01505_);
  nor _52565_ (_01507_, _01506_, _01504_);
  and _52566_ (_01508_, _01507_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _52567_ (_01509_, _01502_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _52568_ (_01510_, _01509_, _01503_);
  and _52569_ (_01511_, _01510_, _01508_);
  nor _52570_ (_01512_, _01511_, _01503_);
  not _52571_ (_01513_, _01512_);
  nor _52572_ (_01514_, _01497_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _52573_ (_01515_, _01514_, _01498_);
  and _52574_ (_01516_, _01515_, _01513_);
  nor _52575_ (_01517_, _01516_, _01498_);
  nor _52576_ (_01518_, _01517_, _01493_);
  or _52577_ (_01519_, _01518_, _01492_);
  or _52578_ (_01520_, _01486_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _52579_ (_01521_, _01520_, _01487_);
  nand _52580_ (_01522_, _01521_, _01519_);
  and _52581_ (_01523_, _01522_, _01487_);
  nor _52582_ (_01524_, _01523_, _01482_);
  or _52583_ (_01525_, _01524_, _01481_);
  and _52584_ (_01526_, _01525_, _01476_);
  nor _52585_ (_01527_, _01526_, _01474_);
  nor _52586_ (_01528_, _01527_, _01469_);
  or _52587_ (_01529_, _01528_, _01468_);
  and _52588_ (_01530_, _01529_, _01467_);
  and _52589_ (_01531_, _01530_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _52590_ (_01532_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _52591_ (_01533_, _01532_, _01531_);
  nor _52592_ (_01534_, _01533_, _01465_);
  not _52593_ (_01535_, _01465_);
  nor _52594_ (_01536_, _01529_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _52595_ (_01537_, _01536_, _38558_);
  and _52596_ (_01538_, _01537_, _38563_);
  and _52597_ (_01539_, _01538_, _38548_);
  nor _52598_ (_01540_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _52599_ (_01541_, _01540_, _01539_);
  nor _52600_ (_01542_, _01541_, _01535_);
  nor _52601_ (_01543_, _01542_, _01534_);
  or _52602_ (_01544_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _52603_ (_01545_, _01465_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _52604_ (_01546_, _01545_, _01544_);
  and _52605_ (_01547_, _01546_, _01543_);
  nand _52606_ (_01548_, _01547_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or _52607_ (_01549_, _01547_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not _52608_ (_01550_, _38247_);
  and _52609_ (_01551_, _01388_, _01550_);
  and _52610_ (_01552_, _01551_, _01423_);
  and _52611_ (_01553_, _01552_, _01451_);
  nor _52612_ (_01554_, _01553_, _42317_);
  nor _52613_ (_01555_, _01554_, _01457_);
  and _52614_ (_01556_, _38224_, _38243_);
  nor _52615_ (_01557_, _01556_, _01385_);
  not _52616_ (_01558_, _01557_);
  and _52617_ (_01559_, _01558_, _01461_);
  nor _52618_ (_01560_, _01559_, _01555_);
  and _52619_ (_01561_, _01560_, _01549_);
  and _52620_ (_01562_, _01561_, _01548_);
  nor _52621_ (_01563_, _01345_, _30603_);
  not _52622_ (_01564_, _38621_);
  and _52623_ (_01565_, _01556_, _01564_);
  and _52624_ (_01566_, _01559_, _01555_);
  and _52625_ (_01567_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _52626_ (_01568_, _01567_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _52627_ (_01569_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _52628_ (_01570_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _52629_ (_01571_, _01570_, _01569_);
  and _52630_ (_01572_, _01571_, _01568_);
  and _52631_ (_01573_, _01572_, _01467_);
  and _52632_ (_01574_, _01573_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _52633_ (_01575_, _01574_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _52634_ (_01576_, _01575_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand _52635_ (_01577_, _01576_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _52636_ (_01578_, _01577_, _38536_);
  or _52637_ (_01579_, _01577_, _38536_);
  and _52638_ (_01580_, _01579_, _01578_);
  and _52639_ (_01581_, _01580_, _01566_);
  and _52640_ (_01582_, _01454_, _42267_);
  or _52641_ (_01583_, _01582_, _01581_);
  and _52642_ (_01584_, _01557_, _01461_);
  and _52643_ (_01585_, _01584_, _01555_);
  and _52644_ (_01586_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _52645_ (_01587_, _01586_, _01583_);
  nor _52646_ (_01588_, _01587_, _01565_);
  nand _52647_ (_01589_, _01588_, _01449_);
  or _52648_ (_01590_, _01589_, _01563_);
  or _52649_ (_01591_, _01590_, _01562_);
  nor _52650_ (_01592_, _36537_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _52651_ (_01593_, _01592_, _42250_);
  nor _52652_ (_01594_, _01593_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _52653_ (_01595_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _52654_ (_01596_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _52655_ (_01597_, _01596_, _01595_);
  not _52656_ (_01598_, _01597_);
  nor _52657_ (_01599_, _01598_, _01594_);
  and _52658_ (_01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _52659_ (_01601_, _01600_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _52660_ (_01602_, _01601_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _52661_ (_01603_, _01602_, _01599_);
  and _52662_ (_01604_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _52663_ (_01605_, _01604_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _52664_ (_01606_, _01605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _52665_ (_01607_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _52666_ (_01608_, _01607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _52667_ (_01609_, _01608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand _52668_ (_01610_, _01608_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _52669_ (_01611_, _01610_, _01609_);
  or _52670_ (_01612_, _01611_, _01449_);
  and _52671_ (_01613_, _01612_, _42882_);
  and _52672_ (_39064_, _01613_, _01591_);
  and _52673_ (_01614_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _42882_);
  and _52674_ (_01615_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _52675_ (_01616_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _52676_ (_01617_, _36450_, _01616_);
  not _52677_ (_01618_, _01617_);
  not _52678_ (_01619_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _52679_ (_01620_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _52680_ (_01621_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not _52681_ (_01622_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _52682_ (_01623_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _52683_ (_01624_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _52684_ (_01625_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _52685_ (_01626_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor _52686_ (_01627_, _01626_, _01624_);
  and _52687_ (_01629_, _01627_, _01625_);
  nor _52688_ (_01630_, _01629_, _01624_);
  nor _52689_ (_01632_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _52690_ (_01633_, _01632_, _01623_);
  not _52691_ (_01635_, _01633_);
  nor _52692_ (_01636_, _01635_, _01630_);
  nor _52693_ (_01638_, _01636_, _01623_);
  not _52694_ (_01639_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _52695_ (_01641_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9], \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _52696_ (_01642_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _52697_ (_01644_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _52698_ (_01645_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _52699_ (_01647_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _52700_ (_01648_, _01647_, _01645_);
  and _52701_ (_01650_, _01648_, _01644_);
  and _52702_ (_01651_, _01650_, _01642_);
  and _52703_ (_01653_, _01651_, _01641_);
  and _52704_ (_01654_, _01653_, _01639_);
  and _52705_ (_01656_, _01654_, _01638_);
  and _52706_ (_01657_, _01656_, _01622_);
  and _52707_ (_01659_, _01657_, _01621_);
  and _52708_ (_01660_, _01659_, _01620_);
  and _52709_ (_01661_, _01660_, _01619_);
  nor _52710_ (_01662_, _01661_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _52711_ (_01663_, _01661_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _52712_ (_01664_, _01663_, _01662_);
  not _52713_ (_01665_, _01664_);
  nor _52714_ (_01666_, _01660_, _01619_);
  nor _52715_ (_01667_, _01666_, _01661_);
  not _52716_ (_01668_, _01667_);
  nor _52717_ (_01669_, _01659_, _01620_);
  or _52718_ (_01670_, _01669_, _01660_);
  nor _52719_ (_01671_, _01657_, _01621_);
  nor _52720_ (_01672_, _01671_, _01659_);
  not _52721_ (_01673_, _01672_);
  nor _52722_ (_01674_, _01656_, _01622_);
  nor _52723_ (_01675_, _01674_, _01657_);
  not _52724_ (_01676_, _01675_);
  and _52725_ (_01677_, _01653_, _01638_);
  nor _52726_ (_01678_, _01677_, _01639_);
  nor _52727_ (_01679_, _01678_, _01656_);
  not _52728_ (_01680_, _01679_);
  not _52729_ (_01681_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _52730_ (_01682_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _52731_ (_01683_, _01651_, _01638_);
  and _52732_ (_01684_, _01683_, _01682_);
  nor _52733_ (_01685_, _01684_, _01681_);
  nor _52734_ (_01686_, _01685_, _01677_);
  not _52735_ (_01687_, _01686_);
  and _52736_ (_01688_, _01648_, _01638_);
  and _52737_ (_01689_, _01688_, _01644_);
  nor _52738_ (_01690_, _01689_, _01642_);
  or _52739_ (_01691_, _01690_, _01683_);
  nor _52740_ (_01692_, _01688_, _01644_);
  or _52741_ (_01693_, _01692_, _01689_);
  and _52742_ (_01694_, _01647_, _01638_);
  nor _52743_ (_01695_, _01694_, _01645_);
  nor _52744_ (_01696_, _01695_, _01688_);
  not _52745_ (_01697_, _01696_);
  not _52746_ (_01698_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _52747_ (_01699_, _01638_, _01698_);
  nor _52748_ (_01700_, _01638_, _01698_);
  nor _52749_ (_01701_, _01700_, _01699_);
  not _52750_ (_01702_, _01701_);
  and _52751_ (_01703_, _00706_, _00635_);
  and _52752_ (_01704_, _01703_, _00708_);
  not _52753_ (_01705_, _01704_);
  or _52754_ (_01706_, _00711_, _00658_);
  and _52755_ (_01707_, _01706_, _00708_);
  not _52756_ (_01708_, _00708_);
  and _52757_ (_01709_, _00651_, _00644_);
  nor _52758_ (_01710_, _01709_, _00683_);
  nor _52759_ (_01711_, _01710_, _01708_);
  nor _52760_ (_01712_, _01711_, _01707_);
  and _52761_ (_01713_, _01712_, _01705_);
  and _52762_ (_01714_, _00713_, _00704_);
  and _52763_ (_01715_, _00708_, _00661_);
  nor _52764_ (_01716_, _01715_, _01714_);
  not _52765_ (_01717_, _00660_);
  nor _52766_ (_01718_, _00658_, _00707_);
  nor _52767_ (_01719_, _01718_, _01717_);
  not _52768_ (_01720_, _00667_);
  and _52769_ (_01721_, _00678_, _00635_);
  nor _52770_ (_01722_, _01721_, _00645_);
  nor _52771_ (_01723_, _01722_, _01720_);
  nor _52772_ (_01724_, _01723_, _01719_);
  and _52773_ (_01725_, _01724_, _01716_);
  and _52774_ (_01726_, _01725_, _01713_);
  and _52775_ (_01727_, _01726_, _00688_);
  not _52776_ (_01728_, _00673_);
  and _52777_ (_01729_, _00703_, _00658_);
  nor _52778_ (_01730_, _01729_, _00646_);
  and _52779_ (_01731_, _00657_, _00689_);
  and _52780_ (_01732_, _00694_, _01731_);
  and _52781_ (_01733_, _00635_, _00642_);
  and _52782_ (_01734_, _00649_, _38185_);
  and _52783_ (_01735_, _01734_, _01733_);
  nor _52784_ (_01736_, _01735_, _01732_);
  and _52785_ (_01737_, _01736_, _01730_);
  and _52786_ (_01738_, _01737_, _01728_);
  and _52787_ (_01739_, _00672_, _00635_);
  nor _52788_ (_01740_, _00650_, _00639_);
  and _52789_ (_01741_, _00683_, _37905_);
  nor _52790_ (_01742_, _01741_, _00679_);
  nor _52791_ (_01743_, _01742_, _01740_);
  nor _52792_ (_01744_, _01743_, _01739_);
  and _52793_ (_01745_, _01744_, _01738_);
  and _52794_ (_01746_, _00683_, _00640_);
  and _52795_ (_01747_, _00678_, _00644_);
  and _52796_ (_01748_, _01747_, _00708_);
  nor _52797_ (_01749_, _01748_, _01746_);
  and _52798_ (_01750_, _00711_, _00660_);
  not _52799_ (_01751_, _00703_);
  nor _52800_ (_01752_, _01703_, _00685_);
  nor _52801_ (_01753_, _01752_, _01751_);
  nor _52802_ (_01754_, _01753_, _01750_);
  and _52803_ (_01755_, _01754_, _01749_);
  nor _52804_ (_01756_, _00712_, _00663_);
  nor _52805_ (_01757_, _01733_, _00658_);
  nor _52806_ (_01758_, _01757_, _38210_);
  nor _52807_ (_01759_, _01758_, _00699_);
  and _52808_ (_01760_, _01759_, _01756_);
  and _52809_ (_01761_, _01760_, _01755_);
  and _52810_ (_01762_, _01761_, _01745_);
  not _52811_ (_01763_, _00653_);
  not _52812_ (_01764_, _00671_);
  and _52813_ (_01765_, _00657_, _00706_);
  and _52814_ (_01766_, _01765_, _00640_);
  nor _52815_ (_01767_, _01766_, _00709_);
  and _52816_ (_01768_, _01767_, _01764_);
  and _52817_ (_01769_, _01768_, _01763_);
  and _52818_ (_01770_, _00670_, _00635_);
  nor _52819_ (_01771_, _01770_, _00652_);
  nor _52820_ (_01772_, _01771_, _01717_);
  not _52821_ (_01773_, _01772_);
  not _52822_ (_01774_, _01765_);
  nor _52823_ (_01775_, _00660_, _00650_);
  nor _52824_ (_01776_, _01775_, _01774_);
  and _52825_ (_01777_, _00669_, _00644_);
  not _52826_ (_01778_, _01777_);
  nor _52827_ (_01779_, _00708_, _00660_);
  nor _52828_ (_01780_, _01779_, _01778_);
  nor _52829_ (_01781_, _01780_, _01776_);
  and _52830_ (_01782_, _01781_, _01773_);
  and _52831_ (_01783_, _01782_, _01769_);
  and _52832_ (_01784_, _01783_, _01762_);
  and _52833_ (_01785_, _01784_, _01727_);
  not _52834_ (_01786_, _01785_);
  nor _52835_ (_01787_, _01627_, _01625_);
  nor _52836_ (_01788_, _01787_, _01629_);
  nand _52837_ (_01789_, _01788_, _01786_);
  and _52838_ (_01790_, _00657_, _00642_);
  and _52839_ (_01791_, _01790_, _00640_);
  and _52840_ (_01792_, _01703_, _00667_);
  or _52841_ (_01793_, _01792_, _01707_);
  or _52842_ (_01794_, _00686_, _00663_);
  or _52843_ (_01795_, _01794_, _01793_);
  or _52844_ (_01796_, _01795_, _01791_);
  not _52845_ (_01797_, _00699_);
  nand _52846_ (_01798_, _01769_, _01797_);
  or _52847_ (_01799_, _01798_, _01796_);
  nor _52848_ (_01800_, _01799_, _01785_);
  not _52849_ (_01801_, _01800_);
  nor _52850_ (_01802_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _52851_ (_01803_, _01802_, _01625_);
  and _52852_ (_01804_, _01803_, _01801_);
  or _52853_ (_01805_, _01788_, _01786_);
  and _52854_ (_01806_, _01805_, _01789_);
  nand _52855_ (_01807_, _01806_, _01804_);
  and _52856_ (_01808_, _01807_, _01789_);
  not _52857_ (_01809_, _01808_);
  and _52858_ (_01810_, _01635_, _01630_);
  nor _52859_ (_01811_, _01810_, _01636_);
  and _52860_ (_01812_, _01811_, _01809_);
  and _52861_ (_01813_, _01812_, _01702_);
  not _52862_ (_01814_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _52863_ (_01815_, _01699_, _01814_);
  or _52864_ (_01816_, _01815_, _01694_);
  and _52865_ (_01817_, _01816_, _01813_);
  and _52866_ (_01818_, _01817_, _01697_);
  and _52867_ (_01819_, _01818_, _01693_);
  and _52868_ (_01820_, _01819_, _01691_);
  nor _52869_ (_01821_, _01683_, _01682_);
  or _52870_ (_01822_, _01821_, _01684_);
  and _52871_ (_01823_, _01822_, _01820_);
  and _52872_ (_01824_, _01823_, _01687_);
  and _52873_ (_01825_, _01824_, _01680_);
  and _52874_ (_01826_, _01825_, _01676_);
  and _52875_ (_01827_, _01826_, _01673_);
  and _52876_ (_01828_, _01827_, _01670_);
  nand _52877_ (_01829_, _01828_, _01668_);
  nand _52878_ (_01830_, _01829_, _01665_);
  or _52879_ (_01831_, _01829_, _01665_);
  and _52880_ (_01832_, _01831_, _01830_);
  or _52881_ (_01833_, _01832_, _01618_);
  or _52882_ (_01834_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor _52883_ (_01835_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  and _52884_ (_01836_, _01835_, _01834_);
  and _52885_ (_01837_, _01836_, _01833_);
  or _52886_ (_39066_, _01837_, _01615_);
  nor _52887_ (_01838_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _52888_ (_39067_, _01838_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _52889_ (_39068_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _42882_);
  not _52890_ (_01839_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor _52891_ (_01840_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _52892_ (_01841_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _52893_ (_01842_, _01841_, _01840_);
  not _52894_ (_01843_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor _52895_ (_01844_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _52896_ (_01845_, _01844_, _01843_);
  and _52897_ (_01846_, _01845_, _01842_);
  and _52898_ (_01847_, _01846_, _01839_);
  and _52899_ (_01848_, \oc8051_top_1.oc8051_rom1.ea_int , _36418_);
  nand _52900_ (_01849_, _01848_, _36450_);
  nand _52901_ (_01850_, _01849_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand _52902_ (_01851_, _01850_, _01847_);
  and _52903_ (_39069_, _01851_, _42882_);
  and _52904_ (_01852_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _52905_ (_01853_, _01852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _52906_ (_39071_, _01853_, _42882_);
  nor _52907_ (_01854_, _01594_, _42250_);
  or _52908_ (_01855_, _01785_, _36646_);
  nor _52909_ (_01856_, _01800_, _36570_);
  nand _52910_ (_01857_, _01785_, _36646_);
  and _52911_ (_01858_, _01857_, _01855_);
  nand _52912_ (_01859_, _01858_, _01856_);
  and _52913_ (_01860_, _01859_, _01855_);
  nor _52914_ (_01861_, _01860_, _42250_);
  and _52915_ (_01862_, _01861_, _36494_);
  nor _52916_ (_01863_, _01861_, _36494_);
  nor _52917_ (_01864_, _01863_, _01862_);
  nor _52918_ (_01865_, _01864_, _01854_);
  and _52919_ (_01866_, _36657_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and _52920_ (_01867_, _01866_, _01854_);
  and _52921_ (_01868_, _01867_, _01799_);
  or _52922_ (_01869_, _01868_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _52923_ (_01870_, _01869_, _01865_);
  and _52924_ (_39072_, _01870_, _42882_);
  nor _52925_ (_01871_, _38179_, _36767_);
  and _52926_ (_01872_, _37313_, _37062_);
  and _52927_ (_01873_, _01872_, _01871_);
  nand _52928_ (_01874_, _01342_, _38101_);
  nor _52929_ (_01875_, _01874_, _37861_);
  not _52930_ (_01876_, _38206_);
  and _52931_ (_01877_, _01876_, _37586_);
  and _52932_ (_01878_, _01877_, _01875_);
  and _52933_ (_39075_, _01878_, _01873_);
  nor _52934_ (_01879_, \oc8051_top_1.oc8051_memory_interface1.istb_t , rst);
  and _52935_ (_01880_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  and _52936_ (_01881_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [7]);
  and _52937_ (_39078_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _42882_);
  and _52938_ (_01882_, _39078_, _01881_);
  or _52939_ (_39076_, _01882_, _01880_);
  not _52940_ (_01883_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and _52941_ (_01884_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _52942_ (_01885_, _01884_, _01883_);
  and _52943_ (_01886_, _01884_, _01883_);
  nor _52944_ (_01887_, _01886_, _01885_);
  not _52945_ (_01888_, _01887_);
  and _52946_ (_01889_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _52947_ (_01890_, _01889_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _52948_ (_01891_, _01889_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _52949_ (_01892_, _01891_, _01890_);
  or _52950_ (_01893_, _01892_, _01884_);
  and _52951_ (_01894_, _01893_, _01888_);
  nor _52952_ (_01895_, _01885_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _52953_ (_01896_, _01885_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _52954_ (_01897_, _01896_, _01895_);
  or _52955_ (_01898_, _01890_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _52956_ (_39080_, _01898_, _42882_);
  and _52957_ (_01899_, _39080_, _01897_);
  and _52958_ (_39079_, _01899_, _01894_);
  not _52959_ (_01900_, \oc8051_top_1.oc8051_rom1.ea_int );
  nor _52960_ (_01901_, _01594_, _01900_);
  and _52961_ (_01902_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  not _52962_ (_01903_, _01901_);
  and _52963_ (_01904_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or _52964_ (_01905_, _01904_, _01902_);
  and _52965_ (_39081_, _01905_, _42882_);
  and _52966_ (_01906_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _52967_ (_01907_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or _52968_ (_01908_, _01907_, _01906_);
  and _52969_ (_39082_, _01908_, _42882_);
  and _52970_ (_01909_, \oc8051_top_1.oc8051_decoder1.mem_act [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  not _52971_ (_01910_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52972_ (_01911_, \oc8051_top_1.oc8051_decoder1.mem_act [0], _01910_);
  and _52973_ (_01912_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _52974_ (_01913_, _01912_, _01909_);
  and _52975_ (_39083_, _01913_, _42882_);
  and _52976_ (_01914_, \oc8051_top_1.oc8051_memory_interface1.dwe_o , \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52977_ (_01915_, _01914_, _01911_);
  and _52978_ (_39084_, _01915_, _42882_);
  or _52979_ (_01916_, _01910_, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  and _52980_ (_39086_, _01916_, _42882_);
  not _52981_ (_01917_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _52982_ (_01918_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _52983_ (_01919_, _01918_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _52984_ (_01920_, _01910_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  and _52985_ (_01921_, _01920_, _42882_);
  and _52986_ (_39087_, _01921_, _01919_);
  or _52987_ (_01922_, _01910_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  and _52988_ (_39088_, _01922_, _42882_);
  nor _52989_ (_01923_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  and _52990_ (_01924_, _01923_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _52991_ (_01925_, _01924_, _42882_);
  and _52992_ (_01926_, _39078_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _52993_ (_39089_, _01926_, _01925_);
  and _52994_ (_01927_, _01900_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _52995_ (_01928_, _01927_, _01924_);
  and _52996_ (_39090_, _01928_, _42882_);
  nand _52997_ (_01929_, _01924_, _38621_);
  or _52998_ (_01930_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [15]);
  and _52999_ (_01931_, _01930_, _42882_);
  and _53000_ (_39091_, _01931_, _01929_);
  nand _53001_ (_01932_, _38257_, _42882_);
  nor _53002_ (_39092_, _01932_, _38398_);
  or _53003_ (_01933_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _53004_ (_01934_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _53005_ (_01935_, _01934_, _42882_);
  and _53006_ (_39128_, _01935_, _01933_);
  or _53007_ (_01936_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _53008_ (_01937_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand _53009_ (_01938_, _01336_, _01937_);
  and _53010_ (_01939_, _01938_, _42882_);
  and _53011_ (_39129_, _01939_, _01936_);
  or _53012_ (_01940_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _53013_ (_01941_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _53014_ (_01942_, _01336_, _01941_);
  and _53015_ (_01943_, _01942_, _42882_);
  and _53016_ (_39130_, _01943_, _01940_);
  or _53017_ (_01944_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _53018_ (_01945_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand _53019_ (_01946_, _01336_, _01945_);
  and _53020_ (_01947_, _01946_, _42882_);
  and _53021_ (_39131_, _01947_, _01944_);
  or _53022_ (_01948_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not _53023_ (_01949_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand _53024_ (_01950_, _01336_, _01949_);
  and _53025_ (_01951_, _01950_, _42882_);
  and _53026_ (_39132_, _01951_, _01948_);
  or _53027_ (_01952_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not _53028_ (_01953_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand _53029_ (_01954_, _01336_, _01953_);
  and _53030_ (_01955_, _01954_, _42882_);
  and _53031_ (_39134_, _01955_, _01952_);
  or _53032_ (_01956_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  or _53033_ (_01957_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _53034_ (_01958_, _01957_, _42882_);
  and _53035_ (_39135_, _01958_, _01956_);
  or _53036_ (_01959_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  not _53037_ (_01960_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand _53038_ (_01961_, _01336_, _01960_);
  and _53039_ (_01962_, _01961_, _42882_);
  and _53040_ (_39136_, _01962_, _01959_);
  or _53041_ (_01963_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _53042_ (_01964_, _01336_, _38552_);
  and _53043_ (_01965_, _01964_, _42882_);
  and _53044_ (_39137_, _01965_, _01963_);
  or _53045_ (_01966_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _53046_ (_01967_, _01336_, _38558_);
  and _53047_ (_01968_, _01967_, _42882_);
  and _53048_ (_39138_, _01968_, _01966_);
  or _53049_ (_01969_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _53050_ (_01970_, _01336_, _38563_);
  and _53051_ (_01971_, _01970_, _42882_);
  and _53052_ (_39139_, _01971_, _01969_);
  or _53053_ (_01972_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _53054_ (_01973_, _01336_, _38548_);
  and _53055_ (_01974_, _01973_, _42882_);
  and _53056_ (_39140_, _01974_, _01972_);
  or _53057_ (_01975_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _53058_ (_01976_, _01336_, _38569_);
  and _53059_ (_01977_, _01976_, _42882_);
  and _53060_ (_39141_, _01977_, _01975_);
  or _53061_ (_01978_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _53062_ (_01979_, _01336_, _38544_);
  and _53063_ (_01980_, _01979_, _42882_);
  and _53064_ (_39142_, _01980_, _01978_);
  or _53065_ (_01981_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _53066_ (_01982_, _01336_, _38540_);
  and _53067_ (_01983_, _01982_, _42882_);
  and _53068_ (_39143_, _01983_, _01981_);
  and _53069_ (_01984_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _53070_ (_01985_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _53071_ (_01986_, _01985_, _01984_);
  and _53072_ (_39148_, _01986_, _42882_);
  and _53073_ (_01987_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _53074_ (_01988_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  or _53075_ (_01989_, _01988_, _01987_);
  and _53076_ (_39149_, _01989_, _42882_);
  and _53077_ (_01990_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _53078_ (_01991_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  or _53079_ (_01992_, _01991_, _01990_);
  and _53080_ (_39150_, _01992_, _42882_);
  and _53081_ (_01993_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _53082_ (_01994_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _53083_ (_01995_, _01994_, _01993_);
  and _53084_ (_39151_, _01995_, _42882_);
  and _53085_ (_01996_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _53086_ (_01997_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or _53087_ (_01998_, _01997_, _01996_);
  and _53088_ (_39152_, _01998_, _42882_);
  and _53089_ (_01999_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _53090_ (_02000_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  or _53091_ (_02001_, _02000_, _01999_);
  and _53092_ (_39153_, _02001_, _42882_);
  and _53093_ (_02002_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  and _53094_ (_02003_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  or _53095_ (_02004_, _02003_, _02002_);
  and _53096_ (_39154_, _02004_, _42882_);
  and _53097_ (_02005_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _53098_ (_02006_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  or _53099_ (_02007_, _02006_, _02005_);
  and _53100_ (_39155_, _02007_, _42882_);
  and _53101_ (_02008_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _53102_ (_02009_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  or _53103_ (_02010_, _02009_, _02008_);
  and _53104_ (_39156_, _02010_, _42882_);
  and _53105_ (_02011_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _53106_ (_02012_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  or _53107_ (_02013_, _02012_, _02011_);
  and _53108_ (_39157_, _02013_, _42882_);
  and _53109_ (_02014_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _53110_ (_02015_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  or _53111_ (_02016_, _02015_, _02014_);
  and _53112_ (_39159_, _02016_, _42882_);
  and _53113_ (_02017_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _53114_ (_02018_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or _53115_ (_02019_, _02018_, _02017_);
  and _53116_ (_39160_, _02019_, _42882_);
  and _53117_ (_02020_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _53118_ (_02021_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  or _53119_ (_02022_, _02021_, _02020_);
  and _53120_ (_39161_, _02022_, _42882_);
  and _53121_ (_02023_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _53122_ (_02024_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or _53123_ (_02025_, _02024_, _02023_);
  and _53124_ (_39162_, _02025_, _42882_);
  and _53125_ (_02026_, _01336_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _53126_ (_02027_, _01340_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or _53127_ (_02028_, _02027_, _02026_);
  and _53128_ (_39163_, _02028_, _42882_);
  and _53129_ (_39339_, _37960_, _42882_);
  and _53130_ (_39340_, _38190_, _42882_);
  and _53131_ (_39341_, _38167_, _42882_);
  nor _53132_ (_39342_, _42273_, rst);
  and _53133_ (_02029_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _53134_ (_02030_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  or _53135_ (_02031_, _02030_, _02029_);
  and _53136_ (_39343_, _02031_, _42882_);
  and _53137_ (_02032_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _53138_ (_02033_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [1]);
  and _53139_ (_02034_, _02033_, _01901_);
  or _53140_ (_02035_, _02034_, _02032_);
  and _53141_ (_39344_, _02035_, _42882_);
  and _53142_ (_02036_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _53143_ (_02037_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _53144_ (_02038_, _02037_, _02036_);
  and _53145_ (_39345_, _02038_, _42882_);
  and _53146_ (_02039_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _53147_ (_02040_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  or _53148_ (_02041_, _02040_, _02039_);
  and _53149_ (_39346_, _02041_, _42882_);
  and _53150_ (_02042_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _53151_ (_02043_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  or _53152_ (_02044_, _02043_, _02042_);
  and _53153_ (_39348_, _02044_, _42882_);
  and _53154_ (_02045_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _53155_ (_02046_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  or _53156_ (_02047_, _02046_, _02045_);
  and _53157_ (_39349_, _02047_, _42882_);
  and _53158_ (_02048_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _53159_ (_02049_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or _53160_ (_02050_, _02049_, _02048_);
  and _53161_ (_39350_, _02050_, _42882_);
  and _53162_ (_02051_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _53163_ (_02052_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  or _53164_ (_02053_, _02052_, _02051_);
  and _53165_ (_39351_, _02053_, _42882_);
  and _53166_ (_02054_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  and _53167_ (_02055_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  or _53168_ (_02056_, _02055_, _02054_);
  and _53169_ (_39352_, _02056_, _42882_);
  and _53170_ (_02057_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  and _53171_ (_02058_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or _53172_ (_02059_, _02058_, _02057_);
  and _53173_ (_39353_, _02059_, _42882_);
  and _53174_ (_02060_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  and _53175_ (_02061_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _53176_ (_02062_, _02061_, _02060_);
  and _53177_ (_39354_, _02062_, _42882_);
  and _53178_ (_02063_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  and _53179_ (_02064_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or _53180_ (_02065_, _02064_, _02063_);
  and _53181_ (_39355_, _02065_, _42882_);
  and _53182_ (_02066_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  and _53183_ (_02067_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _53184_ (_02068_, _02067_, _02066_);
  and _53185_ (_39356_, _02068_, _42882_);
  and _53186_ (_02069_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  and _53187_ (_02070_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or _53188_ (_02071_, _02070_, _02069_);
  and _53189_ (_39357_, _02071_, _42882_);
  and _53190_ (_02072_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  and _53191_ (_02073_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or _53192_ (_02074_, _02073_, _02072_);
  and _53193_ (_39359_, _02074_, _42882_);
  and _53194_ (_02075_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  and _53195_ (_02076_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or _53196_ (_02077_, _02076_, _02075_);
  and _53197_ (_39360_, _02077_, _42882_);
  and _53198_ (_02078_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  and _53199_ (_02079_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or _53200_ (_02080_, _02079_, _02078_);
  and _53201_ (_39361_, _02080_, _42882_);
  and _53202_ (_02081_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  and _53203_ (_02082_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or _53204_ (_02083_, _02082_, _02081_);
  and _53205_ (_39362_, _02083_, _42882_);
  and _53206_ (_02084_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  and _53207_ (_02085_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  or _53208_ (_02086_, _02085_, _02084_);
  and _53209_ (_39363_, _02086_, _42882_);
  and _53210_ (_02087_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  and _53211_ (_02088_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  or _53212_ (_02089_, _02088_, _02087_);
  and _53213_ (_39364_, _02089_, _42882_);
  and _53214_ (_02090_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  and _53215_ (_02091_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or _53216_ (_02092_, _02091_, _02090_);
  and _53217_ (_39365_, _02092_, _42882_);
  and _53218_ (_02093_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  and _53219_ (_02094_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or _53220_ (_02095_, _02094_, _02093_);
  and _53221_ (_39366_, _02095_, _42882_);
  and _53222_ (_02096_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  and _53223_ (_02097_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or _53224_ (_02098_, _02097_, _02096_);
  and _53225_ (_39367_, _02098_, _42882_);
  and _53226_ (_02099_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  and _53227_ (_02100_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  or _53228_ (_02101_, _02100_, _02099_);
  and _53229_ (_39368_, _02101_, _42882_);
  and _53230_ (_02102_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  and _53231_ (_02103_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _53232_ (_02104_, _02103_, _02102_);
  and _53233_ (_39370_, _02104_, _42882_);
  and _53234_ (_02105_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  and _53235_ (_02106_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or _53236_ (_02107_, _02106_, _02105_);
  and _53237_ (_39371_, _02107_, _42882_);
  and _53238_ (_02110_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  and _53239_ (_02112_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or _53240_ (_02114_, _02112_, _02110_);
  and _53241_ (_39372_, _02114_, _42882_);
  and _53242_ (_02117_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  and _53243_ (_02119_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or _53244_ (_02121_, _02119_, _02117_);
  and _53245_ (_39373_, _02121_, _42882_);
  and _53246_ (_02124_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  and _53247_ (_02126_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or _53248_ (_02128_, _02126_, _02124_);
  and _53249_ (_39374_, _02128_, _42882_);
  and _53250_ (_02131_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  and _53251_ (_02133_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  or _53252_ (_02135_, _02133_, _02131_);
  and _53253_ (_39375_, _02135_, _42882_);
  and _53254_ (_02138_, _01901_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  and _53255_ (_02140_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or _53256_ (_02142_, _02140_, _02138_);
  and _53257_ (_39376_, _02142_, _42882_);
  nor _53258_ (_39377_, _42476_, rst);
  and _53259_ (_39379_, _42398_, _42882_);
  nor _53260_ (_39380_, _42602_, rst);
  nor _53261_ (_39381_, _42444_, rst);
  nor _53262_ (_39382_, _42356_, rst);
  nor _53263_ (_39383_, _42564_, rst);
  and _53264_ (_39385_, _42505_, _42882_);
  and _53265_ (_39401_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _42882_);
  and _53266_ (_39402_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _42882_);
  and _53267_ (_39403_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _42882_);
  and _53268_ (_39404_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _42882_);
  and _53269_ (_39405_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _42882_);
  and _53270_ (_39407_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _42882_);
  and _53271_ (_39408_, \oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _42882_);
  not _53272_ (_02158_, _01450_);
  and _53273_ (_02159_, _02158_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _53274_ (_02160_, _01566_, _42465_);
  and _53275_ (_02161_, _01454_, _01505_);
  or _53276_ (_02162_, _02161_, _02160_);
  or _53277_ (_02163_, _01507_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _53278_ (_02164_, _01508_);
  and _53279_ (_02165_, _01560_, _02164_);
  and _53280_ (_02166_, _02165_, _02163_);
  or _53281_ (_02167_, _02166_, _02162_);
  or _53282_ (_02168_, _01585_, _01556_);
  and _53283_ (_02169_, _02168_, _31783_);
  or _53284_ (_02170_, _02169_, _02167_);
  and _53285_ (_02171_, _02170_, _01449_);
  or _53286_ (_02172_, _02171_, _02159_);
  and _53287_ (_39409_, _02172_, _42882_);
  and _53288_ (_02173_, _02158_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _53289_ (_02174_, _01566_, _42385_);
  and _53290_ (_02175_, _01454_, _01500_);
  or _53291_ (_02176_, _02175_, _02174_);
  or _53292_ (_02177_, _01510_, _01508_);
  not _53293_ (_02178_, _01511_);
  and _53294_ (_02179_, _01560_, _02178_);
  and _53295_ (_02180_, _02179_, _02177_);
  or _53296_ (_02181_, _02180_, _02176_);
  and _53297_ (_02182_, _02168_, _32469_);
  or _53298_ (_02183_, _02182_, _02181_);
  and _53299_ (_02184_, _02183_, _01449_);
  or _53300_ (_02185_, _02184_, _02173_);
  and _53301_ (_39410_, _02185_, _42882_);
  and _53302_ (_02186_, _02168_, _33165_);
  or _53303_ (_02187_, _01515_, _01513_);
  not _53304_ (_02188_, _01516_);
  and _53305_ (_02189_, _01560_, _02188_);
  nand _53306_ (_02190_, _02189_, _02187_);
  and _53307_ (_02191_, _01566_, _42590_);
  and _53308_ (_02192_, _01454_, _01495_);
  and _53309_ (_02193_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _53310_ (_02194_, _02193_, _02192_);
  nor _53311_ (_02195_, _02194_, _02191_);
  and _53312_ (_02196_, _02195_, _02190_);
  nand _53313_ (_02197_, _02196_, _01449_);
  or _53314_ (_02198_, _02197_, _02186_);
  not _53315_ (_02199_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _53316_ (_02200_, _01594_, _02199_);
  and _53317_ (_02201_, _01594_, _02199_);
  nor _53318_ (_02202_, _02201_, _02200_);
  or _53319_ (_02203_, _02202_, _01449_);
  and _53320_ (_02204_, _02203_, _42882_);
  and _53321_ (_39411_, _02204_, _02198_);
  and _53322_ (_02205_, _02168_, _33916_);
  or _53323_ (_02206_, _01493_, _01492_);
  or _53324_ (_02207_, _02206_, _01517_);
  nand _53325_ (_02208_, _02206_, _01517_);
  and _53326_ (_02209_, _02208_, _01560_);
  nand _53327_ (_02210_, _02209_, _02207_);
  and _53328_ (_02211_, _01566_, _42430_);
  and _53329_ (_02212_, _01454_, _01489_);
  and _53330_ (_02213_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _53331_ (_02214_, _02213_, _02212_);
  nor _53332_ (_02215_, _02214_, _02211_);
  and _53333_ (_02216_, _02215_, _02210_);
  nand _53334_ (_02217_, _02216_, _01449_);
  or _53335_ (_02218_, _02217_, _02205_);
  and _53336_ (_02219_, _02200_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _53337_ (_02220_, _02200_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _53338_ (_02221_, _02220_, _02219_);
  or _53339_ (_02222_, _02221_, _01449_);
  and _53340_ (_02223_, _02222_, _42882_);
  and _53341_ (_39412_, _02223_, _02218_);
  and _53342_ (_02224_, _02168_, _34678_);
  or _53343_ (_02225_, _01521_, _01519_);
  and _53344_ (_02226_, _01560_, _01522_);
  and _53345_ (_02227_, _02226_, _02225_);
  and _53346_ (_02228_, _01566_, _42337_);
  and _53347_ (_02229_, _01454_, _01484_);
  and _53348_ (_02230_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _53349_ (_02231_, _02230_, _02229_);
  or _53350_ (_02232_, _02231_, _02228_);
  nor _53351_ (_02233_, _02232_, _02227_);
  nand _53352_ (_02234_, _02233_, _01449_);
  or _53353_ (_02235_, _02234_, _02224_);
  and _53354_ (_02236_, _02219_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _53355_ (_02237_, _02219_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _53356_ (_02238_, _02237_, _02236_);
  or _53357_ (_02239_, _02238_, _01449_);
  and _53358_ (_02240_, _02239_, _42882_);
  and _53359_ (_39413_, _02240_, _02235_);
  and _53360_ (_02241_, _02168_, _35472_);
  or _53361_ (_02242_, _01482_, _01481_);
  nand _53362_ (_02243_, _02242_, _01523_);
  or _53363_ (_02244_, _02242_, _01523_);
  and _53364_ (_02245_, _02244_, _01560_);
  nand _53365_ (_02246_, _02245_, _02243_);
  and _53366_ (_02247_, _01566_, _42552_);
  and _53367_ (_02248_, _01454_, _01478_);
  and _53368_ (_02249_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _53369_ (_02250_, _02249_, _02248_);
  nor _53370_ (_02251_, _02250_, _02247_);
  and _53371_ (_02252_, _02251_, _02246_);
  nand _53372_ (_02253_, _02252_, _01449_);
  or _53373_ (_02254_, _02253_, _02241_);
  nor _53374_ (_02255_, _02236_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _53375_ (_02256_, _02255_, _01599_);
  or _53376_ (_02257_, _02256_, _01449_);
  and _53377_ (_02258_, _02257_, _42882_);
  and _53378_ (_39414_, _02258_, _02254_);
  nor _53379_ (_02259_, _01599_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _53380_ (_02260_, _01599_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _53381_ (_02261_, _02260_, _02259_);
  or _53382_ (_02262_, _02261_, _01449_);
  and _53383_ (_02263_, _02262_, _42882_);
  and _53384_ (_02264_, _02168_, _36190_);
  and _53385_ (_02265_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _53386_ (_02266_, _01454_, _01471_);
  and _53387_ (_02267_, _01566_, _42524_);
  or _53388_ (_02268_, _02267_, _02266_);
  or _53389_ (_02269_, _02268_, _02265_);
  or _53390_ (_02270_, _01525_, _01476_);
  not _53391_ (_02271_, _01526_);
  and _53392_ (_02272_, _01560_, _02271_);
  and _53393_ (_02273_, _02272_, _02270_);
  nor _53394_ (_02274_, _02273_, _02269_);
  nand _53395_ (_02275_, _02274_, _01449_);
  or _53396_ (_02276_, _02275_, _02264_);
  and _53397_ (_39415_, _02276_, _02263_);
  and _53398_ (_02277_, _02168_, _30614_);
  or _53399_ (_02278_, _01468_, _01469_);
  or _53400_ (_02279_, _02278_, _01527_);
  nand _53401_ (_02280_, _02278_, _01527_);
  and _53402_ (_02281_, _02280_, _01560_);
  and _53403_ (_02282_, _02281_, _02279_);
  and _53404_ (_02283_, _01454_, _01463_);
  and _53405_ (_02284_, _01566_, _42267_);
  and _53406_ (_02285_, _38352_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _53407_ (_02286_, _02285_, _02284_);
  nor _53408_ (_02287_, _02286_, _02283_);
  nand _53409_ (_02288_, _02287_, _01449_);
  or _53410_ (_02289_, _02288_, _02282_);
  or _53411_ (_02290_, _02289_, _02277_);
  nor _53412_ (_02291_, _02260_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _53413_ (_02292_, _02260_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _53414_ (_02293_, _02292_, _02291_);
  or _53415_ (_02294_, _02293_, _01449_);
  and _53416_ (_02295_, _02294_, _42882_);
  and _53417_ (_39416_, _02295_, _02290_);
  nor _53418_ (_02296_, _01345_, _31782_);
  not _53419_ (_02297_, _38660_);
  and _53420_ (_02298_, _01556_, _02297_);
  and _53421_ (_02299_, _01529_, _38552_);
  nor _53422_ (_02300_, _01529_, _38552_);
  nor _53423_ (_02301_, _02300_, _02299_);
  nand _53424_ (_02302_, _02301_, _01535_);
  or _53425_ (_02303_, _02301_, _01535_);
  and _53426_ (_02304_, _02303_, _01560_);
  and _53427_ (_02305_, _02304_, _02302_);
  and _53428_ (_02306_, _01566_, _00689_);
  and _53429_ (_02307_, _01454_, _42465_);
  or _53430_ (_02308_, _02307_, _02306_);
  and _53431_ (_02309_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _53432_ (_02310_, _02309_, _02308_);
  nand _53433_ (_02311_, _02310_, _01449_);
  or _53434_ (_02312_, _02311_, _02305_);
  or _53435_ (_02313_, _02312_, _02298_);
  or _53436_ (_02314_, _02313_, _02296_);
  or _53437_ (_02315_, _02292_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand _53438_ (_02316_, _01601_, _01599_);
  and _53439_ (_02317_, _02316_, _02315_);
  or _53440_ (_02318_, _02317_, _01449_);
  and _53441_ (_02319_, _02318_, _42882_);
  and _53442_ (_39418_, _02319_, _02314_);
  nor _53443_ (_02320_, _01345_, _32458_);
  and _53444_ (_02321_, _01529_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _53445_ (_02322_, _02321_, _01535_);
  and _53446_ (_02323_, _01536_, _01465_);
  nor _53447_ (_02324_, _02323_, _02322_);
  nand _53448_ (_02325_, _02324_, _38558_);
  or _53449_ (_02326_, _02324_, _38558_);
  and _53450_ (_02327_, _02326_, _01560_);
  and _53451_ (_02328_, _02327_, _02325_);
  not _53452_ (_02329_, _38693_);
  nand _53453_ (_02330_, _01556_, _02329_);
  and _53454_ (_02331_, _01566_, _00656_);
  and _53455_ (_02332_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _53456_ (_02333_, _01454_, _42385_);
  or _53457_ (_02334_, _02333_, _02332_);
  nor _53458_ (_02335_, _02334_, _02331_);
  and _53459_ (_02336_, _02335_, _02330_);
  nand _53460_ (_02337_, _02336_, _01449_);
  or _53461_ (_02338_, _02337_, _02328_);
  or _53462_ (_02339_, _02338_, _02320_);
  nand _53463_ (_02340_, _02316_, _01681_);
  or _53464_ (_02341_, _02316_, _01681_);
  and _53465_ (_02342_, _02341_, _02340_);
  or _53466_ (_02343_, _02342_, _01449_);
  and _53467_ (_02344_, _02343_, _42882_);
  and _53468_ (_39419_, _02344_, _02339_);
  nor _53469_ (_02345_, _01345_, _33154_);
  and _53470_ (_02346_, _01537_, _01465_);
  and _53471_ (_02347_, _02322_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _53472_ (_02348_, _02347_, _02346_);
  nand _53473_ (_02349_, _02348_, _38563_);
  or _53474_ (_02350_, _02348_, _38563_);
  and _53475_ (_02351_, _02350_, _01560_);
  and _53476_ (_02352_, _02351_, _02349_);
  not _53477_ (_02353_, _38724_);
  and _53478_ (_02354_, _01556_, _02353_);
  and _53479_ (_02355_, _01566_, _00634_);
  and _53480_ (_02357_, _01454_, _42590_);
  or _53481_ (_02358_, _02357_, _02355_);
  and _53482_ (_02359_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _53483_ (_02360_, _02359_, _02358_);
  nor _53484_ (_02361_, _02360_, _02354_);
  nand _53485_ (_02362_, _02361_, _01449_);
  or _53486_ (_02363_, _02362_, _02352_);
  or _53487_ (_02364_, _02363_, _02345_);
  nor _53488_ (_02365_, _01603_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _53489_ (_02366_, _02365_, _01604_);
  or _53490_ (_02367_, _02366_, _01449_);
  and _53491_ (_02368_, _02367_, _42882_);
  and _53492_ (_39420_, _02368_, _02364_);
  nor _53493_ (_02369_, _01345_, _33906_);
  and _53494_ (_02370_, _01530_, _01535_);
  and _53495_ (_02371_, _01538_, _01465_);
  nor _53496_ (_02372_, _02371_, _02370_);
  nand _53497_ (_02373_, _02372_, _38548_);
  or _53498_ (_02374_, _02372_, _38548_);
  and _53499_ (_02375_, _02374_, _01560_);
  and _53500_ (_02376_, _02375_, _02373_);
  not _53501_ (_02377_, _38756_);
  and _53502_ (_02378_, _01556_, _02377_);
  and _53503_ (_02379_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _53504_ (_02380_, _01573_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _53505_ (_02381_, _02380_, _01574_);
  and _53506_ (_02382_, _02381_, _01566_);
  and _53507_ (_02383_, _01454_, _42430_);
  or _53508_ (_02384_, _02383_, _02382_);
  or _53509_ (_02385_, _02384_, _02379_);
  nor _53510_ (_02386_, _02385_, _02378_);
  nand _53511_ (_02387_, _02386_, _01449_);
  or _53512_ (_02388_, _02387_, _02376_);
  or _53513_ (_02389_, _02388_, _02369_);
  nor _53514_ (_02390_, _01604_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor _53515_ (_02391_, _02390_, _01605_);
  or _53516_ (_02392_, _02391_, _01449_);
  and _53517_ (_02393_, _02392_, _42882_);
  and _53518_ (_39421_, _02393_, _02389_);
  nor _53519_ (_02394_, _01345_, _34667_);
  and _53520_ (_02395_, _01531_, _01535_);
  and _53521_ (_02396_, _01539_, _01465_);
  nor _53522_ (_02397_, _02396_, _02395_);
  nand _53523_ (_02398_, _02397_, _38569_);
  or _53524_ (_02399_, _02397_, _38569_);
  and _53525_ (_02400_, _02399_, _01560_);
  and _53526_ (_02401_, _02400_, _02398_);
  not _53527_ (_02402_, _38787_);
  nand _53528_ (_02403_, _01556_, _02402_);
  and _53529_ (_02404_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _53530_ (_02405_, _01574_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _53531_ (_02406_, _02405_, _01575_);
  and _53532_ (_02407_, _02406_, _01566_);
  and _53533_ (_02408_, _01454_, _42337_);
  or _53534_ (_02409_, _02408_, _02407_);
  nor _53535_ (_02410_, _02409_, _02404_);
  and _53536_ (_02411_, _02410_, _02403_);
  nand _53537_ (_02412_, _02411_, _01449_);
  or _53538_ (_02413_, _02412_, _02401_);
  or _53539_ (_02414_, _02413_, _02394_);
  nor _53540_ (_02415_, _01605_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _53541_ (_02416_, _02415_, _01606_);
  or _53542_ (_02417_, _02416_, _01449_);
  and _53543_ (_02418_, _02417_, _42882_);
  and _53544_ (_39422_, _02418_, _02414_);
  nor _53545_ (_02419_, _01345_, _35461_);
  and _53546_ (_02420_, _02395_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _53547_ (_02421_, _02396_, _38569_);
  nor _53548_ (_02422_, _02421_, _02420_);
  nand _53549_ (_02423_, _02422_, _38544_);
  or _53550_ (_02424_, _02422_, _38544_);
  and _53551_ (_02425_, _02424_, _01560_);
  and _53552_ (_02426_, _02425_, _02423_);
  not _53553_ (_02427_, _38821_);
  nand _53554_ (_02428_, _01556_, _02427_);
  and _53555_ (_02429_, _01454_, _42552_);
  nor _53556_ (_02430_, _01575_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor _53557_ (_02431_, _02430_, _01576_);
  and _53558_ (_02432_, _02431_, _01566_);
  and _53559_ (_02433_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _53560_ (_02434_, _02433_, _02432_);
  nor _53561_ (_02435_, _02434_, _02429_);
  and _53562_ (_02436_, _02435_, _02428_);
  nand _53563_ (_02437_, _02436_, _01449_);
  or _53564_ (_02438_, _02437_, _02426_);
  or _53565_ (_02439_, _02438_, _02419_);
  nor _53566_ (_02440_, _01606_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _53567_ (_02441_, _02440_, _01607_);
  or _53568_ (_02442_, _02441_, _01449_);
  and _53569_ (_02443_, _02442_, _42882_);
  and _53570_ (_39423_, _02443_, _02439_);
  nor _53571_ (_02444_, _01345_, _36179_);
  nor _53572_ (_02445_, _01543_, _38540_);
  and _53573_ (_02446_, _01543_, _38540_);
  or _53574_ (_02447_, _02446_, _02445_);
  and _53575_ (_02448_, _02447_, _01560_);
  and _53576_ (_02449_, _01556_, _38847_);
  or _53577_ (_02450_, _01576_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _53578_ (_02451_, _02450_, _01577_);
  and _53579_ (_02452_, _02451_, _01566_);
  and _53580_ (_02453_, _01585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and _53581_ (_02454_, _01454_, _42524_);
  or _53582_ (_02455_, _02454_, _02453_);
  or _53583_ (_02456_, _02455_, _02452_);
  nor _53584_ (_02457_, _02456_, _02449_);
  nand _53585_ (_02458_, _02457_, _01449_);
  or _53586_ (_02459_, _02458_, _02448_);
  or _53587_ (_02460_, _02459_, _02444_);
  nor _53588_ (_02461_, _01607_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _53589_ (_02462_, _02461_, _01608_);
  or _53590_ (_02463_, _02462_, _01449_);
  and _53591_ (_02464_, _02463_, _42882_);
  and _53592_ (_39424_, _02464_, _02460_);
  and _53593_ (_02465_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor _53594_ (_02466_, _01803_, _01801_);
  nor _53595_ (_02467_, _02466_, _01804_);
  or _53596_ (_02468_, _02467_, _01618_);
  or _53597_ (_02469_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _53598_ (_02470_, _02469_, _01835_);
  and _53599_ (_02471_, _02470_, _02468_);
  or _53600_ (_39425_, _02471_, _02465_);
  or _53601_ (_02472_, _01806_, _01804_);
  and _53602_ (_02473_, _02472_, _01807_);
  or _53603_ (_02474_, _02473_, _01618_);
  or _53604_ (_02475_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _53605_ (_02476_, _02475_, _01835_);
  and _53606_ (_02477_, _02476_, _02474_);
  and _53607_ (_02478_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _53608_ (_39426_, _02478_, _02477_);
  or _53609_ (_02479_, _01811_, _01809_);
  nor _53610_ (_02480_, _01812_, _01618_);
  and _53611_ (_02481_, _02480_, _02479_);
  nor _53612_ (_02482_, _01617_, _01941_);
  or _53613_ (_02483_, _02482_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _53614_ (_02484_, _02483_, _02481_);
  or _53615_ (_02485_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _36418_);
  and _53616_ (_02486_, _02485_, _42882_);
  and _53617_ (_39427_, _02486_, _02484_);
  and _53618_ (_02487_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _53619_ (_02488_, _01812_, _01702_);
  nor _53620_ (_02489_, _02488_, _01813_);
  or _53621_ (_02490_, _02489_, _01618_);
  or _53622_ (_02491_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _53623_ (_02492_, _02491_, _01835_);
  and _53624_ (_02493_, _02492_, _02490_);
  or _53625_ (_39429_, _02493_, _02487_);
  and _53626_ (_02494_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _53627_ (_02495_, _01816_, _01813_);
  nor _53628_ (_02496_, _02495_, _01817_);
  or _53629_ (_02497_, _02496_, _01618_);
  or _53630_ (_02498_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _53631_ (_02499_, _02498_, _01835_);
  and _53632_ (_02500_, _02499_, _02497_);
  or _53633_ (_39430_, _02500_, _02494_);
  and _53634_ (_02501_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _53635_ (_02502_, _01817_, _01697_);
  nor _53636_ (_02503_, _02502_, _01818_);
  or _53637_ (_02504_, _02503_, _01618_);
  or _53638_ (_02505_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _53639_ (_02506_, _02505_, _01835_);
  and _53640_ (_02507_, _02506_, _02504_);
  or _53641_ (_39431_, _02507_, _02501_);
  nor _53642_ (_02508_, _01818_, _01693_);
  nor _53643_ (_02509_, _02508_, _01819_);
  or _53644_ (_02510_, _02509_, _01618_);
  or _53645_ (_02511_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _53646_ (_02512_, _02511_, _01835_);
  and _53647_ (_02513_, _02512_, _02510_);
  and _53648_ (_02514_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _53649_ (_39432_, _02514_, _02513_);
  nor _53650_ (_02515_, _01819_, _01691_);
  nor _53651_ (_02516_, _02515_, _01820_);
  or _53652_ (_02517_, _02516_, _01618_);
  or _53653_ (_02518_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _53654_ (_02519_, _02518_, _01835_);
  and _53655_ (_02520_, _02519_, _02517_);
  and _53656_ (_02521_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _53657_ (_39433_, _02521_, _02520_);
  and _53658_ (_02522_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _53659_ (_02523_, _01822_, _01820_);
  nor _53660_ (_02524_, _02523_, _01823_);
  or _53661_ (_02525_, _02524_, _01618_);
  or _53662_ (_02526_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _53663_ (_02527_, _02526_, _01835_);
  and _53664_ (_02528_, _02527_, _02525_);
  or _53665_ (_39434_, _02528_, _02522_);
  and _53666_ (_02529_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _53667_ (_02530_, _01823_, _01687_);
  nor _53668_ (_02531_, _02530_, _01824_);
  or _53669_ (_02532_, _02531_, _01618_);
  or _53670_ (_02533_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _53671_ (_02534_, _02533_, _01835_);
  and _53672_ (_02535_, _02534_, _02532_);
  or _53673_ (_39435_, _02535_, _02529_);
  nor _53674_ (_02536_, _01824_, _01680_);
  nor _53675_ (_02537_, _02536_, _01825_);
  or _53676_ (_02538_, _02537_, _01618_);
  or _53677_ (_02539_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _53678_ (_02540_, _02539_, _01835_);
  and _53679_ (_02541_, _02540_, _02538_);
  and _53680_ (_02543_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _53681_ (_39436_, _02543_, _02541_);
  nor _53682_ (_02544_, _01825_, _01676_);
  nor _53683_ (_02545_, _02544_, _01826_);
  or _53684_ (_02546_, _02545_, _01618_);
  or _53685_ (_02547_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _53686_ (_02548_, _02547_, _01835_);
  and _53687_ (_02549_, _02548_, _02546_);
  and _53688_ (_02550_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _53689_ (_39437_, _02550_, _02549_);
  nor _53690_ (_02551_, _01826_, _01673_);
  nor _53691_ (_02552_, _02551_, _01827_);
  or _53692_ (_02553_, _02552_, _01618_);
  or _53693_ (_02554_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _53694_ (_02555_, _02554_, _01835_);
  and _53695_ (_02556_, _02555_, _02553_);
  and _53696_ (_02557_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _53697_ (_39438_, _02557_, _02556_);
  and _53698_ (_02558_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _53699_ (_02559_, _01827_, _01670_);
  nor _53700_ (_02560_, _02559_, _01828_);
  or _53701_ (_02561_, _02560_, _01618_);
  or _53702_ (_02562_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _53703_ (_02564_, _02562_, _01835_);
  and _53704_ (_02565_, _02564_, _02561_);
  or _53705_ (_39440_, _02565_, _02558_);
  or _53706_ (_02566_, _01828_, _01668_);
  and _53707_ (_02567_, _02566_, _01829_);
  or _53708_ (_02568_, _02567_, _01618_);
  or _53709_ (_02569_, _01617_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _53710_ (_02570_, _02569_, _01835_);
  and _53711_ (_02571_, _02570_, _02568_);
  and _53712_ (_02572_, _01614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _53713_ (_39441_, _02572_, _02571_);
  and _53714_ (_02574_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _53715_ (_02575_, _02574_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _53716_ (_39442_, _02575_, _42882_);
  and _53717_ (_02576_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _53718_ (_02577_, _02576_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _53719_ (_39443_, _02577_, _42882_);
  and _53720_ (_02578_, _01846_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  or _53721_ (_02579_, _02578_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _53722_ (_39444_, _02579_, _42882_);
  and _53723_ (_02580_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _53724_ (_02581_, _02580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _53725_ (_39445_, _02581_, _42882_);
  and _53726_ (_02582_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _53727_ (_02583_, _02582_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _53728_ (_39446_, _02583_, _42882_);
  and _53729_ (_02584_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _53730_ (_02585_, _02584_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _53731_ (_39447_, _02585_, _42882_);
  and _53732_ (_02586_, _01847_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or _53733_ (_02587_, _02586_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _53734_ (_39448_, _02587_, _42882_);
  nor _53735_ (_02588_, _01800_, _42250_);
  nand _53736_ (_02589_, _02588_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or _53737_ (_02590_, _02588_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _53738_ (_02591_, _02590_, _01835_);
  and _53739_ (_39449_, _02591_, _02589_);
  or _53740_ (_02592_, _01858_, _01856_);
  and _53741_ (_02593_, _02592_, _01859_);
  or _53742_ (_02594_, _02593_, _42250_);
  or _53743_ (_02595_, _36450_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _53744_ (_02596_, _02595_, _01835_);
  and _53745_ (_39450_, _02596_, _02594_);
  and _53746_ (_02597_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  and _53747_ (_02598_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [0]);
  and _53748_ (_02599_, _02598_, _39078_);
  or _53749_ (_39466_, _02599_, _02597_);
  and _53750_ (_02600_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  and _53751_ (_02601_, _02033_, _39078_);
  or _53752_ (_39467_, _02601_, _02600_);
  and _53753_ (_02602_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  and _53754_ (_02603_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [2]);
  and _53755_ (_02604_, _02603_, _39078_);
  or _53756_ (_39468_, _02604_, _02602_);
  and _53757_ (_02605_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  and _53758_ (_02606_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [3]);
  and _53759_ (_02607_, _02606_, _39078_);
  or _53760_ (_39469_, _02607_, _02605_);
  and _53761_ (_02608_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [4]);
  and _53762_ (_02609_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [4]);
  and _53763_ (_02610_, _02609_, _39078_);
  or _53764_ (_39470_, _02610_, _02608_);
  and _53765_ (_02611_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _53766_ (_02612_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [5]);
  and _53767_ (_02613_, _02612_, _39078_);
  or _53768_ (_39472_, _02613_, _02611_);
  and _53769_ (_02614_, _01879_, \oc8051_top_1.oc8051_memory_interface1.cdata [6]);
  and _53770_ (_02615_, \oc8051_top_1.oc8051_rom1.ea_int , \oc8051_top_1.oc8051_rom1.data_o [6]);
  and _53771_ (_02616_, _02615_, _39078_);
  or _53772_ (_39473_, _02616_, _02614_);
  and _53773_ (_39474_, _01887_, _42882_);
  nor _53774_ (_39475_, _01897_, rst);
  and _53775_ (_39476_, _01893_, _42882_);
  and _53776_ (_02617_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _53777_ (_02618_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  or _53778_ (_02619_, _02618_, _02617_);
  and _53779_ (_39477_, _02619_, _42882_);
  and _53780_ (_02620_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _53781_ (_02621_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  or _53782_ (_02622_, _02621_, _02620_);
  and _53783_ (_39478_, _02622_, _42882_);
  and _53784_ (_02623_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _53785_ (_02624_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  or _53786_ (_02625_, _02624_, _02623_);
  and _53787_ (_39479_, _02625_, _42882_);
  and _53788_ (_02626_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _53789_ (_02627_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  or _53790_ (_02628_, _02627_, _02626_);
  and _53791_ (_39480_, _02628_, _42882_);
  and _53792_ (_02629_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _53793_ (_02630_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  or _53794_ (_02631_, _02630_, _02629_);
  and _53795_ (_39481_, _02631_, _42882_);
  and _53796_ (_02632_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _53797_ (_02633_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  or _53798_ (_02634_, _02633_, _02632_);
  and _53799_ (_39483_, _02634_, _42882_);
  and _53800_ (_02635_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _53801_ (_02636_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  or _53802_ (_02637_, _02636_, _02635_);
  and _53803_ (_39484_, _02637_, _42882_);
  and _53804_ (_02638_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _53805_ (_02639_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  or _53806_ (_02640_, _02639_, _02638_);
  and _53807_ (_39485_, _02640_, _42882_);
  and _53808_ (_02641_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _53809_ (_02642_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  or _53810_ (_02643_, _02642_, _02641_);
  and _53811_ (_39486_, _02643_, _42882_);
  and _53812_ (_02644_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _53813_ (_02645_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  or _53814_ (_02646_, _02645_, _02644_);
  and _53815_ (_39487_, _02646_, _42882_);
  and _53816_ (_02647_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _53817_ (_02648_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  or _53818_ (_02649_, _02648_, _02647_);
  and _53819_ (_39488_, _02649_, _42882_);
  and _53820_ (_02650_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _53821_ (_02651_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  or _53822_ (_02652_, _02651_, _02650_);
  and _53823_ (_39489_, _02652_, _42882_);
  and _53824_ (_02653_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _53825_ (_02654_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  or _53826_ (_02655_, _02654_, _02653_);
  and _53827_ (_39490_, _02655_, _42882_);
  and _53828_ (_02656_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _53829_ (_02657_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  or _53830_ (_02658_, _02657_, _02656_);
  and _53831_ (_39491_, _02658_, _42882_);
  and _53832_ (_02659_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and _53833_ (_02660_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or _53834_ (_02661_, _02660_, _02659_);
  and _53835_ (_39492_, _02661_, _42882_);
  and _53836_ (_02662_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _53837_ (_02663_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  or _53838_ (_02664_, _02663_, _02662_);
  and _53839_ (_39494_, _02664_, _42882_);
  and _53840_ (_02665_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _53841_ (_02666_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  or _53842_ (_02667_, _02666_, _02665_);
  and _53843_ (_39495_, _02667_, _42882_);
  and _53844_ (_02668_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _53845_ (_02669_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or _53846_ (_02670_, _02669_, _02668_);
  and _53847_ (_39496_, _02670_, _42882_);
  and _53848_ (_02671_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _53849_ (_02672_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or _53850_ (_02673_, _02672_, _02671_);
  and _53851_ (_39497_, _02673_, _42882_);
  and _53852_ (_02674_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _53853_ (_02675_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or _53854_ (_02676_, _02675_, _02674_);
  and _53855_ (_39498_, _02676_, _42882_);
  and _53856_ (_02677_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _53857_ (_02678_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or _53858_ (_02679_, _02678_, _02677_);
  and _53859_ (_39499_, _02679_, _42882_);
  and _53860_ (_02680_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _53861_ (_02681_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or _53862_ (_02682_, _02681_, _02680_);
  and _53863_ (_39500_, _02682_, _42882_);
  and _53864_ (_02683_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _53865_ (_02684_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or _53866_ (_02685_, _02684_, _02683_);
  and _53867_ (_39501_, _02685_, _42882_);
  and _53868_ (_02686_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _53869_ (_02687_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or _53870_ (_02688_, _02687_, _02686_);
  and _53871_ (_39502_, _02688_, _42882_);
  and _53872_ (_02689_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _53873_ (_02690_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  or _53874_ (_02691_, _02690_, _02689_);
  and _53875_ (_39503_, _02691_, _42882_);
  and _53876_ (_02692_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _53877_ (_02693_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or _53878_ (_02694_, _02693_, _02692_);
  and _53879_ (_39505_, _02694_, _42882_);
  and _53880_ (_02696_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _53881_ (_02697_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or _53882_ (_02698_, _02697_, _02696_);
  and _53883_ (_39506_, _02698_, _42882_);
  and _53884_ (_02699_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _53885_ (_02700_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or _53886_ (_02701_, _02700_, _02699_);
  and _53887_ (_39507_, _02701_, _42882_);
  and _53888_ (_02702_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _53889_ (_02703_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or _53890_ (_02704_, _02703_, _02702_);
  and _53891_ (_39508_, _02704_, _42882_);
  and _53892_ (_02705_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _53893_ (_02706_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or _53894_ (_02707_, _02706_, _02705_);
  and _53895_ (_39509_, _02707_, _42882_);
  and _53896_ (_02708_, _01901_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _53897_ (_02709_, _01903_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or _53898_ (_02710_, _02709_, _02708_);
  and _53899_ (_39510_, _02710_, _42882_);
  and _53900_ (_02711_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53901_ (_02712_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _53902_ (_02713_, _02712_, _02711_);
  and _53903_ (_39511_, _02713_, _42882_);
  and _53904_ (_02714_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53905_ (_02715_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _53906_ (_02716_, _02715_, _02714_);
  and _53907_ (_39512_, _02716_, _42882_);
  and _53908_ (_02717_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53909_ (_02718_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _53910_ (_02719_, _02718_, _02717_);
  and _53911_ (_39513_, _02719_, _42882_);
  and _53912_ (_02720_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53913_ (_02721_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _53914_ (_02722_, _02721_, _02720_);
  and _53915_ (_39514_, _02722_, _42882_);
  and _53916_ (_02723_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53917_ (_02724_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _53918_ (_02725_, _02724_, _02723_);
  and _53919_ (_39516_, _02725_, _42882_);
  and _53920_ (_02726_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53921_ (_02727_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _53922_ (_02728_, _02727_, _02726_);
  and _53923_ (_39517_, _02728_, _42882_);
  and _53924_ (_02729_, \oc8051_top_1.oc8051_memory_interface1.ddat_o [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _53925_ (_02730_, _01911_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _53926_ (_02731_, _02730_, _02729_);
  and _53927_ (_39518_, _02731_, _42882_);
  and _53928_ (_02732_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53929_ (_02733_, _42476_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53930_ (_02734_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _53931_ (_02735_, _02734_, _01910_);
  and _53932_ (_02736_, _02735_, _02733_);
  or _53933_ (_02737_, _02736_, _02732_);
  and _53934_ (_39519_, _02737_, _42882_);
  and _53935_ (_02738_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53936_ (_02739_, _42398_, _01917_);
  or _53937_ (_02740_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _53938_ (_02741_, _02740_, _01910_);
  and _53939_ (_02742_, _02741_, _02739_);
  or _53940_ (_02743_, _02742_, _02738_);
  and _53941_ (_39520_, _02743_, _42882_);
  and _53942_ (_02744_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53943_ (_02745_, _42602_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53944_ (_02746_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _53945_ (_02747_, _02746_, _01910_);
  and _53946_ (_02748_, _02747_, _02745_);
  or _53947_ (_02749_, _02748_, _02744_);
  and _53948_ (_39521_, _02749_, _42882_);
  and _53949_ (_02750_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53950_ (_02751_, _42444_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53951_ (_02752_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _53952_ (_02753_, _02752_, _01910_);
  and _53953_ (_02754_, _02753_, _02751_);
  or _53954_ (_02755_, _02754_, _02750_);
  and _53955_ (_39522_, _02755_, _42882_);
  and _53956_ (_02756_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53957_ (_02757_, _42356_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53958_ (_02758_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _53959_ (_02759_, _02758_, _01910_);
  and _53960_ (_02760_, _02759_, _02757_);
  or _53961_ (_02761_, _02760_, _02756_);
  and _53962_ (_39523_, _02761_, _42882_);
  and _53963_ (_02762_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nand _53964_ (_02763_, _42564_, \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  or _53965_ (_02764_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _53966_ (_02765_, _02764_, _01910_);
  and _53967_ (_02766_, _02765_, _02763_);
  or _53968_ (_02767_, _02766_, _02762_);
  and _53969_ (_39524_, _02767_, _42882_);
  and _53970_ (_02768_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53971_ (_02769_, _42505_, _01917_);
  or _53972_ (_02770_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _53973_ (_02771_, _02770_, _01910_);
  and _53974_ (_02772_, _02771_, _02769_);
  or _53975_ (_02773_, _02772_, _02768_);
  and _53976_ (_39525_, _02773_, _42882_);
  and _53977_ (_02774_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53978_ (_02775_, _42300_, _01917_);
  or _53979_ (_02776_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _53980_ (_02777_, _02776_, _01910_);
  and _53981_ (_02778_, _02777_, _02775_);
  or _53982_ (_02779_, _02778_, _02774_);
  and _53983_ (_39527_, _02779_, _42882_);
  and _53984_ (_02780_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _53985_ (_02781_, _02780_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53986_ (_02782_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _01910_);
  and _53987_ (_02783_, _02782_, _42882_);
  and _53988_ (_39528_, _02783_, _02781_);
  and _53989_ (_02784_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _53990_ (_02785_, _02784_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53991_ (_02786_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _01910_);
  and _53992_ (_02787_, _02786_, _42882_);
  and _53993_ (_39529_, _02787_, _02785_);
  and _53994_ (_02788_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _53995_ (_02789_, _02788_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _53996_ (_02790_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _01910_);
  and _53997_ (_02791_, _02790_, _42882_);
  and _53998_ (_39530_, _02791_, _02789_);
  and _53999_ (_02792_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _54000_ (_02793_, _02792_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54001_ (_02794_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _01910_);
  and _54002_ (_02795_, _02794_, _42882_);
  and _54003_ (_39531_, _02795_, _02793_);
  and _54004_ (_02797_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _54005_ (_02798_, _02797_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54006_ (_02799_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _01910_);
  and _54007_ (_02800_, _02799_, _42882_);
  and _54008_ (_39532_, _02800_, _02798_);
  and _54009_ (_02802_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _54010_ (_02803_, _02802_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54011_ (_02804_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _01910_);
  and _54012_ (_02805_, _02804_, _42882_);
  and _54013_ (_39533_, _02805_, _02803_);
  and _54014_ (_02807_, _01917_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _54015_ (_02808_, _02807_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  or _54016_ (_02809_, \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _01910_);
  and _54017_ (_02810_, _02809_, _42882_);
  and _54018_ (_39534_, _02810_, _02808_);
  nand _54019_ (_02812_, _01924_, _31782_);
  or _54020_ (_02813_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _54021_ (_02814_, _02813_, _42882_);
  and _54022_ (_39535_, _02814_, _02812_);
  nand _54023_ (_02816_, _01924_, _32458_);
  or _54024_ (_02817_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _54025_ (_02818_, _02817_, _42882_);
  and _54026_ (_39536_, _02818_, _02816_);
  nand _54027_ (_02819_, _01924_, _33154_);
  or _54028_ (_02821_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _54029_ (_02822_, _02821_, _42882_);
  and _54030_ (_39538_, _02822_, _02819_);
  nand _54031_ (_02823_, _01924_, _33906_);
  or _54032_ (_02824_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _54033_ (_02826_, _02824_, _42882_);
  and _54034_ (_39539_, _02826_, _02823_);
  nand _54035_ (_02828_, _01924_, _34667_);
  or _54036_ (_02829_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [4]);
  and _54037_ (_02830_, _02829_, _42882_);
  and _54038_ (_39540_, _02830_, _02828_);
  nand _54039_ (_02831_, _01924_, _35461_);
  or _54040_ (_02833_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [5]);
  and _54041_ (_02834_, _02833_, _42882_);
  and _54042_ (_39541_, _02834_, _02831_);
  nand _54043_ (_02836_, _01924_, _36179_);
  or _54044_ (_02837_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [6]);
  and _54045_ (_02839_, _02837_, _42882_);
  and _54046_ (_39542_, _02839_, _02836_);
  nand _54047_ (_02840_, _01924_, _30603_);
  or _54048_ (_02842_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [7]);
  and _54049_ (_02843_, _02842_, _42882_);
  and _54050_ (_39543_, _02843_, _02840_);
  nand _54051_ (_02846_, _01924_, _38660_);
  or _54052_ (_02847_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [8]);
  and _54053_ (_02848_, _02847_, _42882_);
  and _54054_ (_39544_, _02848_, _02846_);
  nand _54055_ (_02850_, _01924_, _38693_);
  or _54056_ (_02851_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [9]);
  and _54057_ (_02853_, _02851_, _42882_);
  and _54058_ (_39545_, _02853_, _02850_);
  nand _54059_ (_02854_, _01924_, _38724_);
  or _54060_ (_02856_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [10]);
  and _54061_ (_02857_, _02856_, _42882_);
  and _54062_ (_39546_, _02857_, _02854_);
  nand _54063_ (_02859_, _01924_, _38756_);
  or _54064_ (_02860_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [11]);
  and _54065_ (_02861_, _02860_, _42882_);
  and _54066_ (_39547_, _02861_, _02859_);
  nand _54067_ (_02862_, _01924_, _38787_);
  or _54068_ (_02863_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [12]);
  and _54069_ (_02865_, _02863_, _42882_);
  and _54070_ (_39549_, _02865_, _02862_);
  nand _54071_ (_02867_, _01924_, _38821_);
  or _54072_ (_02869_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [13]);
  and _54073_ (_02870_, _02869_, _42882_);
  and _54074_ (_39550_, _02870_, _02867_);
  not _54075_ (_02872_, _01924_);
  or _54076_ (_02873_, _02872_, _38847_);
  or _54077_ (_02874_, _01924_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [14]);
  and _54078_ (_02876_, _02874_, _42882_);
  and _54079_ (_39551_, _02876_, _02873_);
  nor _54080_ (_39760_, _42319_, rst);
  and _54081_ (_02879_, _42275_, _39022_);
  nand _54082_ (_02880_, _02879_, _38485_);
  or _54083_ (_02881_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _54084_ (_02883_, _02881_, _42882_);
  and _54085_ (_39762_, _02883_, _02880_);
  and _54086_ (_02884_, _42275_, _39280_);
  nand _54087_ (_02886_, _02884_, _38485_);
  or _54088_ (_02887_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _54089_ (_02889_, _02887_, _42882_);
  and _54090_ (_39763_, _02889_, _02886_);
  and _54091_ (_02891_, _42275_, _27045_);
  nor _54092_ (_02892_, _02884_, _02891_);
  and _54093_ (_02893_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _54094_ (_02895_, _27045_, _27714_);
  not _54095_ (_02896_, _02895_);
  nor _54096_ (_02897_, _02896_, _38485_);
  and _54097_ (_02899_, _33329_, _27703_);
  and _54098_ (_02900_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  or _54099_ (_02901_, _02900_, _02897_);
  and _54100_ (_02903_, _02901_, _42275_);
  or _54101_ (_02904_, _02903_, _02893_);
  and _54102_ (_39764_, _02904_, _42882_);
  and _54103_ (_02906_, _42275_, _41396_);
  nand _54104_ (_02907_, _02906_, _38485_);
  or _54105_ (_02908_, _02906_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _54106_ (_02910_, _02908_, _42882_);
  and _54107_ (_39765_, _02910_, _02907_);
  nand _54108_ (_02911_, _02879_, _38464_);
  or _54109_ (_02913_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _54110_ (_02915_, _02913_, _42882_);
  and _54111_ (_39792_, _02915_, _02911_);
  nand _54112_ (_02917_, _02879_, _38456_);
  or _54113_ (_02918_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _54114_ (_02920_, _02918_, _42882_);
  and _54115_ (_39793_, _02920_, _02917_);
  nand _54116_ (_02921_, _02879_, _38449_);
  or _54117_ (_02922_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _54118_ (_02923_, _02922_, _42882_);
  and _54119_ (_39794_, _02923_, _02921_);
  nand _54120_ (_02925_, _02879_, _38442_);
  or _54121_ (_02927_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _54122_ (_02928_, _02927_, _42882_);
  and _54123_ (_39795_, _02928_, _02925_);
  nand _54124_ (_02930_, _02879_, _38434_);
  or _54125_ (_02931_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _54126_ (_02932_, _02931_, _42882_);
  and _54127_ (_39796_, _02932_, _02930_);
  nand _54128_ (_02934_, _02879_, _38428_);
  or _54129_ (_02935_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _54130_ (_02938_, _02935_, _42882_);
  and _54131_ (_39797_, _02938_, _02934_);
  nand _54132_ (_02939_, _02879_, _38420_);
  or _54133_ (_02941_, _02879_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _54134_ (_02942_, _02941_, _42882_);
  and _54135_ (_39798_, _02942_, _02939_);
  nand _54136_ (_02944_, _02884_, _38464_);
  or _54137_ (_02945_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _54138_ (_02946_, _02945_, _42882_);
  and _54139_ (_39799_, _02946_, _02944_);
  nand _54140_ (_02949_, _02884_, _38456_);
  or _54141_ (_02951_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _54142_ (_02952_, _02951_, _42882_);
  and _54143_ (_39800_, _02952_, _02949_);
  nand _54144_ (_02953_, _02884_, _38449_);
  or _54145_ (_02955_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _54146_ (_02956_, _02955_, _42882_);
  and _54147_ (_39801_, _02956_, _02953_);
  nand _54148_ (_02958_, _02884_, _38442_);
  or _54149_ (_02959_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _54150_ (_02961_, _02959_, _42882_);
  and _54151_ (_39803_, _02961_, _02958_);
  nand _54152_ (_02963_, _02884_, _38434_);
  or _54153_ (_02964_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _54154_ (_02966_, _02964_, _42882_);
  and _54155_ (_39804_, _02966_, _02963_);
  nand _54156_ (_02967_, _02884_, _38428_);
  or _54157_ (_02969_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _54158_ (_02970_, _02969_, _42882_);
  and _54159_ (_39805_, _02970_, _02967_);
  nand _54160_ (_02973_, _02884_, _38420_);
  or _54161_ (_02974_, _02884_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _54162_ (_02975_, _02974_, _42882_);
  and _54163_ (_39806_, _02975_, _02973_);
  not _54164_ (_02977_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _54165_ (_02979_, _42275_, _02895_);
  nor _54166_ (_02980_, _02979_, _02977_);
  and _54167_ (_02981_, _02979_, _38465_);
  or _54168_ (_02982_, _02981_, _02980_);
  and _54169_ (_39807_, _02982_, _42882_);
  and _54170_ (_02985_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _54171_ (_02986_, _02896_, _38456_);
  and _54172_ (_02988_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or _54173_ (_02989_, _02988_, _02986_);
  and _54174_ (_02990_, _02989_, _42275_);
  or _54175_ (_02992_, _02990_, _02985_);
  and _54176_ (_39808_, _02992_, _42882_);
  and _54177_ (_02993_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor _54178_ (_02995_, _02896_, _38449_);
  and _54179_ (_02996_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or _54180_ (_02998_, _02996_, _02995_);
  and _54181_ (_03000_, _02998_, _42275_);
  or _54182_ (_03001_, _03000_, _02993_);
  and _54183_ (_39809_, _03001_, _42882_);
  and _54184_ (_03003_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor _54185_ (_03004_, _02896_, _38442_);
  and _54186_ (_03005_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or _54187_ (_03007_, _03005_, _03004_);
  and _54188_ (_03008_, _03007_, _42275_);
  or _54189_ (_03010_, _03008_, _03003_);
  and _54190_ (_39810_, _03010_, _42882_);
  and _54191_ (_03012_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor _54192_ (_03013_, _02896_, _38434_);
  and _54193_ (_03015_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or _54194_ (_03016_, _03015_, _03013_);
  and _54195_ (_03017_, _03016_, _42275_);
  or _54196_ (_03019_, _03017_, _03012_);
  and _54197_ (_39811_, _03019_, _42882_);
  and _54198_ (_03020_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor _54199_ (_03022_, _02896_, _38428_);
  and _54200_ (_03023_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or _54201_ (_03024_, _03023_, _03022_);
  and _54202_ (_03026_, _03024_, _42275_);
  or _54203_ (_03027_, _03026_, _03020_);
  and _54204_ (_39812_, _03027_, _42882_);
  and _54205_ (_03029_, _02892_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor _54206_ (_03030_, _02896_, _38420_);
  and _54207_ (_03031_, _02899_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _54208_ (_03033_, _03031_, _03030_);
  and _54209_ (_03034_, _03033_, _42275_);
  or _54210_ (_03035_, _03034_, _03029_);
  and _54211_ (_39814_, _03035_, _42882_);
  not _54212_ (_03037_, _02906_);
  nor _54213_ (_03039_, _03037_, _38464_);
  and _54214_ (_03040_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or _54215_ (_03041_, _03040_, _03039_);
  and _54216_ (_39815_, _03041_, _42882_);
  nor _54217_ (_03042_, _03037_, _38456_);
  and _54218_ (_03043_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or _54219_ (_03044_, _03043_, _03042_);
  and _54220_ (_39816_, _03044_, _42882_);
  nand _54221_ (_03046_, _02906_, _38449_);
  or _54222_ (_03047_, _02906_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _54223_ (_03049_, _03047_, _42882_);
  and _54224_ (_39817_, _03049_, _03046_);
  nor _54225_ (_03050_, _03037_, _38442_);
  and _54226_ (_03052_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or _54227_ (_03053_, _03052_, _03050_);
  and _54228_ (_39818_, _03053_, _42882_);
  nand _54229_ (_03055_, _02906_, _38434_);
  or _54230_ (_03056_, _02906_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and _54231_ (_03057_, _03056_, _42882_);
  and _54232_ (_39819_, _03057_, _03055_);
  nand _54233_ (_03059_, _02906_, _38428_);
  or _54234_ (_03060_, _02906_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and _54235_ (_03062_, _03060_, _42882_);
  and _54236_ (_39820_, _03062_, _03059_);
  nor _54237_ (_03063_, _03037_, _38420_);
  and _54238_ (_03065_, _03037_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  or _54239_ (_03066_, _03065_, _03063_);
  and _54240_ (_39821_, _03066_, _42882_);
  not _54241_ (_03068_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _54242_ (_03069_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and _54243_ (_03070_, _03069_, _03068_);
  and _54244_ (_03072_, \oc8051_top_1.oc8051_sfr1.prescaler [3], _42882_);
  and _54245_ (_39849_, _03072_, _03070_);
  nor _54246_ (_03073_, _03070_, rst);
  nand _54247_ (_03075_, _03069_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  or _54248_ (_03076_, _03069_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _54249_ (_03077_, _03076_, _03075_);
  and _54250_ (_39850_, _03077_, _03073_);
  nor _54251_ (_03079_, _42527_, _42573_);
  not _54252_ (_03080_, _42304_);
  and _54253_ (_03082_, _42365_, _03080_);
  and _54254_ (_03083_, _03082_, _03079_);
  and _54255_ (_03084_, _03083_, _42448_);
  and _54256_ (_03086_, _03084_, _39021_);
  nor _54257_ (_03087_, _03086_, _01364_);
  not _54258_ (_03088_, _42527_);
  and _54259_ (_03090_, _03088_, _42573_);
  nor _54260_ (_03091_, _42365_, _42304_);
  and _54261_ (_03092_, _03091_, _42448_);
  and _54262_ (_03094_, _03092_, _03090_);
  not _54263_ (_03095_, _42610_);
  and _54264_ (_03097_, _39113_, _39100_);
  nor _54265_ (_03098_, _39113_, _39100_);
  or _54266_ (_03099_, _03098_, _03097_);
  nor _54267_ (_03100_, _39169_, _39125_);
  and _54268_ (_03102_, _39169_, _39125_);
  nor _54269_ (_03103_, _03102_, _03100_);
  nor _54270_ (_03104_, _03103_, _03099_);
  and _54271_ (_03106_, _03103_, _03099_);
  nor _54272_ (_03107_, _03106_, _03104_);
  and _54273_ (_03108_, _39193_, _39181_);
  nor _54274_ (_03110_, _39193_, _39181_);
  nor _54275_ (_03111_, _03110_, _03108_);
  nor _54276_ (_03112_, _39204_, _39045_);
  and _54277_ (_03114_, _39204_, _39045_);
  nor _54278_ (_03115_, _03114_, _03112_);
  or _54279_ (_03116_, _03115_, _03111_);
  nand _54280_ (_03119_, _03115_, _03111_);
  and _54281_ (_03120_, _03119_, _03116_);
  or _54282_ (_03121_, _03120_, _03107_);
  nand _54283_ (_03123_, _03120_, _03107_);
  and _54284_ (_03124_, _03123_, _03121_);
  or _54285_ (_03125_, _03124_, _03095_);
  and _54286_ (_03127_, _42484_, _42402_);
  or _54287_ (_03128_, _42610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _54288_ (_03130_, _03128_, _03127_);
  and _54289_ (_03131_, _03130_, _03125_);
  nor _54290_ (_03132_, _42484_, _42402_);
  nor _54291_ (_03133_, _42610_, _38889_);
  and _54292_ (_03135_, _42610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _54293_ (_03136_, _03135_, _03133_);
  and _54294_ (_03137_, _03136_, _03132_);
  or _54295_ (_03139_, _42610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  not _54296_ (_03140_, _42484_);
  and _54297_ (_03141_, _03140_, _42402_);
  nand _54298_ (_03143_, _42610_, _38905_);
  and _54299_ (_03144_, _03143_, _03141_);
  and _54300_ (_03145_, _03144_, _03139_);
  or _54301_ (_03147_, _03145_, _03137_);
  or _54302_ (_03148_, _03095_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nor _54303_ (_03149_, _03140_, _42402_);
  or _54304_ (_03151_, _42610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _54305_ (_03152_, _03151_, _03149_);
  and _54306_ (_03153_, _03152_, _03148_);
  or _54307_ (_03155_, _03153_, _03147_);
  or _54308_ (_03156_, _03155_, _03131_);
  and _54309_ (_03157_, _03156_, _03094_);
  and _54310_ (_03159_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _54311_ (_03160_, _03159_, _42610_);
  and _54312_ (_03162_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _54313_ (_03163_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _54314_ (_03164_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _54315_ (_03165_, _03164_, _03163_);
  or _54316_ (_03166_, _03165_, _03162_);
  or _54317_ (_03168_, _03166_, _03160_);
  and _54318_ (_03169_, _42527_, _42573_);
  and _54319_ (_03170_, _03091_, _42449_);
  and _54320_ (_03172_, _03170_, _03169_);
  and _54321_ (_03173_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _54322_ (_03174_, _03173_, _03095_);
  and _54323_ (_03176_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and _54324_ (_03177_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _54325_ (_03178_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _54326_ (_03180_, _03178_, _03177_);
  or _54327_ (_03181_, _03180_, _03176_);
  or _54328_ (_03182_, _03181_, _03174_);
  and _54329_ (_03184_, _03182_, _03172_);
  and _54330_ (_03185_, _03184_, _03168_);
  and _54331_ (_03186_, _38244_, _38271_);
  nor _54332_ (_03188_, _03186_, _38369_);
  not _54333_ (_03189_, _38288_);
  and _54334_ (_03190_, _00836_, _03189_);
  and _54335_ (_03192_, _03190_, _03188_);
  and _54336_ (_03193_, _38265_, _38260_);
  or _54337_ (_03195_, _00921_, _00768_);
  or _54338_ (_03196_, _03195_, _00834_);
  or _54339_ (_03197_, _03196_, _38300_);
  or _54340_ (_03198_, _03197_, _00766_);
  nor _54341_ (_03200_, _03198_, _03193_);
  and _54342_ (_03201_, _03200_, _38324_);
  and _54343_ (_03202_, _03201_, _03192_);
  and _54344_ (_03204_, _03202_, _01110_);
  nor _54345_ (_03205_, _03204_, _36407_);
  or _54346_ (_03206_, _03205_, p3_in[0]);
  not _54347_ (_03208_, _03205_);
  or _54348_ (_03209_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _54349_ (_03210_, _03209_, _03206_);
  and _54350_ (_03212_, _03210_, _03127_);
  or _54351_ (_03213_, _03212_, _03095_);
  or _54352_ (_03214_, _03205_, p3_in[3]);
  or _54353_ (_03216_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _54354_ (_03217_, _03216_, _03214_);
  and _54355_ (_03218_, _03217_, _03132_);
  or _54356_ (_03220_, _03205_, p3_in[2]);
  or _54357_ (_03221_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _54358_ (_03222_, _03221_, _03220_);
  and _54359_ (_03224_, _03222_, _03149_);
  or _54360_ (_03225_, _03205_, p3_in[1]);
  or _54361_ (_03227_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _54362_ (_03228_, _03227_, _03225_);
  and _54363_ (_03229_, _03228_, _03141_);
  or _54364_ (_03230_, _03229_, _03224_);
  or _54365_ (_03232_, _03230_, _03218_);
  or _54366_ (_03233_, _03232_, _03213_);
  and _54367_ (_03234_, _03092_, _42574_);
  and _54368_ (_03236_, _03234_, _42527_);
  or _54369_ (_03237_, _03205_, p3_in[4]);
  or _54370_ (_03238_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _54371_ (_03240_, _03238_, _03237_);
  and _54372_ (_03241_, _03240_, _03127_);
  or _54373_ (_03242_, _03241_, _42610_);
  or _54374_ (_03244_, _03205_, p3_in[7]);
  or _54375_ (_03245_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _54376_ (_03246_, _03245_, _03244_);
  and _54377_ (_03248_, _03246_, _03132_);
  or _54378_ (_03249_, _03205_, p3_in[6]);
  or _54379_ (_03250_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _54380_ (_03252_, _03250_, _03249_);
  and _54381_ (_03253_, _03252_, _03149_);
  or _54382_ (_03254_, _03205_, p3_in[5]);
  or _54383_ (_03256_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _54384_ (_03257_, _03256_, _03254_);
  and _54385_ (_03259_, _03257_, _03141_);
  or _54386_ (_03260_, _03259_, _03253_);
  or _54387_ (_03261_, _03260_, _03248_);
  or _54388_ (_03262_, _03261_, _03242_);
  and _54389_ (_03264_, _03262_, _03236_);
  and _54390_ (_03265_, _03264_, _03233_);
  or _54391_ (_03266_, _03265_, _03185_);
  or _54392_ (_03268_, _03205_, p0_in[1]);
  or _54393_ (_03269_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _54394_ (_03270_, _03269_, _03268_);
  and _54395_ (_03272_, _03270_, _03141_);
  or _54396_ (_03273_, _03272_, _03095_);
  or _54397_ (_03274_, _03205_, p0_in[3]);
  or _54398_ (_03276_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _54399_ (_03277_, _03276_, _03274_);
  and _54400_ (_03278_, _03277_, _03132_);
  or _54401_ (_03280_, _03205_, p0_in[0]);
  or _54402_ (_03281_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _54403_ (_03282_, _03281_, _03280_);
  and _54404_ (_03284_, _03282_, _03127_);
  or _54405_ (_03285_, _03205_, p0_in[2]);
  or _54406_ (_03286_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _54407_ (_03288_, _03286_, _03285_);
  and _54408_ (_03289_, _03288_, _03149_);
  or _54409_ (_03290_, _03289_, _03284_);
  or _54410_ (_03291_, _03290_, _03278_);
  or _54411_ (_03292_, _03291_, _03273_);
  and _54412_ (_03293_, _03169_, _03082_);
  and _54413_ (_03294_, _03293_, _42448_);
  or _54414_ (_03295_, _03205_, p0_in[5]);
  or _54415_ (_03296_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _54416_ (_03297_, _03296_, _03295_);
  and _54417_ (_03298_, _03297_, _03141_);
  or _54418_ (_03299_, _03298_, _42610_);
  or _54419_ (_03300_, _03205_, p0_in[7]);
  or _54420_ (_03301_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _54421_ (_03302_, _03301_, _03300_);
  and _54422_ (_03303_, _03302_, _03132_);
  or _54423_ (_03304_, _03205_, p0_in[4]);
  or _54424_ (_03305_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _54425_ (_03306_, _03305_, _03304_);
  and _54426_ (_03307_, _03306_, _03127_);
  or _54427_ (_03308_, _03205_, p0_in[6]);
  or _54428_ (_03309_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _54429_ (_03310_, _03309_, _03308_);
  and _54430_ (_03311_, _03310_, _03149_);
  or _54431_ (_03312_, _03311_, _03307_);
  or _54432_ (_03313_, _03312_, _03303_);
  or _54433_ (_03314_, _03313_, _03299_);
  and _54434_ (_03315_, _03314_, _03294_);
  and _54435_ (_03316_, _03315_, _03292_);
  and _54436_ (_03317_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _54437_ (_03318_, _03317_, _03095_);
  and _54438_ (_03319_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _54439_ (_03320_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _54440_ (_03321_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _54441_ (_03322_, _03321_, _03320_);
  or _54442_ (_03323_, _03322_, _03319_);
  or _54443_ (_03324_, _03323_, _03318_);
  and _54444_ (_03325_, _42527_, _42574_);
  and _54445_ (_03326_, _03325_, _03170_);
  and _54446_ (_03327_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _54447_ (_03328_, _03327_, _42610_);
  and _54448_ (_03329_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _54449_ (_03330_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and _54450_ (_03331_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _54451_ (_03332_, _03331_, _03330_);
  or _54452_ (_03333_, _03332_, _03329_);
  or _54453_ (_03334_, _03333_, _03328_);
  and _54454_ (_03335_, _03334_, _03326_);
  and _54455_ (_03336_, _03335_, _03324_);
  or _54456_ (_03337_, _03336_, _03316_);
  or _54457_ (_03338_, _03337_, _03266_);
  and _54458_ (_03339_, _01379_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or _54459_ (_03340_, _03205_, p2_in[1]);
  or _54460_ (_03341_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _54461_ (_03342_, _03341_, _03340_);
  and _54462_ (_03343_, _03342_, _03141_);
  or _54463_ (_03344_, _03343_, _03095_);
  or _54464_ (_03345_, _03205_, p2_in[3]);
  or _54465_ (_03346_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _54466_ (_03347_, _03346_, _03345_);
  and _54467_ (_03348_, _03347_, _03132_);
  or _54468_ (_03349_, _03205_, p2_in[0]);
  or _54469_ (_03350_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _54470_ (_03351_, _03350_, _03349_);
  and _54471_ (_03352_, _03351_, _03127_);
  or _54472_ (_03353_, _03205_, p2_in[2]);
  or _54473_ (_03354_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _54474_ (_03355_, _03354_, _03353_);
  and _54475_ (_03356_, _03355_, _03149_);
  or _54476_ (_03357_, _03356_, _03352_);
  or _54477_ (_03358_, _03357_, _03348_);
  or _54478_ (_03359_, _03358_, _03344_);
  and _54479_ (_03360_, _03325_, _03082_);
  and _54480_ (_03362_, _03360_, _42448_);
  or _54481_ (_03363_, _03205_, p2_in[5]);
  or _54482_ (_03364_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _54483_ (_03365_, _03364_, _03363_);
  and _54484_ (_03366_, _03365_, _03141_);
  or _54485_ (_03367_, _03366_, _42610_);
  or _54486_ (_03368_, _03205_, p2_in[7]);
  or _54487_ (_03369_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _54488_ (_03370_, _03369_, _03368_);
  and _54489_ (_03371_, _03370_, _03132_);
  or _54490_ (_03372_, _03205_, p2_in[4]);
  or _54491_ (_03373_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _54492_ (_03374_, _03373_, _03372_);
  and _54493_ (_03375_, _03374_, _03127_);
  or _54494_ (_03376_, _03205_, p2_in[6]);
  or _54495_ (_03377_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _54496_ (_03378_, _03377_, _03376_);
  and _54497_ (_03379_, _03378_, _03149_);
  or _54498_ (_03380_, _03379_, _03375_);
  or _54499_ (_03381_, _03380_, _03371_);
  or _54500_ (_03382_, _03381_, _03367_);
  and _54501_ (_03383_, _03382_, _03362_);
  and _54502_ (_03384_, _03383_, _03359_);
  or _54503_ (_03385_, _03384_, _03339_);
  and _54504_ (_03386_, _42527_, _03080_);
  nand _54505_ (_03387_, _03386_, _42449_);
  nor _54506_ (_03388_, _03092_, _28613_);
  and _54507_ (_03389_, _03388_, _03387_);
  nor _54508_ (_03390_, _03362_, _03084_);
  and _54509_ (_03391_, _03090_, _03082_);
  and _54510_ (_03392_, _03391_, _42449_);
  nor _54511_ (_03393_, _03392_, _03294_);
  and _54512_ (_03394_, _03393_, _03390_);
  and _54513_ (_03395_, _03394_, _03389_);
  and _54514_ (_03396_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _54515_ (_03397_, _03396_, _42610_);
  and _54516_ (_03398_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _54517_ (_03399_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _54518_ (_03400_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _54519_ (_03401_, _03400_, _03399_);
  or _54520_ (_03402_, _03401_, _03398_);
  or _54521_ (_03403_, _03402_, _03397_);
  and _54522_ (_03404_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _54523_ (_03405_, _03404_, _03095_);
  and _54524_ (_03406_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _54525_ (_03407_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _54526_ (_03408_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _54527_ (_03409_, _03408_, _03407_);
  or _54528_ (_03410_, _03409_, _03406_);
  or _54529_ (_03411_, _03410_, _03405_);
  and _54530_ (_03412_, _03411_, _03084_);
  and _54531_ (_03413_, _03412_, _03403_);
  or _54532_ (_03414_, _03413_, _03395_);
  or _54533_ (_03415_, _03414_, _03385_);
  or _54534_ (_03416_, _03415_, _03338_);
  and _54535_ (_03417_, _03082_, _42449_);
  and _54536_ (_03418_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _54537_ (_03419_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or _54538_ (_03420_, _03419_, _03418_);
  and _54539_ (_03421_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _54540_ (_03422_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _54541_ (_03423_, _03422_, _03421_);
  or _54542_ (_03424_, _03423_, _03420_);
  and _54543_ (_03425_, _03424_, _42610_);
  and _54544_ (_03426_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _54545_ (_03427_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _54546_ (_03428_, _03427_, _03426_);
  and _54547_ (_03429_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _54548_ (_03430_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  or _54549_ (_03431_, _03430_, _03429_);
  or _54550_ (_03432_, _03431_, _03428_);
  and _54551_ (_03433_, _03432_, _03095_);
  or _54552_ (_03434_, _03433_, _03425_);
  and _54553_ (_03435_, _03434_, _03325_);
  and _54554_ (_03436_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _54555_ (_03437_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _54556_ (_03438_, _03437_, _03436_);
  and _54557_ (_03439_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _54558_ (_03440_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _54559_ (_03441_, _03440_, _03439_);
  or _54560_ (_03442_, _03441_, _03438_);
  and _54561_ (_03443_, _03442_, _03095_);
  and _54562_ (_03444_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _54563_ (_03445_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or _54564_ (_03446_, _03445_, _03444_);
  and _54565_ (_03447_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _54566_ (_03448_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _54567_ (_03449_, _03448_, _03447_);
  or _54568_ (_03450_, _03449_, _03446_);
  and _54569_ (_03451_, _03450_, _42610_);
  or _54570_ (_03452_, _03451_, _03443_);
  and _54571_ (_03453_, _03452_, _03169_);
  or _54572_ (_03454_, _03453_, _03435_);
  and _54573_ (_03455_, _03454_, _03417_);
  or _54574_ (_03456_, _03205_, p1_in[4]);
  or _54575_ (_03457_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _54576_ (_03458_, _03457_, _03456_);
  and _54577_ (_03459_, _03458_, _03127_);
  or _54578_ (_03460_, _03459_, _42610_);
  or _54579_ (_03461_, _03205_, p1_in[7]);
  or _54580_ (_03462_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _54581_ (_03463_, _03462_, _03461_);
  and _54582_ (_03464_, _03463_, _03132_);
  or _54583_ (_03465_, _03205_, p1_in[6]);
  or _54584_ (_03466_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _54585_ (_03467_, _03466_, _03465_);
  and _54586_ (_03468_, _03467_, _03149_);
  or _54587_ (_03469_, _03205_, p1_in[5]);
  or _54588_ (_03470_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _54589_ (_03471_, _03470_, _03469_);
  and _54590_ (_03472_, _03471_, _03141_);
  or _54591_ (_03473_, _03472_, _03468_);
  or _54592_ (_03474_, _03473_, _03464_);
  or _54593_ (_03475_, _03474_, _03460_);
  and _54594_ (_03476_, _03169_, _03092_);
  or _54595_ (_03477_, _03205_, p1_in[0]);
  or _54596_ (_03478_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _54597_ (_03479_, _03478_, _03477_);
  and _54598_ (_03480_, _03479_, _03127_);
  or _54599_ (_03481_, _03480_, _03095_);
  or _54600_ (_03482_, _03205_, p1_in[3]);
  or _54601_ (_03483_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _54602_ (_03484_, _03483_, _03482_);
  and _54603_ (_03485_, _03484_, _03132_);
  or _54604_ (_03486_, _03205_, p1_in[2]);
  or _54605_ (_03487_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _54606_ (_03488_, _03487_, _03486_);
  and _54607_ (_03489_, _03488_, _03149_);
  or _54608_ (_03490_, _03205_, p1_in[1]);
  or _54609_ (_03491_, _03208_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _54610_ (_03492_, _03491_, _03490_);
  and _54611_ (_03493_, _03492_, _03141_);
  or _54612_ (_03494_, _03493_, _03489_);
  or _54613_ (_03495_, _03494_, _03485_);
  or _54614_ (_03496_, _03495_, _03481_);
  and _54615_ (_03497_, _03496_, _03476_);
  and _54616_ (_03498_, _03497_, _03475_);
  and _54617_ (_03499_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or _54618_ (_03500_, _03499_, _42610_);
  and _54619_ (_03501_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _54620_ (_03502_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _54621_ (_03503_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or _54622_ (_03504_, _03503_, _03502_);
  or _54623_ (_03505_, _03504_, _03501_);
  or _54624_ (_03506_, _03505_, _03500_);
  and _54625_ (_03507_, _03234_, _03088_);
  and _54626_ (_03508_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _54627_ (_03509_, _03508_, _03095_);
  and _54628_ (_03510_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _54629_ (_03511_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _54630_ (_03512_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _54631_ (_03513_, _03512_, _03511_);
  or _54632_ (_03514_, _03513_, _03510_);
  or _54633_ (_03515_, _03514_, _03509_);
  and _54634_ (_03516_, _03515_, _03507_);
  and _54635_ (_03517_, _03516_, _03506_);
  and _54636_ (_03518_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _54637_ (_03519_, _03518_, _03095_);
  and _54638_ (_03520_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _54639_ (_03521_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _54640_ (_03522_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _54641_ (_03523_, _03522_, _03521_);
  or _54642_ (_03524_, _03523_, _03520_);
  or _54643_ (_03525_, _03524_, _03519_);
  and _54644_ (_03526_, _03149_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _54645_ (_03527_, _03526_, _42610_);
  and _54646_ (_03528_, _03132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and _54647_ (_03529_, _03127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _54648_ (_03530_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or _54649_ (_03531_, _03530_, _03529_);
  or _54650_ (_03532_, _03531_, _03528_);
  or _54651_ (_03533_, _03532_, _03527_);
  and _54652_ (_03534_, _03533_, _03392_);
  and _54653_ (_03535_, _03534_, _03525_);
  or _54654_ (_03536_, _03535_, _03517_);
  or _54655_ (_03537_, _03536_, _03498_);
  or _54656_ (_03538_, _03537_, _03455_);
  or _54657_ (_03539_, _03538_, _03416_);
  or _54658_ (_03540_, _03539_, _03157_);
  nand _54659_ (_03541_, _03339_, _31282_);
  nand _54660_ (_03542_, _03541_, _03540_);
  nand _54661_ (_03543_, _03542_, _03087_);
  nand _54662_ (_03544_, _42610_, _38456_);
  nand _54663_ (_03545_, _03095_, _38428_);
  and _54664_ (_03546_, _03545_, _03141_);
  and _54665_ (_03547_, _03546_, _03544_);
  and _54666_ (_03548_, _42610_, _42600_);
  nor _54667_ (_03549_, _42610_, _38420_);
  or _54668_ (_03550_, _03549_, _03548_);
  and _54669_ (_03551_, _03550_, _03149_);
  nor _54670_ (_03552_, _42610_, _38434_);
  and _54671_ (_03553_, _42610_, _38465_);
  or _54672_ (_03554_, _03553_, _03552_);
  and _54673_ (_03555_, _03554_, _03127_);
  nand _54674_ (_03556_, _42610_, _38442_);
  nand _54675_ (_03557_, _03095_, _38485_);
  and _54676_ (_03558_, _03557_, _03132_);
  and _54677_ (_03559_, _03558_, _03556_);
  or _54678_ (_03560_, _03559_, _03555_);
  or _54679_ (_03561_, _03560_, _03551_);
  or _54680_ (_03563_, _03561_, _03547_);
  or _54681_ (_03564_, _03563_, _03087_);
  and _54682_ (_03565_, _03564_, _42882_);
  and _54683_ (_39851_, _03565_, _03543_);
  nor _54684_ (_03566_, _42365_, _42574_);
  nor _54685_ (_03567_, _42527_, _42304_);
  and _54686_ (_03568_, _42448_, _42610_);
  and _54687_ (_03569_, _03568_, _03127_);
  and _54688_ (_03570_, _03569_, _03567_);
  and _54689_ (_03571_, _03570_, _03566_);
  and _54690_ (_03572_, _03571_, _01438_);
  and _54691_ (_03573_, _03569_, _03083_);
  and _54692_ (_03574_, _03573_, _39018_);
  nor _54693_ (_03575_, _03574_, _03572_);
  and _54694_ (_03576_, _03568_, _03132_);
  and _54695_ (_03577_, _03576_, _03293_);
  nand _54696_ (_03578_, _03577_, _38533_);
  and _54697_ (_03579_, _03578_, _03575_);
  nor _54698_ (_03580_, _03579_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _54699_ (_03581_, _03580_);
  not _54700_ (_03582_, _39031_);
  and _54701_ (_03583_, _03132_, _03095_);
  nor _54702_ (_03584_, _03583_, _03582_);
  and _54703_ (_03585_, _03584_, _01362_);
  and _54704_ (_03586_, _03573_, _39021_);
  nor _54705_ (_03587_, _03586_, _03585_);
  and _54706_ (_03588_, _03587_, _01382_);
  and _54707_ (_03589_, _03588_, _03581_);
  and _54708_ (_03590_, _03293_, _03149_);
  and _54709_ (_03591_, _03590_, _03568_);
  and _54710_ (_03592_, _03591_, _38533_);
  or _54711_ (_03593_, _03592_, rst);
  nor _54712_ (_39853_, _03593_, _03589_);
  nand _54713_ (_03594_, _03592_, _30603_);
  and _54714_ (_03595_, _42449_, _42610_);
  and _54715_ (_03596_, _03595_, _03127_);
  and _54716_ (_03597_, _03596_, _03391_);
  and _54717_ (_03598_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor _54718_ (_03599_, _42448_, _42610_);
  and _54719_ (_03600_, _03599_, _03127_);
  and _54720_ (_03601_, _03600_, _03391_);
  and _54721_ (_03602_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _54722_ (_03603_, _03602_, _03598_);
  and _54723_ (_03604_, _03595_, _03149_);
  and _54724_ (_03605_, _03604_, _03391_);
  and _54725_ (_03606_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and _54726_ (_03607_, _03599_, _03141_);
  and _54727_ (_03608_, _03607_, _03391_);
  and _54728_ (_03609_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _54729_ (_03610_, _03609_, _03606_);
  or _54730_ (_03611_, _03610_, _03603_);
  and _54731_ (_03612_, _03596_, _03293_);
  and _54732_ (_03613_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _54733_ (_03614_, _03595_, _03132_);
  and _54734_ (_03615_, _03614_, _03391_);
  and _54735_ (_03616_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or _54736_ (_03617_, _03616_, _03613_);
  and _54737_ (_03618_, _03596_, _03360_);
  and _54738_ (_03619_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _54739_ (_03620_, _03583_, _42448_);
  nor _54740_ (_03621_, _42365_, _42573_);
  and _54741_ (_03622_, _03621_, _03386_);
  and _54742_ (_03623_, _03622_, _03620_);
  and _54743_ (_03624_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or _54744_ (_03625_, _03624_, _03619_);
  or _54745_ (_03626_, _03625_, _03617_);
  or _54746_ (_03627_, _03626_, _03611_);
  and _54747_ (_03628_, _03614_, _03293_);
  and _54748_ (_03629_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _54749_ (_03630_, _03595_, _03141_);
  and _54750_ (_03631_, _03630_, _03293_);
  and _54751_ (_03632_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or _54752_ (_03633_, _03632_, _03629_);
  and _54753_ (_03634_, _03607_, _03293_);
  and _54754_ (_03635_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _54755_ (_03636_, _03604_, _03293_);
  and _54756_ (_03637_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _54757_ (_03638_, _03637_, _03635_);
  or _54758_ (_03639_, _03638_, _03633_);
  and _54759_ (_03640_, _03169_, _03091_);
  and _54760_ (_03641_, _03640_, _03630_);
  and _54761_ (_03642_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _54762_ (_03643_, _03596_, _03640_);
  and _54763_ (_03644_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _54764_ (_03645_, _03644_, _03642_);
  and _54765_ (_03646_, _03600_, _03293_);
  and _54766_ (_03647_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _54767_ (_03648_, _03583_, _03294_);
  and _54768_ (_03649_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _54769_ (_03650_, _03649_, _03647_);
  or _54770_ (_03651_, _03650_, _03645_);
  or _54771_ (_03652_, _03651_, _03639_);
  or _54772_ (_03653_, _03652_, _03627_);
  and _54773_ (_03654_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _54774_ (_03655_, _03293_, _03132_);
  and _54775_ (_03656_, _03655_, _03568_);
  and _54776_ (_03657_, _03656_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or _54777_ (_03658_, _03657_, _03654_);
  and _54778_ (_03659_, _03621_, _03570_);
  and _54779_ (_03660_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _54780_ (_03661_, _03293_, _03141_);
  and _54781_ (_03662_, _03661_, _03568_);
  and _54782_ (_03663_, _03662_, _42245_);
  or _54783_ (_03664_, _03663_, _03660_);
  or _54784_ (_03665_, _03664_, _03658_);
  and _54785_ (_03666_, _03569_, _03360_);
  and _54786_ (_03667_, _03666_, _03370_);
  and _54787_ (_03668_, _03622_, _03569_);
  and _54788_ (_03669_, _03668_, _03246_);
  or _54789_ (_03670_, _03669_, _03667_);
  and _54790_ (_03671_, _03569_, _03293_);
  and _54791_ (_03672_, _03671_, _03302_);
  and _54792_ (_03673_, _03640_, _03569_);
  and _54793_ (_03674_, _03673_, _03463_);
  or _54794_ (_03675_, _03674_, _03672_);
  or _54795_ (_03676_, _03675_, _03670_);
  or _54796_ (_03677_, _03676_, _03665_);
  and _54797_ (_03678_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and _54798_ (_03679_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _54799_ (_03680_, _03679_, _03678_);
  or _54800_ (_03681_, _03680_, _03677_);
  or _54801_ (_03682_, _03681_, _03653_);
  and _54802_ (_03683_, _03682_, _03589_);
  and _54803_ (_03684_, _03569_, _03386_);
  or _54804_ (_03685_, _03659_, _03684_);
  or _54805_ (_03686_, _03685_, _03662_);
  and _54806_ (_03687_, _03595_, _03655_);
  or _54807_ (_03688_, _03646_, _03641_);
  or _54808_ (_03689_, _03634_, _03643_);
  or _54809_ (_03690_, _03689_, _03688_);
  or _54810_ (_03691_, _03690_, _03687_);
  or _54811_ (_03692_, _03691_, _03686_);
  or _54812_ (_03693_, _03623_, _03573_);
  or _54813_ (_03694_, _03648_, _03571_);
  or _54814_ (_03695_, _03694_, _03693_);
  or _54815_ (_03696_, _03615_, _03605_);
  or _54816_ (_03697_, _03608_, _03612_);
  or _54817_ (_03698_, _03697_, _03696_);
  or _54818_ (_03699_, _03698_, _03656_);
  or _54819_ (_03700_, _03699_, _03695_);
  and _54820_ (_03701_, _03595_, _03590_);
  or _54821_ (_03702_, _03631_, _03618_);
  or _54822_ (_03703_, _03702_, _03701_);
  and _54823_ (_03704_, _03392_, _03127_);
  or _54824_ (_03705_, _03704_, _03591_);
  or _54825_ (_03706_, _03705_, _03703_);
  or _54826_ (_03707_, _03706_, _03700_);
  or _54827_ (_03708_, _03707_, _03692_);
  nand _54828_ (_03709_, _03708_, _03589_);
  and _54829_ (_03710_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or _54830_ (_03711_, _03710_, _03683_);
  or _54831_ (_03712_, _03711_, _03592_);
  and _54832_ (_03713_, _03712_, _42882_);
  and _54833_ (_39854_, _03713_, _03594_);
  nor _54834_ (_39935_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or _54835_ (_03714_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor _54836_ (_03715_, _03069_, rst);
  and _54837_ (_39936_, _03715_, _03714_);
  nor _54838_ (_03716_, _03069_, _03068_);
  or _54839_ (_03717_, _03716_, _03070_);
  and _54840_ (_03718_, _03075_, _42882_);
  and _54841_ (_39937_, _03718_, _03717_);
  and _54842_ (_03719_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _54843_ (_03720_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or _54844_ (_03721_, _03720_, _03719_);
  and _54845_ (_03722_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _54846_ (_03723_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _54847_ (_03724_, _03723_, _03722_);
  or _54848_ (_03725_, _03724_, _03721_);
  and _54849_ (_03726_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _54850_ (_03727_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or _54851_ (_03728_, _03727_, _03726_);
  and _54852_ (_03729_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _54853_ (_03730_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _54854_ (_03731_, _03730_, _03729_);
  or _54855_ (_03732_, _03731_, _03728_);
  or _54856_ (_03733_, _03732_, _03725_);
  and _54857_ (_03734_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _54858_ (_03735_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or _54859_ (_03736_, _03735_, _03734_);
  and _54860_ (_03737_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _54861_ (_03738_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or _54862_ (_03739_, _03738_, _03737_);
  or _54863_ (_03740_, _03739_, _03736_);
  and _54864_ (_03741_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and _54865_ (_03742_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _54866_ (_03743_, _03742_, _03741_);
  and _54867_ (_03744_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _54868_ (_03745_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  or _54869_ (_03746_, _03745_, _03744_);
  or _54870_ (_03747_, _03746_, _03743_);
  or _54871_ (_03748_, _03747_, _03740_);
  or _54872_ (_03749_, _03748_, _03733_);
  and _54873_ (_03750_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and _54874_ (_03751_, _03662_, _42480_);
  or _54875_ (_03752_, _03751_, _03750_);
  and _54876_ (_03753_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _54877_ (_03754_, _03577_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or _54878_ (_03755_, _03754_, _03753_);
  or _54879_ (_03756_, _03755_, _03752_);
  and _54880_ (_03758_, _03666_, _03351_);
  and _54881_ (_03759_, _03668_, _03210_);
  or _54882_ (_03760_, _03759_, _03758_);
  and _54883_ (_03761_, _03671_, _03282_);
  and _54884_ (_03762_, _03673_, _03479_);
  or _54885_ (_03763_, _03762_, _03761_);
  or _54886_ (_03764_, _03763_, _03760_);
  or _54887_ (_03765_, _03764_, _03756_);
  and _54888_ (_03766_, _03571_, _03124_);
  and _54889_ (_03767_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _54890_ (_03768_, _03767_, _03766_);
  or _54891_ (_03769_, _03768_, _03765_);
  or _54892_ (_03770_, _03769_, _03749_);
  and _54893_ (_03771_, _03770_, _03589_);
  and _54894_ (_03772_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or _54895_ (_03773_, _03772_, _03592_);
  or _54896_ (_03774_, _03773_, _03771_);
  nand _54897_ (_03775_, _03592_, _31782_);
  and _54898_ (_03776_, _03775_, _42882_);
  and _54899_ (_39938_, _03776_, _03774_);
  and _54900_ (_03777_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _54901_ (_03778_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _54902_ (_03779_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _54903_ (_03780_, _03779_, _03778_);
  and _54904_ (_03781_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _54905_ (_03782_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _54906_ (_03783_, _03782_, _03781_);
  or _54907_ (_03784_, _03783_, _03780_);
  and _54908_ (_03785_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _54909_ (_03786_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _54910_ (_03787_, _03786_, _03785_);
  and _54911_ (_03788_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _54912_ (_03789_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _54913_ (_03790_, _03789_, _03788_);
  or _54914_ (_03791_, _03790_, _03787_);
  or _54915_ (_03792_, _03791_, _03784_);
  and _54916_ (_03793_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _54917_ (_03794_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _54918_ (_03795_, _03794_, _03793_);
  and _54919_ (_03796_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _54920_ (_03797_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _54921_ (_03798_, _03797_, _03796_);
  or _54922_ (_03799_, _03798_, _03795_);
  and _54923_ (_03800_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and _54924_ (_03801_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _54925_ (_03802_, _03801_, _03800_);
  and _54926_ (_03803_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _54927_ (_03804_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or _54928_ (_03805_, _03804_, _03803_);
  or _54929_ (_03806_, _03805_, _03802_);
  or _54930_ (_03807_, _03806_, _03799_);
  or _54931_ (_03808_, _03807_, _03792_);
  and _54932_ (_03809_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _54933_ (_03810_, _03662_, _42387_);
  or _54934_ (_03811_, _03810_, _03809_);
  and _54935_ (_03812_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _54936_ (_03813_, _03577_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _54937_ (_03814_, _03813_, _03812_);
  or _54938_ (_03815_, _03814_, _03811_);
  and _54939_ (_03816_, _03666_, _03342_);
  and _54940_ (_03817_, _03668_, _03228_);
  or _54941_ (_03818_, _03817_, _03816_);
  and _54942_ (_03819_, _03671_, _03270_);
  and _54943_ (_03820_, _03673_, _03492_);
  or _54944_ (_03821_, _03820_, _03819_);
  or _54945_ (_03822_, _03821_, _03818_);
  or _54946_ (_03823_, _03822_, _03815_);
  and _54947_ (_03824_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _54948_ (_03825_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _54949_ (_03826_, _03825_, _03824_);
  or _54950_ (_03827_, _03826_, _03823_);
  or _54951_ (_03828_, _03827_, _03808_);
  and _54952_ (_03829_, _03828_, _03589_);
  or _54953_ (_03830_, _03829_, _03592_);
  or _54954_ (_03831_, _03830_, _03777_);
  nand _54955_ (_03832_, _03592_, _32458_);
  and _54956_ (_03833_, _03832_, _42882_);
  and _54957_ (_39939_, _03833_, _03831_);
  and _54958_ (_03834_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and _54959_ (_03835_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _54960_ (_03836_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _54961_ (_03837_, _03836_, _03835_);
  and _54962_ (_03838_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _54963_ (_03839_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _54964_ (_03840_, _03839_, _03838_);
  or _54965_ (_03841_, _03840_, _03837_);
  and _54966_ (_03842_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _54967_ (_03843_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _54968_ (_03844_, _03843_, _03842_);
  and _54969_ (_03845_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _54970_ (_03846_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _54971_ (_03847_, _03846_, _03845_);
  or _54972_ (_03848_, _03847_, _03844_);
  or _54973_ (_03849_, _03848_, _03841_);
  and _54974_ (_03850_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _54975_ (_03851_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _54976_ (_03852_, _03851_, _03850_);
  and _54977_ (_03853_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _54978_ (_03854_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or _54979_ (_03855_, _03854_, _03853_);
  or _54980_ (_03856_, _03855_, _03852_);
  and _54981_ (_03857_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and _54982_ (_03858_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  or _54983_ (_03859_, _03858_, _03857_);
  and _54984_ (_03860_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _54985_ (_03861_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _54986_ (_03862_, _03861_, _03860_);
  or _54987_ (_03863_, _03862_, _03859_);
  or _54988_ (_03864_, _03863_, _03856_);
  or _54989_ (_03865_, _03864_, _03849_);
  and _54990_ (_03866_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _54991_ (_03867_, _03656_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _54992_ (_03868_, _03867_, _03866_);
  and _54993_ (_03869_, _03662_, _42606_);
  and _54994_ (_03870_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _54995_ (_03871_, _03870_, _03869_);
  or _54996_ (_03872_, _03871_, _03868_);
  and _54997_ (_03873_, _03666_, _03355_);
  and _54998_ (_03874_, _03668_, _03222_);
  or _54999_ (_03875_, _03874_, _03873_);
  and _55000_ (_03876_, _03671_, _03288_);
  and _55001_ (_03877_, _03673_, _03488_);
  or _55002_ (_03878_, _03877_, _03876_);
  or _55003_ (_03879_, _03878_, _03875_);
  or _55004_ (_03880_, _03879_, _03872_);
  and _55005_ (_03881_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _55006_ (_03882_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _55007_ (_03883_, _03882_, _03881_);
  or _55008_ (_03884_, _03883_, _03880_);
  or _55009_ (_03885_, _03884_, _03865_);
  and _55010_ (_03886_, _03885_, _03589_);
  or _55011_ (_03887_, _03886_, _03592_);
  or _55012_ (_03888_, _03887_, _03834_);
  nand _55013_ (_03889_, _03592_, _33154_);
  and _55014_ (_03890_, _03889_, _42882_);
  and _55015_ (_39940_, _03890_, _03888_);
  nand _55016_ (_03891_, _03592_, _33906_);
  and _55017_ (_03892_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _55018_ (_03893_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _55019_ (_03894_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _55020_ (_03895_, _03894_, _03893_);
  and _55021_ (_03896_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _55022_ (_03897_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _55023_ (_03898_, _03897_, _03896_);
  or _55024_ (_03899_, _03898_, _03895_);
  and _55025_ (_03900_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _55026_ (_03901_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or _55027_ (_03902_, _03901_, _03900_);
  and _55028_ (_03903_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _55029_ (_03904_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _55030_ (_03905_, _03904_, _03903_);
  or _55031_ (_03906_, _03905_, _03902_);
  or _55032_ (_03907_, _03906_, _03899_);
  and _55033_ (_03908_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _55034_ (_03909_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or _55035_ (_03910_, _03909_, _03908_);
  and _55036_ (_03911_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _55037_ (_03912_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _55038_ (_03913_, _03912_, _03911_);
  or _55039_ (_03914_, _03913_, _03910_);
  and _55040_ (_03915_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and _55041_ (_03916_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or _55042_ (_03917_, _03916_, _03915_);
  and _55043_ (_03918_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _55044_ (_03919_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or _55045_ (_03920_, _03919_, _03918_);
  or _55046_ (_03921_, _03920_, _03917_);
  or _55047_ (_03922_, _03921_, _03914_);
  or _55048_ (_03923_, _03922_, _03907_);
  and _55049_ (_03924_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _55050_ (_03925_, _03656_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _55051_ (_03926_, _03925_, _03924_);
  and _55052_ (_03927_, _03662_, _42433_);
  and _55053_ (_03928_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _55054_ (_03929_, _03928_, _03927_);
  or _55055_ (_03930_, _03929_, _03926_);
  and _55056_ (_03931_, _03666_, _03347_);
  and _55057_ (_03932_, _03668_, _03217_);
  or _55058_ (_03933_, _03932_, _03931_);
  and _55059_ (_03934_, _03671_, _03277_);
  and _55060_ (_03935_, _03673_, _03484_);
  or _55061_ (_03936_, _03935_, _03934_);
  or _55062_ (_03937_, _03936_, _03933_);
  or _55063_ (_03938_, _03937_, _03930_);
  and _55064_ (_03939_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _55065_ (_03940_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _55066_ (_03941_, _03940_, _03939_);
  or _55067_ (_03942_, _03941_, _03938_);
  or _55068_ (_03943_, _03942_, _03923_);
  and _55069_ (_03944_, _03943_, _03589_);
  or _55070_ (_03945_, _03944_, _03892_);
  or _55071_ (_03946_, _03945_, _03592_);
  and _55072_ (_03947_, _03946_, _42882_);
  and _55073_ (_39941_, _03947_, _03891_);
  nand _55074_ (_03948_, _03592_, _34667_);
  and _55075_ (_03949_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and _55076_ (_03950_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _55077_ (_03951_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _55078_ (_03952_, _03951_, _03950_);
  and _55079_ (_03953_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _55080_ (_03955_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _55081_ (_03956_, _03955_, _03953_);
  or _55082_ (_03957_, _03956_, _03952_);
  and _55083_ (_03958_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _55084_ (_03959_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  or _55085_ (_03960_, _03959_, _03958_);
  and _55086_ (_03961_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and _55087_ (_03962_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or _55088_ (_03963_, _03962_, _03961_);
  or _55089_ (_03964_, _03963_, _03960_);
  or _55090_ (_03965_, _03964_, _03957_);
  and _55091_ (_03966_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _55092_ (_03967_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or _55093_ (_03968_, _03967_, _03966_);
  and _55094_ (_03969_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _55095_ (_03970_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or _55096_ (_03971_, _03970_, _03969_);
  or _55097_ (_03972_, _03971_, _03968_);
  and _55098_ (_03973_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and _55099_ (_03974_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _55100_ (_03975_, _03974_, _03973_);
  and _55101_ (_03976_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _55102_ (_03977_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or _55103_ (_03978_, _03977_, _03976_);
  or _55104_ (_03979_, _03978_, _03975_);
  or _55105_ (_03980_, _03979_, _03972_);
  or _55106_ (_03981_, _03980_, _03965_);
  and _55107_ (_03982_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _55108_ (_03983_, _03662_, _42360_);
  or _55109_ (_03984_, _03983_, _03982_);
  and _55110_ (_03985_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _55111_ (_03986_, _03577_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or _55112_ (_03987_, _03986_, _03985_);
  or _55113_ (_03988_, _03987_, _03984_);
  and _55114_ (_03989_, _03666_, _03374_);
  and _55115_ (_03990_, _03668_, _03240_);
  or _55116_ (_03991_, _03990_, _03989_);
  and _55117_ (_03992_, _03671_, _03306_);
  and _55118_ (_03993_, _03673_, _03458_);
  or _55119_ (_03994_, _03993_, _03992_);
  or _55120_ (_03995_, _03994_, _03991_);
  or _55121_ (_03996_, _03995_, _03988_);
  and _55122_ (_03997_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _55123_ (_03998_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or _55124_ (_03999_, _03998_, _03997_);
  or _55125_ (_04000_, _03999_, _03996_);
  or _55126_ (_04001_, _04000_, _03981_);
  and _55127_ (_04002_, _04001_, _03589_);
  or _55128_ (_04003_, _04002_, _03949_);
  or _55129_ (_04004_, _04003_, _03592_);
  and _55130_ (_04005_, _04004_, _42882_);
  and _55131_ (_39943_, _04005_, _03948_);
  nand _55132_ (_04006_, _03592_, _35461_);
  and _55133_ (_04007_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and _55134_ (_04008_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _55135_ (_04009_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _55136_ (_04010_, _04009_, _04008_);
  and _55137_ (_04011_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and _55138_ (_04012_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _55139_ (_04013_, _04012_, _04011_);
  or _55140_ (_04014_, _04013_, _04010_);
  and _55141_ (_04015_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _55142_ (_04016_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _55143_ (_04017_, _04016_, _04015_);
  and _55144_ (_04018_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _55145_ (_04019_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or _55146_ (_04020_, _04019_, _04018_);
  or _55147_ (_04021_, _04020_, _04017_);
  or _55148_ (_04022_, _04021_, _04014_);
  and _55149_ (_04023_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _55150_ (_04024_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _55151_ (_04025_, _04024_, _04023_);
  and _55152_ (_04026_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _55153_ (_04027_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _55154_ (_04028_, _04027_, _04026_);
  or _55155_ (_04029_, _04028_, _04025_);
  and _55156_ (_04030_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _55157_ (_04031_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _55158_ (_04032_, _04031_, _04030_);
  and _55159_ (_04033_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _55160_ (_04034_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or _55161_ (_04035_, _04034_, _04033_);
  or _55162_ (_04036_, _04035_, _04032_);
  or _55163_ (_04037_, _04036_, _04029_);
  or _55164_ (_04038_, _04037_, _04022_);
  not _55165_ (_04039_, _38525_);
  and _55166_ (_04040_, _03662_, _04039_);
  and _55167_ (_04041_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or _55168_ (_04042_, _04041_, _04040_);
  and _55169_ (_04043_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _55170_ (_04044_, _03577_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or _55171_ (_04045_, _04044_, _04043_);
  or _55172_ (_04046_, _04045_, _04042_);
  and _55173_ (_04047_, _03666_, _03365_);
  and _55174_ (_04048_, _03668_, _03257_);
  or _55175_ (_04049_, _04048_, _04047_);
  and _55176_ (_04050_, _03671_, _03297_);
  and _55177_ (_04051_, _03673_, _03471_);
  or _55178_ (_04052_, _04051_, _04050_);
  or _55179_ (_04053_, _04052_, _04049_);
  or _55180_ (_04055_, _04053_, _04046_);
  and _55181_ (_04056_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _55182_ (_04057_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _55183_ (_04058_, _04057_, _04056_);
  or _55184_ (_04059_, _04058_, _04055_);
  or _55185_ (_04060_, _04059_, _04038_);
  and _55186_ (_04061_, _04060_, _03589_);
  or _55187_ (_04062_, _04061_, _04007_);
  or _55188_ (_04063_, _04062_, _03592_);
  and _55189_ (_04064_, _04063_, _42882_);
  and _55190_ (_39944_, _04064_, _04006_);
  and _55191_ (_04065_, _03597_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and _55192_ (_04066_, _03601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or _55193_ (_04067_, _04066_, _04065_);
  and _55194_ (_04068_, _03605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _55195_ (_04069_, _03608_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _55196_ (_04070_, _04069_, _04068_);
  or _55197_ (_04071_, _04070_, _04067_);
  and _55198_ (_04072_, _03615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _55199_ (_04073_, _03612_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _55200_ (_04074_, _04073_, _04072_);
  and _55201_ (_04075_, _03618_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _55202_ (_04076_, _03623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _55203_ (_04077_, _04076_, _04075_);
  or _55204_ (_04078_, _04077_, _04074_);
  or _55205_ (_04079_, _04078_, _04071_);
  and _55206_ (_04080_, _03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _55207_ (_04081_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _55208_ (_04082_, _04081_, _04080_);
  and _55209_ (_04083_, _03634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _55210_ (_04084_, _03636_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _55211_ (_04085_, _04084_, _04083_);
  or _55212_ (_04086_, _04085_, _04082_);
  and _55213_ (_04087_, _03641_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and _55214_ (_04088_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _55215_ (_04089_, _04088_, _04087_);
  and _55216_ (_04090_, _03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _55217_ (_04091_, _03648_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or _55218_ (_04092_, _04091_, _04090_);
  or _55219_ (_04093_, _04092_, _04089_);
  or _55220_ (_04094_, _04093_, _04086_);
  or _55221_ (_04095_, _04094_, _04079_);
  and _55222_ (_04096_, _03591_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _55223_ (_04097_, _03656_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _55224_ (_04098_, _04097_, _04096_);
  and _55225_ (_04099_, _03659_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _55226_ (_04100_, _03662_, _42508_);
  or _55227_ (_04101_, _04100_, _04099_);
  or _55228_ (_04102_, _04101_, _04098_);
  and _55229_ (_04103_, _03666_, _03378_);
  and _55230_ (_04104_, _03668_, _03252_);
  or _55231_ (_04105_, _04104_, _04103_);
  and _55232_ (_04106_, _03671_, _03310_);
  and _55233_ (_04107_, _03673_, _03467_);
  or _55234_ (_04108_, _04107_, _04106_);
  or _55235_ (_04109_, _04108_, _04105_);
  or _55236_ (_04110_, _04109_, _04102_);
  and _55237_ (_04111_, _03571_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _55238_ (_04112_, _03573_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _55239_ (_04113_, _04112_, _04111_);
  or _55240_ (_04114_, _04113_, _04110_);
  or _55241_ (_04115_, _04114_, _04095_);
  and _55242_ (_04116_, _04115_, _03589_);
  and _55243_ (_04117_, _03709_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  or _55244_ (_04118_, _04117_, _04116_);
  or _55245_ (_04119_, _04118_, _03592_);
  nand _55246_ (_04120_, _03592_, _36179_);
  and _55247_ (_04121_, _04120_, _42882_);
  and _55248_ (_39945_, _04121_, _04119_);
  and _55249_ (_40015_, _42648_, _42882_);
  nor _55250_ (_40019_, _42610_, rst);
  and _55251_ (_40041_, _42794_, _42882_);
  nor _55252_ (_40044_, _42484_, rst);
  nor _55253_ (_40045_, _42402_, rst);
  not _55254_ (_04122_, _00317_);
  nor _55255_ (_04123_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _55256_ (_04124_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55257_ (_04125_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _04124_);
  nor _55258_ (_04126_, _04125_, _04123_);
  nor _55259_ (_04127_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55260_ (_04128_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _04124_);
  nor _55261_ (_04129_, _04128_, _04127_);
  nor _55262_ (_04130_, _04129_, _04126_);
  and _55263_ (_04131_, _04129_, _04126_);
  nor _55264_ (_04132_, _02202_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55265_ (_04133_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _04124_);
  nor _55266_ (_04134_, _04133_, _04132_);
  and _55267_ (_04135_, _04134_, _04131_);
  nor _55268_ (_04136_, _04134_, _04131_);
  nor _55269_ (_04137_, _04136_, _04135_);
  not _55270_ (_04138_, _04137_);
  nor _55271_ (_04139_, _02221_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _55272_ (_04140_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _04124_);
  nor _55273_ (_04141_, _04140_, _04139_);
  and _55274_ (_04142_, _04141_, _04135_);
  nor _55275_ (_04143_, _04141_, _04135_);
  nor _55276_ (_04144_, _04143_, _04142_);
  and _55277_ (_04145_, _04144_, _04138_);
  and _55278_ (_04146_, _04145_, _04130_);
  and _55279_ (_04148_, _04146_, _04122_);
  not _55280_ (_04149_, _00358_);
  not _55281_ (_04150_, _04129_);
  and _55282_ (_04151_, _04150_, _04126_);
  and _55283_ (_04152_, _04145_, _04151_);
  and _55284_ (_04153_, _04152_, _04149_);
  or _55285_ (_04154_, _04153_, _04148_);
  not _55286_ (_04155_, _00399_);
  nor _55287_ (_04156_, _04150_, _04126_);
  and _55288_ (_04157_, _04145_, _04156_);
  and _55289_ (_04158_, _04157_, _04155_);
  not _55290_ (_04159_, _00040_);
  nor _55291_ (_04160_, _04144_, _04137_);
  and _55292_ (_04161_, _04160_, _04156_);
  and _55293_ (_04162_, _04161_, _04159_);
  or _55294_ (_04163_, _04162_, _04158_);
  or _55295_ (_04164_, _04163_, _04154_);
  not _55296_ (_04165_, _43768_);
  and _55297_ (_04166_, _04160_, _04130_);
  and _55298_ (_04167_, _04166_, _04165_);
  not _55299_ (_04168_, _43809_);
  and _55300_ (_04169_, _04160_, _04151_);
  and _55301_ (_04170_, _04169_, _04168_);
  or _55302_ (_04171_, _04170_, _04167_);
  not _55303_ (_04172_, _00481_);
  and _55304_ (_04173_, _04141_, _04137_);
  and _55305_ (_04174_, _04173_, _04130_);
  and _55306_ (_04175_, _04174_, _04172_);
  not _55307_ (_04176_, _00522_);
  and _55308_ (_04177_, _04173_, _04151_);
  and _55309_ (_04178_, _04177_, _04176_);
  or _55310_ (_04179_, _04178_, _04175_);
  not _55311_ (_04180_, _00122_);
  not _55312_ (_04181_, _04141_);
  and _55313_ (_04182_, _04181_, _04137_);
  and _55314_ (_04183_, _04182_, _04130_);
  and _55315_ (_04184_, _04183_, _04180_);
  not _55316_ (_04185_, _00194_);
  and _55317_ (_04186_, _04182_, _04151_);
  and _55318_ (_04187_, _04186_, _04185_);
  or _55319_ (_04188_, _04187_, _04184_);
  or _55320_ (_04189_, _04188_, _04179_);
  not _55321_ (_04190_, _00081_);
  and _55322_ (_04191_, _04143_, _04131_);
  and _55323_ (_04192_, _04191_, _04190_);
  not _55324_ (_04193_, _00576_);
  and _55325_ (_04194_, _04134_, _04156_);
  and _55326_ (_04195_, _04194_, _04141_);
  and _55327_ (_04196_, _04195_, _04193_);
  not _55328_ (_04197_, _00276_);
  and _55329_ (_04198_, _04181_, _04135_);
  and _55330_ (_04199_, _04198_, _04197_);
  not _55331_ (_04200_, _43727_);
  and _55332_ (_04201_, _04142_, _04200_);
  or _55333_ (_04202_, _04201_, _04199_);
  or _55334_ (_04203_, _04202_, _04196_);
  or _55335_ (_04204_, _04203_, _04192_);
  not _55336_ (_04205_, _00440_);
  and _55337_ (_04206_, _04173_, _04131_);
  and _55338_ (_04207_, _04206_, _04205_);
  not _55339_ (_04208_, _00235_);
  and _55340_ (_04209_, _04182_, _04156_);
  and _55341_ (_04210_, _04209_, _04208_);
  or _55342_ (_04211_, _04210_, _04207_);
  or _55343_ (_04212_, _04211_, _04204_);
  or _55344_ (_04213_, _04212_, _04189_);
  or _55345_ (_04214_, _04213_, _04171_);
  or _55346_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], _04214_, _04164_);
  and _55347_ (_04215_, _04157_, _04205_);
  and _55348_ (_04216_, _04152_, _04155_);
  or _55349_ (_04217_, _04216_, _04215_);
  and _55350_ (_04218_, _04146_, _04149_);
  and _55351_ (_04219_, _04161_, _04190_);
  or _55352_ (_04220_, _04219_, _04218_);
  or _55353_ (_04221_, _04220_, _04217_);
  and _55354_ (_04222_, _04186_, _04208_);
  and _55355_ (_04223_, _04183_, _04185_);
  or _55356_ (_04224_, _04223_, _04222_);
  and _55357_ (_04225_, _04174_, _04176_);
  and _55358_ (_04226_, _04209_, _04197_);
  or _55359_ (_04227_, _04226_, _04225_);
  or _55360_ (_04228_, _04227_, _04224_);
  and _55361_ (_04229_, _04191_, _04180_);
  and _55362_ (_04230_, _04142_, _04165_);
  and _55363_ (_04231_, _04198_, _04122_);
  and _55364_ (_04232_, _04195_, _04200_);
  or _55365_ (_04233_, _04232_, _04231_);
  or _55366_ (_04234_, _04233_, _04230_);
  or _55367_ (_04235_, _04234_, _04229_);
  and _55368_ (_04236_, _04177_, _04193_);
  and _55369_ (_04237_, _04206_, _04172_);
  or _55370_ (_04238_, _04237_, _04236_);
  or _55371_ (_04239_, _04238_, _04235_);
  or _55372_ (_04240_, _04239_, _04228_);
  and _55373_ (_04241_, _04169_, _04159_);
  and _55374_ (_04242_, _04166_, _04168_);
  or _55375_ (_04243_, _04242_, _04241_);
  or _55376_ (_04244_, _04243_, _04240_);
  or _55377_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], _04244_, _04221_);
  and _55378_ (_04245_, _04146_, _04155_);
  and _55379_ (_04247_, _04152_, _04205_);
  or _55380_ (_04248_, _04247_, _04245_);
  and _55381_ (_04249_, _04157_, _04172_);
  and _55382_ (_04250_, _04161_, _04180_);
  or _55383_ (_04251_, _04250_, _04249_);
  or _55384_ (_04252_, _04251_, _04248_);
  and _55385_ (_04253_, _04169_, _04190_);
  and _55386_ (_04254_, _04166_, _04159_);
  or _55387_ (_04255_, _04254_, _04253_);
  and _55388_ (_04256_, _04209_, _04122_);
  and _55389_ (_04257_, _04186_, _04197_);
  or _55390_ (_04258_, _04257_, _04256_);
  and _55391_ (_04259_, _04183_, _04208_);
  and _55392_ (_04260_, _04177_, _04200_);
  or _55393_ (_04261_, _04260_, _04259_);
  or _55394_ (_04262_, _04261_, _04258_);
  and _55395_ (_04263_, _04191_, _04185_);
  and _55396_ (_04264_, _04142_, _04168_);
  and _55397_ (_04265_, _04198_, _04149_);
  and _55398_ (_04266_, _04195_, _04165_);
  or _55399_ (_04267_, _04266_, _04265_);
  or _55400_ (_04268_, _04267_, _04264_);
  or _55401_ (_04269_, _04268_, _04263_);
  and _55402_ (_04270_, _04174_, _04193_);
  and _55403_ (_04271_, _04206_, _04176_);
  or _55404_ (_04272_, _04271_, _04270_);
  or _55405_ (_04273_, _04272_, _04269_);
  or _55406_ (_04274_, _04273_, _04262_);
  or _55407_ (_04275_, _04274_, _04255_);
  or _55408_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], _04275_, _04252_);
  and _55409_ (_04276_, _04142_, _04193_);
  and _55410_ (_04277_, _04161_, _04168_);
  and _55411_ (_04278_, _04166_, _04200_);
  or _55412_ (_04279_, _04278_, _04277_);
  and _55413_ (_04280_, _04169_, _04165_);
  and _55414_ (_04281_, _04209_, _04185_);
  and _55415_ (_04282_, _04186_, _04180_);
  or _55416_ (_04283_, _04282_, _04281_);
  and _55417_ (_04284_, _04183_, _04190_);
  and _55418_ (_04285_, _04191_, _04159_);
  or _55419_ (_04286_, _04285_, _04284_);
  or _55420_ (_04287_, _04286_, _04283_);
  or _55421_ (_04288_, _04287_, _04280_);
  or _55422_ (_04289_, _04288_, _04279_);
  and _55423_ (_04290_, _04177_, _04172_);
  and _55424_ (_04291_, _04195_, _04176_);
  or _55425_ (_04292_, _04291_, _04290_);
  and _55426_ (_04293_, _04206_, _04155_);
  and _55427_ (_04294_, _04174_, _04205_);
  or _55428_ (_04295_, _04294_, _04293_);
  or _55429_ (_04296_, _04295_, _04292_);
  and _55430_ (_04297_, _04157_, _04149_);
  and _55431_ (_04298_, _04152_, _04122_);
  or _55432_ (_04299_, _04298_, _04297_);
  and _55433_ (_04300_, _04146_, _04197_);
  and _55434_ (_04301_, _04198_, _04208_);
  or _55435_ (_04302_, _04301_, _04300_);
  or _55436_ (_04303_, _04302_, _04299_);
  or _55437_ (_04304_, _04303_, _04296_);
  or _55438_ (_04305_, _04304_, _04289_);
  or _55439_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], _04305_, _04276_);
  not _55440_ (_04306_, _00404_);
  and _55441_ (_04307_, _04146_, _04306_);
  not _55442_ (_04308_, _00127_);
  and _55443_ (_04309_, _04161_, _04308_);
  or _55444_ (_04310_, _04309_, _04307_);
  not _55445_ (_04311_, _00445_);
  and _55446_ (_04312_, _04152_, _04311_);
  not _55447_ (_04313_, _00486_);
  and _55448_ (_04314_, _04157_, _04313_);
  or _55449_ (_04315_, _04314_, _04312_);
  or _55450_ (_04316_, _04315_, _04310_);
  not _55451_ (_04317_, _00045_);
  and _55452_ (_04318_, _04166_, _04317_);
  not _55453_ (_04319_, _00086_);
  and _55454_ (_04320_, _04169_, _04319_);
  or _55455_ (_04321_, _04320_, _04318_);
  not _55456_ (_04322_, _00584_);
  and _55457_ (_04323_, _04174_, _04322_);
  not _55458_ (_04324_, _00322_);
  and _55459_ (_04325_, _04209_, _04324_);
  or _55460_ (_04326_, _04325_, _04323_);
  not _55461_ (_04327_, _00527_);
  and _55462_ (_04328_, _04206_, _04327_);
  not _55463_ (_04329_, _00240_);
  and _55464_ (_04330_, _04183_, _04329_);
  or _55465_ (_04331_, _04330_, _04328_);
  or _55466_ (_04332_, _04331_, _04326_);
  not _55467_ (_04333_, _00199_);
  and _55468_ (_04334_, _04191_, _04333_);
  not _55469_ (_04335_, _43773_);
  and _55470_ (_04336_, _04195_, _04335_);
  not _55471_ (_04337_, _00363_);
  and _55472_ (_04338_, _04198_, _04337_);
  not _55473_ (_04339_, _00004_);
  and _55474_ (_04340_, _04142_, _04339_);
  or _55475_ (_04341_, _04340_, _04338_);
  or _55476_ (_04342_, _04341_, _04336_);
  or _55477_ (_04343_, _04342_, _04334_);
  not _55478_ (_04344_, _00281_);
  and _55479_ (_04346_, _04186_, _04344_);
  not _55480_ (_04347_, _43732_);
  and _55481_ (_04348_, _04177_, _04347_);
  or _55482_ (_04349_, _04348_, _04346_);
  or _55483_ (_04350_, _04349_, _04343_);
  or _55484_ (_04351_, _04350_, _04332_);
  or _55485_ (_04352_, _04351_, _04321_);
  or _55486_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], _04352_, _04316_);
  not _55487_ (_04353_, _00409_);
  and _55488_ (_04354_, _04146_, _04353_);
  not _55489_ (_04355_, _00135_);
  and _55490_ (_04356_, _04161_, _04355_);
  or _55491_ (_04357_, _04356_, _04354_);
  not _55492_ (_04358_, _00450_);
  and _55493_ (_04359_, _04152_, _04358_);
  not _55494_ (_04360_, _00491_);
  and _55495_ (_04361_, _04157_, _04360_);
  or _55496_ (_04362_, _04361_, _04359_);
  or _55497_ (_04363_, _04362_, _04357_);
  not _55498_ (_04364_, _00050_);
  and _55499_ (_04365_, _04166_, _04364_);
  not _55500_ (_04366_, _00091_);
  and _55501_ (_04367_, _04169_, _04366_);
  or _55502_ (_04368_, _04367_, _04365_);
  not _55503_ (_04369_, _00592_);
  and _55504_ (_04370_, _04174_, _04369_);
  not _55505_ (_04371_, _00327_);
  and _55506_ (_04372_, _04209_, _04371_);
  or _55507_ (_04373_, _04372_, _04370_);
  not _55508_ (_04374_, _00532_);
  and _55509_ (_04375_, _04206_, _04374_);
  not _55510_ (_04376_, _00245_);
  and _55511_ (_04377_, _04183_, _04376_);
  or _55512_ (_04378_, _04377_, _04375_);
  or _55513_ (_04379_, _04378_, _04373_);
  not _55514_ (_04380_, _00204_);
  and _55515_ (_04381_, _04191_, _04380_);
  not _55516_ (_04382_, _43778_);
  and _55517_ (_04383_, _04195_, _04382_);
  not _55518_ (_04384_, _00368_);
  and _55519_ (_04385_, _04198_, _04384_);
  not _55520_ (_04386_, _00009_);
  and _55521_ (_04387_, _04142_, _04386_);
  or _55522_ (_04388_, _04387_, _04385_);
  or _55523_ (_04389_, _04388_, _04383_);
  or _55524_ (_04390_, _04389_, _04381_);
  not _55525_ (_04391_, _00286_);
  and _55526_ (_04392_, _04186_, _04391_);
  not _55527_ (_04393_, _43737_);
  and _55528_ (_04394_, _04177_, _04393_);
  or _55529_ (_04395_, _04394_, _04392_);
  or _55530_ (_04396_, _04395_, _04390_);
  or _55531_ (_04397_, _04396_, _04379_);
  or _55532_ (_04398_, _04397_, _04368_);
  or _55533_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], _04398_, _04363_);
  not _55534_ (_04399_, _00455_);
  and _55535_ (_04400_, _04152_, _04399_);
  not _55536_ (_04401_, _00146_);
  and _55537_ (_04402_, _04161_, _04401_);
  or _55538_ (_04403_, _04402_, _04400_);
  not _55539_ (_04404_, _00496_);
  and _55540_ (_04405_, _04157_, _04404_);
  not _55541_ (_04406_, _00414_);
  and _55542_ (_04407_, _04146_, _04406_);
  or _55543_ (_04408_, _04407_, _04405_);
  or _55544_ (_04409_, _04408_, _04403_);
  not _55545_ (_04410_, _00096_);
  and _55546_ (_04411_, _04169_, _04410_);
  not _55547_ (_04412_, _00055_);
  and _55548_ (_04413_, _04166_, _04412_);
  or _55549_ (_04414_, _04413_, _04411_);
  not _55550_ (_04415_, _00537_);
  and _55551_ (_04416_, _04206_, _04415_);
  not _55552_ (_04417_, _43742_);
  and _55553_ (_04418_, _04177_, _04417_);
  or _55554_ (_04419_, _04418_, _04416_);
  not _55555_ (_04420_, _00332_);
  and _55556_ (_04421_, _04209_, _04420_);
  not _55557_ (_04422_, _00250_);
  and _55558_ (_04423_, _04183_, _04422_);
  or _55559_ (_04424_, _04423_, _04421_);
  or _55560_ (_04425_, _04424_, _04419_);
  not _55561_ (_04426_, _00209_);
  and _55562_ (_04427_, _04191_, _04426_);
  not _55563_ (_04428_, _00373_);
  and _55564_ (_04429_, _04198_, _04428_);
  not _55565_ (_04430_, _43783_);
  and _55566_ (_04431_, _04195_, _04430_);
  not _55567_ (_04432_, _00014_);
  and _55568_ (_04433_, _04142_, _04432_);
  or _55569_ (_04434_, _04433_, _04431_);
  or _55570_ (_04435_, _04434_, _04429_);
  or _55571_ (_04436_, _04435_, _04427_);
  not _55572_ (_04437_, _00597_);
  and _55573_ (_04438_, _04174_, _04437_);
  not _55574_ (_04439_, _00291_);
  and _55575_ (_04440_, _04186_, _04439_);
  or _55576_ (_04441_, _04440_, _04438_);
  or _55577_ (_04442_, _04441_, _04436_);
  or _55578_ (_04443_, _04442_, _04425_);
  or _55579_ (_04445_, _04443_, _04414_);
  or _55580_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], _04445_, _04409_);
  not _55581_ (_04446_, _00419_);
  and _55582_ (_04447_, _04146_, _04446_);
  not _55583_ (_04448_, _00157_);
  and _55584_ (_04449_, _04161_, _04448_);
  or _55585_ (_04450_, _04449_, _04447_);
  not _55586_ (_04451_, _00460_);
  and _55587_ (_04452_, _04152_, _04451_);
  not _55588_ (_04453_, _00501_);
  and _55589_ (_04454_, _04157_, _04453_);
  or _55590_ (_04455_, _04454_, _04452_);
  or _55591_ (_04456_, _04455_, _04450_);
  not _55592_ (_04457_, _00060_);
  and _55593_ (_04458_, _04166_, _04457_);
  not _55594_ (_04459_, _00101_);
  and _55595_ (_04460_, _04169_, _04459_);
  or _55596_ (_04461_, _04460_, _04458_);
  not _55597_ (_04462_, _00602_);
  and _55598_ (_04463_, _04174_, _04462_);
  not _55599_ (_04464_, _00337_);
  and _55600_ (_04465_, _04209_, _04464_);
  or _55601_ (_04466_, _04465_, _04463_);
  not _55602_ (_04467_, _00542_);
  and _55603_ (_04468_, _04206_, _04467_);
  not _55604_ (_04469_, _00255_);
  and _55605_ (_04470_, _04183_, _04469_);
  or _55606_ (_04471_, _04470_, _04468_);
  or _55607_ (_04472_, _04471_, _04466_);
  not _55608_ (_04473_, _00214_);
  and _55609_ (_04474_, _04191_, _04473_);
  not _55610_ (_04475_, _43788_);
  and _55611_ (_04476_, _04195_, _04475_);
  not _55612_ (_04477_, _00378_);
  and _55613_ (_04478_, _04198_, _04477_);
  not _55614_ (_04479_, _00019_);
  and _55615_ (_04480_, _04142_, _04479_);
  or _55616_ (_04481_, _04480_, _04478_);
  or _55617_ (_04482_, _04481_, _04476_);
  or _55618_ (_04483_, _04482_, _04474_);
  not _55619_ (_04484_, _00296_);
  and _55620_ (_04485_, _04186_, _04484_);
  not _55621_ (_04486_, _43747_);
  and _55622_ (_04487_, _04177_, _04486_);
  or _55623_ (_04488_, _04487_, _04485_);
  or _55624_ (_04489_, _04488_, _04483_);
  or _55625_ (_04490_, _04489_, _04472_);
  or _55626_ (_04491_, _04490_, _04461_);
  or _55627_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], _04491_, _04456_);
  not _55628_ (_04492_, _00424_);
  and _55629_ (_04493_, _04146_, _04492_);
  not _55630_ (_04494_, _00168_);
  and _55631_ (_04495_, _04161_, _04494_);
  or _55632_ (_04496_, _04495_, _04493_);
  not _55633_ (_04497_, _00465_);
  and _55634_ (_04498_, _04152_, _04497_);
  not _55635_ (_04499_, _00506_);
  and _55636_ (_04500_, _04157_, _04499_);
  or _55637_ (_04501_, _04500_, _04498_);
  or _55638_ (_04502_, _04501_, _04496_);
  not _55639_ (_04503_, _00065_);
  and _55640_ (_04504_, _04166_, _04503_);
  not _55641_ (_04505_, _00106_);
  and _55642_ (_04506_, _04169_, _04505_);
  or _55643_ (_04507_, _04506_, _04504_);
  not _55644_ (_04508_, _00607_);
  and _55645_ (_04509_, _04174_, _04508_);
  not _55646_ (_04510_, _00342_);
  and _55647_ (_04511_, _04209_, _04510_);
  or _55648_ (_04512_, _04511_, _04509_);
  not _55649_ (_04513_, _00550_);
  and _55650_ (_04514_, _04206_, _04513_);
  not _55651_ (_04515_, _00260_);
  and _55652_ (_04516_, _04183_, _04515_);
  or _55653_ (_04517_, _04516_, _04514_);
  or _55654_ (_04518_, _04517_, _04512_);
  not _55655_ (_04519_, _00219_);
  and _55656_ (_04520_, _04191_, _04519_);
  not _55657_ (_04521_, _43793_);
  and _55658_ (_04522_, _04195_, _04521_);
  not _55659_ (_04523_, _00383_);
  and _55660_ (_04524_, _04198_, _04523_);
  not _55661_ (_04525_, _00024_);
  and _55662_ (_04526_, _04142_, _04525_);
  or _55663_ (_04527_, _04526_, _04524_);
  or _55664_ (_04528_, _04527_, _04522_);
  or _55665_ (_04529_, _04528_, _04520_);
  not _55666_ (_04530_, _00301_);
  and _55667_ (_04531_, _04186_, _04530_);
  not _55668_ (_04532_, _43752_);
  and _55669_ (_04533_, _04177_, _04532_);
  or _55670_ (_04534_, _04533_, _04531_);
  or _55671_ (_04535_, _04534_, _04529_);
  or _55672_ (_04536_, _04535_, _04518_);
  or _55673_ (_04537_, _04536_, _04507_);
  or _55674_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], _04537_, _04502_);
  not _55675_ (_04538_, _00511_);
  and _55676_ (_04539_, _04157_, _04538_);
  not _55677_ (_04540_, _00429_);
  and _55678_ (_04541_, _04146_, _04540_);
  or _55679_ (_04543_, _04541_, _04539_);
  not _55680_ (_04544_, _00470_);
  and _55681_ (_04545_, _04152_, _04544_);
  not _55682_ (_04546_, _00179_);
  and _55683_ (_04547_, _04161_, _04546_);
  or _55684_ (_04548_, _04547_, _04545_);
  or _55685_ (_04549_, _04548_, _04543_);
  not _55686_ (_04550_, _00111_);
  and _55687_ (_04551_, _04169_, _04550_);
  not _55688_ (_04552_, _00070_);
  and _55689_ (_04553_, _04166_, _04552_);
  or _55690_ (_04554_, _04553_, _04551_);
  not _55691_ (_04555_, _00347_);
  and _55692_ (_04556_, _04209_, _04555_);
  not _55693_ (_04557_, _00306_);
  and _55694_ (_04558_, _04186_, _04557_);
  or _55695_ (_04559_, _04558_, _04556_);
  not _55696_ (_04560_, _00265_);
  and _55697_ (_04561_, _04183_, _04560_);
  not _55698_ (_04562_, _43757_);
  and _55699_ (_04563_, _04177_, _04562_);
  or _55700_ (_04564_, _04563_, _04561_);
  or _55701_ (_04565_, _04564_, _04559_);
  not _55702_ (_04566_, _00224_);
  and _55703_ (_04567_, _04191_, _04566_);
  not _55704_ (_04568_, _00029_);
  and _55705_ (_04569_, _04142_, _04568_);
  not _55706_ (_04570_, _00388_);
  and _55707_ (_04571_, _04198_, _04570_);
  not _55708_ (_04572_, _43798_);
  and _55709_ (_04573_, _04195_, _04572_);
  or _55710_ (_04574_, _04573_, _04571_);
  or _55711_ (_04575_, _04574_, _04569_);
  or _55712_ (_04576_, _04575_, _04567_);
  not _55713_ (_04577_, _00612_);
  and _55714_ (_04578_, _04174_, _04577_);
  not _55715_ (_04579_, _00558_);
  and _55716_ (_04580_, _04206_, _04579_);
  or _55717_ (_04581_, _04580_, _04578_);
  or _55718_ (_04582_, _04581_, _04576_);
  or _55719_ (_04583_, _04582_, _04565_);
  or _55720_ (_04584_, _04583_, _04554_);
  or _55721_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], _04584_, _04549_);
  not _55722_ (_04585_, _00434_);
  and _55723_ (_04586_, _04146_, _04585_);
  not _55724_ (_04587_, _00475_);
  and _55725_ (_04588_, _04152_, _04587_);
  or _55726_ (_04589_, _04588_, _04586_);
  not _55727_ (_04590_, _00516_);
  and _55728_ (_04591_, _04157_, _04590_);
  not _55729_ (_04592_, _00188_);
  and _55730_ (_04593_, _04161_, _04592_);
  or _55731_ (_04594_, _04593_, _04591_);
  or _55732_ (_04595_, _04594_, _04589_);
  not _55733_ (_04596_, _00116_);
  and _55734_ (_04597_, _04169_, _04596_);
  not _55735_ (_04598_, _00075_);
  and _55736_ (_04599_, _04166_, _04598_);
  or _55737_ (_04600_, _04599_, _04597_);
  not _55738_ (_04601_, _00352_);
  and _55739_ (_04602_, _04209_, _04601_);
  not _55740_ (_04603_, _00311_);
  and _55741_ (_04604_, _04186_, _04603_);
  or _55742_ (_04605_, _04604_, _04602_);
  not _55743_ (_04606_, _00270_);
  and _55744_ (_04607_, _04183_, _04606_);
  not _55745_ (_04608_, _43762_);
  and _55746_ (_04609_, _04177_, _04608_);
  or _55747_ (_04610_, _04609_, _04607_);
  or _55748_ (_04611_, _04610_, _04605_);
  not _55749_ (_04612_, _00229_);
  and _55750_ (_04613_, _04191_, _04612_);
  not _55751_ (_04614_, _00034_);
  and _55752_ (_04615_, _04142_, _04614_);
  not _55753_ (_04616_, _00393_);
  and _55754_ (_04617_, _04198_, _04616_);
  not _55755_ (_04618_, _43803_);
  and _55756_ (_04619_, _04195_, _04618_);
  or _55757_ (_04620_, _04619_, _04617_);
  or _55758_ (_04621_, _04620_, _04615_);
  or _55759_ (_04622_, _04621_, _04613_);
  not _55760_ (_04623_, _00617_);
  and _55761_ (_04624_, _04174_, _04623_);
  not _55762_ (_04625_, _00566_);
  and _55763_ (_04626_, _04206_, _04625_);
  or _55764_ (_04627_, _04626_, _04624_);
  or _55765_ (_04628_, _04627_, _04622_);
  or _55766_ (_04629_, _04628_, _04611_);
  or _55767_ (_04630_, _04629_, _04600_);
  or _55768_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], _04630_, _04595_);
  and _55769_ (_04631_, _04157_, _04311_);
  and _55770_ (_04632_, _04161_, _04319_);
  or _55771_ (_04633_, _04632_, _04631_);
  and _55772_ (_04634_, _04152_, _04306_);
  and _55773_ (_04635_, _04146_, _04337_);
  or _55774_ (_04636_, _04635_, _04634_);
  or _55775_ (_04637_, _04636_, _04633_);
  and _55776_ (_04638_, _04209_, _04344_);
  and _55777_ (_04639_, _04183_, _04333_);
  or _55778_ (_04640_, _04639_, _04638_);
  and _55779_ (_04642_, _04206_, _04313_);
  and _55780_ (_04643_, _04186_, _04329_);
  or _55781_ (_04644_, _04643_, _04642_);
  or _55782_ (_04645_, _04644_, _04640_);
  and _55783_ (_04646_, _04191_, _04308_);
  and _55784_ (_04647_, _04198_, _04324_);
  and _55785_ (_04648_, _04195_, _04347_);
  and _55786_ (_04649_, _04142_, _04335_);
  or _55787_ (_04650_, _04649_, _04648_);
  or _55788_ (_04651_, _04650_, _04647_);
  or _55789_ (_04652_, _04651_, _04646_);
  and _55790_ (_04653_, _04177_, _04322_);
  and _55791_ (_04654_, _04174_, _04327_);
  or _55792_ (_04655_, _04654_, _04653_);
  or _55793_ (_04656_, _04655_, _04652_);
  or _55794_ (_04657_, _04656_, _04645_);
  and _55795_ (_04658_, _04169_, _04317_);
  and _55796_ (_04659_, _04166_, _04339_);
  or _55797_ (_04660_, _04659_, _04658_);
  or _55798_ (_04661_, _04660_, _04657_);
  or _55799_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], _04661_, _04637_);
  and _55800_ (_04662_, _04157_, _04358_);
  and _55801_ (_04663_, _04152_, _04353_);
  or _55802_ (_04664_, _04663_, _04662_);
  and _55803_ (_04665_, _04146_, _04384_);
  and _55804_ (_04666_, _04161_, _04366_);
  or _55805_ (_04667_, _04666_, _04665_);
  or _55806_ (_04668_, _04667_, _04664_);
  and _55807_ (_04669_, _04186_, _04376_);
  and _55808_ (_04670_, _04183_, _04380_);
  or _55809_ (_04671_, _04670_, _04669_);
  and _55810_ (_04672_, _04174_, _04374_);
  and _55811_ (_04673_, _04209_, _04391_);
  or _55812_ (_04674_, _04673_, _04672_);
  or _55813_ (_04675_, _04674_, _04671_);
  and _55814_ (_04676_, _04191_, _04355_);
  and _55815_ (_04677_, _04142_, _04382_);
  and _55816_ (_04678_, _04198_, _04371_);
  and _55817_ (_04679_, _04195_, _04393_);
  or _55818_ (_04680_, _04679_, _04678_);
  or _55819_ (_04681_, _04680_, _04677_);
  or _55820_ (_04682_, _04681_, _04676_);
  and _55821_ (_04683_, _04177_, _04369_);
  and _55822_ (_04684_, _04206_, _04360_);
  or _55823_ (_04685_, _04684_, _04683_);
  or _55824_ (_04686_, _04685_, _04682_);
  or _55825_ (_04687_, _04686_, _04675_);
  and _55826_ (_04688_, _04169_, _04364_);
  and _55827_ (_04689_, _04166_, _04386_);
  or _55828_ (_04690_, _04689_, _04688_);
  or _55829_ (_04691_, _04690_, _04687_);
  or _55830_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], _04691_, _04668_);
  and _55831_ (_04692_, _04157_, _04399_);
  and _55832_ (_04693_, _04161_, _04410_);
  or _55833_ (_04694_, _04693_, _04692_);
  and _55834_ (_04695_, _04152_, _04406_);
  and _55835_ (_04696_, _04146_, _04428_);
  or _55836_ (_04697_, _04696_, _04695_);
  or _55837_ (_04698_, _04697_, _04694_);
  and _55838_ (_04699_, _04177_, _04437_);
  and _55839_ (_04700_, _04174_, _04415_);
  or _55840_ (_04701_, _04700_, _04699_);
  and _55841_ (_04702_, _04209_, _04439_);
  and _55842_ (_04703_, _04183_, _04426_);
  or _55843_ (_04704_, _04703_, _04702_);
  or _55844_ (_04705_, _04704_, _04701_);
  and _55845_ (_04706_, _04191_, _04401_);
  and _55846_ (_04707_, _04198_, _04420_);
  and _55847_ (_04708_, _04195_, _04417_);
  and _55848_ (_04709_, _04142_, _04430_);
  or _55849_ (_04710_, _04709_, _04708_);
  or _55850_ (_04711_, _04710_, _04707_);
  or _55851_ (_04712_, _04711_, _04706_);
  and _55852_ (_04713_, _04206_, _04404_);
  and _55853_ (_04714_, _04186_, _04422_);
  or _55854_ (_04715_, _04714_, _04713_);
  or _55855_ (_04716_, _04715_, _04712_);
  or _55856_ (_04717_, _04716_, _04705_);
  and _55857_ (_04718_, _04169_, _04412_);
  and _55858_ (_04719_, _04166_, _04432_);
  or _55859_ (_04720_, _04719_, _04718_);
  or _55860_ (_04721_, _04720_, _04717_);
  or _55861_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], _04721_, _04698_);
  and _55862_ (_04722_, _04152_, _04446_);
  and _55863_ (_04723_, _04157_, _04451_);
  or _55864_ (_04724_, _04723_, _04722_);
  and _55865_ (_04725_, _04146_, _04477_);
  and _55866_ (_04726_, _04161_, _04459_);
  or _55867_ (_04727_, _04726_, _04725_);
  or _55868_ (_04728_, _04727_, _04724_);
  and _55869_ (_04729_, _04186_, _04469_);
  and _55870_ (_04730_, _04183_, _04473_);
  or _55871_ (_04731_, _04730_, _04729_);
  and _55872_ (_04732_, _04177_, _04462_);
  and _55873_ (_04733_, _04206_, _04453_);
  or _55874_ (_04734_, _04733_, _04732_);
  or _55875_ (_04735_, _04734_, _04731_);
  and _55876_ (_04736_, _04191_, _04448_);
  and _55877_ (_04737_, _04195_, _04486_);
  and _55878_ (_04738_, _04198_, _04464_);
  and _55879_ (_04739_, _04142_, _04475_);
  or _55880_ (_04740_, _04739_, _04738_);
  or _55881_ (_04741_, _04740_, _04737_);
  or _55882_ (_04742_, _04741_, _04736_);
  and _55883_ (_04743_, _04174_, _04467_);
  and _55884_ (_04744_, _04209_, _04484_);
  or _55885_ (_04745_, _04744_, _04743_);
  or _55886_ (_04746_, _04745_, _04742_);
  or _55887_ (_04747_, _04746_, _04735_);
  and _55888_ (_04748_, _04169_, _04457_);
  and _55889_ (_04749_, _04166_, _04479_);
  or _55890_ (_04750_, _04749_, _04748_);
  or _55891_ (_04751_, _04750_, _04747_);
  or _55892_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], _04751_, _04728_);
  and _55893_ (_04752_, _04157_, _04497_);
  and _55894_ (_04753_, _04146_, _04523_);
  or _55895_ (_04754_, _04753_, _04752_);
  and _55896_ (_04755_, _04152_, _04492_);
  and _55897_ (_04756_, _04161_, _04505_);
  or _55898_ (_04757_, _04756_, _04755_);
  or _55899_ (_04758_, _04757_, _04754_);
  and _55900_ (_04759_, _04186_, _04515_);
  and _55901_ (_04760_, _04183_, _04519_);
  or _55902_ (_04761_, _04760_, _04759_);
  and _55903_ (_04762_, _04174_, _04513_);
  and _55904_ (_04763_, _04209_, _04530_);
  or _55905_ (_04764_, _04763_, _04762_);
  or _55906_ (_04765_, _04764_, _04761_);
  and _55907_ (_04766_, _04191_, _04494_);
  and _55908_ (_04767_, _04142_, _04521_);
  and _55909_ (_04768_, _04198_, _04510_);
  and _55910_ (_04769_, _04195_, _04532_);
  or _55911_ (_04770_, _04769_, _04768_);
  or _55912_ (_04771_, _04770_, _04767_);
  or _55913_ (_04772_, _04771_, _04766_);
  and _55914_ (_04773_, _04177_, _04508_);
  and _55915_ (_04774_, _04206_, _04499_);
  or _55916_ (_04775_, _04774_, _04773_);
  or _55917_ (_04776_, _04775_, _04772_);
  or _55918_ (_04777_, _04776_, _04765_);
  and _55919_ (_04778_, _04169_, _04503_);
  and _55920_ (_04779_, _04166_, _04525_);
  or _55921_ (_04780_, _04779_, _04778_);
  or _55922_ (_04781_, _04780_, _04777_);
  or _55923_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], _04781_, _04758_);
  and _55924_ (_04782_, _04152_, _04540_);
  and _55925_ (_04783_, _04157_, _04544_);
  or _55926_ (_04784_, _04783_, _04782_);
  and _55927_ (_04785_, _04146_, _04570_);
  and _55928_ (_04786_, _04161_, _04550_);
  or _55929_ (_04787_, _04786_, _04785_);
  or _55930_ (_04788_, _04787_, _04784_);
  and _55931_ (_04789_, _04186_, _04560_);
  and _55932_ (_04790_, _04183_, _04566_);
  or _55933_ (_04791_, _04790_, _04789_);
  and _55934_ (_04792_, _04177_, _04577_);
  and _55935_ (_04793_, _04206_, _04538_);
  or _55936_ (_04794_, _04793_, _04792_);
  or _55937_ (_04795_, _04794_, _04791_);
  and _55938_ (_04796_, _04191_, _04546_);
  and _55939_ (_04797_, _04195_, _04562_);
  and _55940_ (_04798_, _04198_, _04555_);
  and _55941_ (_04799_, _04142_, _04572_);
  or _55942_ (_04800_, _04799_, _04798_);
  or _55943_ (_04801_, _04800_, _04797_);
  or _55944_ (_04802_, _04801_, _04796_);
  and _55945_ (_04803_, _04174_, _04579_);
  and _55946_ (_04804_, _04209_, _04557_);
  or _55947_ (_04805_, _04804_, _04803_);
  or _55948_ (_04806_, _04805_, _04802_);
  or _55949_ (_04807_, _04806_, _04795_);
  and _55950_ (_04808_, _04169_, _04552_);
  and _55951_ (_04809_, _04166_, _04568_);
  or _55952_ (_04810_, _04809_, _04808_);
  or _55953_ (_04811_, _04810_, _04807_);
  or _55954_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], _04811_, _04788_);
  and _55955_ (_04812_, _04157_, _04587_);
  and _55956_ (_04813_, _04146_, _04616_);
  or _55957_ (_04814_, _04813_, _04812_);
  and _55958_ (_04815_, _04152_, _04585_);
  and _55959_ (_04816_, _04161_, _04596_);
  or _55960_ (_04817_, _04816_, _04815_);
  or _55961_ (_04818_, _04817_, _04814_);
  and _55962_ (_04819_, _04186_, _04606_);
  and _55963_ (_04820_, _04183_, _04612_);
  or _55964_ (_04821_, _04820_, _04819_);
  and _55965_ (_04822_, _04174_, _04625_);
  and _55966_ (_04823_, _04209_, _04603_);
  or _55967_ (_04824_, _04823_, _04822_);
  or _55968_ (_04825_, _04824_, _04821_);
  and _55969_ (_04826_, _04191_, _04592_);
  and _55970_ (_04827_, _04142_, _04618_);
  and _55971_ (_04828_, _04198_, _04601_);
  and _55972_ (_04829_, _04195_, _04608_);
  or _55973_ (_04830_, _04829_, _04828_);
  or _55974_ (_04831_, _04830_, _04827_);
  or _55975_ (_04832_, _04831_, _04826_);
  and _55976_ (_04833_, _04177_, _04623_);
  and _55977_ (_04834_, _04206_, _04590_);
  or _55978_ (_04835_, _04834_, _04833_);
  or _55979_ (_04836_, _04835_, _04832_);
  or _55980_ (_04837_, _04836_, _04825_);
  and _55981_ (_04838_, _04169_, _04598_);
  and _55982_ (_04839_, _04166_, _04614_);
  or _55983_ (_04840_, _04839_, _04838_);
  or _55984_ (_04841_, _04840_, _04837_);
  or _55985_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], _04841_, _04818_);
  and _55986_ (_04842_, _04161_, _04339_);
  and _55987_ (_04843_, _04157_, _04337_);
  or _55988_ (_04844_, _04843_, _04842_);
  and _55989_ (_04845_, _04152_, _04324_);
  and _55990_ (_04846_, _04146_, _04344_);
  or _55991_ (_04847_, _04846_, _04845_);
  or _55992_ (_04848_, _04847_, _04844_);
  and _55993_ (_04849_, _04183_, _04319_);
  and _55994_ (_04850_, _04177_, _04313_);
  or _55995_ (_04851_, _04850_, _04849_);
  and _55996_ (_04852_, _04209_, _04333_);
  and _55997_ (_04853_, _04206_, _04306_);
  or _55998_ (_04854_, _04853_, _04852_);
  or _55999_ (_04855_, _04854_, _04851_);
  and _56000_ (_04856_, _04191_, _04317_);
  and _56001_ (_04857_, _04198_, _04329_);
  and _56002_ (_04858_, _04142_, _04322_);
  and _56003_ (_04859_, _04195_, _04327_);
  or _56004_ (_04860_, _04859_, _04858_);
  or _56005_ (_04861_, _04860_, _04857_);
  or _56006_ (_04862_, _04861_, _04856_);
  and _56007_ (_04863_, _04186_, _04308_);
  and _56008_ (_04864_, _04174_, _04311_);
  or _56009_ (_04865_, _04864_, _04863_);
  or _56010_ (_04866_, _04865_, _04862_);
  or _56011_ (_04867_, _04866_, _04855_);
  and _56012_ (_04868_, _04166_, _04347_);
  and _56013_ (_04869_, _04169_, _04335_);
  or _56014_ (_04870_, _04869_, _04868_);
  or _56015_ (_04871_, _04870_, _04867_);
  or _56016_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], _04871_, _04848_);
  and _56017_ (_04872_, _04152_, _04371_);
  and _56018_ (_04873_, _04157_, _04384_);
  or _56019_ (_04874_, _04873_, _04872_);
  and _56020_ (_04875_, _04146_, _04391_);
  and _56021_ (_04876_, _04161_, _04386_);
  or _56022_ (_04877_, _04876_, _04875_);
  or _56023_ (_04878_, _04877_, _04874_);
  and _56024_ (_04879_, _04177_, _04360_);
  and _56025_ (_04880_, _04183_, _04366_);
  or _56026_ (_04881_, _04880_, _04879_);
  and _56027_ (_04882_, _04206_, _04353_);
  and _56028_ (_04883_, _04209_, _04380_);
  or _56029_ (_04884_, _04883_, _04882_);
  or _56030_ (_04885_, _04884_, _04881_);
  and _56031_ (_04886_, _04191_, _04364_);
  and _56032_ (_04887_, _04142_, _04369_);
  and _56033_ (_04888_, _04195_, _04374_);
  and _56034_ (_04889_, _04198_, _04376_);
  or _56035_ (_04890_, _04889_, _04888_);
  or _56036_ (_04891_, _04890_, _04887_);
  or _56037_ (_04892_, _04891_, _04886_);
  and _56038_ (_04893_, _04174_, _04358_);
  and _56039_ (_04894_, _04186_, _04355_);
  or _56040_ (_04895_, _04894_, _04893_);
  or _56041_ (_04896_, _04895_, _04892_);
  or _56042_ (_04897_, _04896_, _04885_);
  and _56043_ (_04898_, _04166_, _04393_);
  and _56044_ (_04899_, _04169_, _04382_);
  or _56045_ (_04900_, _04899_, _04898_);
  or _56046_ (_04901_, _04900_, _04897_);
  or _56047_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], _04901_, _04878_);
  and _56048_ (_04902_, _04142_, _04437_);
  and _56049_ (_04903_, _04161_, _04432_);
  and _56050_ (_04904_, _04166_, _04417_);
  or _56051_ (_04905_, _04904_, _04903_);
  and _56052_ (_04906_, _04169_, _04430_);
  and _56053_ (_04907_, _04209_, _04426_);
  and _56054_ (_04908_, _04186_, _04401_);
  or _56055_ (_04909_, _04908_, _04907_);
  and _56056_ (_04910_, _04183_, _04410_);
  and _56057_ (_04911_, _04191_, _04412_);
  or _56058_ (_04912_, _04911_, _04910_);
  or _56059_ (_04913_, _04912_, _04909_);
  or _56060_ (_04914_, _04913_, _04906_);
  or _56061_ (_04915_, _04914_, _04905_);
  and _56062_ (_04916_, _04177_, _04404_);
  and _56063_ (_04917_, _04195_, _04415_);
  or _56064_ (_04918_, _04917_, _04916_);
  and _56065_ (_04919_, _04206_, _04406_);
  and _56066_ (_04920_, _04174_, _04399_);
  or _56067_ (_04921_, _04920_, _04919_);
  or _56068_ (_04922_, _04921_, _04918_);
  and _56069_ (_04923_, _04157_, _04428_);
  and _56070_ (_04924_, _04152_, _04420_);
  or _56071_ (_04925_, _04924_, _04923_);
  and _56072_ (_04926_, _04146_, _04439_);
  and _56073_ (_04927_, _04198_, _04422_);
  or _56074_ (_04928_, _04927_, _04926_);
  or _56075_ (_04929_, _04928_, _04925_);
  or _56076_ (_04930_, _04929_, _04922_);
  or _56077_ (_04931_, _04930_, _04915_);
  or _56078_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], _04931_, _04902_);
  and _56079_ (_04932_, _04142_, _04462_);
  and _56080_ (_04933_, _04161_, _04479_);
  and _56081_ (_04934_, _04166_, _04486_);
  or _56082_ (_04935_, _04934_, _04933_);
  and _56083_ (_04936_, _04169_, _04475_);
  and _56084_ (_04937_, _04209_, _04473_);
  and _56085_ (_04938_, _04186_, _04448_);
  or _56086_ (_04939_, _04938_, _04937_);
  and _56087_ (_04940_, _04183_, _04459_);
  and _56088_ (_04941_, _04191_, _04457_);
  or _56089_ (_04942_, _04941_, _04940_);
  or _56090_ (_04943_, _04942_, _04939_);
  or _56091_ (_04944_, _04943_, _04936_);
  or _56092_ (_04945_, _04944_, _04935_);
  and _56093_ (_04946_, _04177_, _04453_);
  and _56094_ (_04947_, _04195_, _04467_);
  or _56095_ (_04948_, _04947_, _04946_);
  and _56096_ (_04949_, _04206_, _04446_);
  and _56097_ (_04950_, _04174_, _04451_);
  or _56098_ (_04951_, _04950_, _04949_);
  or _56099_ (_04952_, _04951_, _04948_);
  and _56100_ (_04953_, _04157_, _04477_);
  and _56101_ (_04954_, _04152_, _04464_);
  or _56102_ (_04955_, _04954_, _04953_);
  and _56103_ (_04956_, _04146_, _04484_);
  and _56104_ (_04957_, _04198_, _04469_);
  or _56105_ (_04958_, _04957_, _04956_);
  or _56106_ (_04959_, _04958_, _04955_);
  or _56107_ (_04960_, _04959_, _04952_);
  or _56108_ (_04961_, _04960_, _04945_);
  or _56109_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], _04961_, _04932_);
  and _56110_ (_04962_, _04152_, _04510_);
  and _56111_ (_04963_, _04161_, _04525_);
  or _56112_ (_04964_, _04963_, _04962_);
  and _56113_ (_04965_, _04157_, _04523_);
  and _56114_ (_04966_, _04146_, _04530_);
  or _56115_ (_04967_, _04966_, _04965_);
  or _56116_ (_04968_, _04967_, _04964_);
  and _56117_ (_04969_, _04177_, _04499_);
  and _56118_ (_04970_, _04183_, _04505_);
  or _56119_ (_04971_, _04970_, _04969_);
  and _56120_ (_04972_, _04206_, _04492_);
  and _56121_ (_04973_, _04209_, _04519_);
  or _56122_ (_04974_, _04973_, _04972_);
  or _56123_ (_04975_, _04974_, _04971_);
  and _56124_ (_04976_, _04191_, _04503_);
  and _56125_ (_04977_, _04142_, _04508_);
  and _56126_ (_04978_, _04195_, _04513_);
  and _56127_ (_04979_, _04198_, _04515_);
  or _56128_ (_04980_, _04979_, _04978_);
  or _56129_ (_04981_, _04980_, _04977_);
  or _56130_ (_04982_, _04981_, _04976_);
  and _56131_ (_04983_, _04174_, _04497_);
  and _56132_ (_04984_, _04186_, _04494_);
  or _56133_ (_04985_, _04984_, _04983_);
  or _56134_ (_04986_, _04985_, _04982_);
  or _56135_ (_04987_, _04986_, _04975_);
  and _56136_ (_04988_, _04166_, _04532_);
  and _56137_ (_04989_, _04169_, _04521_);
  or _56138_ (_04990_, _04989_, _04988_);
  or _56139_ (_04991_, _04990_, _04987_);
  or _56140_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], _04991_, _04968_);
  and _56141_ (_04992_, _04152_, _04555_);
  and _56142_ (_04993_, _04157_, _04570_);
  or _56143_ (_04994_, _04993_, _04992_);
  and _56144_ (_04995_, _04146_, _04557_);
  and _56145_ (_04996_, _04161_, _04568_);
  or _56146_ (_04997_, _04996_, _04995_);
  or _56147_ (_04998_, _04997_, _04994_);
  and _56148_ (_04999_, _04177_, _04538_);
  and _56149_ (_05000_, _04183_, _04550_);
  or _56150_ (_05001_, _05000_, _04999_);
  and _56151_ (_05002_, _04206_, _04540_);
  and _56152_ (_05003_, _04209_, _04566_);
  or _56153_ (_05004_, _05003_, _05002_);
  or _56154_ (_05005_, _05004_, _05001_);
  and _56155_ (_05006_, _04191_, _04552_);
  and _56156_ (_05007_, _04142_, _04577_);
  and _56157_ (_05008_, _04195_, _04579_);
  and _56158_ (_05009_, _04198_, _04560_);
  or _56159_ (_05010_, _05009_, _05008_);
  or _56160_ (_05011_, _05010_, _05007_);
  or _56161_ (_05012_, _05011_, _05006_);
  and _56162_ (_05013_, _04174_, _04544_);
  and _56163_ (_05014_, _04186_, _04546_);
  or _56164_ (_05015_, _05014_, _05013_);
  or _56165_ (_05016_, _05015_, _05012_);
  or _56166_ (_05017_, _05016_, _05005_);
  and _56167_ (_05018_, _04166_, _04562_);
  and _56168_ (_05019_, _04169_, _04572_);
  or _56169_ (_05020_, _05019_, _05018_);
  or _56170_ (_05021_, _05020_, _05017_);
  or _56171_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], _05021_, _04998_);
  and _56172_ (_05022_, _04142_, _04623_);
  and _56173_ (_05023_, _04161_, _04614_);
  and _56174_ (_05024_, _04166_, _04608_);
  or _56175_ (_05025_, _05024_, _05023_);
  and _56176_ (_05026_, _04169_, _04618_);
  and _56177_ (_05027_, _04209_, _04612_);
  and _56178_ (_05028_, _04186_, _04592_);
  or _56179_ (_05029_, _05028_, _05027_);
  and _56180_ (_05030_, _04183_, _04596_);
  and _56181_ (_05031_, _04191_, _04598_);
  or _56182_ (_05032_, _05031_, _05030_);
  or _56183_ (_05033_, _05032_, _05029_);
  or _56184_ (_05034_, _05033_, _05026_);
  or _56185_ (_05035_, _05034_, _05025_);
  and _56186_ (_05036_, _04177_, _04590_);
  and _56187_ (_05037_, _04195_, _04625_);
  or _56188_ (_05038_, _05037_, _05036_);
  and _56189_ (_05039_, _04206_, _04585_);
  and _56190_ (_05040_, _04174_, _04587_);
  or _56191_ (_05041_, _05040_, _05039_);
  or _56192_ (_05042_, _05041_, _05038_);
  and _56193_ (_05043_, _04157_, _04616_);
  and _56194_ (_05044_, _04152_, _04601_);
  or _56195_ (_05045_, _05044_, _05043_);
  and _56196_ (_05046_, _04146_, _04603_);
  and _56197_ (_05047_, _04198_, _04606_);
  or _56198_ (_05048_, _05047_, _05046_);
  or _56199_ (_05049_, _05048_, _05045_);
  or _56200_ (_05050_, _05049_, _05042_);
  or _56201_ (_05051_, _05050_, _05035_);
  or _56202_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], _05051_, _05022_);
  and _56203_ (_05052_, _04157_, _04306_);
  and _56204_ (_05053_, _04146_, _04324_);
  or _56205_ (_05054_, _05053_, _05052_);
  and _56206_ (_05055_, _04152_, _04337_);
  and _56207_ (_05056_, _04161_, _04317_);
  or _56208_ (_05057_, _05056_, _05055_);
  or _56209_ (_05058_, _05057_, _05054_);
  and _56210_ (_05059_, _04166_, _04335_);
  and _56211_ (_05060_, _04169_, _04339_);
  or _56212_ (_05061_, _05060_, _05059_);
  and _56213_ (_05062_, _04174_, _04313_);
  and _56214_ (_05063_, _04177_, _04327_);
  or _56215_ (_05064_, _05063_, _05062_);
  and _56216_ (_05065_, _04183_, _04308_);
  and _56217_ (_05066_, _04186_, _04333_);
  or _56218_ (_05067_, _05066_, _05065_);
  or _56219_ (_05068_, _05067_, _05064_);
  and _56220_ (_05069_, _04191_, _04319_);
  and _56221_ (_05070_, _04195_, _04322_);
  and _56222_ (_05071_, _04198_, _04344_);
  and _56223_ (_05072_, _04142_, _04347_);
  or _56224_ (_05073_, _05072_, _05071_);
  or _56225_ (_05074_, _05073_, _05070_);
  or _56226_ (_05075_, _05074_, _05069_);
  and _56227_ (_05076_, _04206_, _04311_);
  and _56228_ (_05077_, _04209_, _04329_);
  or _56229_ (_05078_, _05077_, _05076_);
  or _56230_ (_05079_, _05078_, _05075_);
  or _56231_ (_05080_, _05079_, _05068_);
  or _56232_ (_05082_, _05080_, _05061_);
  or _56233_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], _05082_, _05058_);
  and _56234_ (_05085_, _04157_, _04353_);
  and _56235_ (_05087_, _04146_, _04371_);
  or _56236_ (_05089_, _05087_, _05085_);
  and _56237_ (_05091_, _04152_, _04384_);
  and _56238_ (_05093_, _04161_, _04364_);
  or _56239_ (_05094_, _05093_, _05091_);
  or _56240_ (_05095_, _05094_, _05089_);
  and _56241_ (_05096_, _04166_, _04382_);
  and _56242_ (_05097_, _04169_, _04386_);
  or _56243_ (_05098_, _05097_, _05096_);
  and _56244_ (_05099_, _04183_, _04355_);
  and _56245_ (_05101_, _04186_, _04380_);
  or _56246_ (_05102_, _05101_, _05099_);
  and _56247_ (_05104_, _04174_, _04360_);
  and _56248_ (_05105_, _04209_, _04376_);
  or _56249_ (_05106_, _05105_, _05104_);
  or _56250_ (_05108_, _05106_, _05102_);
  and _56251_ (_05109_, _04191_, _04366_);
  and _56252_ (_05110_, _04142_, _04393_);
  and _56253_ (_05112_, _04195_, _04369_);
  and _56254_ (_05113_, _04198_, _04391_);
  or _56255_ (_05114_, _05113_, _05112_);
  or _56256_ (_05116_, _05114_, _05110_);
  or _56257_ (_05117_, _05116_, _05109_);
  and _56258_ (_05118_, _04177_, _04374_);
  and _56259_ (_05120_, _04206_, _04358_);
  or _56260_ (_05121_, _05120_, _05118_);
  or _56261_ (_05122_, _05121_, _05117_);
  or _56262_ (_05124_, _05122_, _05108_);
  or _56263_ (_05125_, _05124_, _05098_);
  or _56264_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], _05125_, _05095_);
  and _56265_ (_05127_, _04146_, _04420_);
  and _56266_ (_05128_, _04152_, _04428_);
  or _56267_ (_05129_, _05128_, _05127_);
  and _56268_ (_05131_, _04157_, _04406_);
  and _56269_ (_05132_, _04161_, _04412_);
  or _56270_ (_05133_, _05132_, _05131_);
  or _56271_ (_05134_, _05133_, _05129_);
  and _56272_ (_05135_, _04166_, _04430_);
  and _56273_ (_05136_, _04169_, _04432_);
  or _56274_ (_05137_, _05136_, _05135_);
  and _56275_ (_05138_, _04174_, _04404_);
  and _56276_ (_05139_, _04177_, _04415_);
  or _56277_ (_05140_, _05139_, _05138_);
  and _56278_ (_05141_, _04183_, _04401_);
  and _56279_ (_05142_, _04186_, _04426_);
  or _56280_ (_05143_, _05142_, _05141_);
  or _56281_ (_05144_, _05143_, _05140_);
  and _56282_ (_05145_, _04191_, _04410_);
  and _56283_ (_05146_, _04195_, _04437_);
  and _56284_ (_05147_, _04198_, _04439_);
  and _56285_ (_05148_, _04142_, _04417_);
  or _56286_ (_05149_, _05148_, _05147_);
  or _56287_ (_05150_, _05149_, _05146_);
  or _56288_ (_05151_, _05150_, _05145_);
  and _56289_ (_05153_, _04206_, _04399_);
  and _56290_ (_05154_, _04209_, _04422_);
  or _56291_ (_05156_, _05154_, _05153_);
  or _56292_ (_05157_, _05156_, _05151_);
  or _56293_ (_05158_, _05157_, _05144_);
  or _56294_ (_05160_, _05158_, _05137_);
  or _56295_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], _05160_, _05134_);
  and _56296_ (_05161_, _04157_, _04446_);
  and _56297_ (_05163_, _04152_, _04477_);
  or _56298_ (_05164_, _05163_, _05161_);
  and _56299_ (_05165_, _04146_, _04464_);
  and _56300_ (_05167_, _04161_, _04457_);
  or _56301_ (_05168_, _05167_, _05165_);
  or _56302_ (_05169_, _05168_, _05164_);
  and _56303_ (_05171_, _04166_, _04475_);
  and _56304_ (_05172_, _04169_, _04479_);
  or _56305_ (_05173_, _05172_, _05171_);
  and _56306_ (_05175_, _04183_, _04448_);
  and _56307_ (_05176_, _04186_, _04473_);
  or _56308_ (_05177_, _05176_, _05175_);
  and _56309_ (_05179_, _04177_, _04467_);
  and _56310_ (_05180_, _04206_, _04451_);
  or _56311_ (_05181_, _05180_, _05179_);
  or _56312_ (_05183_, _05181_, _05177_);
  and _56313_ (_05184_, _04191_, _04459_);
  and _56314_ (_05185_, _04195_, _04462_);
  and _56315_ (_05186_, _04198_, _04484_);
  and _56316_ (_05187_, _04142_, _04486_);
  or _56317_ (_05188_, _05187_, _05186_);
  or _56318_ (_05189_, _05188_, _05185_);
  or _56319_ (_05190_, _05189_, _05184_);
  and _56320_ (_05191_, _04174_, _04453_);
  and _56321_ (_05192_, _04209_, _04469_);
  or _56322_ (_05193_, _05192_, _05191_);
  or _56323_ (_05194_, _05193_, _05190_);
  or _56324_ (_05195_, _05194_, _05183_);
  or _56325_ (_05196_, _05195_, _05173_);
  or _56326_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], _05196_, _05169_);
  and _56327_ (_05197_, _04146_, _04510_);
  and _56328_ (_05198_, _04152_, _04523_);
  or _56329_ (_05199_, _05198_, _05197_);
  and _56330_ (_05200_, _04157_, _04492_);
  and _56331_ (_05201_, _04161_, _04503_);
  or _56332_ (_05202_, _05201_, _05200_);
  or _56333_ (_05204_, _05202_, _05199_);
  and _56334_ (_05205_, _04166_, _04521_);
  and _56335_ (_05207_, _04169_, _04525_);
  or _56336_ (_05208_, _05207_, _05205_);
  and _56337_ (_05209_, _04174_, _04499_);
  and _56338_ (_05211_, _04177_, _04513_);
  or _56339_ (_05212_, _05211_, _05209_);
  and _56340_ (_05213_, _04183_, _04494_);
  and _56341_ (_05215_, _04186_, _04519_);
  or _56342_ (_05216_, _05215_, _05213_);
  or _56343_ (_05217_, _05216_, _05212_);
  and _56344_ (_05219_, _04191_, _04505_);
  and _56345_ (_05220_, _04195_, _04508_);
  and _56346_ (_05221_, _04198_, _04530_);
  and _56347_ (_05223_, _04142_, _04532_);
  or _56348_ (_05224_, _05223_, _05221_);
  or _56349_ (_05225_, _05224_, _05220_);
  or _56350_ (_05227_, _05225_, _05219_);
  and _56351_ (_05228_, _04206_, _04497_);
  and _56352_ (_05229_, _04209_, _04515_);
  or _56353_ (_05231_, _05229_, _05228_);
  or _56354_ (_05232_, _05231_, _05227_);
  or _56355_ (_05233_, _05232_, _05217_);
  or _56356_ (_05235_, _05233_, _05208_);
  or _56357_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], _05235_, _05204_);
  and _56358_ (_05236_, _04152_, _04570_);
  and _56359_ (_05237_, _04161_, _04552_);
  or _56360_ (_05238_, _05237_, _05236_);
  and _56361_ (_05239_, _04157_, _04540_);
  and _56362_ (_05240_, _04146_, _04555_);
  or _56363_ (_05241_, _05240_, _05239_);
  or _56364_ (_05242_, _05241_, _05238_);
  and _56365_ (_05243_, _04166_, _04572_);
  and _56366_ (_05244_, _04169_, _04568_);
  or _56367_ (_05245_, _05244_, _05243_);
  and _56368_ (_05246_, _04174_, _04538_);
  and _56369_ (_05247_, _04206_, _04544_);
  or _56370_ (_05248_, _05247_, _05246_);
  and _56371_ (_05249_, _04209_, _04560_);
  and _56372_ (_05250_, _04183_, _04546_);
  or _56373_ (_05251_, _05250_, _05249_);
  or _56374_ (_05252_, _05251_, _05248_);
  and _56375_ (_05253_, _04191_, _04550_);
  and _56376_ (_05254_, _04198_, _04557_);
  and _56377_ (_05256_, _04195_, _04577_);
  and _56378_ (_05257_, _04142_, _04562_);
  or _56379_ (_05259_, _05257_, _05256_);
  or _56380_ (_05260_, _05259_, _05254_);
  or _56381_ (_05261_, _05260_, _05253_);
  and _56382_ (_05263_, _04177_, _04579_);
  and _56383_ (_05264_, _04186_, _04566_);
  or _56384_ (_05265_, _05264_, _05263_);
  or _56385_ (_05267_, _05265_, _05261_);
  or _56386_ (_05268_, _05267_, _05252_);
  or _56387_ (_05269_, _05268_, _05245_);
  or _56388_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], _05269_, _05242_);
  and _56389_ (_05271_, _04157_, _04585_);
  and _56390_ (_05272_, _04152_, _04616_);
  or _56391_ (_05274_, _05272_, _05271_);
  and _56392_ (_05275_, _04146_, _04601_);
  and _56393_ (_05276_, _04161_, _04598_);
  or _56394_ (_05278_, _05276_, _05275_);
  or _56395_ (_05279_, _05278_, _05274_);
  and _56396_ (_05280_, _04166_, _04618_);
  and _56397_ (_05282_, _04169_, _04614_);
  or _56398_ (_05283_, _05282_, _05280_);
  and _56399_ (_05284_, _04183_, _04592_);
  and _56400_ (_05286_, _04186_, _04612_);
  or _56401_ (_05287_, _05286_, _05284_);
  and _56402_ (_05288_, _04177_, _04625_);
  and _56403_ (_05289_, _04206_, _04587_);
  or _56404_ (_05290_, _05289_, _05288_);
  or _56405_ (_05291_, _05290_, _05287_);
  and _56406_ (_05292_, _04191_, _04596_);
  and _56407_ (_05293_, _04195_, _04623_);
  and _56408_ (_05294_, _04198_, _04603_);
  and _56409_ (_05295_, _04142_, _04608_);
  or _56410_ (_05296_, _05295_, _05294_);
  or _56411_ (_05297_, _05296_, _05293_);
  or _56412_ (_05298_, _05297_, _05292_);
  and _56413_ (_05299_, _04174_, _04590_);
  and _56414_ (_05300_, _04209_, _04606_);
  or _56415_ (_05301_, _05300_, _05299_);
  or _56416_ (_05302_, _05301_, _05298_);
  or _56417_ (_05303_, _05302_, _05291_);
  or _56418_ (_05304_, _05303_, _05283_);
  or _56419_ (\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], _05304_, _05279_);
  nand _56420_ (_05305_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  not _56421_ (_05307_, \oc8051_golden_model_1.PC [3]);
  or _56422_ (_05308_, \oc8051_golden_model_1.PC [2], _05307_);
  or _56423_ (_05310_, _05308_, _05305_);
  or _56424_ (_05311_, _05310_, _00434_);
  not _56425_ (_05312_, \oc8051_golden_model_1.PC [1]);
  or _56426_ (_05314_, _05312_, \oc8051_golden_model_1.PC [0]);
  or _56427_ (_05315_, _05314_, _05308_);
  or _56428_ (_05316_, _05315_, _00393_);
  and _56429_ (_05318_, _05316_, _05311_);
  not _56430_ (_05319_, \oc8051_golden_model_1.PC [2]);
  or _56431_ (_05320_, _05319_, \oc8051_golden_model_1.PC [3]);
  or _56432_ (_05322_, _05320_, _05305_);
  or _56433_ (_05323_, _05322_, _00270_);
  or _56434_ (_05324_, _05320_, _05314_);
  or _56435_ (_05326_, _05324_, _00229_);
  and _56436_ (_05327_, _05326_, _05323_);
  and _56437_ (_05328_, _05327_, _05318_);
  nand _56438_ (_05330_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _56439_ (_05331_, _05330_, _05305_);
  or _56440_ (_05332_, _05331_, _00617_);
  or _56441_ (_05334_, _05330_, _05314_);
  or _56442_ (_05335_, _05334_, _00566_);
  and _56443_ (_05336_, _05335_, _05332_);
  or _56444_ (_05338_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [3]);
  or _56445_ (_05339_, _05338_, _05305_);
  or _56446_ (_05340_, _05339_, _00075_);
  or _56447_ (_05341_, _05338_, _05314_);
  or _56448_ (_05342_, _05341_, _00034_);
  and _56449_ (_05343_, _05342_, _05340_);
  and _56450_ (_05344_, _05343_, _05336_);
  and _56451_ (_05345_, _05344_, _05328_);
  not _56452_ (_05346_, \oc8051_golden_model_1.PC [0]);
  or _56453_ (_05347_, \oc8051_golden_model_1.PC [1], _05346_);
  or _56454_ (_05348_, _05347_, _05330_);
  or _56455_ (_05349_, _05348_, _00516_);
  or _56456_ (_05350_, \oc8051_golden_model_1.PC [1], \oc8051_golden_model_1.PC [0]);
  or _56457_ (_05351_, _05350_, _05330_);
  or _56458_ (_05352_, _05351_, _00475_);
  and _56459_ (_05353_, _05352_, _05349_);
  or _56460_ (_05354_, _05338_, _05350_);
  or _56461_ (_05355_, _05354_, _43762_);
  or _56462_ (_05356_, _05338_, _05347_);
  or _56463_ (_05357_, _05356_, _43803_);
  and _56464_ (_05358_, _05357_, _05355_);
  and _56465_ (_05360_, _05358_, _05353_);
  or _56466_ (_05361_, _05347_, _05308_);
  or _56467_ (_05363_, _05361_, _00352_);
  or _56468_ (_05364_, _05350_, _05308_);
  or _56469_ (_05365_, _05364_, _00311_);
  and _56470_ (_05367_, _05365_, _05363_);
  or _56471_ (_05368_, _05347_, _05320_);
  or _56472_ (_05369_, _05368_, _00188_);
  or _56473_ (_05371_, _05350_, _05320_);
  or _56474_ (_05372_, _05371_, _00116_);
  and _56475_ (_05373_, _05372_, _05369_);
  and _56476_ (_05375_, _05373_, _05367_);
  and _56477_ (_05376_, _05375_, _05360_);
  and _56478_ (_05377_, _05376_, _05345_);
  or _56479_ (_05379_, _05310_, _00399_);
  or _56480_ (_05380_, _05315_, _00358_);
  and _56481_ (_05381_, _05380_, _05379_);
  or _56482_ (_05383_, _05322_, _00235_);
  or _56483_ (_05384_, _05324_, _00194_);
  and _56484_ (_05385_, _05384_, _05383_);
  and _56485_ (_05387_, _05385_, _05381_);
  or _56486_ (_05388_, _05331_, _00576_);
  or _56487_ (_05389_, _05334_, _00522_);
  and _56488_ (_05391_, _05389_, _05388_);
  or _56489_ (_05392_, _05339_, _00040_);
  or _56490_ (_05393_, _05341_, _43809_);
  and _56491_ (_05394_, _05393_, _05392_);
  and _56492_ (_05395_, _05394_, _05391_);
  and _56493_ (_05396_, _05395_, _05387_);
  or _56494_ (_05397_, _05348_, _00481_);
  or _56495_ (_05398_, _05351_, _00440_);
  and _56496_ (_05399_, _05398_, _05397_);
  or _56497_ (_05400_, _05354_, _43727_);
  or _56498_ (_05401_, _05356_, _43768_);
  and _56499_ (_05402_, _05401_, _05400_);
  and _56500_ (_05403_, _05402_, _05399_);
  or _56501_ (_05404_, _05361_, _00317_);
  or _56502_ (_05405_, _05364_, _00276_);
  and _56503_ (_05406_, _05405_, _05404_);
  or _56504_ (_05407_, _05368_, _00122_);
  or _56505_ (_05408_, _05371_, _00081_);
  and _56506_ (_05409_, _05408_, _05407_);
  and _56507_ (_05410_, _05409_, _05406_);
  and _56508_ (_05411_, _05410_, _05403_);
  and _56509_ (_05413_, _05411_, _05396_);
  and _56510_ (_05414_, _05413_, _05377_);
  or _56511_ (_05416_, _05310_, _00424_);
  or _56512_ (_05417_, _05315_, _00383_);
  and _56513_ (_05418_, _05417_, _05416_);
  or _56514_ (_05420_, _05322_, _00260_);
  or _56515_ (_05421_, _05324_, _00219_);
  and _56516_ (_05422_, _05421_, _05420_);
  and _56517_ (_05424_, _05422_, _05418_);
  or _56518_ (_05425_, _05331_, _00607_);
  or _56519_ (_05426_, _05334_, _00550_);
  and _56520_ (_05428_, _05426_, _05425_);
  or _56521_ (_05429_, _05339_, _00065_);
  or _56522_ (_05430_, _05341_, _00024_);
  and _56523_ (_05432_, _05430_, _05429_);
  and _56524_ (_05433_, _05432_, _05428_);
  and _56525_ (_05434_, _05433_, _05424_);
  or _56526_ (_05436_, _05348_, _00506_);
  or _56527_ (_05437_, _05351_, _00465_);
  and _56528_ (_05438_, _05437_, _05436_);
  or _56529_ (_05440_, _05354_, _43752_);
  or _56530_ (_05441_, _05356_, _43793_);
  and _56531_ (_05442_, _05441_, _05440_);
  and _56532_ (_05444_, _05442_, _05438_);
  or _56533_ (_05445_, _05361_, _00342_);
  or _56534_ (_05446_, _05364_, _00301_);
  and _56535_ (_05447_, _05446_, _05445_);
  or _56536_ (_05448_, _05368_, _00168_);
  or _56537_ (_05449_, _05371_, _00106_);
  and _56538_ (_05450_, _05449_, _05448_);
  and _56539_ (_05451_, _05450_, _05447_);
  and _56540_ (_05452_, _05451_, _05444_);
  nand _56541_ (_05453_, _05452_, _05434_);
  or _56542_ (_05454_, _05310_, _00429_);
  or _56543_ (_05455_, _05315_, _00388_);
  and _56544_ (_05456_, _05455_, _05454_);
  or _56545_ (_05457_, _05322_, _00265_);
  or _56546_ (_05458_, _05324_, _00224_);
  and _56547_ (_05459_, _05458_, _05457_);
  and _56548_ (_05460_, _05459_, _05456_);
  or _56549_ (_05461_, _05331_, _00612_);
  or _56550_ (_05462_, _05334_, _00558_);
  and _56551_ (_05463_, _05462_, _05461_);
  or _56552_ (_05464_, _05339_, _00070_);
  or _56553_ (_05466_, _05341_, _00029_);
  and _56554_ (_05467_, _05466_, _05464_);
  and _56555_ (_05469_, _05467_, _05463_);
  and _56556_ (_05470_, _05469_, _05460_);
  or _56557_ (_05471_, _05348_, _00511_);
  or _56558_ (_05473_, _05351_, _00470_);
  and _56559_ (_05474_, _05473_, _05471_);
  or _56560_ (_05475_, _05354_, _43757_);
  or _56561_ (_05477_, _05356_, _43798_);
  and _56562_ (_05478_, _05477_, _05475_);
  and _56563_ (_05479_, _05478_, _05474_);
  or _56564_ (_05481_, _05361_, _00347_);
  or _56565_ (_05482_, _05364_, _00306_);
  and _56566_ (_05483_, _05482_, _05481_);
  or _56567_ (_05485_, _05368_, _00179_);
  or _56568_ (_05486_, _05371_, _00111_);
  and _56569_ (_05487_, _05486_, _05485_);
  and _56570_ (_05489_, _05487_, _05483_);
  and _56571_ (_05490_, _05489_, _05479_);
  and _56572_ (_05491_, _05490_, _05470_);
  nand _56573_ (_05493_, _05491_, _05453_);
  not _56574_ (_05494_, _05493_);
  and _56575_ (_05495_, _05494_, _05414_);
  or _56576_ (_05497_, _05310_, _00414_);
  or _56577_ (_05498_, _05315_, _00373_);
  and _56578_ (_05499_, _05498_, _05497_);
  or _56579_ (_05500_, _05322_, _00250_);
  or _56580_ (_05501_, _05324_, _00209_);
  and _56581_ (_05502_, _05501_, _05500_);
  and _56582_ (_05503_, _05502_, _05499_);
  or _56583_ (_05504_, _05331_, _00597_);
  or _56584_ (_05505_, _05334_, _00537_);
  and _56585_ (_05506_, _05505_, _05504_);
  or _56586_ (_05507_, _05339_, _00055_);
  or _56587_ (_05508_, _05341_, _00014_);
  and _56588_ (_05509_, _05508_, _05507_);
  and _56589_ (_05510_, _05509_, _05506_);
  and _56590_ (_05511_, _05510_, _05503_);
  or _56591_ (_05512_, _05348_, _00496_);
  or _56592_ (_05513_, _05351_, _00455_);
  and _56593_ (_05514_, _05513_, _05512_);
  or _56594_ (_05515_, _05354_, _43742_);
  or _56595_ (_05516_, _05356_, _43783_);
  and _56596_ (_05517_, _05516_, _05515_);
  and _56597_ (_05519_, _05517_, _05514_);
  or _56598_ (_05520_, _05361_, _00332_);
  or _56599_ (_05522_, _05364_, _00291_);
  and _56600_ (_05523_, _05522_, _05520_);
  or _56601_ (_05524_, _05368_, _00146_);
  or _56602_ (_05526_, _05371_, _00096_);
  and _56603_ (_05527_, _05526_, _05524_);
  and _56604_ (_05528_, _05527_, _05523_);
  and _56605_ (_05530_, _05528_, _05519_);
  nand _56606_ (_05531_, _05530_, _05511_);
  or _56607_ (_05532_, _05310_, _00419_);
  or _56608_ (_05534_, _05315_, _00378_);
  and _56609_ (_05535_, _05534_, _05532_);
  or _56610_ (_05536_, _05322_, _00255_);
  or _56611_ (_05538_, _05324_, _00214_);
  and _56612_ (_05539_, _05538_, _05536_);
  and _56613_ (_05540_, _05539_, _05535_);
  or _56614_ (_05542_, _05331_, _00602_);
  or _56615_ (_05543_, _05334_, _00542_);
  and _56616_ (_05544_, _05543_, _05542_);
  or _56617_ (_05546_, _05339_, _00060_);
  or _56618_ (_05547_, _05341_, _00019_);
  and _56619_ (_05548_, _05547_, _05546_);
  and _56620_ (_05550_, _05548_, _05544_);
  and _56621_ (_05551_, _05550_, _05540_);
  or _56622_ (_05552_, _05348_, _00501_);
  or _56623_ (_05553_, _05351_, _00460_);
  and _56624_ (_05554_, _05553_, _05552_);
  or _56625_ (_05555_, _05354_, _43747_);
  or _56626_ (_05556_, _05356_, _43788_);
  and _56627_ (_05557_, _05556_, _05555_);
  and _56628_ (_05558_, _05557_, _05554_);
  or _56629_ (_05559_, _05361_, _00337_);
  or _56630_ (_05560_, _05364_, _00296_);
  and _56631_ (_05561_, _05560_, _05559_);
  or _56632_ (_05562_, _05368_, _00157_);
  or _56633_ (_05563_, _05371_, _00101_);
  and _56634_ (_05564_, _05563_, _05562_);
  and _56635_ (_05565_, _05564_, _05561_);
  and _56636_ (_05566_, _05565_, _05558_);
  nand _56637_ (_05567_, _05566_, _05551_);
  or _56638_ (_05568_, _05567_, _05531_);
  not _56639_ (_05569_, _05568_);
  or _56640_ (_05570_, _05310_, _00409_);
  or _56641_ (_05572_, _05315_, _00368_);
  and _56642_ (_05573_, _05572_, _05570_);
  or _56643_ (_05575_, _05322_, _00245_);
  or _56644_ (_05576_, _05324_, _00204_);
  and _56645_ (_05577_, _05576_, _05575_);
  and _56646_ (_05579_, _05577_, _05573_);
  or _56647_ (_05580_, _05331_, _00592_);
  or _56648_ (_05581_, _05334_, _00532_);
  and _56649_ (_05583_, _05581_, _05580_);
  or _56650_ (_05584_, _05339_, _00050_);
  or _56651_ (_05585_, _05341_, _00009_);
  and _56652_ (_05587_, _05585_, _05584_);
  and _56653_ (_05588_, _05587_, _05583_);
  and _56654_ (_05589_, _05588_, _05579_);
  or _56655_ (_05591_, _05348_, _00491_);
  or _56656_ (_05592_, _05351_, _00450_);
  and _56657_ (_05593_, _05592_, _05591_);
  or _56658_ (_05595_, _05354_, _43737_);
  or _56659_ (_05596_, _05356_, _43778_);
  and _56660_ (_05597_, _05596_, _05595_);
  and _56661_ (_05599_, _05597_, _05593_);
  or _56662_ (_05600_, _05361_, _00327_);
  or _56663_ (_05601_, _05364_, _00286_);
  and _56664_ (_05603_, _05601_, _05600_);
  or _56665_ (_05604_, _05368_, _00135_);
  or _56666_ (_05605_, _05371_, _00091_);
  and _56667_ (_05606_, _05605_, _05604_);
  and _56668_ (_05607_, _05606_, _05603_);
  and _56669_ (_05608_, _05607_, _05599_);
  nand _56670_ (_05609_, _05608_, _05589_);
  not _56671_ (_05610_, _05609_);
  or _56672_ (_05611_, _05310_, _00404_);
  or _56673_ (_05612_, _05315_, _00363_);
  and _56674_ (_05613_, _05612_, _05611_);
  or _56675_ (_05614_, _05322_, _00240_);
  or _56676_ (_05615_, _05324_, _00199_);
  and _56677_ (_05616_, _05615_, _05614_);
  and _56678_ (_05617_, _05616_, _05613_);
  or _56679_ (_05618_, _05331_, _00584_);
  or _56680_ (_05619_, _05334_, _00527_);
  and _56681_ (_05620_, _05619_, _05618_);
  or _56682_ (_05621_, _05339_, _00045_);
  or _56683_ (_05622_, _05341_, _00004_);
  and _56684_ (_05623_, _05622_, _05621_);
  and _56685_ (_05625_, _05623_, _05620_);
  and _56686_ (_05626_, _05625_, _05617_);
  or _56687_ (_05628_, _05348_, _00486_);
  or _56688_ (_05629_, _05351_, _00445_);
  and _56689_ (_05630_, _05629_, _05628_);
  or _56690_ (_05632_, _05354_, _43732_);
  or _56691_ (_05633_, _05356_, _43773_);
  and _56692_ (_05634_, _05633_, _05632_);
  and _56693_ (_05636_, _05634_, _05630_);
  or _56694_ (_05637_, _05361_, _00322_);
  or _56695_ (_05638_, _05364_, _00281_);
  and _56696_ (_05640_, _05638_, _05637_);
  or _56697_ (_05641_, _05368_, _00127_);
  or _56698_ (_05642_, _05371_, _00086_);
  and _56699_ (_05644_, _05642_, _05641_);
  and _56700_ (_05645_, _05644_, _05640_);
  and _56701_ (_05646_, _05645_, _05636_);
  and _56702_ (_05648_, _05646_, _05626_);
  and _56703_ (_05649_, _05648_, _05610_);
  and _56704_ (_05650_, _05649_, _05569_);
  and _56705_ (_05652_, _05650_, _05495_);
  not _56706_ (_05653_, _05652_);
  and _56707_ (_05654_, _05452_, _05434_);
  nand _56708_ (_05656_, _05491_, _05654_);
  nand _56709_ (_05657_, _05376_, _05345_);
  or _56710_ (_05658_, _05413_, _05657_);
  nor _56711_ (_05659_, _05658_, _05656_);
  not _56712_ (_05660_, _05659_);
  or _56713_ (_05661_, _05648_, _05610_);
  or _56714_ (_05662_, _05661_, _05568_);
  nor _56715_ (_05663_, _05662_, _05660_);
  not _56716_ (_05664_, _05663_);
  or _56717_ (_05665_, _05648_, _05609_);
  not _56718_ (_05666_, _05531_);
  or _56719_ (_05667_, _05567_, _05666_);
  or _56720_ (_05668_, _05667_, _05665_);
  or _56721_ (_05669_, _05668_, _05660_);
  or _56722_ (_05670_, _05665_, _05568_);
  nor _56723_ (_05671_, _05658_, _05493_);
  not _56724_ (_05672_, _05671_);
  or _56725_ (_05673_, _05672_, _05670_);
  and _56726_ (_05674_, _05673_, _05669_);
  or _56727_ (_05675_, _05672_, _05662_);
  not _56728_ (_05676_, _05675_);
  and _56729_ (_05678_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _56730_ (_05679_, \oc8051_golden_model_1.DPL [0], \oc8051_golden_model_1.ACC [0]);
  nor _56731_ (_05681_, _05679_, _05678_);
  nand _56732_ (_05682_, _05681_, _05676_);
  or _56733_ (_05683_, _05491_, _05654_);
  or _56734_ (_05685_, _05683_, _05658_);
  or _56735_ (_05686_, _05685_, _05670_);
  or _56736_ (_05687_, _05413_, _05377_);
  or _56737_ (_05689_, _05687_, _05493_);
  or _56738_ (_05690_, _05689_, _05670_);
  and _56739_ (_05691_, _05690_, _05686_);
  or _56740_ (_05693_, _05687_, _05656_);
  or _56741_ (_05694_, _05693_, _05670_);
  or _56742_ (_05695_, _05491_, _05453_);
  or _56743_ (_05697_, _05695_, _05687_);
  or _56744_ (_05698_, _05697_, _05670_);
  and _56745_ (_05699_, _05698_, _05694_);
  or _56746_ (_05701_, _05695_, _05658_);
  or _56747_ (_05702_, _05701_, _05670_);
  or _56748_ (_05703_, _05687_, _05683_);
  or _56749_ (_05705_, _05703_, _05670_);
  and _56750_ (_05706_, _05705_, _05702_);
  and _56751_ (_05707_, _05706_, _05699_);
  and _56752_ (_05709_, _05707_, _05691_);
  and _56753_ (_05710_, _05675_, _05346_);
  nand _56754_ (_05711_, _05710_, _05709_);
  nand _56755_ (_05712_, _05711_, _05682_);
  nand _56756_ (_05713_, _05712_, _05674_);
  and _56757_ (_05714_, _05709_, _05674_);
  or _56758_ (_05715_, _05714_, _05346_);
  nand _56759_ (_05716_, _05715_, _05713_);
  nand _56760_ (_05717_, _05716_, _05664_);
  not _56761_ (_05718_, _05670_);
  and _56762_ (_05719_, _05718_, _05659_);
  not _56763_ (_05720_, _05719_);
  not _56764_ (_05721_, _05683_);
  and _56765_ (_05722_, _05413_, _05657_);
  and _56766_ (_05723_, _05722_, _05721_);
  and _56767_ (_05724_, _05723_, _05718_);
  not _56768_ (_05725_, _05695_);
  and _56769_ (_05726_, _05722_, _05725_);
  and _56770_ (_05727_, _05726_, _05718_);
  nor _56771_ (_05728_, _05727_, _05724_);
  and _56772_ (_05729_, _05728_, _05720_);
  and _56773_ (_05731_, _05721_, _05414_);
  and _56774_ (_05732_, _05731_, _05718_);
  not _56775_ (_05734_, _05732_);
  and _56776_ (_05735_, _05722_, _05494_);
  and _56777_ (_05736_, _05735_, _05718_);
  not _56778_ (_05738_, _05656_);
  and _56779_ (_05739_, _05722_, _05738_);
  and _56780_ (_05740_, _05739_, _05718_);
  nor _56781_ (_05742_, _05740_, _05736_);
  and _56782_ (_05743_, _05742_, _05734_);
  and _56783_ (_05744_, _05743_, _05729_);
  and _56784_ (_05746_, _05725_, _05414_);
  and _56785_ (_05747_, _05746_, _05718_);
  not _56786_ (_05748_, _05747_);
  and _56787_ (_05750_, _05738_, _05414_);
  and _56788_ (_05751_, _05750_, _05718_);
  and _56789_ (_05752_, _05718_, _05495_);
  nor _56790_ (_05754_, _05752_, _05751_);
  and _56791_ (_05755_, _05754_, _05748_);
  and _56792_ (_05756_, _05755_, _05744_);
  not _56793_ (_05758_, \oc8051_golden_model_1.ACC [0]);
  and _56794_ (_05759_, _05758_, \oc8051_golden_model_1.PC [0]);
  and _56795_ (_05760_, \oc8051_golden_model_1.ACC [0], _05346_);
  or _56796_ (_05762_, _05760_, _05664_);
  or _56797_ (_05763_, _05762_, _05759_);
  and _56798_ (_05764_, _05763_, _05756_);
  nand _56799_ (_05765_, _05764_, _05717_);
  or _56800_ (_05766_, _05756_, \oc8051_golden_model_1.PC [0]);
  and _56801_ (_05767_, _05766_, _05765_);
  and _56802_ (_05768_, _05756_, _05714_);
  or _56803_ (_05769_, _05768_, _05312_);
  and _56804_ (_05770_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor _56805_ (_05771_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.ACC [1]);
  nor _56806_ (_05772_, _05771_, _05770_);
  and _56807_ (_05773_, _05772_, _05678_);
  nor _56808_ (_05774_, _05772_, _05678_);
  nor _56809_ (_05775_, _05774_, _05773_);
  or _56810_ (_05776_, _05775_, _05675_);
  and _56811_ (_05777_, _05347_, _05314_);
  and _56812_ (_05778_, _05777_, _05675_);
  nand _56813_ (_05779_, _05778_, _05709_);
  nand _56814_ (_05780_, _05779_, _05776_);
  and _56815_ (_05781_, _05674_, _05664_);
  and _56816_ (_05782_, _05781_, _05780_);
  not _56817_ (_05784_, \oc8051_golden_model_1.ACC [1]);
  nor _56818_ (_05785_, _05777_, _05784_);
  and _56819_ (_05787_, _05777_, _05784_);
  nor _56820_ (_05788_, _05787_, _05785_);
  and _56821_ (_05789_, _05788_, _05760_);
  nor _56822_ (_05791_, _05788_, _05760_);
  nor _56823_ (_05792_, _05791_, _05789_);
  nor _56824_ (_05793_, _05792_, _05664_);
  or _56825_ (_05795_, _05793_, _05782_);
  nand _56826_ (_05796_, _05795_, _05756_);
  nand _56827_ (_05797_, _05796_, _05769_);
  or _56828_ (_05799_, _05797_, _05767_);
  and _56829_ (_05800_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _56830_ (_05801_, \oc8051_golden_model_1.PC [2], \oc8051_golden_model_1.PC [1]);
  nor _56831_ (_05803_, _05801_, _05800_);
  not _56832_ (_05804_, _05803_);
  nor _56833_ (_05805_, _05804_, _05755_);
  not _56834_ (_05807_, _05805_);
  nor _56835_ (_05808_, _05773_, _05770_);
  and _56836_ (_05809_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor _56837_ (_05811_, \oc8051_golden_model_1.DPL [2], \oc8051_golden_model_1.ACC [2]);
  nor _56838_ (_05812_, _05811_, _05809_);
  not _56839_ (_05813_, _05812_);
  nor _56840_ (_05815_, _05813_, _05808_);
  and _56841_ (_05816_, _05813_, _05808_);
  nor _56842_ (_05817_, _05816_, _05815_);
  not _56843_ (_05818_, _05817_);
  or _56844_ (_05819_, _05818_, _05675_);
  and _56845_ (_05820_, _05819_, _05674_);
  nor _56846_ (_05821_, _05305_, _05319_);
  and _56847_ (_05822_, _05305_, _05319_);
  nor _56848_ (_05823_, _05822_, _05821_);
  not _56849_ (_05824_, _05823_);
  nand _56850_ (_05825_, _05824_, _05709_);
  nand _56851_ (_05826_, _05825_, _05675_);
  nand _56852_ (_05827_, _05826_, _05820_);
  or _56853_ (_05828_, _05803_, _05714_);
  and _56854_ (_05829_, _05828_, _05664_);
  nand _56855_ (_05830_, _05829_, _05827_);
  nor _56856_ (_05831_, _05789_, _05785_);
  and _56857_ (_05832_, _05823_, \oc8051_golden_model_1.ACC [2]);
  nor _56858_ (_05833_, _05823_, \oc8051_golden_model_1.ACC [2]);
  nor _56859_ (_05834_, _05833_, _05832_);
  not _56860_ (_05835_, _05834_);
  and _56861_ (_05837_, _05835_, _05831_);
  nor _56862_ (_05838_, _05835_, _05831_);
  nor _56863_ (_05840_, _05838_, _05837_);
  and _56864_ (_05841_, _05840_, _05663_);
  not _56865_ (_05842_, _05841_);
  and _56866_ (_05844_, _05842_, _05744_);
  nand _56867_ (_05845_, _05844_, _05830_);
  or _56868_ (_05846_, _05803_, _05756_);
  nand _56869_ (_05848_, _05846_, _05845_);
  and _56870_ (_05849_, _05848_, _05807_);
  nor _56871_ (_05850_, _05330_, _05312_);
  nor _56872_ (_05852_, _05800_, \oc8051_golden_model_1.PC [3]);
  nor _56873_ (_05853_, _05852_, _05850_);
  or _56874_ (_05854_, _05853_, _05768_);
  nor _56875_ (_05856_, _05815_, _05809_);
  and _56876_ (_05857_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _56877_ (_05858_, \oc8051_golden_model_1.DPL [3], \oc8051_golden_model_1.ACC [3]);
  nor _56878_ (_05860_, _05858_, _05857_);
  not _56879_ (_05861_, _05860_);
  nor _56880_ (_05862_, _05861_, _05856_);
  and _56881_ (_05864_, _05861_, _05856_);
  nor _56882_ (_05865_, _05864_, _05862_);
  or _56883_ (_05866_, _05865_, _05675_);
  not _56884_ (_05868_, _05322_);
  nor _56885_ (_05869_, _05821_, _05307_);
  nor _56886_ (_05870_, _05869_, _05868_);
  and _56887_ (_05871_, _05675_, _05870_);
  nand _56888_ (_05872_, _05871_, _05709_);
  nand _56889_ (_05873_, _05872_, _05866_);
  and _56890_ (_05874_, _05873_, _05781_);
  nor _56891_ (_05875_, _05838_, _05832_);
  nor _56892_ (_05876_, _05870_, \oc8051_golden_model_1.ACC [3]);
  and _56893_ (_05877_, _05870_, \oc8051_golden_model_1.ACC [3]);
  nor _56894_ (_05878_, _05877_, _05876_);
  and _56895_ (_05879_, _05878_, _05875_);
  nor _56896_ (_05880_, _05878_, _05875_);
  nor _56897_ (_05881_, _05880_, _05879_);
  nor _56898_ (_05882_, _05881_, _05664_);
  or _56899_ (_05883_, _05882_, _05874_);
  nand _56900_ (_05884_, _05883_, _05756_);
  and _56901_ (_05885_, _05884_, _05854_);
  or _56902_ (_05886_, _05885_, _05849_);
  or _56903_ (_05887_, _05886_, _05799_);
  or _56904_ (_05888_, _05887_, _00194_);
  nand _56905_ (_05890_, _05766_, _05765_);
  and _56906_ (_05891_, _05796_, _05769_);
  or _56907_ (_05893_, _05891_, _05890_);
  or _56908_ (_05894_, _05893_, _05886_);
  or _56909_ (_05895_, _05894_, _00122_);
  and _56910_ (_05897_, _05895_, _05888_);
  nand _56911_ (_05898_, _05884_, _05854_);
  or _56912_ (_05899_, _05898_, _05849_);
  or _56913_ (_05901_, _05797_, _05890_);
  or _56914_ (_05902_, _05901_, _05899_);
  or _56915_ (_05903_, _05902_, _00576_);
  nand _56916_ (_05905_, _05848_, _05807_);
  or _56917_ (_05906_, _05898_, _05905_);
  or _56918_ (_05907_, _05906_, _05901_);
  or _56919_ (_05909_, _05907_, _00399_);
  and _56920_ (_05910_, _05909_, _05903_);
  and _56921_ (_05911_, _05910_, _05897_);
  or _56922_ (_05913_, _05906_, _05799_);
  or _56923_ (_05914_, _05913_, _00358_);
  or _56924_ (_05915_, _05906_, _05893_);
  or _56925_ (_05917_, _05915_, _00317_);
  and _56926_ (_05918_, _05917_, _05914_);
  or _56927_ (_05919_, _05899_, _05893_);
  or _56928_ (_05921_, _05919_, _00481_);
  or _56929_ (_05922_, _05891_, _05767_);
  or _56930_ (_05923_, _05922_, _05899_);
  or _56931_ (_05924_, _05923_, _00440_);
  and _56932_ (_05925_, _05924_, _05921_);
  and _56933_ (_05926_, _05925_, _05918_);
  and _56934_ (_05927_, _05926_, _05911_);
  or _56935_ (_05928_, _05885_, _05905_);
  or _56936_ (_05929_, _05928_, _05922_);
  or _56937_ (_05930_, _05929_, _43727_);
  or _56938_ (_05931_, _05928_, _05799_);
  or _56939_ (_05932_, _05931_, _43809_);
  and _56940_ (_05933_, _05932_, _05930_);
  or _56941_ (_05934_, _05901_, _05886_);
  or _56942_ (_05935_, _05934_, _00235_);
  or _56943_ (_05936_, _05922_, _05886_);
  or _56944_ (_05937_, _05936_, _00081_);
  and _56945_ (_05938_, _05937_, _05935_);
  and _56946_ (_05939_, _05938_, _05933_);
  or _56947_ (_05940_, _05899_, _05799_);
  or _56948_ (_05941_, _05940_, _00522_);
  or _56949_ (_05942_, _05906_, _05922_);
  or _56950_ (_05943_, _05942_, _00276_);
  and _56951_ (_05944_, _05943_, _05941_);
  or _56952_ (_05945_, _05928_, _05901_);
  or _56953_ (_05946_, _05945_, _00040_);
  or _56954_ (_05947_, _05928_, _05893_);
  or _56955_ (_05948_, _05947_, _43768_);
  and _56956_ (_05949_, _05948_, _05946_);
  and _56957_ (_05950_, _05949_, _05944_);
  and _56958_ (_05951_, _05950_, _05939_);
  nand _56959_ (_05952_, _05951_, _05927_);
  or _56960_ (_05953_, _05907_, _00419_);
  or _56961_ (_05954_, _05929_, _43747_);
  and _56962_ (_05955_, _05954_, _05953_);
  or _56963_ (_05956_, _05919_, _00501_);
  or _56964_ (_05957_, _05887_, _00214_);
  and _56965_ (_05958_, _05957_, _05956_);
  and _56966_ (_05959_, _05958_, _05955_);
  or _56967_ (_05960_, _05913_, _00378_);
  or _56968_ (_05961_, _05915_, _00337_);
  and _56969_ (_05962_, _05961_, _05960_);
  or _56970_ (_05963_, _05940_, _00542_);
  or _56971_ (_05964_, _05945_, _00060_);
  and _56972_ (_05965_, _05964_, _05963_);
  and _56973_ (_05966_, _05965_, _05962_);
  and _56974_ (_05967_, _05966_, _05959_);
  or _56975_ (_05968_, _05936_, _00101_);
  or _56976_ (_05969_, _05947_, _43788_);
  and _56977_ (_05970_, _05969_, _05968_);
  or _56978_ (_05971_, _05934_, _00255_);
  or _56979_ (_05972_, _05894_, _00157_);
  and _56980_ (_05973_, _05972_, _05971_);
  and _56981_ (_05974_, _05973_, _05970_);
  or _56982_ (_05975_, _05942_, _00296_);
  or _56983_ (_05976_, _05931_, _00019_);
  and _56984_ (_05977_, _05976_, _05975_);
  or _56985_ (_05978_, _05902_, _00602_);
  or _56986_ (_05979_, _05923_, _00460_);
  and _56987_ (_05980_, _05979_, _05978_);
  and _56988_ (_05981_, _05980_, _05977_);
  and _56989_ (_05982_, _05981_, _05974_);
  and _56990_ (_05983_, _05982_, _05967_);
  or _56991_ (_05984_, _05983_, _05952_);
  nor _56992_ (_05985_, _05984_, _05653_);
  or _56993_ (_05986_, _05945_, _00045_);
  or _56994_ (_05987_, _05929_, _43732_);
  and _56995_ (_05988_, _05987_, _05986_);
  or _56996_ (_05989_, _05942_, _00281_);
  or _56997_ (_05990_, _05931_, _00004_);
  and _56998_ (_05991_, _05990_, _05989_);
  and _56999_ (_05992_, _05991_, _05988_);
  or _57000_ (_05993_, _05934_, _00240_);
  or _57001_ (_05994_, _05887_, _00199_);
  and _57002_ (_05995_, _05994_, _05993_);
  or _57003_ (_05996_, _05902_, _00584_);
  or _57004_ (_05997_, _05923_, _00445_);
  and _57005_ (_05998_, _05997_, _05996_);
  and _57006_ (_05999_, _05998_, _05995_);
  and _57007_ (_06000_, _05999_, _05992_);
  or _57008_ (_06001_, _05936_, _00086_);
  or _57009_ (_06002_, _05947_, _43773_);
  and _57010_ (_06003_, _06002_, _06001_);
  or _57011_ (_06004_, _05907_, _00404_);
  or _57012_ (_06005_, _05913_, _00363_);
  and _57013_ (_06006_, _06005_, _06004_);
  and _57014_ (_06007_, _06006_, _06003_);
  or _57015_ (_06008_, _05940_, _00527_);
  or _57016_ (_06009_, _05919_, _00486_);
  and _57017_ (_06010_, _06009_, _06008_);
  or _57018_ (_06011_, _05915_, _00322_);
  or _57019_ (_06012_, _05894_, _00127_);
  and _57020_ (_06013_, _06012_, _06011_);
  and _57021_ (_06014_, _06013_, _06010_);
  and _57022_ (_06015_, _06014_, _06007_);
  and _57023_ (_06016_, _06015_, _06000_);
  not _57024_ (_06017_, _06016_);
  not _57025_ (_06018_, _05668_);
  and _57026_ (_06019_, _05723_, _06018_);
  not _57027_ (_06020_, _06019_);
  nor _57028_ (_06021_, _06020_, _05952_);
  and _57029_ (_06022_, _06021_, _06017_);
  not _57030_ (_06023_, _05673_);
  and _57031_ (_06024_, _05648_, _05609_);
  and _57032_ (_06025_, _06024_, _05569_);
  and _57033_ (_06026_, _06025_, _05671_);
  not _57034_ (_06027_, _06026_);
  nor _57035_ (_06028_, _06027_, _05984_);
  not _57036_ (_06029_, \oc8051_golden_model_1.SP [0]);
  nor _57037_ (_06030_, _05686_, _06029_);
  not _57038_ (_06031_, _05685_);
  and _57039_ (_06032_, _06025_, _06031_);
  not _57040_ (_06033_, _06032_);
  nor _57041_ (_06034_, _06033_, _05984_);
  nor _57042_ (_06035_, _06033_, _05952_);
  not _57043_ (_06036_, _06035_);
  not _57044_ (_06037_, _05693_);
  and _57045_ (_06038_, _06037_, _05650_);
  and _57046_ (_06039_, _06025_, _06037_);
  not _57047_ (_06040_, _06039_);
  nor _57048_ (_06041_, _06040_, _05984_);
  not _57049_ (_06042_, _05689_);
  and _57050_ (_06043_, _06025_, _06042_);
  not _57051_ (_06044_, _06043_);
  or _57052_ (_06045_, _06044_, _05984_);
  not _57053_ (_06046_, _05705_);
  and _57054_ (_06047_, _05750_, _06018_);
  not _57055_ (_06048_, _06047_);
  and _57056_ (_06049_, _06025_, _05746_);
  not _57057_ (_06050_, _06049_);
  and _57058_ (_06051_, _05746_, _06018_);
  not _57059_ (_06052_, _06051_);
  not _57060_ (_06053_, _05952_);
  nor _57061_ (_06054_, _05907_, _00434_);
  nor _57062_ (_06055_, _05934_, _00270_);
  nor _57063_ (_06056_, _06055_, _06054_);
  nor _57064_ (_06057_, _05887_, _00229_);
  nor _57065_ (_06058_, _05929_, _43762_);
  nor _57066_ (_06059_, _06058_, _06057_);
  and _57067_ (_06060_, _06059_, _06056_);
  nor _57068_ (_06061_, _05919_, _00516_);
  nor _57069_ (_06062_, _05940_, _00566_);
  nor _57070_ (_06063_, _06062_, _06061_);
  nor _57071_ (_06064_, _05902_, _00617_);
  nor _57072_ (_06065_, _05945_, _00075_);
  nor _57073_ (_06066_, _06065_, _06064_);
  and _57074_ (_06067_, _06066_, _06063_);
  and _57075_ (_06068_, _06067_, _06060_);
  nor _57076_ (_06069_, _05894_, _00188_);
  nor _57077_ (_06070_, _05936_, _00116_);
  nor _57078_ (_06071_, _06070_, _06069_);
  nor _57079_ (_06072_, _05923_, _00475_);
  nor _57080_ (_06073_, _05947_, _43803_);
  nor _57081_ (_06074_, _06073_, _06072_);
  and _57082_ (_06075_, _06074_, _06071_);
  nor _57083_ (_06076_, _05913_, _00393_);
  nor _57084_ (_06077_, _05931_, _00034_);
  nor _57085_ (_06078_, _06077_, _06076_);
  nor _57086_ (_06079_, _05915_, _00352_);
  nor _57087_ (_06080_, _05942_, _00311_);
  nor _57088_ (_06081_, _06080_, _06079_);
  and _57089_ (_06082_, _06081_, _06078_);
  and _57090_ (_06083_, _06082_, _06075_);
  and _57091_ (_06084_, _06083_, _06068_);
  and _57092_ (_06085_, _06084_, _06053_);
  and _57093_ (_06086_, _05983_, _05952_);
  nor _57094_ (_06087_, _06086_, _06085_);
  and _57095_ (_06088_, _06025_, _05723_);
  and _57096_ (_06089_, _06025_, _05659_);
  nor _57097_ (_06090_, _06089_, _06088_);
  nor _57098_ (_06091_, _06090_, _06087_);
  not _57099_ (_06092_, _05661_);
  and _57100_ (_06093_, _05567_, _05531_);
  and _57101_ (_06094_, _06093_, _06092_);
  and _57102_ (_06095_, _05567_, _05666_);
  and _57103_ (_06096_, _06095_, _05649_);
  not _57104_ (_06097_, _05665_);
  and _57105_ (_06098_, _06093_, _06097_);
  or _57106_ (_06099_, _06098_, _06096_);
  nor _57107_ (_06100_, _06099_, _06094_);
  or _57108_ (_06101_, _06100_, _05685_);
  nor _57109_ (_06102_, _05689_, _05668_);
  nor _57110_ (_06103_, _05667_, _05610_);
  and _57111_ (_06104_, _06103_, _06031_);
  nor _57112_ (_06105_, _06104_, _06102_);
  and _57113_ (_06106_, _06105_, _06101_);
  not _57114_ (_06107_, _05662_);
  and _57115_ (_06108_, _05735_, _06107_);
  nor _57116_ (_06109_, _06108_, _06019_);
  and _57117_ (_06110_, _05671_, _05650_);
  not _57118_ (_06111_, _06110_);
  and _57119_ (_06112_, _05726_, _06107_);
  not _57120_ (_06113_, _05667_);
  and _57121_ (_06114_, _06113_, _05649_);
  and _57122_ (_06115_, _06114_, _06031_);
  nor _57123_ (_06116_, _06115_, _06112_);
  and _57124_ (_06117_, _06116_, _06111_);
  and _57125_ (_06118_, _06117_, _06109_);
  and _57126_ (_06119_, _06025_, _05750_);
  nor _57127_ (_06120_, _06119_, _05652_);
  nor _57128_ (_06121_, _05685_, _05668_);
  and _57129_ (_06122_, _06093_, _06024_);
  and _57130_ (_06123_, _06122_, _06031_);
  nor _57131_ (_06124_, _06123_, _06121_);
  and _57132_ (_06125_, _06124_, _06120_);
  and _57133_ (_06126_, _05746_, _05650_);
  and _57134_ (_06127_, _06025_, _05495_);
  nor _57135_ (_06128_, _06127_, _06126_);
  and _57136_ (_06129_, _05731_, _05650_);
  and _57137_ (_06130_, _05739_, _06107_);
  nor _57138_ (_06131_, _06130_, _06129_);
  and _57139_ (_06132_, _06131_, _06128_);
  and _57140_ (_06133_, _06095_, _06097_);
  and _57141_ (_06134_, _06133_, _06031_);
  and _57142_ (_06135_, _06095_, _05609_);
  and _57143_ (_06136_, _06093_, _05649_);
  nor _57144_ (_06137_, _06136_, _06135_);
  nor _57145_ (_06138_, _06137_, _05685_);
  or _57146_ (_06139_, _06138_, _06134_);
  not _57147_ (_06140_, _06139_);
  and _57148_ (_06141_, _06140_, _06132_);
  and _57149_ (_06142_, _06141_, _06125_);
  and _57150_ (_06143_, _06142_, _06118_);
  and _57151_ (_06144_, _06143_, _06106_);
  nor _57152_ (_06145_, _06144_, _05803_);
  and _57153_ (_06146_, _06144_, _05824_);
  nor _57154_ (_06147_, _06146_, _06145_);
  not _57155_ (_06148_, _05853_);
  nor _57156_ (_06149_, _06144_, _06148_);
  not _57157_ (_06150_, _05870_);
  and _57158_ (_06151_, _06144_, _06150_);
  nor _57159_ (_06152_, _06151_, _06149_);
  nor _57160_ (_06153_, _06152_, _06147_);
  and _57161_ (_06154_, _06144_, _05346_);
  nor _57162_ (_06155_, _06154_, \oc8051_golden_model_1.PC [1]);
  and _57163_ (_06156_, _06154_, \oc8051_golden_model_1.PC [1]);
  nor _57164_ (_06157_, _06156_, _06155_);
  nor _57165_ (_06158_, _06144_, _05346_);
  nor _57166_ (_06159_, _06158_, _06154_);
  nor _57167_ (_06160_, _06159_, _06157_);
  and _57168_ (_06161_, _06160_, _06153_);
  and _57169_ (_06162_, _06161_, _04446_);
  and _57170_ (_06163_, _06159_, _06157_);
  not _57171_ (_06164_, _06152_);
  nor _57172_ (_06165_, _06164_, _06147_);
  and _57173_ (_06166_, _06165_, _06163_);
  and _57174_ (_06167_, _06166_, _04486_);
  nor _57175_ (_06168_, _06167_, _06162_);
  and _57176_ (_06169_, _06164_, _06147_);
  and _57177_ (_06170_, _06169_, _06160_);
  and _57178_ (_06171_, _06170_, _04462_);
  not _57179_ (_06172_, _06159_);
  nor _57180_ (_06173_, _06172_, _06157_);
  and _57181_ (_06174_, _06152_, _06147_);
  and _57182_ (_06175_, _06174_, _06173_);
  and _57183_ (_06176_, _06175_, _04473_);
  nor _57184_ (_06177_, _06176_, _06171_);
  and _57185_ (_06178_, _06177_, _06168_);
  and _57186_ (_06179_, _06173_, _06153_);
  and _57187_ (_06180_, _06179_, _04477_);
  and _57188_ (_06181_, _06172_, _06157_);
  and _57189_ (_06182_, _06181_, _06153_);
  and _57190_ (_06183_, _06182_, _04464_);
  nor _57191_ (_06184_, _06183_, _06180_);
  and _57192_ (_06185_, _06173_, _06169_);
  and _57193_ (_06186_, _06185_, _04467_);
  and _57194_ (_06187_, _06165_, _06160_);
  and _57195_ (_06188_, _06187_, _04457_);
  nor _57196_ (_06189_, _06188_, _06186_);
  and _57197_ (_06190_, _06189_, _06184_);
  and _57198_ (_06191_, _06190_, _06178_);
  and _57199_ (_06192_, _06174_, _06163_);
  and _57200_ (_06193_, _06192_, _04459_);
  and _57201_ (_06194_, _06181_, _06165_);
  and _57202_ (_06195_, _06194_, _04475_);
  nor _57203_ (_06196_, _06195_, _06193_);
  and _57204_ (_06197_, _06174_, _06160_);
  and _57205_ (_06198_, _06197_, _04469_);
  and _57206_ (_06199_, _06174_, _06181_);
  and _57207_ (_06200_, _06199_, _04448_);
  nor _57208_ (_06201_, _06200_, _06198_);
  and _57209_ (_06202_, _06201_, _06196_);
  and _57210_ (_06203_, _06163_, _06153_);
  and _57211_ (_06204_, _06203_, _04484_);
  and _57212_ (_06205_, _06173_, _06165_);
  and _57213_ (_06206_, _06205_, _04479_);
  nor _57214_ (_06207_, _06206_, _06204_);
  and _57215_ (_06208_, _06181_, _06169_);
  and _57216_ (_06209_, _06208_, _04453_);
  and _57217_ (_06210_, _06169_, _06163_);
  and _57218_ (_06211_, _06210_, _04451_);
  nor _57219_ (_06212_, _06211_, _06209_);
  and _57220_ (_06213_, _06212_, _06207_);
  and _57221_ (_06214_, _06213_, _06202_);
  and _57222_ (_06215_, _06214_, _06191_);
  nor _57223_ (_06216_, _06215_, _05669_);
  not _57224_ (_06217_, _06090_);
  nor _57225_ (_06218_, _06121_, _06038_);
  nor _57226_ (_06219_, _05693_, _05668_);
  not _57227_ (_06220_, _06219_);
  not _57228_ (_06221_, _05701_);
  and _57229_ (_06222_, _06093_, _06221_);
  not _57230_ (_06223_, _06222_);
  and _57231_ (_06224_, _06096_, _06221_);
  and _57232_ (_06225_, _06133_, _06221_);
  nor _57233_ (_06226_, _06225_, _06224_);
  and _57234_ (_06227_, _06095_, _06024_);
  and _57235_ (_06228_, _06227_, _06221_);
  and _57236_ (_06229_, _06095_, _06092_);
  and _57237_ (_06230_, _06229_, _06221_);
  nor _57238_ (_06231_, _06230_, _06228_);
  and _57239_ (_06232_, _06231_, _06226_);
  and _57240_ (_06233_, _06232_, _06223_);
  and _57241_ (_06234_, _06233_, _06220_);
  and _57242_ (_06235_, _06234_, _06218_);
  or _57243_ (_06236_, _06235_, _05983_);
  nor _57244_ (_06237_, _06044_, _06087_);
  not _57245_ (_06238_, \oc8051_golden_model_1.SP [3]);
  and _57246_ (_06239_, _06042_, _05650_);
  and _57247_ (_06240_, _06239_, _06238_);
  nor _57248_ (_06241_, _05697_, _05668_);
  nor _57249_ (_06242_, _06241_, _06102_);
  or _57250_ (_06243_, _06242_, _05983_);
  nor _57251_ (_06244_, _06239_, _06043_);
  nand _57252_ (_06245_, _06242_, \oc8051_golden_model_1.PSW [3]);
  and _57253_ (_06246_, _06245_, _06244_);
  or _57254_ (_06247_, _06246_, _06219_);
  and _57255_ (_06248_, _06247_, _06243_);
  or _57256_ (_06249_, _06248_, _06240_);
  and _57257_ (_06250_, _06221_, _05650_);
  and _57258_ (_06251_, _06025_, _06221_);
  nor _57259_ (_06252_, _06251_, _06250_);
  and _57260_ (_06253_, _06031_, _05650_);
  nor _57261_ (_06254_, _06032_, _06253_);
  and _57262_ (_06255_, _06254_, _06040_);
  and _57263_ (_06256_, _06255_, _06252_);
  and _57264_ (_06257_, _06256_, _06249_);
  or _57265_ (_06258_, _06257_, _06237_);
  and _57266_ (_06259_, _06258_, _06236_);
  nor _57267_ (_06260_, _06256_, _06087_);
  nor _57268_ (_06261_, _05672_, _05668_);
  nand _57269_ (_06262_, _06233_, _06218_);
  and _57270_ (_06263_, _06262_, _05983_);
  or _57271_ (_06264_, _06263_, _06261_);
  or _57272_ (_06265_, _06264_, _06260_);
  nor _57273_ (_06266_, _06265_, _06259_);
  not _57274_ (_06267_, _06261_);
  nor _57275_ (_06268_, _06267_, _05983_);
  or _57276_ (_06269_, _06268_, _06266_);
  and _57277_ (_06270_, _06269_, _06027_);
  and _57278_ (_06271_, _06087_, _06026_);
  or _57279_ (_06272_, _06271_, _06270_);
  and _57280_ (_06273_, _06272_, _05669_);
  or _57281_ (_06274_, _06273_, _06217_);
  nor _57282_ (_06275_, _06274_, _06216_);
  or _57283_ (_06276_, _06275_, _06091_);
  and _57284_ (_06277_, _06025_, _05735_);
  not _57285_ (_06278_, _06277_);
  and _57286_ (_06279_, _05735_, _06018_);
  nor _57287_ (_06280_, _06279_, _06108_);
  and _57288_ (_06281_, _06280_, _06278_);
  and _57289_ (_06282_, _05726_, _06018_);
  not _57290_ (_06283_, _06282_);
  and _57291_ (_06284_, _06025_, _05726_);
  nor _57292_ (_06285_, _06284_, _06112_);
  and _57293_ (_06286_, _06285_, _06283_);
  and _57294_ (_06287_, _06286_, _06281_);
  and _57295_ (_06288_, _05731_, _06018_);
  not _57296_ (_06289_, _06288_);
  and _57297_ (_06290_, _05739_, _06018_);
  not _57298_ (_06291_, _06290_);
  and _57299_ (_06292_, _06025_, _05739_);
  nor _57300_ (_06293_, _06292_, _06130_);
  and _57301_ (_06294_, _06293_, _06291_);
  and _57302_ (_06295_, _06294_, _06289_);
  and _57303_ (_06296_, _06295_, _06287_);
  nand _57304_ (_06297_, _06296_, _06276_);
  and _57305_ (_06298_, _06025_, _05731_);
  not _57306_ (_06299_, _05983_);
  nor _57307_ (_06300_, _06296_, _06299_);
  nor _57308_ (_06301_, _06300_, _06298_);
  and _57309_ (_06302_, _06301_, _06297_);
  and _57310_ (_06303_, _06298_, \oc8051_golden_model_1.SP [3]);
  or _57311_ (_06304_, _06303_, _06129_);
  nor _57312_ (_06305_, _06304_, _06302_);
  not _57313_ (_06306_, _06129_);
  nor _57314_ (_06307_, _06087_, _06306_);
  or _57315_ (_06308_, _06307_, _06305_);
  and _57316_ (_06309_, _06308_, _06052_);
  and _57317_ (_06310_, _06051_, _05983_);
  or _57318_ (_06311_, _06310_, _06309_);
  nand _57319_ (_06312_, _06311_, _06050_);
  and _57320_ (_06313_, _06049_, _06238_);
  nor _57321_ (_06314_, _06313_, _06126_);
  nand _57322_ (_06315_, _06314_, _06312_);
  and _57323_ (_06316_, _06018_, _05495_);
  and _57324_ (_06317_, _06126_, _06087_);
  nor _57325_ (_06318_, _06317_, _06316_);
  nand _57326_ (_06319_, _06318_, _06315_);
  and _57327_ (_06320_, _06316_, _05983_);
  nor _57328_ (_06321_, _06320_, _05652_);
  and _57329_ (_06322_, _06321_, _06319_);
  and _57330_ (_06323_, _06087_, _05652_);
  or _57331_ (_06324_, _06323_, _06322_);
  nand _57332_ (_06325_, _06324_, _06048_);
  nor _57333_ (_06326_, _06048_, _05983_);
  not _57334_ (_06327_, _06326_);
  and _57335_ (_06328_, _06327_, _06325_);
  nor _57336_ (_06329_, _05902_, _00612_);
  nor _57337_ (_06330_, _05915_, _00347_);
  nor _57338_ (_06331_, _06330_, _06329_);
  nor _57339_ (_06332_, _05913_, _00388_);
  nor _57340_ (_06333_, _05945_, _00070_);
  nor _57341_ (_06334_, _06333_, _06332_);
  and _57342_ (_06335_, _06334_, _06331_);
  nor _57343_ (_06336_, _05934_, _00265_);
  nor _57344_ (_06337_, _05894_, _00179_);
  nor _57345_ (_06338_, _06337_, _06336_);
  nor _57346_ (_06339_, _05940_, _00558_);
  nor _57347_ (_06340_, _05923_, _00470_);
  nor _57348_ (_06341_, _06340_, _06339_);
  and _57349_ (_06342_, _06341_, _06338_);
  and _57350_ (_06343_, _06342_, _06335_);
  nor _57351_ (_06344_, _05936_, _00111_);
  nor _57352_ (_06345_, _05931_, _00029_);
  nor _57353_ (_06346_, _06345_, _06344_);
  nor _57354_ (_06347_, _05929_, _43757_);
  nor _57355_ (_06348_, _05947_, _43798_);
  nor _57356_ (_06349_, _06348_, _06347_);
  and _57357_ (_06350_, _06349_, _06346_);
  nor _57358_ (_06351_, _05919_, _00511_);
  nor _57359_ (_06352_, _05887_, _00224_);
  nor _57360_ (_06353_, _06352_, _06351_);
  nor _57361_ (_06354_, _05907_, _00429_);
  nor _57362_ (_06355_, _05942_, _00306_);
  nor _57363_ (_06356_, _06355_, _06354_);
  and _57364_ (_06357_, _06356_, _06353_);
  and _57365_ (_06358_, _06357_, _06350_);
  and _57366_ (_06359_, _06358_, _06343_);
  nor _57367_ (_06360_, _06359_, _05952_);
  not _57368_ (_06361_, _06360_);
  and _57369_ (_06362_, _06254_, _06252_);
  nor _57370_ (_06363_, _06126_, _06043_);
  and _57371_ (_06364_, _06363_, _06306_);
  nor _57372_ (_06365_, _06026_, _05652_);
  and _57373_ (_06366_, _06365_, _06090_);
  and _57374_ (_06367_, _06366_, _06364_);
  and _57375_ (_06368_, _06367_, _06362_);
  nor _57376_ (_06369_, _06368_, _06361_);
  not _57377_ (_06370_, _06369_);
  and _57378_ (_06371_, _06360_, _06039_);
  not _57379_ (_06372_, _06371_);
  nor _57380_ (_06373_, _05915_, _00332_);
  nor _57381_ (_06374_, _05936_, _00096_);
  nor _57382_ (_06375_, _06374_, _06373_);
  nor _57383_ (_06376_, _05902_, _00597_);
  nor _57384_ (_06377_, _05934_, _00250_);
  nor _57385_ (_06378_, _06377_, _06376_);
  and _57386_ (_06379_, _06378_, _06375_);
  nor _57387_ (_06380_, _05942_, _00291_);
  nor _57388_ (_06381_, _05894_, _00146_);
  nor _57389_ (_06382_, _06381_, _06380_);
  nor _57390_ (_06383_, _05929_, _43742_);
  nor _57391_ (_06384_, _05947_, _43783_);
  nor _57392_ (_06385_, _06384_, _06383_);
  and _57393_ (_06386_, _06385_, _06382_);
  and _57394_ (_06387_, _06386_, _06379_);
  nor _57395_ (_06388_, _05919_, _00496_);
  nor _57396_ (_06389_, _05913_, _00373_);
  nor _57397_ (_06390_, _06389_, _06388_);
  nor _57398_ (_06391_, _05887_, _00209_);
  nor _57399_ (_06392_, _05931_, _00014_);
  nor _57400_ (_06393_, _06392_, _06391_);
  and _57401_ (_06394_, _06393_, _06390_);
  nor _57402_ (_06395_, _05907_, _00414_);
  nor _57403_ (_06396_, _05923_, _00455_);
  nor _57404_ (_06397_, _06396_, _06395_);
  nor _57405_ (_06398_, _05940_, _00537_);
  nor _57406_ (_06399_, _05945_, _00055_);
  nor _57407_ (_06400_, _06399_, _06398_);
  and _57408_ (_06401_, _06400_, _06397_);
  and _57409_ (_06402_, _06401_, _06394_);
  and _57410_ (_06403_, _06402_, _06387_);
  nor _57411_ (_06404_, _06288_, _06261_);
  and _57412_ (_06405_, _06404_, _06218_);
  and _57413_ (_06406_, _06405_, _06242_);
  and _57414_ (_06407_, _06406_, _06234_);
  nor _57415_ (_06408_, _06316_, _06047_);
  and _57416_ (_06409_, _06408_, _06052_);
  and _57417_ (_06410_, _06409_, _06294_);
  and _57418_ (_06411_, _06410_, _06287_);
  and _57419_ (_06412_, _06411_, _06407_);
  nor _57420_ (_06413_, _06412_, _06403_);
  not _57421_ (_06414_, _06413_);
  and _57422_ (_06415_, _06170_, _04437_);
  and _57423_ (_06416_, _06161_, _04406_);
  nor _57424_ (_06417_, _06416_, _06415_);
  and _57425_ (_06418_, _06192_, _04410_);
  and _57426_ (_06419_, _06166_, _04417_);
  nor _57427_ (_06420_, _06419_, _06418_);
  and _57428_ (_06421_, _06420_, _06417_);
  and _57429_ (_06422_, _06185_, _04415_);
  and _57430_ (_06423_, _06210_, _04399_);
  nor _57431_ (_06424_, _06423_, _06422_);
  and _57432_ (_06425_, _06179_, _04428_);
  and _57433_ (_06426_, _06203_, _04439_);
  nor _57434_ (_06427_, _06426_, _06425_);
  and _57435_ (_06428_, _06427_, _06424_);
  and _57436_ (_06429_, _06428_, _06421_);
  and _57437_ (_06430_, _06197_, _04422_);
  and _57438_ (_06431_, _06175_, _04426_);
  nor _57439_ (_06432_, _06431_, _06430_);
  and _57440_ (_06433_, _06199_, _04401_);
  and _57441_ (_06434_, _06187_, _04412_);
  nor _57442_ (_06435_, _06434_, _06433_);
  and _57443_ (_06436_, _06435_, _06432_);
  and _57444_ (_06437_, _06205_, _04432_);
  and _57445_ (_06438_, _06194_, _04430_);
  nor _57446_ (_06439_, _06438_, _06437_);
  and _57447_ (_06440_, _06208_, _04404_);
  and _57448_ (_06441_, _06182_, _04420_);
  nor _57449_ (_06442_, _06441_, _06440_);
  and _57450_ (_06443_, _06442_, _06439_);
  and _57451_ (_06444_, _06443_, _06436_);
  and _57452_ (_06445_, _06444_, _06429_);
  nor _57453_ (_06446_, _06445_, _05669_);
  not _57454_ (_06447_, \oc8051_golden_model_1.SP [2]);
  nor _57455_ (_06448_, _06298_, _06049_);
  nor _57456_ (_06449_, _06448_, _06447_);
  and _57457_ (_06450_, _06093_, _05609_);
  not _57458_ (_06451_, _06450_);
  and _57459_ (_06452_, _05453_, _05414_);
  or _57460_ (_06453_, _06037_, _05659_);
  nor _57461_ (_06454_, _06453_, _06452_);
  nor _57462_ (_06455_, _06454_, _06451_);
  nor _57463_ (_06456_, _06455_, _06449_);
  and _57464_ (_06457_, _06136_, _05495_);
  and _57465_ (_06458_, _06098_, _05495_);
  nor _57466_ (_06459_, _06458_, _06457_);
  and _57467_ (_06460_, _06093_, _05610_);
  and _57468_ (_06461_, _06460_, _06042_);
  not _57469_ (_06462_, _06461_);
  and _57470_ (_06463_, _06460_, _06037_);
  and _57471_ (_06464_, _06093_, _05750_);
  nor _57472_ (_06465_, _06464_, _06463_);
  and _57473_ (_06466_, _06465_, _06462_);
  and _57474_ (_06467_, _06466_, _06459_);
  and _57475_ (_06468_, _06467_, _06456_);
  not _57476_ (_06469_, _06460_);
  nor _57477_ (_06470_, _05731_, _05659_);
  and _57478_ (_06471_, _05697_, _05685_);
  nor _57479_ (_06472_, _05726_, _05671_);
  and _57480_ (_06473_, _06472_, _06471_);
  and _57481_ (_06474_, _06473_, _06470_);
  nor _57482_ (_06475_, _06474_, _06469_);
  not _57483_ (_06476_, _06475_);
  and _57484_ (_06477_, _06093_, _05739_);
  not _57485_ (_06478_, _06477_);
  and _57486_ (_06479_, _06239_, \oc8051_golden_model_1.SP [2]);
  not _57487_ (_06480_, _06479_);
  and _57488_ (_06481_, _06450_, _05746_);
  and _57489_ (_06482_, _06450_, _05735_);
  nor _57490_ (_06483_, _06482_, _06481_);
  and _57491_ (_06484_, _06483_, _06480_);
  and _57492_ (_06485_, _06484_, _06478_);
  and _57493_ (_06486_, _06471_, _05689_);
  nor _57494_ (_06487_, _06486_, _06451_);
  not _57495_ (_06488_, _06487_);
  and _57496_ (_06489_, _06450_, _05726_);
  and _57497_ (_06490_, _06460_, _05735_);
  nor _57498_ (_06491_, _06490_, _06489_);
  and _57499_ (_06492_, _06450_, _05671_);
  and _57500_ (_06493_, _06460_, _05746_);
  nor _57501_ (_06494_, _06493_, _06492_);
  and _57502_ (_06495_, _06494_, _06491_);
  and _57503_ (_06496_, _06495_, _06488_);
  and _57504_ (_06497_, _06496_, _06485_);
  and _57505_ (_06498_, _06497_, _06476_);
  and _57506_ (_06499_, _06498_, _06468_);
  not _57507_ (_06500_, _06499_);
  nor _57508_ (_06501_, _06500_, _06446_);
  and _57509_ (_06502_, _06501_, _06414_);
  and _57510_ (_06503_, _06502_, _06372_);
  and _57511_ (_06504_, _06503_, _06370_);
  not _57512_ (_06505_, \oc8051_golden_model_1.IRAM[0] [0]);
  nor _57513_ (_06506_, _06048_, _06016_);
  not _57514_ (_06507_, _06506_);
  nor _57515_ (_06508_, _06267_, _06016_);
  not _57516_ (_06509_, _06121_);
  nor _57517_ (_06510_, _06509_, _06016_);
  or _57518_ (_06511_, _06220_, _06016_);
  nor _57519_ (_06512_, _06242_, _06016_);
  and _57520_ (_06513_, _06024_, _06113_);
  and _57521_ (_06514_, _06513_, _06042_);
  not _57522_ (_06515_, _06514_);
  and _57523_ (_06516_, _06122_, _06042_);
  not _57524_ (_06517_, _06096_);
  nor _57525_ (_06518_, _06136_, _06227_);
  nand _57526_ (_06519_, _06518_, _06517_);
  and _57527_ (_06520_, _06519_, _06042_);
  nor _57528_ (_06521_, _06520_, _06516_);
  and _57529_ (_06522_, _06521_, _06515_);
  not _57530_ (_06523_, _05697_);
  and _57531_ (_06524_, _06227_, _06523_);
  and _57532_ (_06525_, _06096_, _06523_);
  nor _57533_ (_06526_, _06525_, _06524_);
  and _57534_ (_06527_, _06513_, _06523_);
  or _57535_ (_06528_, _06527_, _06241_);
  not _57536_ (_06529_, _06528_);
  and _57537_ (_06530_, _06122_, _06523_);
  nor _57538_ (_06531_, _06530_, _06102_);
  and _57539_ (_06532_, _06136_, _06523_);
  not _57540_ (_06533_, _05703_);
  and _57541_ (_06534_, _06513_, _06533_);
  nor _57542_ (_06535_, _06534_, _06532_);
  and _57543_ (_06536_, _06535_, _06531_);
  and _57544_ (_06537_, _06536_, _06529_);
  and _57545_ (_06538_, _06537_, _06526_);
  and _57546_ (_06539_, _06538_, _06522_);
  or _57547_ (_06540_, _06539_, _06512_);
  nand _57548_ (_06541_, _06540_, _06044_);
  nand _57549_ (_06542_, _06045_, _06541_);
  and _57550_ (_06543_, _06239_, _06029_);
  nor _57551_ (_06544_, _06543_, _06219_);
  not _57552_ (_06545_, _05648_);
  and _57553_ (_06546_, _06450_, _06037_);
  and _57554_ (_06547_, _06135_, _06037_);
  nor _57555_ (_06548_, _06547_, _06546_);
  nor _57556_ (_06549_, _06548_, _06545_);
  not _57557_ (_06550_, _06549_);
  and _57558_ (_06551_, _06136_, _06037_);
  not _57559_ (_06552_, _06551_);
  and _57560_ (_06553_, _06513_, _06037_);
  and _57561_ (_06554_, _06096_, _06037_);
  nor _57562_ (_06555_, _06554_, _06553_);
  and _57563_ (_06556_, _06555_, _06552_);
  and _57564_ (_06557_, _06556_, _06550_);
  and _57565_ (_06558_, _06557_, _06544_);
  nand _57566_ (_06559_, _06558_, _06542_);
  nand _57567_ (_06560_, _06559_, _06511_);
  and _57568_ (_06561_, _06560_, _06040_);
  or _57569_ (_06562_, _06041_, _06561_);
  and _57570_ (_06563_, _06038_, _06016_);
  nor _57571_ (_06564_, _06122_, _06018_);
  nor _57572_ (_06565_, _06513_, _06096_);
  and _57573_ (_06566_, _06565_, _06564_);
  and _57574_ (_06567_, _06566_, _06518_);
  nor _57575_ (_06568_, _06567_, _05685_);
  nor _57576_ (_06569_, _06568_, _06563_);
  and _57577_ (_06570_, _06569_, _06562_);
  or _57578_ (_06571_, _06570_, _06510_);
  nand _57579_ (_06572_, _06571_, _06254_);
  not _57580_ (_06573_, _06233_);
  nor _57581_ (_06574_, _06254_, _05984_);
  nor _57582_ (_06575_, _06574_, _06573_);
  nand _57583_ (_06576_, _06575_, _06572_);
  and _57584_ (_06577_, _06573_, _06016_);
  not _57585_ (_06578_, _06252_);
  and _57586_ (_06579_, _06513_, _06221_);
  nor _57587_ (_06580_, _06579_, _06578_);
  not _57588_ (_06581_, _06580_);
  nor _57589_ (_06582_, _06581_, _06577_);
  and _57590_ (_06583_, _06582_, _06576_);
  nor _57591_ (_06584_, _06252_, _05984_);
  or _57592_ (_06585_, _06584_, _06583_);
  nor _57593_ (_06586_, _06096_, _06018_);
  and _57594_ (_06587_, _06093_, _05648_);
  not _57595_ (_06588_, _06587_);
  and _57596_ (_06589_, _06588_, _06586_);
  nor _57597_ (_06590_, _06589_, _05672_);
  and _57598_ (_06591_, _06513_, _05671_);
  and _57599_ (_06592_, _06135_, _05671_);
  and _57600_ (_06593_, _06592_, _05648_);
  nor _57601_ (_06594_, _06593_, _06591_);
  not _57602_ (_06595_, _06594_);
  nor _57603_ (_06596_, _06595_, _06590_);
  and _57604_ (_06597_, _06596_, _06585_);
  or _57605_ (_06598_, _06597_, _06508_);
  and _57606_ (_06599_, _06598_, _06027_);
  nor _57607_ (_06600_, _06599_, _06028_);
  nor _57608_ (_06601_, _06567_, _05660_);
  nor _57609_ (_06602_, _06601_, _06600_);
  and _57610_ (_06603_, _06161_, _04306_);
  and _57611_ (_06604_, _06194_, _04335_);
  nor _57612_ (_06605_, _06604_, _06603_);
  and _57613_ (_06606_, _06170_, _04322_);
  and _57614_ (_06607_, _06175_, _04333_);
  nor _57615_ (_06608_, _06607_, _06606_);
  and _57616_ (_06609_, _06608_, _06605_);
  and _57617_ (_06610_, _06179_, _04337_);
  and _57618_ (_06611_, _06182_, _04324_);
  nor _57619_ (_06612_, _06611_, _06610_);
  and _57620_ (_06613_, _06185_, _04327_);
  and _57621_ (_06614_, _06187_, _04317_);
  nor _57622_ (_06615_, _06614_, _06613_);
  and _57623_ (_06616_, _06615_, _06612_);
  and _57624_ (_06617_, _06616_, _06609_);
  and _57625_ (_06618_, _06192_, _04319_);
  and _57626_ (_06619_, _06166_, _04347_);
  nor _57627_ (_06620_, _06619_, _06618_);
  and _57628_ (_06621_, _06197_, _04329_);
  and _57629_ (_06622_, _06199_, _04308_);
  nor _57630_ (_06623_, _06622_, _06621_);
  and _57631_ (_06624_, _06623_, _06620_);
  and _57632_ (_06625_, _06203_, _04344_);
  and _57633_ (_06626_, _06205_, _04339_);
  nor _57634_ (_06627_, _06626_, _06625_);
  and _57635_ (_06628_, _06208_, _04313_);
  and _57636_ (_06629_, _06210_, _04311_);
  nor _57637_ (_06630_, _06629_, _06628_);
  and _57638_ (_06631_, _06630_, _06627_);
  and _57639_ (_06632_, _06631_, _06624_);
  and _57640_ (_06633_, _06632_, _06617_);
  nor _57641_ (_06634_, _06633_, _05669_);
  or _57642_ (_06635_, _06634_, _06602_);
  not _57643_ (_06636_, _06088_);
  and _57644_ (_06637_, _06089_, _05984_);
  and _57645_ (_06638_, _06513_, _05723_);
  nor _57646_ (_06639_, _06638_, _06637_);
  and _57647_ (_06640_, _06639_, _06636_);
  and _57648_ (_06641_, _06640_, _06635_);
  nor _57649_ (_06642_, _06636_, _05984_);
  or _57650_ (_06643_, _06642_, _06641_);
  not _57651_ (_06644_, _05726_);
  nor _57652_ (_06645_, _06518_, _06644_);
  not _57653_ (_06646_, _06645_);
  and _57654_ (_06647_, _06513_, _05726_);
  not _57655_ (_06648_, _06647_);
  and _57656_ (_06649_, _06122_, _05726_);
  and _57657_ (_06650_, _06096_, _05726_);
  nor _57658_ (_06651_, _06650_, _06649_);
  and _57659_ (_06652_, _06651_, _06648_);
  and _57660_ (_06653_, _06652_, _06646_);
  and _57661_ (_06654_, _06653_, _06643_);
  nor _57662_ (_06655_, _06286_, _06017_);
  not _57663_ (_06656_, _05735_);
  not _57664_ (_06657_, _06227_);
  and _57665_ (_06658_, _06565_, _06657_);
  and _57666_ (_06659_, _06588_, _06658_);
  nor _57667_ (_06660_, _06659_, _06656_);
  nor _57668_ (_06661_, _06660_, _06655_);
  and _57669_ (_06663_, _06661_, _06654_);
  nor _57670_ (_06664_, _06281_, _06017_);
  and _57671_ (_06665_, _06227_, _05739_);
  not _57672_ (_06666_, _06665_);
  and _57673_ (_06667_, _06096_, _05739_);
  not _57674_ (_06668_, _06667_);
  and _57675_ (_06669_, _06513_, _05739_);
  and _57676_ (_06670_, _06587_, _05739_);
  nor _57677_ (_06671_, _06670_, _06669_);
  and _57678_ (_06672_, _06671_, _06668_);
  and _57679_ (_06673_, _06672_, _06666_);
  not _57680_ (_06674_, _06673_);
  nor _57681_ (_06675_, _06674_, _06664_);
  and _57682_ (_06676_, _06675_, _06663_);
  nor _57683_ (_06677_, _06294_, _06017_);
  not _57684_ (_06678_, _05731_);
  nor _57685_ (_06679_, _06567_, _06678_);
  nor _57686_ (_06680_, _06679_, _06677_);
  and _57687_ (_06681_, _06680_, _06676_);
  nor _57688_ (_06682_, _06289_, _06016_);
  or _57689_ (_06683_, _06682_, _06681_);
  and _57690_ (_06684_, _06298_, _06029_);
  nor _57691_ (_06685_, _06684_, _06129_);
  and _57692_ (_06686_, _06685_, _06683_);
  nor _57693_ (_06687_, _06306_, _05984_);
  or _57694_ (_06688_, _06687_, _06686_);
  nor _57695_ (_06689_, _06493_, _06481_);
  or _57696_ (_06690_, _06689_, _06545_);
  and _57697_ (_06691_, _06227_, _05746_);
  and _57698_ (_06692_, _06513_, _05746_);
  and _57699_ (_06693_, _06096_, _05746_);
  or _57700_ (_06694_, _06693_, _06051_);
  or _57701_ (_06695_, _06694_, _06692_);
  nor _57702_ (_06696_, _06695_, _06691_);
  and _57703_ (_06697_, _06696_, _06690_);
  and _57704_ (_06698_, _06697_, _06688_);
  nor _57705_ (_06699_, _06052_, _06016_);
  or _57706_ (_06700_, _06699_, _06698_);
  and _57707_ (_06701_, _06049_, _06029_);
  nor _57708_ (_06702_, _06701_, _06126_);
  and _57709_ (_06703_, _06702_, _06700_);
  not _57710_ (_06704_, _06126_);
  nor _57711_ (_06705_, _06704_, _05984_);
  or _57712_ (_06706_, _06705_, _06703_);
  and _57713_ (_06707_, _06227_, _05495_);
  and _57714_ (_06708_, _06096_, _05495_);
  or _57715_ (_06709_, _06708_, _06707_);
  not _57716_ (_06710_, _06709_);
  and _57717_ (_06711_, _06122_, _05495_);
  and _57718_ (_06712_, _06513_, _05495_);
  nor _57719_ (_06713_, _06712_, _06711_);
  nor _57720_ (_06714_, _06457_, _06316_);
  and _57721_ (_06715_, _06714_, _06713_);
  and _57722_ (_06716_, _06715_, _06710_);
  and _57723_ (_06717_, _06716_, _06706_);
  not _57724_ (_06718_, _06316_);
  nor _57725_ (_06719_, _06718_, _06016_);
  or _57726_ (_06720_, _06719_, _06717_);
  and _57727_ (_06721_, _06720_, _05653_);
  nor _57728_ (_06722_, _06721_, _05985_);
  not _57729_ (_06723_, _05750_);
  nor _57730_ (_06724_, _06567_, _06723_);
  or _57731_ (_06725_, _06724_, _06722_);
  nand _57732_ (_06726_, _06725_, _06507_);
  or _57733_ (_06727_, _06726_, _06505_);
  nor _57734_ (_06728_, _05934_, _00260_);
  nor _57735_ (_06729_, _05887_, _00219_);
  nor _57736_ (_06730_, _06729_, _06728_);
  nor _57737_ (_06731_, _05894_, _00168_);
  nor _57738_ (_06732_, _05945_, _00065_);
  nor _57739_ (_06733_, _06732_, _06731_);
  and _57740_ (_06734_, _06733_, _06730_);
  nor _57741_ (_06735_, _05902_, _00607_);
  nor _57742_ (_06736_, _05940_, _00550_);
  nor _57743_ (_06737_, _06736_, _06735_);
  nor _57744_ (_06738_, _05919_, _00506_);
  nor _57745_ (_06739_, _05913_, _00383_);
  nor _57746_ (_06740_, _06739_, _06738_);
  and _57747_ (_06741_, _06740_, _06737_);
  and _57748_ (_06742_, _06741_, _06734_);
  nor _57749_ (_06743_, _05915_, _00342_);
  nor _57750_ (_06744_, _05929_, _43752_);
  nor _57751_ (_06745_, _06744_, _06743_);
  nor _57752_ (_06746_, _05907_, _00424_);
  nor _57753_ (_06747_, _05947_, _43793_);
  nor _57754_ (_06748_, _06747_, _06746_);
  and _57755_ (_06749_, _06748_, _06745_);
  nor _57756_ (_06750_, _05942_, _00301_);
  nor _57757_ (_06751_, _05931_, _00024_);
  nor _57758_ (_06752_, _06751_, _06750_);
  nor _57759_ (_06753_, _05923_, _00465_);
  nor _57760_ (_06754_, _05936_, _00106_);
  nor _57761_ (_06755_, _06754_, _06753_);
  and _57762_ (_06756_, _06755_, _06752_);
  and _57763_ (_06757_, _06756_, _06749_);
  and _57764_ (_06758_, _06757_, _06742_);
  nor _57765_ (_06759_, _06758_, _05952_);
  nor _57766_ (_06760_, _06039_, _05652_);
  and _57767_ (_06761_, _06760_, _06090_);
  and _57768_ (_06762_, _06761_, _06364_);
  and _57769_ (_06763_, _06762_, _06362_);
  not _57770_ (_06764_, _06763_);
  and _57771_ (_06765_, _06764_, _06759_);
  not _57772_ (_06766_, _06765_);
  and _57773_ (_06767_, _06759_, _06026_);
  not _57774_ (_06768_, _06767_);
  nor _57775_ (_06769_, _05907_, _00409_);
  nor _57776_ (_06770_, _05934_, _00245_);
  nor _57777_ (_06771_, _06770_, _06769_);
  nor _57778_ (_06772_, _05887_, _00204_);
  nor _57779_ (_06773_, _05947_, _43778_);
  nor _57780_ (_06774_, _06773_, _06772_);
  and _57781_ (_06775_, _06774_, _06771_);
  nor _57782_ (_06776_, _05902_, _00592_);
  nor _57783_ (_06777_, _05945_, _00050_);
  nor _57784_ (_06778_, _06777_, _06776_);
  nor _57785_ (_06779_, _05940_, _00532_);
  nor _57786_ (_06780_, _05942_, _00286_);
  nor _57787_ (_06781_, _06780_, _06779_);
  and _57788_ (_06782_, _06781_, _06778_);
  and _57789_ (_06783_, _06782_, _06775_);
  nor _57790_ (_06784_, _05894_, _00135_);
  nor _57791_ (_06785_, _05936_, _00091_);
  nor _57792_ (_06786_, _06785_, _06784_);
  nor _57793_ (_06787_, _05913_, _00368_);
  nor _57794_ (_06788_, _05929_, _43737_);
  nor _57795_ (_06789_, _06788_, _06787_);
  and _57796_ (_06790_, _06789_, _06786_);
  nor _57797_ (_06791_, _05919_, _00491_);
  nor _57798_ (_06792_, _05931_, _00009_);
  nor _57799_ (_06793_, _06792_, _06791_);
  nor _57800_ (_06794_, _05923_, _00450_);
  nor _57801_ (_06795_, _05915_, _00327_);
  nor _57802_ (_06796_, _06795_, _06794_);
  and _57803_ (_06797_, _06796_, _06793_);
  and _57804_ (_06798_, _06797_, _06790_);
  and _57805_ (_06799_, _06798_, _06783_);
  nor _57806_ (_06800_, _06799_, _06412_);
  not _57807_ (_06801_, _06800_);
  and _57808_ (_06802_, _06194_, _04382_);
  and _57809_ (_06803_, _06205_, _04386_);
  nor _57810_ (_06804_, _06803_, _06802_);
  and _57811_ (_06805_, _06185_, _04374_);
  and _57812_ (_06806_, _06175_, _04380_);
  nor _57813_ (_06807_, _06806_, _06805_);
  and _57814_ (_06808_, _06807_, _06804_);
  and _57815_ (_06809_, _06161_, _04353_);
  and _57816_ (_06810_, _06203_, _04391_);
  nor _57817_ (_06811_, _06810_, _06809_);
  and _57818_ (_06812_, _06192_, _04366_);
  and _57819_ (_06813_, _06166_, _04393_);
  nor _57820_ (_06814_, _06813_, _06812_);
  and _57821_ (_06815_, _06814_, _06811_);
  and _57822_ (_06816_, _06815_, _06808_);
  and _57823_ (_06817_, _06210_, _04358_);
  and _57824_ (_06818_, _06182_, _04371_);
  nor _57825_ (_06819_, _06818_, _06817_);
  and _57826_ (_06820_, _06170_, _04369_);
  and _57827_ (_06821_, _06208_, _04360_);
  nor _57828_ (_06822_, _06821_, _06820_);
  and _57829_ (_06823_, _06822_, _06819_);
  and _57830_ (_06824_, _06179_, _04384_);
  and _57831_ (_06825_, _06187_, _04364_);
  nor _57832_ (_06826_, _06825_, _06824_);
  and _57833_ (_06827_, _06197_, _04376_);
  and _57834_ (_06828_, _06199_, _04355_);
  nor _57835_ (_06829_, _06828_, _06827_);
  and _57836_ (_06830_, _06829_, _06826_);
  and _57837_ (_06831_, _06830_, _06823_);
  and _57838_ (_06832_, _06831_, _06816_);
  nor _57839_ (_06833_, _06832_, _05669_);
  and _57840_ (_06834_, _06135_, _05739_);
  and _57841_ (_06835_, _06135_, _05735_);
  nor _57842_ (_06836_, _06835_, _06834_);
  and _57843_ (_06837_, _06135_, _06031_);
  nor _57844_ (_06838_, _06592_, _06837_);
  and _57845_ (_06839_, _06838_, _06836_);
  and _57846_ (_06840_, _06839_, _06488_);
  not _57847_ (_06841_, _05746_);
  nor _57848_ (_06842_, _05739_, _05735_);
  and _57849_ (_06843_, _06842_, _06841_);
  nor _57850_ (_06844_, _06843_, _06451_);
  nor _57851_ (_06845_, _06844_, _06455_);
  and _57852_ (_06846_, _06845_, _06840_);
  not _57853_ (_06847_, \oc8051_golden_model_1.SP [1]);
  not _57854_ (_06848_, _06239_);
  and _57855_ (_06849_, _06448_, _06848_);
  nor _57856_ (_06850_, _06849_, _06847_);
  not _57857_ (_06851_, _06850_);
  not _57858_ (_06852_, _06229_);
  nor _57859_ (_06853_, _05746_, _06523_);
  nor _57860_ (_06854_, _06853_, _06852_);
  not _57861_ (_06855_, _06854_);
  nor _57862_ (_06856_, _06450_, _06135_);
  nor _57863_ (_06857_, _05750_, _05726_);
  nor _57864_ (_06858_, _06857_, _06856_);
  not _57865_ (_06859_, _06135_);
  nor _57866_ (_06860_, _06470_, _06859_);
  nor _57867_ (_06861_, _06860_, _06858_);
  and _57868_ (_06862_, _06861_, _06855_);
  and _57869_ (_06863_, _06135_, _06042_);
  not _57870_ (_06864_, _06863_);
  and _57871_ (_06865_, _06229_, _05495_);
  nor _57872_ (_06866_, _06865_, _06707_);
  and _57873_ (_06867_, _06866_, _06864_);
  nor _57874_ (_06868_, _06547_, _06492_);
  and _57875_ (_06869_, _06868_, _06867_);
  nor _57876_ (_06870_, _06691_, _06524_);
  and _57877_ (_06871_, _06870_, _06869_);
  and _57878_ (_06872_, _06871_, _06862_);
  and _57879_ (_06873_, _06872_, _06851_);
  and _57880_ (_06874_, _06873_, _06846_);
  not _57881_ (_06875_, _06874_);
  nor _57882_ (_06876_, _06875_, _06833_);
  and _57883_ (_06877_, _06876_, _06801_);
  and _57884_ (_06878_, _06877_, _06768_);
  and _57885_ (_06879_, _06878_, _06766_);
  not _57886_ (_06880_, \oc8051_golden_model_1.IRAM[1] [0]);
  and _57887_ (_06881_, _06725_, _06507_);
  or _57888_ (_06882_, _06881_, _06880_);
  and _57889_ (_06883_, _06882_, _06879_);
  nand _57890_ (_06884_, _06883_, _06727_);
  not _57891_ (_06885_, \oc8051_golden_model_1.IRAM[3] [0]);
  or _57892_ (_06886_, _06881_, _06885_);
  not _57893_ (_06887_, _06879_);
  not _57894_ (_06888_, \oc8051_golden_model_1.IRAM[2] [0]);
  or _57895_ (_06889_, _06726_, _06888_);
  and _57896_ (_06890_, _06889_, _06887_);
  nand _57897_ (_06891_, _06890_, _06886_);
  nand _57898_ (_06892_, _06891_, _06884_);
  nand _57899_ (_06893_, _06892_, _06504_);
  not _57900_ (_06894_, _06504_);
  not _57901_ (_06895_, \oc8051_golden_model_1.IRAM[7] [0]);
  or _57902_ (_06896_, _06881_, _06895_);
  nand _57903_ (_06897_, _06881_, \oc8051_golden_model_1.IRAM[6] [0]);
  and _57904_ (_06898_, _06897_, _06887_);
  nand _57905_ (_06899_, _06898_, _06896_);
  nand _57906_ (_06900_, _06881_, \oc8051_golden_model_1.IRAM[4] [0]);
  nand _57907_ (_06901_, _06726_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _57908_ (_06902_, _06901_, _06879_);
  nand _57909_ (_06903_, _06902_, _06900_);
  nand _57910_ (_06904_, _06903_, _06899_);
  nand _57911_ (_06905_, _06904_, _06894_);
  nand _57912_ (_06906_, _06905_, _06893_);
  nand _57913_ (_06907_, _06906_, _06328_);
  not _57914_ (_06908_, _06328_);
  nand _57915_ (_06909_, _06726_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand _57916_ (_06910_, _06881_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _57917_ (_06911_, _06910_, _06887_);
  nand _57918_ (_06912_, _06911_, _06909_);
  nand _57919_ (_06913_, _06881_, \oc8051_golden_model_1.IRAM[8] [0]);
  nand _57920_ (_06914_, _06726_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _57921_ (_06915_, _06914_, _06879_);
  nand _57922_ (_06916_, _06915_, _06913_);
  nand _57923_ (_06917_, _06916_, _06912_);
  nand _57924_ (_06918_, _06917_, _06504_);
  nand _57925_ (_06919_, _06726_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand _57926_ (_06920_, _06881_, \oc8051_golden_model_1.IRAM[14] [0]);
  and _57927_ (_06921_, _06920_, _06887_);
  nand _57928_ (_06922_, _06921_, _06919_);
  nand _57929_ (_06923_, _06881_, \oc8051_golden_model_1.IRAM[12] [0]);
  nand _57930_ (_06924_, _06726_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _57931_ (_06925_, _06924_, _06879_);
  nand _57932_ (_06926_, _06925_, _06923_);
  nand _57933_ (_06927_, _06926_, _06922_);
  nand _57934_ (_06928_, _06927_, _06894_);
  nand _57935_ (_06929_, _06928_, _06918_);
  nand _57936_ (_06930_, _06929_, _06908_);
  and _57937_ (_06931_, _06930_, _06907_);
  and _57938_ (_06932_, _06931_, _06046_);
  nor _57939_ (_06933_, _06114_, _05718_);
  and _57940_ (_06934_, _06933_, _06565_);
  nor _57941_ (_06935_, _06934_, _05703_);
  not _57942_ (_06936_, _06935_);
  nor _57943_ (_06937_, _06936_, _06932_);
  and _57944_ (_06938_, _06094_, _06523_);
  not _57945_ (_06939_, _06938_);
  nor _57946_ (_06940_, _06939_, _05952_);
  and _57947_ (_06941_, _06940_, _06016_);
  nor _57948_ (_06942_, _06941_, _06937_);
  and _57949_ (_06943_, _06098_, _06523_);
  and _57950_ (_06944_, _06943_, \oc8051_golden_model_1.SP [0]);
  not _57951_ (_06945_, _06944_);
  and _57952_ (_06946_, _06945_, _06521_);
  and _57953_ (_06947_, _06946_, _06942_);
  and _57954_ (_06948_, _06103_, _06042_);
  not _57955_ (_06949_, _06948_);
  nor _57956_ (_06950_, _06949_, _06931_);
  not _57957_ (_06951_, _06950_);
  and _57958_ (_06952_, _06951_, _06947_);
  nor _57959_ (_06953_, _06044_, _05952_);
  not _57960_ (_06954_, _06102_);
  nor _57961_ (_06955_, _06954_, _05952_);
  and _57962_ (_06956_, _06955_, _06016_);
  nor _57963_ (_06957_, _06956_, _06953_);
  and _57964_ (_06958_, _06957_, _06952_);
  not _57965_ (_06959_, _06958_);
  and _57966_ (_06960_, _06959_, _06045_);
  nor _57967_ (_06961_, _05690_, _06029_);
  nor _57968_ (_06962_, _06961_, _06960_);
  nor _57969_ (_06963_, _06848_, _05952_);
  and _57970_ (_06964_, _06963_, _06016_);
  or _57971_ (_06965_, _06554_, _06551_);
  nor _57972_ (_06966_, _06965_, _06549_);
  not _57973_ (_06967_, _06966_);
  nor _57974_ (_06968_, _06967_, _06964_);
  and _57975_ (_06969_, _06968_, _06962_);
  and _57976_ (_06970_, _06103_, _06037_);
  not _57977_ (_06971_, _06970_);
  nor _57978_ (_06972_, _06971_, _06931_);
  not _57979_ (_06973_, _06972_);
  and _57980_ (_06974_, _06973_, _06969_);
  nor _57981_ (_06975_, _06040_, _05952_);
  nor _57982_ (_06976_, _06220_, _05952_);
  and _57983_ (_06977_, _06976_, _06016_);
  nor _57984_ (_06978_, _06977_, _06975_);
  and _57985_ (_06979_, _06978_, _06974_);
  nor _57986_ (_06980_, _06979_, _06041_);
  or _57987_ (_06981_, _06980_, _06038_);
  nand _57988_ (_06982_, _06038_, _06029_);
  nand _57989_ (_06983_, _06982_, _06981_);
  and _57990_ (_06984_, _06983_, _06036_);
  nor _57991_ (_06985_, _06984_, _06034_);
  or _57992_ (_06986_, _06228_, _06224_);
  and _57993_ (_06987_, _06587_, _06221_);
  or _57994_ (_06988_, _06987_, _06986_);
  or _57995_ (_06989_, _06988_, _06985_);
  nor _57996_ (_06990_, _06989_, _06030_);
  nor _57997_ (_06991_, _06027_, _05952_);
  and _57998_ (_06992_, _06103_, _06221_);
  not _57999_ (_06993_, _06992_);
  nor _58000_ (_06994_, _06993_, _06931_);
  nor _58001_ (_06995_, _06994_, _06991_);
  and _58002_ (_06996_, _06995_, _06990_);
  nor _58003_ (_06997_, _06996_, _06028_);
  nor _58004_ (_06998_, _06997_, _06023_);
  nor _58005_ (_06999_, _05673_, \oc8051_golden_model_1.SP [0]);
  nor _58006_ (_07000_, _06999_, _06998_);
  nor _58007_ (_07001_, _05952_, _05660_);
  and _58008_ (_07002_, _06095_, _05610_);
  or _58009_ (_07003_, _07002_, _06136_);
  and _58010_ (_07004_, _07003_, _07001_);
  or _58011_ (_07005_, _06450_, _06098_);
  nor _58012_ (_07006_, _07005_, _06135_);
  not _58013_ (_07007_, _07006_);
  and _58014_ (_07008_, _07007_, _07001_);
  nor _58015_ (_07009_, _07008_, _07004_);
  nor _58016_ (_07010_, _05952_, _05669_);
  and _58017_ (_07011_, _06103_, _05659_);
  not _58018_ (_07012_, _07011_);
  nor _58019_ (_07013_, _07012_, _05952_);
  nor _58020_ (_07014_, _07013_, _07010_);
  and _58021_ (_07015_, _07014_, _07009_);
  nor _58022_ (_07016_, _07015_, _06017_);
  and _58023_ (_07017_, _05648_, _05567_);
  and _58024_ (_07018_, _07017_, _05723_);
  nor _58025_ (_07019_, _07018_, _07016_);
  not _58026_ (_07020_, _07019_);
  nor _58027_ (_07021_, _07020_, _07000_);
  not _58028_ (_07022_, _06931_);
  and _58029_ (_07023_, _06103_, _05723_);
  and _58030_ (_07024_, _07023_, _07022_);
  nor _58031_ (_07025_, _07024_, _06021_);
  and _58032_ (_07026_, _07025_, _07021_);
  nor _58033_ (_07027_, _07026_, _06022_);
  nor _58034_ (_07028_, _07027_, _05724_);
  and _58035_ (_07029_, _05724_, _06029_);
  nor _58036_ (_07030_, _07029_, _07028_);
  nor _58037_ (_07031_, _06278_, _05952_);
  not _58038_ (_07032_, _06108_);
  and _58039_ (_07033_, _06285_, _07032_);
  nor _58040_ (_07034_, _07033_, _05952_);
  nor _58041_ (_07035_, _07034_, _07031_);
  nor _58042_ (_07036_, _07035_, _06017_);
  nor _58043_ (_07037_, _07036_, _05736_);
  not _58044_ (_07038_, _07037_);
  nor _58045_ (_07039_, _07038_, _07030_);
  and _58046_ (_07040_, _05736_, _06029_);
  nor _58047_ (_07041_, _07040_, _07039_);
  nor _58048_ (_07042_, _06293_, _05952_);
  and _58049_ (_07043_, _07042_, _06016_);
  nor _58050_ (_07044_, _07043_, _07041_);
  and _58051_ (_07045_, _05732_, \oc8051_golden_model_1.SP [0]);
  and _58052_ (_07046_, _06587_, _05495_);
  nor _58053_ (_07047_, _07046_, _07045_);
  and _58054_ (_07048_, _07047_, _06710_);
  and _58055_ (_07049_, _07048_, _07044_);
  nor _58056_ (_07050_, _06718_, _05952_);
  and _58057_ (_07051_, _06103_, _05495_);
  not _58058_ (_07052_, _07051_);
  nor _58059_ (_07053_, _07052_, _06931_);
  nor _58060_ (_07054_, _07053_, _07050_);
  and _58061_ (_07055_, _07054_, _07049_);
  and _58062_ (_07056_, _07050_, _06017_);
  nor _58063_ (_07057_, _07056_, _07055_);
  nor _58064_ (_07058_, _05952_, _05653_);
  nor _58065_ (_07059_, _06127_, _05752_);
  nor _58066_ (_07060_, _07059_, _06029_);
  nor _58067_ (_07061_, _07060_, _07058_);
  not _58068_ (_07062_, _07061_);
  nor _58069_ (_07063_, _07062_, _07057_);
  nor _58070_ (_07064_, _07063_, _05985_);
  and _58071_ (_07065_, _07017_, _05750_);
  nor _58072_ (_07066_, _07065_, _07064_);
  nor _58073_ (_07067_, _06048_, _05952_);
  and _58074_ (_07068_, _06103_, _05750_);
  not _58075_ (_07069_, _07068_);
  nor _58076_ (_07070_, _07069_, _06931_);
  nor _58077_ (_07071_, _07070_, _07067_);
  and _58078_ (_07072_, _07071_, _07066_);
  and _58079_ (_07073_, _07067_, _06017_);
  nor _58080_ (_07074_, _07073_, _07072_);
  not _58081_ (_07075_, _07074_);
  not _58082_ (_07076_, _06799_);
  and _58083_ (_07077_, _07067_, _07076_);
  and _58084_ (_07078_, _06460_, _05750_);
  and _58085_ (_07079_, _06759_, _05652_);
  and _58086_ (_07080_, _06847_, \oc8051_golden_model_1.SP [0]);
  and _58087_ (_07081_, \oc8051_golden_model_1.SP [1], _06029_);
  nor _58088_ (_07082_, _07081_, _07080_);
  not _58089_ (_07083_, _07082_);
  nor _58090_ (_07084_, _07083_, _07059_);
  and _58091_ (_07085_, _07083_, _05732_);
  and _58092_ (_07086_, _07076_, _06021_);
  and _58093_ (_07087_, _06103_, _06533_);
  nand _58094_ (_07088_, _06881_, \oc8051_golden_model_1.IRAM[0] [1]);
  nand _58095_ (_07089_, _06726_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _58096_ (_07090_, _07089_, _06879_);
  nand _58097_ (_07091_, _07090_, _07088_);
  nand _58098_ (_07092_, _06726_, \oc8051_golden_model_1.IRAM[3] [1]);
  nand _58099_ (_07093_, _06881_, \oc8051_golden_model_1.IRAM[2] [1]);
  and _58100_ (_07094_, _07093_, _06887_);
  nand _58101_ (_07095_, _07094_, _07092_);
  nand _58102_ (_07096_, _07095_, _07091_);
  nand _58103_ (_07097_, _07096_, _06504_);
  nand _58104_ (_07098_, _06726_, \oc8051_golden_model_1.IRAM[7] [1]);
  nand _58105_ (_07099_, _06881_, \oc8051_golden_model_1.IRAM[6] [1]);
  and _58106_ (_07100_, _07099_, _06887_);
  nand _58107_ (_07101_, _07100_, _07098_);
  nand _58108_ (_07102_, _06881_, \oc8051_golden_model_1.IRAM[4] [1]);
  nand _58109_ (_07103_, _06726_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _58110_ (_07104_, _07103_, _06879_);
  nand _58111_ (_07105_, _07104_, _07102_);
  nand _58112_ (_07106_, _07105_, _07101_);
  nand _58113_ (_07107_, _07106_, _06894_);
  nand _58114_ (_07108_, _07107_, _07097_);
  nand _58115_ (_07109_, _07108_, _06328_);
  nand _58116_ (_07110_, _06726_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand _58117_ (_07111_, _06881_, \oc8051_golden_model_1.IRAM[10] [1]);
  and _58118_ (_07112_, _07111_, _06887_);
  nand _58119_ (_07113_, _07112_, _07110_);
  nand _58120_ (_07114_, _06881_, \oc8051_golden_model_1.IRAM[8] [1]);
  nand _58121_ (_07115_, _06726_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _58122_ (_07116_, _07115_, _06879_);
  nand _58123_ (_07117_, _07116_, _07114_);
  nand _58124_ (_07118_, _07117_, _07113_);
  nand _58125_ (_07119_, _07118_, _06504_);
  nand _58126_ (_07120_, _06726_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand _58127_ (_07121_, _06881_, \oc8051_golden_model_1.IRAM[14] [1]);
  and _58128_ (_07122_, _07121_, _06887_);
  nand _58129_ (_07123_, _07122_, _07120_);
  nand _58130_ (_07124_, _06881_, \oc8051_golden_model_1.IRAM[12] [1]);
  nand _58131_ (_07125_, _06726_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _58132_ (_07126_, _07125_, _06879_);
  nand _58133_ (_07127_, _07126_, _07124_);
  nand _58134_ (_07128_, _07127_, _07123_);
  nand _58135_ (_07129_, _07128_, _06894_);
  nand _58136_ (_07130_, _07129_, _07119_);
  nand _58137_ (_07131_, _07130_, _06908_);
  nand _58138_ (_07132_, _07131_, _07109_);
  and _58139_ (_07133_, _07132_, _06046_);
  or _58140_ (_07134_, _07133_, _07087_);
  and _58141_ (_07135_, _06940_, _06799_);
  or _58142_ (_07136_, _07135_, _07134_);
  and _58143_ (_07137_, _07082_, _06943_);
  not _58144_ (_07138_, _07137_);
  and _58145_ (_07139_, _07002_, _06042_);
  nor _58146_ (_07140_, _07139_, _06461_);
  and _58147_ (_07141_, _07140_, _07138_);
  not _58148_ (_07142_, _07141_);
  nor _58149_ (_07143_, _07142_, _07136_);
  and _58150_ (_07144_, _07132_, _06948_);
  nor _58151_ (_07145_, _07144_, _06955_);
  and _58152_ (_07146_, _07145_, _07143_);
  and _58153_ (_07147_, _06955_, _07076_);
  nor _58154_ (_07148_, _07147_, _07146_);
  and _58155_ (_07149_, _06758_, _06953_);
  nor _58156_ (_07150_, _07149_, _07148_);
  or _58157_ (_07151_, _07083_, _05690_);
  nand _58158_ (_07152_, _07151_, _07150_);
  and _58159_ (_07153_, _06963_, _06799_);
  and _58160_ (_07154_, _07002_, _06037_);
  nor _58161_ (_07155_, _07154_, _06463_);
  not _58162_ (_07156_, _07155_);
  nor _58163_ (_07157_, _07156_, _07153_);
  not _58164_ (_07158_, _07157_);
  nor _58165_ (_07159_, _07158_, _07152_);
  and _58166_ (_07160_, _07132_, _06970_);
  nor _58167_ (_07161_, _07160_, _06976_);
  and _58168_ (_07162_, _07161_, _07159_);
  and _58169_ (_07163_, _06976_, _07076_);
  nor _58170_ (_07164_, _07163_, _07162_);
  and _58171_ (_07165_, _06758_, _06975_);
  nor _58172_ (_07166_, _07165_, _06038_);
  not _58173_ (_07167_, _07166_);
  nor _58174_ (_07168_, _07167_, _07164_);
  and _58175_ (_07169_, _07083_, _06038_);
  nor _58176_ (_07170_, _07169_, _07168_);
  and _58177_ (_07171_, _06035_, _06758_);
  nor _58178_ (_07172_, _07171_, _07170_);
  nand _58179_ (_07173_, _06222_, _05610_);
  and _58180_ (_07174_, _07002_, _06221_);
  nor _58181_ (_07175_, _07083_, _05686_);
  nor _58182_ (_07176_, _07175_, _07174_);
  and _58183_ (_07177_, _07176_, _07173_);
  and _58184_ (_07178_, _07177_, _07172_);
  and _58185_ (_07179_, _07132_, _06992_);
  nor _58186_ (_07180_, _07179_, _06991_);
  and _58187_ (_07181_, _07180_, _07178_);
  nor _58188_ (_07182_, _07181_, _06767_);
  nor _58189_ (_07183_, _07182_, _06023_);
  nor _58190_ (_07184_, _07082_, _05673_);
  nor _58191_ (_07185_, _07184_, _07183_);
  nor _58192_ (_07186_, _07015_, _07076_);
  and _58193_ (_07187_, _05723_, _05610_);
  and _58194_ (_07188_, _07187_, _05567_);
  nor _58195_ (_07189_, _07188_, _07186_);
  not _58196_ (_07190_, _07189_);
  nor _58197_ (_07191_, _07190_, _07185_);
  and _58198_ (_07192_, _07132_, _07023_);
  nor _58199_ (_07193_, _07192_, _06021_);
  and _58200_ (_07194_, _07193_, _07191_);
  nor _58201_ (_07195_, _07194_, _07086_);
  nor _58202_ (_07196_, _07195_, _05724_);
  and _58203_ (_07197_, _07083_, _05724_);
  nor _58204_ (_07198_, _07197_, _07196_);
  nor _58205_ (_07199_, _07035_, _07076_);
  nor _58206_ (_07200_, _07199_, _05736_);
  not _58207_ (_07201_, _07200_);
  nor _58208_ (_07202_, _07201_, _07198_);
  and _58209_ (_07203_, _07083_, _05736_);
  nor _58210_ (_07204_, _07203_, _07202_);
  and _58211_ (_07205_, _07042_, _06799_);
  nor _58212_ (_07206_, _07205_, _05732_);
  not _58213_ (_07207_, _07206_);
  nor _58214_ (_07208_, _07207_, _07204_);
  nor _58215_ (_07209_, _07208_, _07085_);
  and _58216_ (_07210_, _07002_, _05495_);
  not _58217_ (_07211_, _07210_);
  and _58218_ (_07212_, _07211_, _06459_);
  not _58219_ (_07213_, _07212_);
  nor _58220_ (_07214_, _07213_, _07209_);
  and _58221_ (_07215_, _07132_, _07051_);
  nor _58222_ (_07216_, _07215_, _07050_);
  and _58223_ (_07217_, _07216_, _07214_);
  and _58224_ (_07218_, _07050_, _07076_);
  nor _58225_ (_07219_, _07218_, _07217_);
  or _58226_ (_07220_, _07219_, _07058_);
  nor _58227_ (_07221_, _07220_, _07084_);
  nor _58228_ (_07222_, _07221_, _07079_);
  and _58229_ (_07223_, _07002_, _05750_);
  or _58230_ (_07224_, _07223_, _07222_);
  nor _58231_ (_07225_, _07224_, _07078_);
  and _58232_ (_07226_, _07132_, _07068_);
  nor _58233_ (_07227_, _07226_, _07067_);
  and _58234_ (_07228_, _07227_, _07225_);
  nor _58235_ (_07229_, _07228_, _07077_);
  not _58236_ (_07230_, _00000_);
  not _58237_ (_07231_, _07013_);
  not _58238_ (_07232_, _07067_);
  not _58239_ (_07233_, _06943_);
  and _58240_ (_07234_, _07059_, _07233_);
  nor _58241_ (_07235_, _05736_, _05732_);
  and _58242_ (_07236_, _06867_, _07235_);
  and _58243_ (_07237_, _07236_, _07234_);
  and _58244_ (_07238_, _06450_, _06042_);
  nor _58245_ (_07239_, _06948_, _07238_);
  and _58246_ (_07240_, _07239_, _06548_);
  nor _58247_ (_07241_, _06554_, _06038_);
  nor _58248_ (_07242_, _07051_, _06992_);
  and _58249_ (_07243_, _07242_, _07241_);
  and _58250_ (_07244_, _07243_, _07240_);
  and _58251_ (_07245_, _07244_, _07237_);
  nand _58252_ (_07246_, _06933_, _05668_);
  and _58253_ (_07247_, _07246_, _06533_);
  nor _58254_ (_07248_, _07002_, _06103_);
  nor _58255_ (_07249_, _07248_, _05703_);
  or _58256_ (_07250_, _07249_, _07247_);
  not _58257_ (_07251_, _07250_);
  and _58258_ (_07252_, _06095_, _05723_);
  not _58259_ (_07253_, _07252_);
  and _58260_ (_07254_, _06094_, _05723_);
  and _58261_ (_07255_, _06222_, _06545_);
  nor _58262_ (_07256_, _07255_, _07254_);
  and _58263_ (_07257_, _07256_, _07253_);
  and _58264_ (_07258_, _07257_, _07251_);
  and _58265_ (_07259_, _07258_, _07245_);
  and _58266_ (_07260_, _07069_, _06467_);
  and _58267_ (_07261_, _06133_, _06037_);
  nor _58268_ (_07262_, _07261_, _07139_);
  nor _58269_ (_07263_, _07210_, _07174_);
  and _58270_ (_07264_, _07263_, _07262_);
  nor _58271_ (_07265_, _06987_, _06970_);
  and _58272_ (_07266_, _06093_, _05661_);
  and _58273_ (_07267_, _07266_, _05723_);
  nor _58274_ (_07268_, _07267_, _07023_);
  and _58275_ (_07269_, _07268_, _07265_);
  and _58276_ (_07270_, _07269_, _07264_);
  and _58277_ (_07271_, _05686_, _05673_);
  not _58278_ (_07272_, _05690_);
  nor _58279_ (_07273_, _05724_, _07272_);
  and _58280_ (_07274_, _07273_, _07271_);
  and _58281_ (_07275_, _06135_, _06221_);
  and _58282_ (_07276_, _06135_, _05750_);
  nor _58283_ (_07277_, _07276_, _07275_);
  and _58284_ (_07278_, _06450_, _05495_);
  nor _58285_ (_07279_, _07223_, _07278_);
  and _58286_ (_07280_, _07279_, _07277_);
  and _58287_ (_07281_, _07280_, _07274_);
  and _58288_ (_07282_, _07281_, _07270_);
  and _58289_ (_07283_, _07282_, _07260_);
  and _58290_ (_07284_, _07283_, _07259_);
  and _58291_ (_07285_, _07284_, _07232_);
  and _58292_ (_07286_, _07285_, _07231_);
  and _58293_ (_07287_, _07286_, _07009_);
  nor _58294_ (_07288_, _06976_, _06963_);
  nor _58295_ (_07289_, _06955_, _06940_);
  and _58296_ (_07290_, _07289_, _07288_);
  nor _58297_ (_07291_, _07042_, _06021_);
  nor _58298_ (_07292_, _07010_, _06975_);
  and _58299_ (_07293_, _07292_, _07291_);
  and _58300_ (_07294_, _07293_, _07290_);
  not _58301_ (_07295_, _07058_);
  nor _58302_ (_07296_, _07050_, _07034_);
  and _58303_ (_07297_, _07296_, _07295_);
  nor _58304_ (_07298_, _06035_, _06953_);
  nor _58305_ (_07299_, _07031_, _06991_);
  and _58306_ (_07300_, _07299_, _07298_);
  and _58307_ (_07301_, _07300_, _07297_);
  and _58308_ (_07302_, _07301_, _07294_);
  and _58309_ (_07303_, _07302_, _07287_);
  nor _58310_ (_07304_, _07303_, _07230_);
  not _58311_ (_07305_, _07304_);
  nor _58312_ (_07306_, _07305_, _07229_);
  and _58313_ (_07307_, _07306_, _07075_);
  not _58314_ (_07308_, _06991_);
  nand _58315_ (_07309_, _06881_, \oc8051_golden_model_1.IRAM[0] [3]);
  nand _58316_ (_07310_, _06726_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _58317_ (_07311_, _07310_, _06879_);
  nand _58318_ (_07312_, _07311_, _07309_);
  nand _58319_ (_07313_, _06726_, \oc8051_golden_model_1.IRAM[3] [3]);
  nand _58320_ (_07314_, _06881_, \oc8051_golden_model_1.IRAM[2] [3]);
  and _58321_ (_07315_, _07314_, _06887_);
  nand _58322_ (_07316_, _07315_, _07313_);
  nand _58323_ (_07317_, _07316_, _07312_);
  nand _58324_ (_07318_, _07317_, _06504_);
  nand _58325_ (_07319_, _06726_, \oc8051_golden_model_1.IRAM[7] [3]);
  nand _58326_ (_07320_, _06881_, \oc8051_golden_model_1.IRAM[6] [3]);
  and _58327_ (_07321_, _07320_, _06887_);
  nand _58328_ (_07322_, _07321_, _07319_);
  nand _58329_ (_07323_, _06881_, \oc8051_golden_model_1.IRAM[4] [3]);
  nand _58330_ (_07324_, _06726_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _58331_ (_07325_, _07324_, _06879_);
  nand _58332_ (_07326_, _07325_, _07323_);
  nand _58333_ (_07327_, _07326_, _07322_);
  nand _58334_ (_07328_, _07327_, _06894_);
  nand _58335_ (_07329_, _07328_, _07318_);
  nand _58336_ (_07330_, _07329_, _06328_);
  nand _58337_ (_07331_, _06726_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _58338_ (_07332_, _06881_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _58339_ (_07333_, _07332_, _06887_);
  nand _58340_ (_07334_, _07333_, _07331_);
  nand _58341_ (_07335_, _06881_, \oc8051_golden_model_1.IRAM[8] [3]);
  nand _58342_ (_07336_, _06726_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _58343_ (_07337_, _07336_, _06879_);
  nand _58344_ (_07338_, _07337_, _07335_);
  nand _58345_ (_07339_, _07338_, _07334_);
  nand _58346_ (_07340_, _07339_, _06504_);
  nand _58347_ (_07341_, _06726_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _58348_ (_07342_, _06881_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _58349_ (_07343_, _07342_, _06887_);
  nand _58350_ (_07344_, _07343_, _07341_);
  nand _58351_ (_07345_, _06881_, \oc8051_golden_model_1.IRAM[12] [3]);
  nand _58352_ (_07346_, _06726_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _58353_ (_07347_, _07346_, _06879_);
  nand _58354_ (_07348_, _07347_, _07345_);
  nand _58355_ (_07349_, _07348_, _07344_);
  nand _58356_ (_07350_, _07349_, _06894_);
  nand _58357_ (_07351_, _07350_, _07340_);
  nand _58358_ (_07352_, _07351_, _06908_);
  nand _58359_ (_07353_, _07352_, _07330_);
  and _58360_ (_07354_, _07353_, _06992_);
  not _58361_ (_07355_, _05686_);
  and _58362_ (_07356_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _58363_ (_07357_, _07356_, \oc8051_golden_model_1.SP [2]);
  nor _58364_ (_07358_, _07357_, \oc8051_golden_model_1.SP [3]);
  and _58365_ (_07359_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _58366_ (_07360_, _07359_, \oc8051_golden_model_1.SP [3]);
  and _58367_ (_07361_, _07360_, \oc8051_golden_model_1.SP [0]);
  nor _58368_ (_07362_, _07361_, _07358_);
  and _58369_ (_07363_, _07362_, _07355_);
  not _58370_ (_07364_, _06038_);
  and _58371_ (_07365_, _06953_, _06084_);
  and _58372_ (_07366_, _07353_, _06948_);
  and _58373_ (_07367_, _07362_, _06943_);
  and _58374_ (_07368_, _07353_, _06046_);
  not _58375_ (_07369_, \oc8051_golden_model_1.PSW [3]);
  and _58376_ (_07370_, _05705_, _07369_);
  nor _58377_ (_07371_, _07370_, _06940_);
  not _58378_ (_07372_, _07371_);
  nor _58379_ (_07373_, _07372_, _07368_);
  and _58380_ (_07374_, _06940_, _06299_);
  nor _58381_ (_07375_, _07374_, _07373_);
  nor _58382_ (_07376_, _07375_, _06943_);
  or _58383_ (_07377_, _07376_, _06948_);
  nor _58384_ (_07378_, _07377_, _07367_);
  or _58385_ (_07379_, _07378_, _06955_);
  nor _58386_ (_07380_, _07379_, _07366_);
  and _58387_ (_07381_, _06955_, _06299_);
  or _58388_ (_07382_, _07381_, _06953_);
  nor _58389_ (_07383_, _07382_, _07380_);
  nor _58390_ (_07384_, _07383_, _07365_);
  nor _58391_ (_07385_, _07384_, _07272_);
  nor _58392_ (_07386_, _07362_, _05690_);
  nor _58393_ (_07387_, _07386_, _06963_);
  not _58394_ (_07388_, _07387_);
  nor _58395_ (_07389_, _07388_, _07385_);
  and _58396_ (_07390_, _06963_, _06299_);
  nor _58397_ (_07391_, _07390_, _06970_);
  not _58398_ (_07392_, _07391_);
  nor _58399_ (_07393_, _07392_, _07389_);
  and _58400_ (_07394_, _07353_, _06970_);
  nor _58401_ (_07395_, _07394_, _06976_);
  not _58402_ (_07396_, _07395_);
  nor _58403_ (_07397_, _07396_, _07393_);
  and _58404_ (_07398_, _06976_, _06299_);
  or _58405_ (_07399_, _07398_, _06975_);
  nor _58406_ (_07400_, _07399_, _07397_);
  and _58407_ (_07401_, _06084_, _06975_);
  nor _58408_ (_07402_, _07401_, _07400_);
  and _58409_ (_07403_, _07402_, _07364_);
  and _58410_ (_07404_, _07362_, _06038_);
  or _58411_ (_07405_, _07404_, _06035_);
  nor _58412_ (_07406_, _07405_, _07403_);
  and _58413_ (_07407_, _06032_, _06085_);
  or _58414_ (_07408_, _07407_, _07355_);
  nor _58415_ (_07409_, _07408_, _07406_);
  or _58416_ (_07410_, _07409_, _06992_);
  nor _58417_ (_07411_, _07410_, _07363_);
  nor _58418_ (_07412_, _07411_, _07354_);
  and _58419_ (_07413_, _07412_, _07308_);
  not _58420_ (_07414_, _06084_);
  and _58421_ (_07415_, _06991_, _07414_);
  or _58422_ (_07416_, _07415_, _07413_);
  and _58423_ (_07417_, _07416_, _05673_);
  and _58424_ (_07418_, _07362_, _06023_);
  not _58425_ (_07419_, _07418_);
  and _58426_ (_07420_, _07419_, _07015_);
  not _58427_ (_07421_, _07420_);
  nor _58428_ (_07422_, _07421_, _07417_);
  nor _58429_ (_07423_, _07015_, _06299_);
  nor _58430_ (_07424_, _07423_, _07422_);
  nor _58431_ (_07425_, _07424_, _07023_);
  and _58432_ (_07426_, _07353_, _07023_);
  nor _58433_ (_07427_, _07426_, _06021_);
  not _58434_ (_07428_, _07427_);
  nor _58435_ (_07429_, _07428_, _07425_);
  nor _58436_ (_07430_, _06020_, _05984_);
  nor _58437_ (_07431_, _07430_, _07429_);
  nor _58438_ (_07432_, _07431_, _05724_);
  and _58439_ (_07433_, _07362_, _05724_);
  not _58440_ (_07434_, _07433_);
  and _58441_ (_07435_, _07434_, _07035_);
  not _58442_ (_07436_, _07435_);
  nor _58443_ (_07437_, _07436_, _07432_);
  nor _58444_ (_07438_, _07035_, _06299_);
  nor _58445_ (_07439_, _07438_, _05736_);
  not _58446_ (_07440_, _07439_);
  nor _58447_ (_07441_, _07440_, _07437_);
  and _58448_ (_07442_, _07362_, _05736_);
  nor _58449_ (_07443_, _07442_, _07042_);
  not _58450_ (_07444_, _07443_);
  nor _58451_ (_07445_, _07444_, _07441_);
  and _58452_ (_07446_, _07042_, _05983_);
  nor _58453_ (_07447_, _07446_, _05732_);
  not _58454_ (_07448_, _07447_);
  nor _58455_ (_07449_, _07448_, _07445_);
  and _58456_ (_07450_, _07362_, _05732_);
  nor _58457_ (_07451_, _07450_, _07051_);
  not _58458_ (_07452_, _07451_);
  nor _58459_ (_07453_, _07452_, _07449_);
  and _58460_ (_07454_, _07353_, _07051_);
  nor _58461_ (_07455_, _07454_, _07050_);
  not _58462_ (_07456_, _07455_);
  nor _58463_ (_07457_, _07456_, _07453_);
  not _58464_ (_07458_, _07059_);
  and _58465_ (_07459_, _07050_, _06299_);
  nor _58466_ (_07460_, _07459_, _07458_);
  not _58467_ (_07461_, _07460_);
  nor _58468_ (_07462_, _07461_, _07457_);
  nor _58469_ (_07463_, _07362_, _07059_);
  nor _58470_ (_07464_, _07463_, _07058_);
  not _58471_ (_07465_, _07464_);
  nor _58472_ (_07466_, _07465_, _07462_);
  and _58473_ (_07467_, _07058_, _07414_);
  nor _58474_ (_07468_, _07467_, _07068_);
  not _58475_ (_07469_, _07468_);
  nor _58476_ (_07470_, _07469_, _07466_);
  and _58477_ (_07471_, _07353_, _07068_);
  nor _58478_ (_07472_, _07471_, _07067_);
  not _58479_ (_07473_, _07472_);
  nor _58480_ (_07474_, _07473_, _07470_);
  nor _58481_ (_07475_, _06048_, _05984_);
  nor _58482_ (_07476_, _07475_, _07474_);
  not _58483_ (_07477_, _06403_);
  and _58484_ (_07478_, _07067_, _07477_);
  and _58485_ (_07479_, _06360_, _05652_);
  nor _58486_ (_07480_, _07356_, \oc8051_golden_model_1.SP [2]);
  nor _58487_ (_07481_, _07480_, _07357_);
  and _58488_ (_07482_, _07481_, _05732_);
  and _58489_ (_07483_, _07477_, _06021_);
  nor _58490_ (_07484_, _07481_, _05686_);
  and _58491_ (_07485_, _06976_, _07477_);
  nand _58492_ (_07486_, _06881_, \oc8051_golden_model_1.IRAM[0] [2]);
  nand _58493_ (_07487_, _06726_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _58494_ (_07488_, _07487_, _06879_);
  nand _58495_ (_07489_, _07488_, _07486_);
  nand _58496_ (_07490_, _06726_, \oc8051_golden_model_1.IRAM[3] [2]);
  nand _58497_ (_07491_, _06881_, \oc8051_golden_model_1.IRAM[2] [2]);
  and _58498_ (_07492_, _07491_, _06887_);
  nand _58499_ (_07493_, _07492_, _07490_);
  nand _58500_ (_07494_, _07493_, _07489_);
  nand _58501_ (_07495_, _07494_, _06504_);
  nand _58502_ (_07496_, _06726_, \oc8051_golden_model_1.IRAM[7] [2]);
  nand _58503_ (_07497_, _06881_, \oc8051_golden_model_1.IRAM[6] [2]);
  and _58504_ (_07498_, _07497_, _06887_);
  nand _58505_ (_07499_, _07498_, _07496_);
  nand _58506_ (_07500_, _06881_, \oc8051_golden_model_1.IRAM[4] [2]);
  nand _58507_ (_07501_, _06726_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _58508_ (_07502_, _07501_, _06879_);
  nand _58509_ (_07503_, _07502_, _07500_);
  nand _58510_ (_07504_, _07503_, _07499_);
  nand _58511_ (_07505_, _07504_, _06894_);
  nand _58512_ (_07506_, _07505_, _07495_);
  nand _58513_ (_07507_, _07506_, _06328_);
  nand _58514_ (_07508_, _06726_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand _58515_ (_07509_, _06881_, \oc8051_golden_model_1.IRAM[10] [2]);
  and _58516_ (_07510_, _07509_, _06887_);
  nand _58517_ (_07511_, _07510_, _07508_);
  nand _58518_ (_07512_, _06881_, \oc8051_golden_model_1.IRAM[8] [2]);
  nand _58519_ (_07513_, _06726_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _58520_ (_07514_, _07513_, _06879_);
  nand _58521_ (_07515_, _07514_, _07512_);
  nand _58522_ (_07516_, _07515_, _07511_);
  nand _58523_ (_07517_, _07516_, _06504_);
  nand _58524_ (_07518_, _06726_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand _58525_ (_07519_, _06881_, \oc8051_golden_model_1.IRAM[14] [2]);
  and _58526_ (_07520_, _07519_, _06887_);
  nand _58527_ (_07521_, _07520_, _07518_);
  nand _58528_ (_07522_, _06881_, \oc8051_golden_model_1.IRAM[12] [2]);
  nand _58529_ (_07523_, _06726_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _58530_ (_07524_, _07523_, _06879_);
  nand _58531_ (_07525_, _07524_, _07522_);
  nand _58532_ (_07526_, _07525_, _07521_);
  nand _58533_ (_07527_, _07526_, _06894_);
  nand _58534_ (_07528_, _07527_, _07517_);
  nand _58535_ (_07529_, _07528_, _06908_);
  nand _58536_ (_07530_, _07529_, _07507_);
  or _58537_ (_07531_, _07530_, _05670_);
  and _58538_ (_07532_, _07531_, _07247_);
  and _58539_ (_07533_, _06940_, _06403_);
  nor _58540_ (_07534_, _07533_, _07532_);
  not _58541_ (_07535_, _07481_);
  and _58542_ (_07536_, _07535_, _06943_);
  and _58543_ (_07537_, _06095_, _06042_);
  nor _58544_ (_07538_, _07537_, _07536_);
  and _58545_ (_07539_, _07538_, _07534_);
  and _58546_ (_07540_, _07530_, _06948_);
  nor _58547_ (_07541_, _07540_, _06955_);
  and _58548_ (_07542_, _07541_, _07539_);
  and _58549_ (_07543_, _06955_, _07477_);
  nor _58550_ (_07544_, _07543_, _07542_);
  and _58551_ (_07545_, _06953_, _06359_);
  nor _58552_ (_07546_, _07545_, _07544_);
  or _58553_ (_07547_, _07481_, _05690_);
  nand _58554_ (_07548_, _07547_, _07546_);
  and _58555_ (_07549_, _06095_, _06037_);
  and _58556_ (_07550_, _06963_, _06403_);
  nor _58557_ (_07551_, _07550_, _07549_);
  not _58558_ (_07552_, _07551_);
  nor _58559_ (_07553_, _07552_, _07548_);
  and _58560_ (_07554_, _07530_, _06970_);
  nor _58561_ (_07555_, _07554_, _06976_);
  and _58562_ (_07556_, _07555_, _07553_);
  nor _58563_ (_07557_, _07556_, _07485_);
  nor _58564_ (_07558_, _07557_, _06975_);
  nor _58565_ (_07559_, _07558_, _06371_);
  nor _58566_ (_07560_, _07559_, _06038_);
  and _58567_ (_07561_, _07481_, _06038_);
  nor _58568_ (_07562_, _07561_, _07560_);
  and _58569_ (_07563_, _06035_, _06359_);
  nor _58570_ (_07564_, _07563_, _07562_);
  nand _58571_ (_07565_, _07564_, _06232_);
  nor _58572_ (_07566_, _07565_, _07484_);
  and _58573_ (_07567_, _07530_, _06992_);
  not _58574_ (_07568_, _07567_);
  and _58575_ (_07569_, _07568_, _07566_);
  and _58576_ (_07570_, _06991_, _06359_);
  nor _58577_ (_07571_, _07570_, _06023_);
  and _58578_ (_07572_, _07571_, _07569_);
  nor _58579_ (_07573_, _07535_, _05673_);
  nor _58580_ (_07574_, _07573_, _07572_);
  nor _58581_ (_07575_, _07015_, _07477_);
  nor _58582_ (_07576_, _07575_, _07252_);
  not _58583_ (_07577_, _07576_);
  nor _58584_ (_07578_, _07577_, _07574_);
  and _58585_ (_07579_, _07530_, _07023_);
  nor _58586_ (_07580_, _07579_, _06021_);
  and _58587_ (_07581_, _07580_, _07578_);
  nor _58588_ (_07582_, _07581_, _07483_);
  nor _58589_ (_07583_, _07582_, _05724_);
  and _58590_ (_07584_, _07481_, _05724_);
  nor _58591_ (_07585_, _07584_, _07583_);
  nor _58592_ (_07586_, _07035_, _07477_);
  nor _58593_ (_07587_, _07586_, _05736_);
  not _58594_ (_07588_, _07587_);
  nor _58595_ (_07589_, _07588_, _07585_);
  and _58596_ (_07590_, _07481_, _05736_);
  nor _58597_ (_07591_, _07590_, _07589_);
  and _58598_ (_07592_, _07042_, _06403_);
  nor _58599_ (_07593_, _07592_, _05732_);
  not _58600_ (_07594_, _07593_);
  nor _58601_ (_07595_, _07594_, _07591_);
  nor _58602_ (_07596_, _07595_, _07482_);
  and _58603_ (_07597_, _06095_, _05495_);
  nor _58604_ (_07598_, _07597_, _07596_);
  and _58605_ (_07599_, _07530_, _07051_);
  nor _58606_ (_07600_, _07599_, _07050_);
  and _58607_ (_07601_, _07600_, _07598_);
  and _58608_ (_07602_, _07050_, _07477_);
  nor _58609_ (_07603_, _07602_, _07601_);
  nor _58610_ (_07604_, _07481_, _07059_);
  nor _58611_ (_07605_, _07604_, _07058_);
  not _58612_ (_07606_, _07605_);
  nor _58613_ (_07607_, _07606_, _07603_);
  nor _58614_ (_07608_, _07607_, _07479_);
  and _58615_ (_07609_, _06095_, _05750_);
  nor _58616_ (_07610_, _07609_, _07608_);
  and _58617_ (_07611_, _07530_, _07068_);
  nor _58618_ (_07612_, _07611_, _07067_);
  and _58619_ (_07613_, _07612_, _07610_);
  nor _58620_ (_07614_, _07613_, _07478_);
  nor _58621_ (_07615_, _07614_, _07305_);
  not _58622_ (_07616_, _07615_);
  nor _58623_ (_07617_, _07616_, _07476_);
  and _58624_ (_07618_, _07617_, _07307_);
  or _58625_ (_07619_, _07618_, \oc8051_golden_model_1.IRAM[15] [7]);
  and _58626_ (_07620_, _07359_, _06029_);
  nor _58627_ (_07621_, _07481_, _07081_);
  nor _58628_ (_07622_, _07621_, _07620_);
  and _58629_ (_07623_, _07360_, _06029_);
  nor _58630_ (_07624_, _07620_, _07362_);
  nor _58631_ (_07625_, _07624_, _07623_);
  and _58632_ (_07626_, _07234_, _07235_);
  and _58633_ (_07627_, _07626_, _07274_);
  nor _58634_ (_07628_, _07627_, _07230_);
  and _58635_ (_07629_, _07628_, _07625_);
  and _58636_ (_07630_, _07629_, _07622_);
  and _58637_ (_07631_, _07630_, _07080_);
  not _58638_ (_07632_, _07631_);
  and _58639_ (_07633_, _07632_, _07619_);
  not _58640_ (_07634_, _07618_);
  and _58641_ (_07635_, _06084_, _05952_);
  and _58642_ (_07636_, _07635_, _06359_);
  and _58643_ (_07637_, _07636_, _06758_);
  and _58644_ (_07638_, _07637_, _05983_);
  nor _58645_ (_07639_, _06799_, _06016_);
  and _58646_ (_07640_, _07639_, _07477_);
  and _58647_ (_07641_, _07640_, _07638_);
  and _58648_ (_07642_, _07641_, \oc8051_golden_model_1.PCON [7]);
  not _58649_ (_07643_, _07642_);
  and _58650_ (_07644_, _06799_, _06016_);
  not _58651_ (_07645_, _07644_);
  nand _58652_ (_07646_, _06403_, _06299_);
  nor _58653_ (_07647_, _07646_, _07645_);
  and _58654_ (_07648_, _07647_, _07637_);
  and _58655_ (_07649_, _07648_, \oc8051_golden_model_1.TCON [7]);
  and _58656_ (_07650_, _06799_, _06017_);
  not _58657_ (_07651_, _07650_);
  nor _58658_ (_07652_, _07651_, _07646_);
  and _58659_ (_07653_, _07652_, _07637_);
  and _58660_ (_07654_, _07653_, \oc8051_golden_model_1.TMOD [7]);
  not _58661_ (_07655_, _07637_);
  nor _58662_ (_07656_, _06799_, _06017_);
  not _58663_ (_07657_, _07656_);
  or _58664_ (_07658_, _07657_, _07646_);
  nor _58665_ (_07659_, _07658_, _07655_);
  and _58666_ (_07660_, _07659_, \oc8051_golden_model_1.TL0 [7]);
  or _58667_ (_07661_, _06403_, _05983_);
  or _58668_ (_07662_, _07661_, _07645_);
  nor _58669_ (_07663_, _07662_, _07655_);
  and _58670_ (_07664_, _07663_, \oc8051_golden_model_1.TH0 [7]);
  not _58671_ (_07665_, _07639_);
  or _58672_ (_07666_, _07665_, _07646_);
  nor _58673_ (_07667_, _07666_, _07655_);
  and _58674_ (_07668_, _07667_, \oc8051_golden_model_1.TL1 [7]);
  or _58675_ (_07669_, _07661_, _07651_);
  nor _58676_ (_07670_, _07669_, _07655_);
  and _58677_ (_07671_, _07670_, \oc8051_golden_model_1.TH1 [7]);
  nand _58678_ (_07672_, _06403_, _05983_);
  nor _58679_ (_07673_, _07672_, _07645_);
  not _58680_ (_07674_, _06758_);
  and _58681_ (_07675_, _07674_, _06359_);
  and _58682_ (_07676_, _07675_, _07635_);
  and _58683_ (_07677_, _07676_, _07673_);
  and _58684_ (_07678_, _07677_, \oc8051_golden_model_1.P1 [7]);
  and _58685_ (_07679_, _07676_, _07647_);
  and _58686_ (_07680_, _07679_, \oc8051_golden_model_1.SCON [7]);
  and _58687_ (_07681_, _07652_, _07676_);
  and _58688_ (_07682_, _07681_, \oc8051_golden_model_1.SBUF [7]);
  not _58689_ (_07683_, _06359_);
  and _58690_ (_07684_, _06758_, _07683_);
  and _58691_ (_07685_, _07635_, _07684_);
  and _58692_ (_07686_, _07685_, _07673_);
  and _58693_ (_07687_, _07686_, \oc8051_golden_model_1.P2 [7]);
  and _58694_ (_07688_, _07647_, _07685_);
  and _58695_ (_07689_, _07688_, \oc8051_golden_model_1.IE [7]);
  nor _58696_ (_07690_, _06758_, _06359_);
  and _58697_ (_07691_, _07635_, _07690_);
  and _58698_ (_07692_, _07691_, _07673_);
  and _58699_ (_07693_, _07692_, \oc8051_golden_model_1.P3 [7]);
  and _58700_ (_07694_, _07647_, _07691_);
  and _58701_ (_07695_, _07694_, \oc8051_golden_model_1.IP [7]);
  nor _58702_ (_07696_, _06084_, _06053_);
  and _58703_ (_07697_, _07696_, _07690_);
  and _58704_ (_07698_, _07697_, _07673_);
  and _58705_ (_07699_, _07698_, \oc8051_golden_model_1.B [7]);
  and _58706_ (_07700_, _07684_, _07696_);
  and _58707_ (_07701_, _07700_, _07673_);
  and _58708_ (_07702_, _07701_, \oc8051_golden_model_1.ACC [7]);
  nor _58709_ (_07703_, _07702_, _07699_);
  and _58710_ (_07704_, _07675_, _07696_);
  and _58711_ (_07705_, _07704_, _07673_);
  and _58712_ (_07706_, _07705_, \oc8051_golden_model_1.PSW [7]);
  not _58713_ (_07707_, _07706_);
  nand _58714_ (_07708_, _07707_, _07703_);
  or _58715_ (_07709_, _07708_, _07695_);
  or _58716_ (_07710_, _07709_, _07693_);
  or _58717_ (_07711_, _07710_, _07689_);
  or _58718_ (_07712_, _07711_, _07687_);
  or _58719_ (_07713_, _07712_, _07682_);
  or _58720_ (_07714_, _07713_, _07680_);
  or _58721_ (_07715_, _07714_, _07678_);
  or _58722_ (_07716_, _07715_, _07671_);
  or _58723_ (_07717_, _07716_, _07668_);
  or _58724_ (_07718_, _07717_, _07664_);
  or _58725_ (_07719_, _07718_, _07660_);
  or _58726_ (_07720_, _07719_, _07654_);
  nor _58727_ (_07721_, _07720_, _07649_);
  and _58728_ (_07722_, _07721_, _07643_);
  and _58729_ (_07723_, _07639_, _06403_);
  and _58730_ (_07724_, _07723_, _07638_);
  and _58731_ (_07725_, _07724_, \oc8051_golden_model_1.DPH [7]);
  and _58732_ (_07726_, _07650_, _06403_);
  and _58733_ (_07727_, _07726_, _07638_);
  and _58734_ (_07728_, _07727_, \oc8051_golden_model_1.SP [7]);
  nor _58735_ (_07729_, _07728_, _07725_);
  and _58736_ (_07730_, _07637_, _07673_);
  and _58737_ (_07731_, _07730_, \oc8051_golden_model_1.P0 [7]);
  and _58738_ (_07732_, _07656_, _06403_);
  and _58739_ (_07733_, _07732_, _07638_);
  and _58740_ (_07734_, _07733_, \oc8051_golden_model_1.DPL [7]);
  nor _58741_ (_07735_, _07734_, _07731_);
  and _58742_ (_07736_, _07735_, _07729_);
  and _58743_ (_07737_, _07736_, _07722_);
  not _58744_ (_07738_, \oc8051_golden_model_1.IRAM[0] [7]);
  or _58745_ (_07739_, _06726_, _07738_);
  not _58746_ (_07740_, \oc8051_golden_model_1.IRAM[1] [7]);
  or _58747_ (_07741_, _06881_, _07740_);
  and _58748_ (_07742_, _07741_, _06879_);
  nand _58749_ (_07743_, _07742_, _07739_);
  nand _58750_ (_07744_, _06726_, \oc8051_golden_model_1.IRAM[3] [7]);
  nand _58751_ (_07745_, _06881_, \oc8051_golden_model_1.IRAM[2] [7]);
  and _58752_ (_07746_, _07745_, _06887_);
  nand _58753_ (_07747_, _07746_, _07744_);
  nand _58754_ (_07748_, _07747_, _07743_);
  nand _58755_ (_07749_, _07748_, _06504_);
  nand _58756_ (_07750_, _06726_, \oc8051_golden_model_1.IRAM[7] [7]);
  not _58757_ (_07751_, \oc8051_golden_model_1.IRAM[6] [7]);
  or _58758_ (_07752_, _06726_, _07751_);
  and _58759_ (_07753_, _07752_, _06887_);
  nand _58760_ (_07754_, _07753_, _07750_);
  nand _58761_ (_07755_, _06881_, \oc8051_golden_model_1.IRAM[4] [7]);
  nand _58762_ (_07756_, _06726_, \oc8051_golden_model_1.IRAM[5] [7]);
  and _58763_ (_07757_, _07756_, _06879_);
  nand _58764_ (_07758_, _07757_, _07755_);
  nand _58765_ (_07759_, _07758_, _07754_);
  nand _58766_ (_07760_, _07759_, _06894_);
  nand _58767_ (_07761_, _07760_, _07749_);
  nand _58768_ (_07762_, _07761_, _06328_);
  nand _58769_ (_07763_, _06726_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand _58770_ (_07764_, _06881_, \oc8051_golden_model_1.IRAM[10] [7]);
  and _58771_ (_07765_, _07764_, _06887_);
  nand _58772_ (_07766_, _07765_, _07763_);
  nand _58773_ (_07767_, _06881_, \oc8051_golden_model_1.IRAM[8] [7]);
  nand _58774_ (_07768_, _06726_, \oc8051_golden_model_1.IRAM[9] [7]);
  and _58775_ (_07769_, _07768_, _06879_);
  nand _58776_ (_07770_, _07769_, _07767_);
  nand _58777_ (_07771_, _07770_, _07766_);
  nand _58778_ (_07772_, _07771_, _06504_);
  nand _58779_ (_07773_, _06726_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand _58780_ (_07774_, _06881_, \oc8051_golden_model_1.IRAM[14] [7]);
  and _58781_ (_07775_, _07774_, _06887_);
  nand _58782_ (_07776_, _07775_, _07773_);
  nand _58783_ (_07777_, _06881_, \oc8051_golden_model_1.IRAM[12] [7]);
  nand _58784_ (_07778_, _06726_, \oc8051_golden_model_1.IRAM[13] [7]);
  and _58785_ (_07779_, _07778_, _06879_);
  nand _58786_ (_07780_, _07779_, _07777_);
  nand _58787_ (_07781_, _07780_, _07776_);
  nand _58788_ (_07782_, _07781_, _06894_);
  nand _58789_ (_07783_, _07782_, _07772_);
  nand _58790_ (_07784_, _07783_, _06908_);
  nand _58791_ (_07785_, _07784_, _07762_);
  or _58792_ (_07786_, _07785_, _05952_);
  and _58793_ (_07787_, _07786_, _07737_);
  not _58794_ (_07788_, _07787_);
  and _58795_ (_07789_, _07686_, \oc8051_golden_model_1.P2 [6]);
  not _58796_ (_07790_, _07789_);
  and _58797_ (_07791_, _07681_, \oc8051_golden_model_1.SBUF [6]);
  not _58798_ (_07792_, _07791_);
  and _58799_ (_07793_, _07688_, \oc8051_golden_model_1.IE [6]);
  and _58800_ (_07794_, _07692_, \oc8051_golden_model_1.P3 [6]);
  nor _58801_ (_07795_, _07794_, _07793_);
  and _58802_ (_07796_, _07795_, _07792_);
  and _58803_ (_07797_, _07796_, _07790_);
  and _58804_ (_07798_, _07730_, \oc8051_golden_model_1.P0 [6]);
  not _58805_ (_07799_, _07798_);
  and _58806_ (_07800_, _07733_, \oc8051_golden_model_1.DPL [6]);
  nor _58807_ (_07801_, _07665_, _07672_);
  and _58808_ (_07802_, _07801_, _07637_);
  and _58809_ (_07803_, _07802_, \oc8051_golden_model_1.DPH [6]);
  nor _58810_ (_07804_, _07803_, _07800_);
  and _58811_ (_07805_, _07804_, _07799_);
  and _58812_ (_07806_, _07667_, \oc8051_golden_model_1.TL1 [6]);
  and _58813_ (_07807_, _07670_, \oc8051_golden_model_1.TH1 [6]);
  nor _58814_ (_07808_, _07807_, _07806_);
  and _58815_ (_07809_, _07679_, \oc8051_golden_model_1.SCON [6]);
  and _58816_ (_07810_, _07677_, \oc8051_golden_model_1.P1 [6]);
  nor _58817_ (_07811_, _07810_, _07809_);
  and _58818_ (_07812_, _07811_, _07808_);
  and _58819_ (_07813_, _07812_, _07805_);
  and _58820_ (_07814_, _07813_, _07797_);
  and _58821_ (_07815_, _07694_, \oc8051_golden_model_1.IP [6]);
  not _58822_ (_07816_, _07815_);
  and _58823_ (_07817_, _07698_, \oc8051_golden_model_1.B [6]);
  and _58824_ (_07818_, _07701_, \oc8051_golden_model_1.ACC [6]);
  nor _58825_ (_07819_, _07818_, _07817_);
  and _58826_ (_07820_, _07819_, _07816_);
  and _58827_ (_07821_, _07641_, \oc8051_golden_model_1.PCON [6]);
  and _58828_ (_07822_, _07705_, \oc8051_golden_model_1.PSW [6]);
  nor _58829_ (_07823_, _07822_, _07821_);
  and _58830_ (_07824_, _07823_, _07820_);
  and _58831_ (_07825_, _07653_, \oc8051_golden_model_1.TMOD [6]);
  not _58832_ (_07826_, _07825_);
  and _58833_ (_07827_, _07659_, \oc8051_golden_model_1.TL0 [6]);
  and _58834_ (_07828_, _07663_, \oc8051_golden_model_1.TH0 [6]);
  nor _58835_ (_07829_, _07828_, _07827_);
  and _58836_ (_07830_, _07829_, _07826_);
  and _58837_ (_07831_, _07648_, \oc8051_golden_model_1.TCON [6]);
  or _58838_ (_07832_, _07651_, _07672_);
  nor _58839_ (_07833_, _07832_, _07655_);
  and _58840_ (_07834_, _07833_, \oc8051_golden_model_1.SP [6]);
  nor _58841_ (_07835_, _07834_, _07831_);
  and _58842_ (_07836_, _07835_, _07830_);
  and _58843_ (_07837_, _07836_, _07824_);
  and _58844_ (_07838_, _07837_, _07814_);
  nand _58845_ (_07839_, _06881_, \oc8051_golden_model_1.IRAM[0] [6]);
  nand _58846_ (_07840_, _06726_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _58847_ (_07841_, _07840_, _06879_);
  nand _58848_ (_07842_, _07841_, _07839_);
  nand _58849_ (_07843_, _06726_, \oc8051_golden_model_1.IRAM[3] [6]);
  nand _58850_ (_07844_, _06881_, \oc8051_golden_model_1.IRAM[2] [6]);
  and _58851_ (_07845_, _07844_, _06887_);
  nand _58852_ (_07846_, _07845_, _07843_);
  nand _58853_ (_07847_, _07846_, _07842_);
  nand _58854_ (_07848_, _07847_, _06504_);
  nand _58855_ (_07849_, _06726_, \oc8051_golden_model_1.IRAM[7] [6]);
  nand _58856_ (_07850_, _06881_, \oc8051_golden_model_1.IRAM[6] [6]);
  and _58857_ (_07851_, _07850_, _06887_);
  nand _58858_ (_07852_, _07851_, _07849_);
  nand _58859_ (_07853_, _06881_, \oc8051_golden_model_1.IRAM[4] [6]);
  nand _58860_ (_07854_, _06726_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _58861_ (_07855_, _07854_, _06879_);
  nand _58862_ (_07856_, _07855_, _07853_);
  nand _58863_ (_07857_, _07856_, _07852_);
  nand _58864_ (_07858_, _07857_, _06894_);
  nand _58865_ (_07859_, _07858_, _07848_);
  nand _58866_ (_07860_, _07859_, _06328_);
  nand _58867_ (_07861_, _06726_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _58868_ (_07862_, _06881_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _58869_ (_07863_, _07862_, _06887_);
  nand _58870_ (_07864_, _07863_, _07861_);
  nand _58871_ (_07865_, _06881_, \oc8051_golden_model_1.IRAM[8] [6]);
  nand _58872_ (_07866_, _06726_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _58873_ (_07867_, _07866_, _06879_);
  nand _58874_ (_07868_, _07867_, _07865_);
  nand _58875_ (_07869_, _07868_, _07864_);
  nand _58876_ (_07870_, _07869_, _06504_);
  nand _58877_ (_07871_, _06726_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _58878_ (_07872_, _06881_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _58879_ (_07873_, _07872_, _06887_);
  nand _58880_ (_07874_, _07873_, _07871_);
  nand _58881_ (_07875_, _06881_, \oc8051_golden_model_1.IRAM[12] [6]);
  nand _58882_ (_07876_, _06726_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _58883_ (_07877_, _07876_, _06879_);
  nand _58884_ (_07878_, _07877_, _07875_);
  nand _58885_ (_07879_, _07878_, _07874_);
  nand _58886_ (_07880_, _07879_, _06894_);
  nand _58887_ (_07881_, _07880_, _07870_);
  nand _58888_ (_07882_, _07881_, _06908_);
  nand _58889_ (_07883_, _07882_, _07860_);
  or _58890_ (_07884_, _07883_, _05952_);
  and _58891_ (_07885_, _07884_, _07838_);
  not _58892_ (_07886_, _07885_);
  and _58893_ (_07887_, _07686_, \oc8051_golden_model_1.P2 [5]);
  not _58894_ (_07888_, _07887_);
  and _58895_ (_07889_, _07681_, \oc8051_golden_model_1.SBUF [5]);
  not _58896_ (_07890_, _07889_);
  and _58897_ (_07891_, _07688_, \oc8051_golden_model_1.IE [5]);
  and _58898_ (_07892_, _07692_, \oc8051_golden_model_1.P3 [5]);
  nor _58899_ (_07893_, _07892_, _07891_);
  and _58900_ (_07894_, _07893_, _07890_);
  and _58901_ (_07895_, _07894_, _07888_);
  and _58902_ (_07896_, _07667_, \oc8051_golden_model_1.TL1 [5]);
  and _58903_ (_07897_, _07670_, \oc8051_golden_model_1.TH1 [5]);
  nor _58904_ (_07898_, _07897_, _07896_);
  and _58905_ (_07899_, _07679_, \oc8051_golden_model_1.SCON [5]);
  and _58906_ (_07900_, _07677_, \oc8051_golden_model_1.P1 [5]);
  nor _58907_ (_07901_, _07900_, _07899_);
  and _58908_ (_07902_, _07901_, _07898_);
  and _58909_ (_07903_, _07902_, _07895_);
  and _58910_ (_07904_, _07694_, \oc8051_golden_model_1.IP [5]);
  not _58911_ (_07905_, _07904_);
  and _58912_ (_07906_, _07698_, \oc8051_golden_model_1.B [5]);
  and _58913_ (_07907_, _07701_, \oc8051_golden_model_1.ACC [5]);
  nor _58914_ (_07908_, _07907_, _07906_);
  and _58915_ (_07909_, _07908_, _07905_);
  and _58916_ (_07910_, _07641_, \oc8051_golden_model_1.PCON [5]);
  and _58917_ (_07911_, _07705_, \oc8051_golden_model_1.PSW [5]);
  nor _58918_ (_07912_, _07911_, _07910_);
  and _58919_ (_07913_, _07912_, _07909_);
  and _58920_ (_07914_, _07648_, \oc8051_golden_model_1.TCON [5]);
  not _58921_ (_07915_, _07914_);
  and _58922_ (_07916_, _07663_, \oc8051_golden_model_1.TH0 [5]);
  and _58923_ (_07917_, _07659_, \oc8051_golden_model_1.TL0 [5]);
  nor _58924_ (_07918_, _07917_, _07916_);
  and _58925_ (_07919_, _07918_, _07915_);
  and _58926_ (_07920_, _07653_, \oc8051_golden_model_1.TMOD [5]);
  not _58927_ (_07921_, _07920_);
  and _58928_ (_07922_, _07733_, \oc8051_golden_model_1.DPL [5]);
  and _58929_ (_07923_, _07802_, \oc8051_golden_model_1.DPH [5]);
  nor _58930_ (_07924_, _07923_, _07922_);
  and _58931_ (_07925_, _07730_, \oc8051_golden_model_1.P0 [5]);
  and _58932_ (_07926_, _07833_, \oc8051_golden_model_1.SP [5]);
  nor _58933_ (_07927_, _07926_, _07925_);
  and _58934_ (_07928_, _07927_, _07924_);
  and _58935_ (_07929_, _07928_, _07921_);
  and _58936_ (_07930_, _07929_, _07919_);
  and _58937_ (_07931_, _07930_, _07913_);
  and _58938_ (_07932_, _07931_, _07903_);
  nand _58939_ (_07933_, _06881_, \oc8051_golden_model_1.IRAM[0] [5]);
  nand _58940_ (_07934_, _06726_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _58941_ (_07935_, _07934_, _06879_);
  nand _58942_ (_07936_, _07935_, _07933_);
  nand _58943_ (_07937_, _06726_, \oc8051_golden_model_1.IRAM[3] [5]);
  nand _58944_ (_07938_, _06881_, \oc8051_golden_model_1.IRAM[2] [5]);
  and _58945_ (_07939_, _07938_, _06887_);
  nand _58946_ (_07940_, _07939_, _07937_);
  nand _58947_ (_07941_, _07940_, _07936_);
  nand _58948_ (_07942_, _07941_, _06504_);
  nand _58949_ (_07943_, _06726_, \oc8051_golden_model_1.IRAM[7] [5]);
  nand _58950_ (_07944_, _06881_, \oc8051_golden_model_1.IRAM[6] [5]);
  and _58951_ (_07945_, _07944_, _06887_);
  nand _58952_ (_07946_, _07945_, _07943_);
  nand _58953_ (_07947_, _06881_, \oc8051_golden_model_1.IRAM[4] [5]);
  nand _58954_ (_07948_, _06726_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _58955_ (_07949_, _07948_, _06879_);
  nand _58956_ (_07950_, _07949_, _07947_);
  nand _58957_ (_07951_, _07950_, _07946_);
  nand _58958_ (_07952_, _07951_, _06894_);
  nand _58959_ (_07953_, _07952_, _07942_);
  nand _58960_ (_07954_, _07953_, _06328_);
  nand _58961_ (_07955_, _06726_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand _58962_ (_07956_, _06881_, \oc8051_golden_model_1.IRAM[10] [5]);
  and _58963_ (_07957_, _07956_, _06887_);
  nand _58964_ (_07958_, _07957_, _07955_);
  nand _58965_ (_07959_, _06881_, \oc8051_golden_model_1.IRAM[8] [5]);
  nand _58966_ (_07960_, _06726_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _58967_ (_07961_, _07960_, _06879_);
  nand _58968_ (_07962_, _07961_, _07959_);
  nand _58969_ (_07963_, _07962_, _07958_);
  nand _58970_ (_07964_, _07963_, _06504_);
  nand _58971_ (_07965_, _06726_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand _58972_ (_07966_, _06881_, \oc8051_golden_model_1.IRAM[14] [5]);
  and _58973_ (_07967_, _07966_, _06887_);
  nand _58974_ (_07968_, _07967_, _07965_);
  nand _58975_ (_07969_, _06881_, \oc8051_golden_model_1.IRAM[12] [5]);
  nand _58976_ (_07970_, _06726_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _58977_ (_07971_, _07970_, _06879_);
  nand _58978_ (_07972_, _07971_, _07969_);
  nand _58979_ (_07973_, _07972_, _07968_);
  nand _58980_ (_07974_, _07973_, _06894_);
  nand _58981_ (_07975_, _07974_, _07964_);
  nand _58982_ (_07976_, _07975_, _06908_);
  nand _58983_ (_07977_, _07976_, _07954_);
  or _58984_ (_07978_, _07977_, _05952_);
  and _58985_ (_07979_, _07978_, _07932_);
  not _58986_ (_07980_, _07979_);
  and _58987_ (_07981_, _07667_, \oc8051_golden_model_1.TL1 [3]);
  not _58988_ (_07982_, _07981_);
  and _58989_ (_07983_, _07677_, \oc8051_golden_model_1.P1 [3]);
  and _58990_ (_07984_, _07679_, \oc8051_golden_model_1.SCON [3]);
  nor _58991_ (_07985_, _07984_, _07983_);
  and _58992_ (_07986_, _07985_, _07982_);
  and _58993_ (_07987_, _07681_, \oc8051_golden_model_1.SBUF [3]);
  not _58994_ (_07988_, _07987_);
  and _58995_ (_07989_, _07692_, \oc8051_golden_model_1.P3 [3]);
  and _58996_ (_07990_, _07688_, \oc8051_golden_model_1.IE [3]);
  nor _58997_ (_07991_, _07990_, _07989_);
  and _58998_ (_07992_, _07991_, _07988_);
  and _58999_ (_07993_, _07686_, \oc8051_golden_model_1.P2 [3]);
  and _59000_ (_07994_, _07670_, \oc8051_golden_model_1.TH1 [3]);
  nor _59001_ (_07995_, _07994_, _07993_);
  and _59002_ (_07996_, _07995_, _07992_);
  and _59003_ (_07997_, _07996_, _07986_);
  and _59004_ (_07998_, _07694_, \oc8051_golden_model_1.IP [3]);
  not _59005_ (_07999_, _07998_);
  and _59006_ (_08000_, _07701_, \oc8051_golden_model_1.ACC [3]);
  and _59007_ (_08001_, _07698_, \oc8051_golden_model_1.B [3]);
  nor _59008_ (_08002_, _08001_, _08000_);
  and _59009_ (_08003_, _08002_, _07999_);
  and _59010_ (_08004_, _07641_, \oc8051_golden_model_1.PCON [3]);
  and _59011_ (_08005_, _07705_, \oc8051_golden_model_1.PSW [3]);
  nor _59012_ (_08006_, _08005_, _08004_);
  and _59013_ (_08007_, _08006_, _08003_);
  and _59014_ (_08008_, _07653_, \oc8051_golden_model_1.TMOD [3]);
  not _59015_ (_08009_, _08008_);
  and _59016_ (_08010_, _07663_, \oc8051_golden_model_1.TH0 [3]);
  and _59017_ (_08011_, _07659_, \oc8051_golden_model_1.TL0 [3]);
  nor _59018_ (_08012_, _08011_, _08010_);
  and _59019_ (_08013_, _08012_, _08009_);
  and _59020_ (_08014_, _07648_, \oc8051_golden_model_1.TCON [3]);
  not _59021_ (_08015_, _08014_);
  and _59022_ (_08016_, _07733_, \oc8051_golden_model_1.DPL [3]);
  and _59023_ (_08017_, _07802_, \oc8051_golden_model_1.DPH [3]);
  nor _59024_ (_08018_, _08017_, _08016_);
  and _59025_ (_08019_, _07730_, \oc8051_golden_model_1.P0 [3]);
  and _59026_ (_08020_, _07833_, \oc8051_golden_model_1.SP [3]);
  nor _59027_ (_08021_, _08020_, _08019_);
  and _59028_ (_08022_, _08021_, _08018_);
  and _59029_ (_08023_, _08022_, _08015_);
  and _59030_ (_08024_, _08023_, _08013_);
  and _59031_ (_08025_, _08024_, _08007_);
  and _59032_ (_08026_, _08025_, _07997_);
  or _59033_ (_08027_, _07353_, _05952_);
  and _59034_ (_08028_, _08027_, _08026_);
  not _59035_ (_08029_, _08028_);
  and _59036_ (_08030_, _07670_, \oc8051_golden_model_1.TH1 [1]);
  not _59037_ (_08031_, _08030_);
  and _59038_ (_08032_, _07679_, \oc8051_golden_model_1.SCON [1]);
  and _59039_ (_08033_, _07677_, \oc8051_golden_model_1.P1 [1]);
  nor _59040_ (_08034_, _08033_, _08032_);
  and _59041_ (_08035_, _08034_, _08031_);
  and _59042_ (_08036_, _07681_, \oc8051_golden_model_1.SBUF [1]);
  not _59043_ (_08037_, _08036_);
  and _59044_ (_08038_, _07692_, \oc8051_golden_model_1.P3 [1]);
  and _59045_ (_08039_, _07688_, \oc8051_golden_model_1.IE [1]);
  nor _59046_ (_08040_, _08039_, _08038_);
  and _59047_ (_08041_, _08040_, _08037_);
  and _59048_ (_08042_, _07686_, \oc8051_golden_model_1.P2 [1]);
  and _59049_ (_08043_, _07667_, \oc8051_golden_model_1.TL1 [1]);
  nor _59050_ (_08044_, _08043_, _08042_);
  and _59051_ (_08045_, _08044_, _08041_);
  and _59052_ (_08046_, _08045_, _08035_);
  and _59053_ (_08047_, _07694_, \oc8051_golden_model_1.IP [1]);
  not _59054_ (_08048_, _08047_);
  and _59055_ (_08049_, _07701_, \oc8051_golden_model_1.ACC [1]);
  and _59056_ (_08050_, _07698_, \oc8051_golden_model_1.B [1]);
  nor _59057_ (_08051_, _08050_, _08049_);
  and _59058_ (_08052_, _08051_, _08048_);
  and _59059_ (_08053_, _07641_, \oc8051_golden_model_1.PCON [1]);
  and _59060_ (_08054_, _07705_, \oc8051_golden_model_1.PSW [1]);
  nor _59061_ (_08055_, _08054_, _08053_);
  and _59062_ (_08056_, _08055_, _08052_);
  and _59063_ (_08057_, _07653_, \oc8051_golden_model_1.TMOD [1]);
  not _59064_ (_08058_, _08057_);
  and _59065_ (_08059_, _07659_, \oc8051_golden_model_1.TL0 [1]);
  and _59066_ (_08060_, _07663_, \oc8051_golden_model_1.TH0 [1]);
  nor _59067_ (_08061_, _08060_, _08059_);
  and _59068_ (_08062_, _08061_, _08058_);
  and _59069_ (_08063_, _07648_, \oc8051_golden_model_1.TCON [1]);
  not _59070_ (_08064_, _08063_);
  and _59071_ (_08065_, _07730_, \oc8051_golden_model_1.P0 [1]);
  and _59072_ (_08066_, _07833_, \oc8051_golden_model_1.SP [1]);
  nor _59073_ (_08067_, _08066_, _08065_);
  and _59074_ (_08068_, _07733_, \oc8051_golden_model_1.DPL [1]);
  and _59075_ (_08069_, _07802_, \oc8051_golden_model_1.DPH [1]);
  nor _59076_ (_08070_, _08069_, _08068_);
  and _59077_ (_08071_, _08070_, _08067_);
  and _59078_ (_08072_, _08071_, _08064_);
  and _59079_ (_08073_, _08072_, _08062_);
  and _59080_ (_08074_, _08073_, _08056_);
  and _59081_ (_08075_, _08074_, _08046_);
  or _59082_ (_08076_, _07132_, _05952_);
  and _59083_ (_08077_, _08076_, _08075_);
  not _59084_ (_08078_, _08077_);
  and _59085_ (_08079_, _07681_, \oc8051_golden_model_1.SBUF [0]);
  not _59086_ (_08080_, _08079_);
  and _59087_ (_08081_, _07686_, \oc8051_golden_model_1.P2 [0]);
  not _59088_ (_08082_, _08081_);
  and _59089_ (_08083_, _07692_, \oc8051_golden_model_1.P3 [0]);
  and _59090_ (_08084_, _07688_, \oc8051_golden_model_1.IE [0]);
  nor _59091_ (_08085_, _08084_, _08083_);
  and _59092_ (_08086_, _08085_, _08082_);
  and _59093_ (_08087_, _08086_, _08080_);
  and _59094_ (_08088_, _07833_, \oc8051_golden_model_1.SP [0]);
  not _59095_ (_08089_, _08088_);
  and _59096_ (_08090_, _07733_, \oc8051_golden_model_1.DPL [0]);
  and _59097_ (_08091_, _07802_, \oc8051_golden_model_1.DPH [0]);
  nor _59098_ (_08092_, _08091_, _08090_);
  and _59099_ (_08093_, _08092_, _08089_);
  and _59100_ (_08094_, _07677_, \oc8051_golden_model_1.P1 [0]);
  and _59101_ (_08095_, _07679_, \oc8051_golden_model_1.SCON [0]);
  nor _59102_ (_08096_, _08095_, _08094_);
  and _59103_ (_08097_, _07670_, \oc8051_golden_model_1.TH1 [0]);
  and _59104_ (_08098_, _07667_, \oc8051_golden_model_1.TL1 [0]);
  nor _59105_ (_08099_, _08098_, _08097_);
  and _59106_ (_08100_, _08099_, _08096_);
  and _59107_ (_08101_, _08100_, _08093_);
  and _59108_ (_08102_, _08101_, _08087_);
  and _59109_ (_08103_, _07705_, \oc8051_golden_model_1.PSW [0]);
  not _59110_ (_08104_, _08103_);
  and _59111_ (_08105_, _07698_, \oc8051_golden_model_1.B [0]);
  and _59112_ (_08106_, _07701_, \oc8051_golden_model_1.ACC [0]);
  nor _59113_ (_08107_, _08106_, _08105_);
  and _59114_ (_08108_, _08107_, _08104_);
  and _59115_ (_08109_, _07641_, \oc8051_golden_model_1.PCON [0]);
  and _59116_ (_08110_, _07694_, \oc8051_golden_model_1.IP [0]);
  nor _59117_ (_08111_, _08110_, _08109_);
  and _59118_ (_08112_, _08111_, _08108_);
  and _59119_ (_08113_, _07653_, \oc8051_golden_model_1.TMOD [0]);
  not _59120_ (_08114_, _08113_);
  and _59121_ (_08115_, _07659_, \oc8051_golden_model_1.TL0 [0]);
  and _59122_ (_08116_, _07663_, \oc8051_golden_model_1.TH0 [0]);
  nor _59123_ (_08117_, _08116_, _08115_);
  and _59124_ (_08118_, _08117_, _08114_);
  and _59125_ (_08119_, _07730_, \oc8051_golden_model_1.P0 [0]);
  and _59126_ (_08120_, _07648_, \oc8051_golden_model_1.TCON [0]);
  nor _59127_ (_08121_, _08120_, _08119_);
  and _59128_ (_08122_, _08121_, _08118_);
  and _59129_ (_08123_, _08122_, _08112_);
  and _59130_ (_08124_, _08123_, _08102_);
  not _59131_ (_08125_, _08124_);
  and _59132_ (_08126_, _06931_, _06053_);
  or _59133_ (_08127_, _08126_, _08125_);
  and _59134_ (_08128_, _08127_, _08078_);
  and _59135_ (_08129_, _07681_, \oc8051_golden_model_1.SBUF [2]);
  not _59136_ (_08130_, _08129_);
  and _59137_ (_08131_, _07692_, \oc8051_golden_model_1.P3 [2]);
  and _59138_ (_08132_, _07688_, \oc8051_golden_model_1.IE [2]);
  nor _59139_ (_08133_, _08132_, _08131_);
  and _59140_ (_08134_, _08133_, _08130_);
  and _59141_ (_08135_, _07686_, \oc8051_golden_model_1.P2 [2]);
  and _59142_ (_08136_, _07667_, \oc8051_golden_model_1.TL1 [2]);
  nor _59143_ (_08137_, _08136_, _08135_);
  and _59144_ (_08138_, _08137_, _08134_);
  and _59145_ (_08139_, _07653_, \oc8051_golden_model_1.TMOD [2]);
  not _59146_ (_08140_, _08139_);
  and _59147_ (_08141_, _07659_, \oc8051_golden_model_1.TL0 [2]);
  and _59148_ (_08142_, _07663_, \oc8051_golden_model_1.TH0 [2]);
  nor _59149_ (_08143_, _08142_, _08141_);
  and _59150_ (_08144_, _08143_, _08140_);
  and _59151_ (_08145_, _07730_, \oc8051_golden_model_1.P0 [2]);
  and _59152_ (_08146_, _07648_, \oc8051_golden_model_1.TCON [2]);
  nor _59153_ (_08147_, _08146_, _08145_);
  and _59154_ (_08148_, _08147_, _08144_);
  and _59155_ (_08149_, _08148_, _08138_);
  and _59156_ (_08150_, _07705_, \oc8051_golden_model_1.PSW [2]);
  not _59157_ (_08151_, _08150_);
  and _59158_ (_08152_, _07698_, \oc8051_golden_model_1.B [2]);
  and _59159_ (_08153_, _07701_, \oc8051_golden_model_1.ACC [2]);
  nor _59160_ (_08154_, _08153_, _08152_);
  and _59161_ (_08155_, _08154_, _08151_);
  and _59162_ (_08156_, _07641_, \oc8051_golden_model_1.PCON [2]);
  and _59163_ (_08157_, _07694_, \oc8051_golden_model_1.IP [2]);
  nor _59164_ (_08158_, _08157_, _08156_);
  and _59165_ (_08159_, _08158_, _08155_);
  and _59166_ (_08160_, _07833_, \oc8051_golden_model_1.SP [2]);
  not _59167_ (_08161_, _08160_);
  and _59168_ (_08162_, _07733_, \oc8051_golden_model_1.DPL [2]);
  and _59169_ (_08163_, _07802_, \oc8051_golden_model_1.DPH [2]);
  nor _59170_ (_08164_, _08163_, _08162_);
  and _59171_ (_08165_, _08164_, _08161_);
  and _59172_ (_08166_, _07670_, \oc8051_golden_model_1.TH1 [2]);
  not _59173_ (_08167_, _08166_);
  and _59174_ (_08168_, _07677_, \oc8051_golden_model_1.P1 [2]);
  and _59175_ (_08169_, _07679_, \oc8051_golden_model_1.SCON [2]);
  nor _59176_ (_08170_, _08169_, _08168_);
  and _59177_ (_08171_, _08170_, _08167_);
  and _59178_ (_08172_, _08171_, _08165_);
  and _59179_ (_08173_, _08172_, _08159_);
  and _59180_ (_08174_, _08173_, _08149_);
  or _59181_ (_08175_, _07530_, _05952_);
  and _59182_ (_08176_, _08175_, _08174_);
  not _59183_ (_08177_, _08176_);
  and _59184_ (_08178_, _08177_, _08128_);
  and _59185_ (_08179_, _08178_, _08029_);
  and _59186_ (_08180_, _07670_, \oc8051_golden_model_1.TH1 [4]);
  not _59187_ (_08181_, _08180_);
  and _59188_ (_08182_, _07679_, \oc8051_golden_model_1.SCON [4]);
  and _59189_ (_08183_, _07677_, \oc8051_golden_model_1.P1 [4]);
  nor _59190_ (_08184_, _08183_, _08182_);
  and _59191_ (_08185_, _08184_, _08181_);
  and _59192_ (_08186_, _07681_, \oc8051_golden_model_1.SBUF [4]);
  not _59193_ (_08187_, _08186_);
  and _59194_ (_08188_, _07688_, \oc8051_golden_model_1.IE [4]);
  and _59195_ (_08189_, _07692_, \oc8051_golden_model_1.P3 [4]);
  nor _59196_ (_08190_, _08189_, _08188_);
  and _59197_ (_08191_, _08190_, _08187_);
  and _59198_ (_08192_, _07686_, \oc8051_golden_model_1.P2 [4]);
  and _59199_ (_08193_, _07667_, \oc8051_golden_model_1.TL1 [4]);
  nor _59200_ (_08194_, _08193_, _08192_);
  and _59201_ (_08195_, _08194_, _08191_);
  and _59202_ (_08196_, _08195_, _08185_);
  and _59203_ (_08197_, _07694_, \oc8051_golden_model_1.IP [4]);
  not _59204_ (_08198_, _08197_);
  and _59205_ (_08199_, _07698_, \oc8051_golden_model_1.B [4]);
  and _59206_ (_08200_, _07701_, \oc8051_golden_model_1.ACC [4]);
  nor _59207_ (_08201_, _08200_, _08199_);
  and _59208_ (_08202_, _08201_, _08198_);
  and _59209_ (_08203_, _07641_, \oc8051_golden_model_1.PCON [4]);
  and _59210_ (_08204_, _07705_, \oc8051_golden_model_1.PSW [4]);
  nor _59211_ (_08205_, _08204_, _08203_);
  and _59212_ (_08206_, _08205_, _08202_);
  and _59213_ (_08207_, _07648_, \oc8051_golden_model_1.TCON [4]);
  not _59214_ (_08208_, _08207_);
  and _59215_ (_08209_, _07659_, \oc8051_golden_model_1.TL0 [4]);
  and _59216_ (_08210_, _07663_, \oc8051_golden_model_1.TH0 [4]);
  nor _59217_ (_08211_, _08210_, _08209_);
  and _59218_ (_08212_, _08211_, _08208_);
  and _59219_ (_08213_, _07653_, \oc8051_golden_model_1.TMOD [4]);
  not _59220_ (_08214_, _08213_);
  and _59221_ (_08215_, _07730_, \oc8051_golden_model_1.P0 [4]);
  and _59222_ (_08216_, _07833_, \oc8051_golden_model_1.SP [4]);
  nor _59223_ (_08217_, _08216_, _08215_);
  and _59224_ (_08218_, _07733_, \oc8051_golden_model_1.DPL [4]);
  and _59225_ (_08219_, _07802_, \oc8051_golden_model_1.DPH [4]);
  nor _59226_ (_08220_, _08219_, _08218_);
  and _59227_ (_08221_, _08220_, _08217_);
  and _59228_ (_08222_, _08221_, _08214_);
  and _59229_ (_08223_, _08222_, _08212_);
  and _59230_ (_08224_, _08223_, _08206_);
  and _59231_ (_08225_, _08224_, _08196_);
  nand _59232_ (_08226_, _06881_, \oc8051_golden_model_1.IRAM[0] [4]);
  nand _59233_ (_08227_, _06726_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _59234_ (_08228_, _08227_, _06879_);
  nand _59235_ (_08229_, _08228_, _08226_);
  nand _59236_ (_08230_, _06726_, \oc8051_golden_model_1.IRAM[3] [4]);
  nand _59237_ (_08231_, _06881_, \oc8051_golden_model_1.IRAM[2] [4]);
  and _59238_ (_08232_, _08231_, _06887_);
  nand _59239_ (_08233_, _08232_, _08230_);
  nand _59240_ (_08234_, _08233_, _08229_);
  nand _59241_ (_08235_, _08234_, _06504_);
  nand _59242_ (_08236_, _06726_, \oc8051_golden_model_1.IRAM[7] [4]);
  nand _59243_ (_08237_, _06881_, \oc8051_golden_model_1.IRAM[6] [4]);
  and _59244_ (_08238_, _08237_, _06887_);
  nand _59245_ (_08239_, _08238_, _08236_);
  nand _59246_ (_08240_, _06881_, \oc8051_golden_model_1.IRAM[4] [4]);
  nand _59247_ (_08241_, _06726_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _59248_ (_08242_, _08241_, _06879_);
  nand _59249_ (_08243_, _08242_, _08240_);
  nand _59250_ (_08244_, _08243_, _08239_);
  nand _59251_ (_08245_, _08244_, _06894_);
  nand _59252_ (_08246_, _08245_, _08235_);
  nand _59253_ (_08247_, _08246_, _06328_);
  nand _59254_ (_08248_, _06726_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand _59255_ (_08249_, _06881_, \oc8051_golden_model_1.IRAM[10] [4]);
  and _59256_ (_08250_, _08249_, _06887_);
  nand _59257_ (_08251_, _08250_, _08248_);
  nand _59258_ (_08252_, _06881_, \oc8051_golden_model_1.IRAM[8] [4]);
  nand _59259_ (_08253_, _06726_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _59260_ (_08254_, _08253_, _06879_);
  nand _59261_ (_08255_, _08254_, _08252_);
  nand _59262_ (_08256_, _08255_, _08251_);
  nand _59263_ (_08257_, _08256_, _06504_);
  nand _59264_ (_08258_, _06726_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand _59265_ (_08259_, _06881_, \oc8051_golden_model_1.IRAM[14] [4]);
  and _59266_ (_08260_, _08259_, _06887_);
  nand _59267_ (_08261_, _08260_, _08258_);
  nand _59268_ (_08262_, _06881_, \oc8051_golden_model_1.IRAM[12] [4]);
  nand _59269_ (_08263_, _06726_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _59270_ (_08264_, _08263_, _06879_);
  nand _59271_ (_08265_, _08264_, _08262_);
  nand _59272_ (_08266_, _08265_, _08261_);
  nand _59273_ (_08267_, _08266_, _06894_);
  nand _59274_ (_08268_, _08267_, _08257_);
  nand _59275_ (_08269_, _08268_, _06908_);
  nand _59276_ (_08270_, _08269_, _08247_);
  or _59277_ (_08271_, _08270_, _05952_);
  and _59278_ (_08272_, _08271_, _08225_);
  not _59279_ (_08273_, _08272_);
  and _59280_ (_08274_, _08273_, _08179_);
  and _59281_ (_08275_, _08274_, _07980_);
  and _59282_ (_08276_, _08275_, _07886_);
  nor _59283_ (_08277_, _08276_, _07788_);
  and _59284_ (_08278_, _08276_, _07788_);
  nor _59285_ (_08279_, _08278_, _08277_);
  and _59286_ (_08280_, _08279_, _07067_);
  nor _59287_ (_08281_, _06137_, _06723_);
  or _59288_ (_08282_, _07278_, _06458_);
  not _59289_ (_08283_, _08282_);
  not _59290_ (_08284_, _06457_);
  and _59291_ (_08285_, _06866_, _08284_);
  and _59292_ (_08286_, _08285_, _08283_);
  and _59293_ (_08287_, _08286_, _07211_);
  not _59294_ (_08288_, _07785_);
  and _59295_ (_08289_, _08270_, _07977_);
  and _59296_ (_08290_, _07530_, _07353_);
  and _59297_ (_08291_, _07132_, _07022_);
  and _59298_ (_08292_, _08291_, _08290_);
  and _59299_ (_08293_, _08292_, _08289_);
  and _59300_ (_08294_, _08293_, _07883_);
  or _59301_ (_08295_, _08294_, _08288_);
  nand _59302_ (_08296_, _08294_, _08288_);
  and _59303_ (_08297_, _08296_, _08295_);
  and _59304_ (_08298_, _08297_, _07211_);
  or _59305_ (_08299_, _08298_, _08287_);
  not _59306_ (_08300_, _07031_);
  nor _59307_ (_08301_, _07032_, _05952_);
  and _59308_ (_08302_, _06166_, _04200_);
  and _59309_ (_08303_, _06205_, _04168_);
  nor _59310_ (_08304_, _08303_, _08302_);
  and _59311_ (_08305_, _06210_, _04205_);
  and _59312_ (_08306_, _06197_, _04208_);
  nor _59313_ (_08307_, _08306_, _08305_);
  and _59314_ (_08308_, _08307_, _08304_);
  and _59315_ (_08309_, _06161_, _04155_);
  and _59316_ (_08310_, _06203_, _04197_);
  nor _59317_ (_08311_, _08310_, _08309_);
  and _59318_ (_08312_, _06199_, _04180_);
  and _59319_ (_08313_, _06187_, _04159_);
  nor _59320_ (_08314_, _08313_, _08312_);
  and _59321_ (_08315_, _08314_, _08311_);
  and _59322_ (_08316_, _08315_, _08308_);
  and _59323_ (_08317_, _06170_, _04193_);
  and _59324_ (_08318_, _06185_, _04176_);
  nor _59325_ (_08319_, _08318_, _08317_);
  and _59326_ (_08320_, _06208_, _04172_);
  and _59327_ (_08321_, _06182_, _04122_);
  nor _59328_ (_08322_, _08321_, _08320_);
  and _59329_ (_08323_, _08322_, _08319_);
  and _59330_ (_08324_, _06179_, _04149_);
  and _59331_ (_08325_, _06194_, _04165_);
  nor _59332_ (_08326_, _08325_, _08324_);
  and _59333_ (_08327_, _06175_, _04185_);
  and _59334_ (_08328_, _06192_, _04190_);
  nor _59335_ (_08329_, _08328_, _08327_);
  and _59336_ (_08330_, _08329_, _08326_);
  and _59337_ (_08331_, _08330_, _08323_);
  and _59338_ (_08332_, _08331_, _08316_);
  nor _59339_ (_08333_, _08332_, _07787_);
  and _59340_ (_08334_, _08333_, _08301_);
  nand _59341_ (_08335_, _08332_, _06021_);
  and _59342_ (_08336_, _07638_, \oc8051_golden_model_1.P0 [7]);
  not _59343_ (_08337_, _05984_);
  nor _59344_ (_08338_, _06759_, _08337_);
  and _59345_ (_08339_, _08338_, _06361_);
  and _59346_ (_08340_, _08339_, _06087_);
  and _59347_ (_08341_, _08340_, _07637_);
  and _59348_ (_08342_, _08341_, \oc8051_golden_model_1.TCON [7]);
  not _59349_ (_08343_, _06087_);
  and _59350_ (_08344_, _08339_, _08343_);
  and _59351_ (_08345_, _08344_, _07676_);
  and _59352_ (_08346_, _08345_, \oc8051_golden_model_1.P1 [7]);
  and _59353_ (_08347_, _08340_, _07676_);
  and _59354_ (_08348_, _08347_, \oc8051_golden_model_1.SCON [7]);
  and _59355_ (_08349_, _08344_, _07685_);
  and _59356_ (_08350_, _08349_, \oc8051_golden_model_1.P2 [7]);
  and _59357_ (_08351_, _08340_, _07685_);
  and _59358_ (_08352_, _08351_, \oc8051_golden_model_1.IE [7]);
  and _59359_ (_08353_, _08344_, _07691_);
  and _59360_ (_08354_, _08353_, \oc8051_golden_model_1.P3 [7]);
  and _59361_ (_08355_, _07704_, _08344_);
  and _59362_ (_08356_, _08355_, \oc8051_golden_model_1.PSW [7]);
  and _59363_ (_08357_, _08340_, _07691_);
  and _59364_ (_08358_, _08357_, \oc8051_golden_model_1.IP [7]);
  and _59365_ (_08359_, _08344_, _07700_);
  and _59366_ (_08360_, _08359_, \oc8051_golden_model_1.ACC [7]);
  and _59367_ (_08361_, _08344_, _07697_);
  and _59368_ (_08362_, _08361_, \oc8051_golden_model_1.B [7]);
  or _59369_ (_08363_, _08362_, _08360_);
  or _59370_ (_08364_, _08363_, _08358_);
  or _59371_ (_08365_, _08364_, _08356_);
  or _59372_ (_08366_, _08365_, _08354_);
  or _59373_ (_08367_, _08366_, _08352_);
  or _59374_ (_08368_, _08367_, _08350_);
  or _59375_ (_08369_, _08368_, _08348_);
  or _59376_ (_08370_, _08369_, _08346_);
  or _59377_ (_08371_, _08370_, _08342_);
  nor _59378_ (_08372_, _08371_, _08336_);
  and _59379_ (_08373_, _08372_, _07786_);
  nor _59380_ (_08374_, _08373_, _07640_);
  and _59381_ (_08375_, _07640_, \oc8051_golden_model_1.PSW [7]);
  or _59382_ (_08376_, _08375_, _08374_);
  and _59383_ (_08377_, _08376_, _06991_);
  not _59384_ (_08378_, _06975_);
  or _59385_ (_08379_, _08374_, _08378_);
  not _59386_ (_08380_, _06953_);
  not _59387_ (_08381_, _06955_);
  not _59388_ (_08382_, _05567_);
  or _59389_ (_08383_, _05689_, _08382_);
  not _59390_ (_08384_, _08383_);
  and _59391_ (_08385_, _08384_, _08297_);
  and _59392_ (_08386_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [4]);
  and _59393_ (_08387_, _08386_, \oc8051_golden_model_1.PC [6]);
  and _59394_ (_08388_, _08387_, _05850_);
  and _59395_ (_08389_, _08388_, \oc8051_golden_model_1.PC [7]);
  nor _59396_ (_08390_, _08388_, \oc8051_golden_model_1.PC [7]);
  nor _59397_ (_08391_, _08390_, _08389_);
  and _59398_ (_08392_, _08391_, _06943_);
  not _59399_ (_08393_, \oc8051_golden_model_1.ACC [7]);
  nor _59400_ (_08394_, _06943_, _08393_);
  or _59401_ (_08395_, _08394_, _08392_);
  and _59402_ (_08396_, _08395_, _08383_);
  or _59403_ (_08397_, _08396_, _08385_);
  and _59404_ (_08398_, _08397_, _06949_);
  nor _59405_ (_08399_, \oc8051_golden_model_1.SP [1], \oc8051_golden_model_1.SP [0]);
  and _59406_ (_08400_, _08399_, _06447_);
  nor _59407_ (_08401_, _08400_, _06238_);
  nor _59408_ (_08402_, \oc8051_golden_model_1.SP [2], \oc8051_golden_model_1.SP [1]);
  and _59409_ (_08403_, _08402_, _06238_);
  and _59410_ (_08404_, _08403_, _06029_);
  nor _59411_ (_08405_, _08404_, _08401_);
  nor _59412_ (_08406_, _08405_, _06448_);
  not _59413_ (_08407_, _08406_);
  nand _59414_ (_08408_, _07353_, _06993_);
  not _59415_ (_08409_, _06448_);
  and _59416_ (_08410_, _06992_, _05983_);
  nor _59417_ (_08411_, _08410_, _08409_);
  nand _59418_ (_08412_, _08411_, _08408_);
  and _59419_ (_08413_, _08412_, _08407_);
  nor _59420_ (_08414_, _08399_, _06447_);
  nor _59421_ (_08415_, _08414_, _08400_);
  nor _59422_ (_08416_, _08415_, _06448_);
  not _59423_ (_08417_, _08416_);
  nand _59424_ (_08418_, _07530_, _06993_);
  and _59425_ (_08419_, _06992_, _06403_);
  nor _59426_ (_08420_, _08419_, _08409_);
  nand _59427_ (_08421_, _08420_, _08418_);
  and _59428_ (_08422_, _08421_, _08417_);
  nor _59429_ (_08423_, _07132_, _06992_);
  nor _59430_ (_08424_, _06993_, _06799_);
  or _59431_ (_08425_, _08424_, _08423_);
  nand _59432_ (_08426_, _08425_, _06448_);
  nor _59433_ (_08427_, _07083_, _06448_);
  not _59434_ (_08428_, _08427_);
  and _59435_ (_08429_, _08428_, _08426_);
  or _59436_ (_08430_, _06992_, _06931_);
  and _59437_ (_08431_, _06992_, _06016_);
  nor _59438_ (_08432_, _08431_, _08409_);
  nand _59439_ (_08433_, _08432_, _08430_);
  nor _59440_ (_08434_, _06448_, \oc8051_golden_model_1.SP [0]);
  not _59441_ (_08435_, _08434_);
  and _59442_ (_08436_, _08435_, _08433_);
  or _59443_ (_08437_, _08436_, _07740_);
  nand _59444_ (_08438_, _08435_, _08433_);
  or _59445_ (_08439_, _08438_, _07738_);
  nand _59446_ (_08440_, _08439_, _08437_);
  and _59447_ (_08441_, _08440_, _08429_);
  or _59448_ (_08442_, _08438_, \oc8051_golden_model_1.IRAM[2] [7]);
  nand _59449_ (_08443_, _08428_, _08426_);
  or _59450_ (_08444_, _08436_, \oc8051_golden_model_1.IRAM[3] [7]);
  and _59451_ (_08445_, _08444_, _08443_);
  and _59452_ (_08446_, _08445_, _08442_);
  nor _59453_ (_08447_, _08446_, _08441_);
  nand _59454_ (_08448_, _08447_, _08422_);
  not _59455_ (_08449_, _08422_);
  or _59456_ (_08450_, _08436_, \oc8051_golden_model_1.IRAM[5] [7]);
  or _59457_ (_08451_, _08438_, \oc8051_golden_model_1.IRAM[4] [7]);
  and _59458_ (_08452_, _08451_, _08429_);
  and _59459_ (_08453_, _08452_, _08450_);
  or _59460_ (_08454_, _08438_, \oc8051_golden_model_1.IRAM[6] [7]);
  or _59461_ (_08455_, _08436_, \oc8051_golden_model_1.IRAM[7] [7]);
  and _59462_ (_08456_, _08455_, _08443_);
  and _59463_ (_08457_, _08456_, _08454_);
  nor _59464_ (_08458_, _08457_, _08453_);
  nand _59465_ (_08459_, _08458_, _08449_);
  nand _59466_ (_08460_, _08459_, _08448_);
  nand _59467_ (_08461_, _08460_, _08413_);
  not _59468_ (_08462_, _08413_);
  or _59469_ (_08463_, _08438_, \oc8051_golden_model_1.IRAM[8] [7]);
  or _59470_ (_08464_, _08436_, \oc8051_golden_model_1.IRAM[9] [7]);
  nand _59471_ (_08465_, _08464_, _08463_);
  nand _59472_ (_08466_, _08465_, _08429_);
  or _59473_ (_08467_, _08438_, \oc8051_golden_model_1.IRAM[10] [7]);
  or _59474_ (_08468_, _08436_, \oc8051_golden_model_1.IRAM[11] [7]);
  nand _59475_ (_08469_, _08468_, _08467_);
  nand _59476_ (_08470_, _08469_, _08443_);
  nand _59477_ (_08471_, _08470_, _08466_);
  nand _59478_ (_08472_, _08471_, _08422_);
  or _59479_ (_08473_, _08438_, \oc8051_golden_model_1.IRAM[12] [7]);
  or _59480_ (_08474_, _08436_, \oc8051_golden_model_1.IRAM[13] [7]);
  nand _59481_ (_08475_, _08474_, _08473_);
  nand _59482_ (_08476_, _08475_, _08429_);
  or _59483_ (_08477_, _08438_, \oc8051_golden_model_1.IRAM[14] [7]);
  or _59484_ (_08478_, _08436_, \oc8051_golden_model_1.IRAM[15] [7]);
  nand _59485_ (_08479_, _08478_, _08477_);
  nand _59486_ (_08480_, _08479_, _08443_);
  nand _59487_ (_08481_, _08480_, _08476_);
  nand _59488_ (_08482_, _08481_, _08449_);
  nand _59489_ (_08483_, _08482_, _08472_);
  nand _59490_ (_08484_, _08483_, _08462_);
  and _59491_ (_08485_, _08484_, _08461_);
  and _59492_ (_08486_, _08485_, _06948_);
  or _59493_ (_08487_, _08486_, _08398_);
  and _59494_ (_08488_, _08487_, _08381_);
  and _59495_ (_08489_, _08272_, _07979_);
  not _59496_ (_08490_, _08127_);
  and _59497_ (_08491_, _08490_, _08077_);
  and _59498_ (_08492_, _08176_, _08028_);
  and _59499_ (_08493_, _08492_, _08491_);
  and _59500_ (_08494_, _08493_, _08489_);
  and _59501_ (_08495_, _08494_, _07885_);
  or _59502_ (_08496_, _08495_, _07788_);
  nand _59503_ (_08497_, _08495_, _07788_);
  and _59504_ (_08498_, _08497_, _08496_);
  and _59505_ (_08499_, _08498_, _06955_);
  or _59506_ (_08500_, _08499_, _08488_);
  and _59507_ (_08501_, _08500_, _08380_);
  not _59508_ (_08502_, _07640_);
  nand _59509_ (_08503_, _08373_, _08502_);
  and _59510_ (_08504_, _08503_, _06953_);
  or _59511_ (_08505_, _08504_, _07272_);
  or _59512_ (_08506_, _08505_, _08501_);
  nor _59513_ (_08507_, _08391_, _05690_);
  nor _59514_ (_08508_, _08507_, _06963_);
  and _59515_ (_08509_, _08508_, _08506_);
  and _59516_ (_08510_, _08288_, _06963_);
  or _59517_ (_08511_, _08510_, _06975_);
  or _59518_ (_08512_, _08511_, _08509_);
  and _59519_ (_08513_, _08512_, _08379_);
  or _59520_ (_08514_, _08513_, _06038_);
  nand _59521_ (_08515_, _07787_, _06038_);
  and _59522_ (_08516_, _08515_, _06036_);
  and _59523_ (_08517_, _08516_, _08514_);
  nor _59524_ (_08518_, _08373_, _08502_);
  not _59525_ (_08519_, _08518_);
  and _59526_ (_08520_, _08519_, _08503_);
  and _59527_ (_08521_, _08520_, _06035_);
  or _59528_ (_08522_, _08521_, _08517_);
  and _59529_ (_08523_, _08522_, _05686_);
  not _59530_ (_08524_, _08391_);
  or _59531_ (_08525_, _08524_, _05686_);
  nand _59532_ (_08526_, _08525_, _06233_);
  or _59533_ (_08527_, _08526_, _08523_);
  nand _59534_ (_08528_, _07787_, _06573_);
  and _59535_ (_08529_, _08528_, _08527_);
  or _59536_ (_08530_, _08529_, _06992_);
  and _59537_ (_08531_, _08485_, _06053_);
  nand _59538_ (_08532_, _07737_, _06992_);
  or _59539_ (_08533_, _08532_, _08531_);
  and _59540_ (_08534_, _08533_, _07308_);
  and _59541_ (_08535_, _08534_, _08530_);
  or _59542_ (_08536_, _08535_, _08377_);
  and _59543_ (_08537_, _08536_, _05673_);
  or _59544_ (_08538_, _08524_, _05673_);
  nand _59545_ (_08539_, _08538_, _07009_);
  or _59546_ (_08540_, _08539_, _08537_);
  not _59547_ (_08541_, _07009_);
  nand _59548_ (_08542_, _07785_, _08541_);
  and _59549_ (_08543_, _08542_, _08540_);
  or _59550_ (_08544_, _08543_, _07013_);
  not _59551_ (_08545_, _07010_);
  or _59552_ (_08546_, _08485_, _07231_);
  and _59553_ (_08547_, _08546_, _08545_);
  and _59554_ (_08548_, _08547_, _08544_);
  not _59555_ (_08549_, _08332_);
  nor _59556_ (_08550_, _08549_, _07785_);
  and _59557_ (_08551_, _06170_, _04508_);
  and _59558_ (_08552_, _06166_, _04532_);
  nor _59559_ (_08553_, _08552_, _08551_);
  and _59560_ (_08554_, _06161_, _04492_);
  and _59561_ (_08555_, _06187_, _04503_);
  nor _59562_ (_08556_, _08555_, _08554_);
  and _59563_ (_08557_, _08556_, _08553_);
  and _59564_ (_08558_, _06182_, _04510_);
  and _59565_ (_08559_, _06205_, _04525_);
  nor _59566_ (_08560_, _08559_, _08558_);
  and _59567_ (_08561_, _06197_, _04515_);
  and _59568_ (_08562_, _06192_, _04505_);
  nor _59569_ (_08563_, _08562_, _08561_);
  and _59570_ (_08564_, _08563_, _08560_);
  and _59571_ (_08565_, _08564_, _08557_);
  and _59572_ (_08566_, _06199_, _04494_);
  and _59573_ (_08567_, _06194_, _04521_);
  nor _59574_ (_08568_, _08567_, _08566_);
  and _59575_ (_08569_, _06185_, _04513_);
  and _59576_ (_08570_, _06179_, _04523_);
  nor _59577_ (_08571_, _08570_, _08569_);
  and _59578_ (_08572_, _08571_, _08568_);
  and _59579_ (_08573_, _06210_, _04497_);
  and _59580_ (_08574_, _06203_, _04530_);
  nor _59581_ (_08575_, _08574_, _08573_);
  and _59582_ (_08576_, _06208_, _04499_);
  and _59583_ (_08577_, _06175_, _04519_);
  nor _59584_ (_08578_, _08577_, _08576_);
  and _59585_ (_08579_, _08578_, _08575_);
  and _59586_ (_08580_, _08579_, _08572_);
  and _59587_ (_08581_, _08580_, _08565_);
  and _59588_ (_08582_, _06185_, _04579_);
  and _59589_ (_08583_, _06208_, _04538_);
  nor _59590_ (_08584_, _08583_, _08582_);
  and _59591_ (_08585_, _06197_, _04560_);
  and _59592_ (_08586_, _06187_, _04552_);
  nor _59593_ (_08587_, _08586_, _08585_);
  and _59594_ (_08588_, _08587_, _08584_);
  and _59595_ (_08589_, _06205_, _04568_);
  and _59596_ (_08590_, _06194_, _04572_);
  nor _59597_ (_08591_, _08590_, _08589_);
  and _59598_ (_08592_, _06175_, _04566_);
  and _59599_ (_08593_, _06192_, _04550_);
  nor _59600_ (_08594_, _08593_, _08592_);
  and _59601_ (_08595_, _08594_, _08591_);
  and _59602_ (_08596_, _08595_, _08588_);
  and _59603_ (_08597_, _06179_, _04570_);
  and _59604_ (_08598_, _06203_, _04557_);
  nor _59605_ (_08599_, _08598_, _08597_);
  and _59606_ (_08600_, _06170_, _04577_);
  and _59607_ (_08601_, _06210_, _04544_);
  nor _59608_ (_08602_, _08601_, _08600_);
  and _59609_ (_08603_, _08602_, _08599_);
  and _59610_ (_08604_, _06199_, _04546_);
  and _59611_ (_08605_, _06166_, _04562_);
  nor _59612_ (_08606_, _08605_, _08604_);
  and _59613_ (_08607_, _06161_, _04540_);
  and _59614_ (_08608_, _06182_, _04555_);
  nor _59615_ (_08609_, _08608_, _08607_);
  and _59616_ (_08610_, _08609_, _08606_);
  and _59617_ (_08611_, _08610_, _08603_);
  and _59618_ (_08612_, _08611_, _08596_);
  nor _59619_ (_08613_, _08612_, _08581_);
  and _59620_ (_08614_, _06832_, _06633_);
  and _59621_ (_08615_, _06445_, _06215_);
  and _59622_ (_08616_, _08615_, _08614_);
  and _59623_ (_08617_, _06170_, _04623_);
  and _59624_ (_08618_, _06203_, _04603_);
  nor _59625_ (_08619_, _08618_, _08617_);
  and _59626_ (_08620_, _06161_, _04585_);
  and _59627_ (_08621_, _06166_, _04608_);
  nor _59628_ (_08622_, _08621_, _08620_);
  and _59629_ (_08623_, _08622_, _08619_);
  and _59630_ (_08624_, _06197_, _04606_);
  and _59631_ (_08625_, _06199_, _04592_);
  nor _59632_ (_08626_, _08625_, _08624_);
  and _59633_ (_08627_, _06185_, _04625_);
  and _59634_ (_08628_, _06210_, _04587_);
  nor _59635_ (_08629_, _08628_, _08627_);
  and _59636_ (_08630_, _08629_, _08626_);
  and _59637_ (_08631_, _08630_, _08623_);
  and _59638_ (_08632_, _06192_, _04596_);
  and _59639_ (_08633_, _06205_, _04614_);
  nor _59640_ (_08634_, _08633_, _08632_);
  and _59641_ (_08635_, _06187_, _04598_);
  and _59642_ (_08636_, _06194_, _04618_);
  nor _59643_ (_08637_, _08636_, _08635_);
  and _59644_ (_08638_, _08637_, _08634_);
  and _59645_ (_08639_, _06182_, _04601_);
  and _59646_ (_08640_, _06179_, _04616_);
  nor _59647_ (_08641_, _08640_, _08639_);
  and _59648_ (_08642_, _06208_, _04590_);
  and _59649_ (_08643_, _06175_, _04612_);
  nor _59650_ (_08644_, _08643_, _08642_);
  and _59651_ (_08645_, _08644_, _08641_);
  and _59652_ (_08646_, _08645_, _08638_);
  and _59653_ (_08647_, _08646_, _08631_);
  nor _59654_ (_08648_, _08647_, _08332_);
  and _59655_ (_08649_, _08648_, _08616_);
  and _59656_ (_08650_, _08649_, _08613_);
  and _59657_ (_08651_, _08650_, \oc8051_golden_model_1.B [7]);
  not _59658_ (_08652_, _08612_);
  and _59659_ (_08653_, _08652_, _08581_);
  and _59660_ (_08654_, _08653_, _08649_);
  and _59661_ (_08655_, _08654_, \oc8051_golden_model_1.ACC [7]);
  or _59662_ (_08656_, _08655_, _08651_);
  and _59663_ (_08657_, _08647_, _08549_);
  and _59664_ (_08658_, _08612_, _08581_);
  and _59665_ (_08659_, _08658_, _08657_);
  and _59666_ (_08660_, _08659_, _08616_);
  and _59667_ (_08661_, _08660_, \oc8051_golden_model_1.P0 [7]);
  not _59668_ (_08662_, _06215_);
  and _59669_ (_08663_, _06445_, _08662_);
  and _59670_ (_08664_, _08663_, _08614_);
  not _59671_ (_08665_, _08581_);
  and _59672_ (_08666_, _08612_, _08665_);
  and _59673_ (_08667_, _08666_, _08657_);
  and _59674_ (_08668_, _08667_, _08664_);
  and _59675_ (_08669_, _08668_, \oc8051_golden_model_1.SCON [7]);
  or _59676_ (_08670_, _08669_, _08661_);
  or _59677_ (_08671_, _08670_, _08656_);
  not _59678_ (_08672_, _06633_);
  and _59679_ (_08673_, _06832_, _08672_);
  and _59680_ (_08674_, _08673_, _08663_);
  and _59681_ (_08675_, _08674_, _08659_);
  and _59682_ (_08676_, _08675_, \oc8051_golden_model_1.TMOD [7]);
  and _59683_ (_08677_, _08674_, _08667_);
  and _59684_ (_08678_, _08677_, \oc8051_golden_model_1.SBUF [7]);
  or _59685_ (_08679_, _08678_, _08676_);
  and _59686_ (_08680_, _08664_, _08659_);
  and _59687_ (_08681_, _08680_, \oc8051_golden_model_1.TCON [7]);
  and _59688_ (_08682_, _08667_, _08616_);
  and _59689_ (_08683_, _08682_, \oc8051_golden_model_1.P1 [7]);
  or _59690_ (_08684_, _08683_, _08681_);
  or _59691_ (_08685_, _08684_, _08679_);
  and _59692_ (_08686_, _08657_, _08653_);
  and _59693_ (_08687_, _08686_, _08616_);
  and _59694_ (_08688_, _08687_, \oc8051_golden_model_1.P2 [7]);
  and _59695_ (_08689_, _08657_, _08613_);
  and _59696_ (_08690_, _08689_, _08664_);
  and _59697_ (_08691_, _08690_, \oc8051_golden_model_1.IP [7]);
  or _59698_ (_08692_, _08691_, _08688_);
  and _59699_ (_08693_, _08686_, _08664_);
  and _59700_ (_08694_, _08693_, \oc8051_golden_model_1.IE [7]);
  and _59701_ (_08695_, _08689_, _08616_);
  and _59702_ (_08696_, _08695_, \oc8051_golden_model_1.P3 [7]);
  or _59703_ (_08697_, _08696_, _08694_);
  or _59704_ (_08698_, _08697_, _08692_);
  not _59705_ (_08699_, _06832_);
  and _59706_ (_08700_, _08699_, _06633_);
  and _59707_ (_08701_, _08700_, _08663_);
  and _59708_ (_08702_, _08701_, _08659_);
  and _59709_ (_08703_, _08702_, \oc8051_golden_model_1.TL0 [7]);
  and _59710_ (_08704_, _08666_, _08649_);
  and _59711_ (_08705_, _08704_, \oc8051_golden_model_1.PSW [7]);
  or _59712_ (_08706_, _08705_, _08703_);
  or _59713_ (_08707_, _08706_, _08698_);
  or _59714_ (_08708_, _08707_, _08685_);
  or _59715_ (_08709_, _08708_, _08671_);
  nor _59716_ (_08710_, _06445_, _06215_);
  and _59717_ (_08711_, _08710_, _08659_);
  and _59718_ (_08712_, _08711_, _08614_);
  and _59719_ (_08713_, _08712_, \oc8051_golden_model_1.TH0 [7]);
  nor _59720_ (_08714_, _06832_, _06633_);
  and _59721_ (_08715_, _08714_, _08659_);
  and _59722_ (_08716_, _08715_, _08663_);
  and _59723_ (_08717_, _08716_, \oc8051_golden_model_1.TL1 [7]);
  and _59724_ (_08718_, _08659_, _08615_);
  and _59725_ (_08719_, _08673_, _08718_);
  and _59726_ (_08720_, _08719_, \oc8051_golden_model_1.SP [7]);
  or _59727_ (_08721_, _08720_, _08717_);
  or _59728_ (_08722_, _08721_, _08713_);
  and _59729_ (_08723_, _08715_, _08615_);
  and _59730_ (_08724_, _08723_, \oc8051_golden_model_1.DPH [7]);
  and _59731_ (_08725_, _08711_, _08673_);
  and _59732_ (_08726_, _08725_, \oc8051_golden_model_1.TH1 [7]);
  or _59733_ (_08727_, _08726_, _08724_);
  and _59734_ (_08728_, _08700_, _08718_);
  and _59735_ (_08729_, _08728_, \oc8051_golden_model_1.DPL [7]);
  not _59736_ (_08730_, _06445_);
  and _59737_ (_08731_, _08730_, _06215_);
  and _59738_ (_08732_, _08731_, _08715_);
  and _59739_ (_08733_, _08732_, \oc8051_golden_model_1.PCON [7]);
  or _59740_ (_08734_, _08733_, _08729_);
  or _59741_ (_08735_, _08734_, _08727_);
  or _59742_ (_08736_, _08735_, _08722_);
  or _59743_ (_08737_, _08736_, _08709_);
  or _59744_ (_08738_, _08737_, _08550_);
  and _59745_ (_08739_, _08738_, _07010_);
  nor _59746_ (_08740_, _07267_, _07254_);
  nor _59747_ (_08741_, _07023_, _07252_);
  and _59748_ (_08742_, _08741_, _08740_);
  not _59749_ (_08743_, _08742_);
  or _59750_ (_08744_, _08743_, _08739_);
  or _59751_ (_08745_, _08744_, _08548_);
  or _59752_ (_08746_, _08742_, _05952_);
  and _59753_ (_08747_, _08746_, _08745_);
  or _59754_ (_08748_, _08747_, _06021_);
  and _59755_ (_08749_, _08748_, _08335_);
  or _59756_ (_08750_, _08749_, _05724_);
  not _59757_ (_08751_, _06112_);
  nor _59758_ (_08752_, _08751_, _05952_);
  and _59759_ (_08753_, _08524_, _05724_);
  nor _59760_ (_08754_, _08753_, _08752_);
  and _59761_ (_08755_, _08754_, _08750_);
  not _59762_ (_08756_, _06284_);
  nor _59763_ (_08757_, _08756_, _05952_);
  not _59764_ (_08758_, _08333_);
  nand _59765_ (_08759_, _08332_, _07787_);
  and _59766_ (_08760_, _08759_, _08758_);
  and _59767_ (_08761_, _08760_, _08752_);
  or _59768_ (_08762_, _08761_, _08757_);
  or _59769_ (_08763_, _08762_, _08755_);
  not _59770_ (_08764_, _08301_);
  not _59771_ (_08765_, _08757_);
  nor _59772_ (_08766_, _07787_, _08393_);
  and _59773_ (_08767_, _07787_, _08393_);
  nor _59774_ (_08768_, _08767_, _08766_);
  or _59775_ (_08769_, _08768_, _08765_);
  and _59776_ (_08770_, _08769_, _08764_);
  and _59777_ (_08771_, _08770_, _08763_);
  or _59778_ (_08772_, _08771_, _08334_);
  and _59779_ (_08773_, _08772_, _08300_);
  and _59780_ (_08774_, _08766_, _07031_);
  or _59781_ (_08775_, _08774_, _05736_);
  or _59782_ (_08776_, _08775_, _08773_);
  not _59783_ (_08777_, _06130_);
  nor _59784_ (_08778_, _08777_, _05952_);
  and _59785_ (_08779_, _08524_, _05736_);
  nor _59786_ (_08780_, _08779_, _08778_);
  and _59787_ (_08781_, _08780_, _08776_);
  not _59788_ (_08782_, _06292_);
  nor _59789_ (_08783_, _08782_, _05952_);
  and _59790_ (_08784_, _08759_, _08778_);
  or _59791_ (_08785_, _08784_, _08783_);
  or _59792_ (_08786_, _08785_, _08781_);
  nand _59793_ (_08787_, _08767_, _08783_);
  and _59794_ (_08788_, _08787_, _05734_);
  and _59795_ (_08789_, _08788_, _08786_);
  nand _59796_ (_08790_, _08391_, _05732_);
  nand _59797_ (_08791_, _08790_, _08286_);
  or _59798_ (_08792_, _08791_, _08789_);
  and _59799_ (_08793_, _08792_, _08299_);
  and _59800_ (_08794_, _08297_, _07210_);
  or _59801_ (_08795_, _08794_, _07051_);
  or _59802_ (_08796_, _08795_, _08793_);
  not _59803_ (_08797_, _07050_);
  nand _59804_ (_08798_, _08484_, _08461_);
  or _59805_ (_08799_, _08436_, \oc8051_golden_model_1.IRAM[1] [6]);
  or _59806_ (_08800_, _08438_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _59807_ (_08801_, _08800_, _08429_);
  and _59808_ (_08802_, _08801_, _08799_);
  or _59809_ (_08803_, _08438_, \oc8051_golden_model_1.IRAM[2] [6]);
  or _59810_ (_08804_, _08436_, \oc8051_golden_model_1.IRAM[3] [6]);
  and _59811_ (_08805_, _08804_, _08443_);
  and _59812_ (_08806_, _08805_, _08803_);
  nor _59813_ (_08807_, _08806_, _08802_);
  nand _59814_ (_08808_, _08807_, _08422_);
  or _59815_ (_08809_, _08436_, \oc8051_golden_model_1.IRAM[5] [6]);
  or _59816_ (_08810_, _08438_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _59817_ (_08811_, _08810_, _08429_);
  and _59818_ (_08812_, _08811_, _08809_);
  or _59819_ (_08813_, _08438_, \oc8051_golden_model_1.IRAM[6] [6]);
  or _59820_ (_08814_, _08436_, \oc8051_golden_model_1.IRAM[7] [6]);
  and _59821_ (_08815_, _08814_, _08443_);
  and _59822_ (_08816_, _08815_, _08813_);
  nor _59823_ (_08817_, _08816_, _08812_);
  nand _59824_ (_08818_, _08817_, _08449_);
  nand _59825_ (_08819_, _08818_, _08808_);
  nand _59826_ (_08820_, _08819_, _08413_);
  or _59827_ (_08821_, _08438_, \oc8051_golden_model_1.IRAM[8] [6]);
  or _59828_ (_08822_, _08436_, \oc8051_golden_model_1.IRAM[9] [6]);
  nand _59829_ (_08823_, _08822_, _08821_);
  nand _59830_ (_08824_, _08823_, _08429_);
  or _59831_ (_08825_, _08438_, \oc8051_golden_model_1.IRAM[10] [6]);
  or _59832_ (_08826_, _08436_, \oc8051_golden_model_1.IRAM[11] [6]);
  nand _59833_ (_08827_, _08826_, _08825_);
  nand _59834_ (_08828_, _08827_, _08443_);
  nand _59835_ (_08829_, _08828_, _08824_);
  nand _59836_ (_08830_, _08829_, _08422_);
  or _59837_ (_08831_, _08438_, \oc8051_golden_model_1.IRAM[12] [6]);
  or _59838_ (_08832_, _08436_, \oc8051_golden_model_1.IRAM[13] [6]);
  nand _59839_ (_08833_, _08832_, _08831_);
  nand _59840_ (_08834_, _08833_, _08429_);
  or _59841_ (_08835_, _08438_, \oc8051_golden_model_1.IRAM[14] [6]);
  or _59842_ (_08836_, _08436_, \oc8051_golden_model_1.IRAM[15] [6]);
  nand _59843_ (_08837_, _08836_, _08835_);
  nand _59844_ (_08838_, _08837_, _08443_);
  nand _59845_ (_08839_, _08838_, _08834_);
  nand _59846_ (_08840_, _08839_, _08449_);
  nand _59847_ (_08841_, _08840_, _08830_);
  nand _59848_ (_08842_, _08841_, _08462_);
  nand _59849_ (_08843_, _08842_, _08820_);
  or _59850_ (_08844_, _08436_, \oc8051_golden_model_1.IRAM[1] [5]);
  or _59851_ (_08845_, _08438_, \oc8051_golden_model_1.IRAM[0] [5]);
  and _59852_ (_08846_, _08845_, _08429_);
  and _59853_ (_08847_, _08846_, _08844_);
  or _59854_ (_08848_, _08438_, \oc8051_golden_model_1.IRAM[2] [5]);
  or _59855_ (_08849_, _08436_, \oc8051_golden_model_1.IRAM[3] [5]);
  and _59856_ (_08850_, _08849_, _08443_);
  and _59857_ (_08851_, _08850_, _08848_);
  nor _59858_ (_08852_, _08851_, _08847_);
  nand _59859_ (_08853_, _08852_, _08422_);
  or _59860_ (_08854_, _08436_, \oc8051_golden_model_1.IRAM[5] [5]);
  or _59861_ (_08855_, _08438_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _59862_ (_08856_, _08855_, _08429_);
  and _59863_ (_08857_, _08856_, _08854_);
  or _59864_ (_08858_, _08438_, \oc8051_golden_model_1.IRAM[6] [5]);
  or _59865_ (_08859_, _08436_, \oc8051_golden_model_1.IRAM[7] [5]);
  and _59866_ (_08860_, _08859_, _08443_);
  and _59867_ (_08861_, _08860_, _08858_);
  nor _59868_ (_08862_, _08861_, _08857_);
  nand _59869_ (_08863_, _08862_, _08449_);
  nand _59870_ (_08864_, _08863_, _08853_);
  nand _59871_ (_08865_, _08864_, _08413_);
  or _59872_ (_08866_, _08438_, \oc8051_golden_model_1.IRAM[8] [5]);
  or _59873_ (_08867_, _08436_, \oc8051_golden_model_1.IRAM[9] [5]);
  nand _59874_ (_08868_, _08867_, _08866_);
  nand _59875_ (_08869_, _08868_, _08429_);
  or _59876_ (_08870_, _08438_, \oc8051_golden_model_1.IRAM[10] [5]);
  or _59877_ (_08871_, _08436_, \oc8051_golden_model_1.IRAM[11] [5]);
  nand _59878_ (_08872_, _08871_, _08870_);
  nand _59879_ (_08873_, _08872_, _08443_);
  nand _59880_ (_08874_, _08873_, _08869_);
  nand _59881_ (_08875_, _08874_, _08422_);
  or _59882_ (_08876_, _08438_, \oc8051_golden_model_1.IRAM[12] [5]);
  or _59883_ (_08877_, _08436_, \oc8051_golden_model_1.IRAM[13] [5]);
  nand _59884_ (_08878_, _08877_, _08876_);
  nand _59885_ (_08879_, _08878_, _08429_);
  or _59886_ (_08880_, _08438_, \oc8051_golden_model_1.IRAM[14] [5]);
  or _59887_ (_08881_, _08436_, \oc8051_golden_model_1.IRAM[15] [5]);
  nand _59888_ (_08882_, _08881_, _08880_);
  nand _59889_ (_08883_, _08882_, _08443_);
  nand _59890_ (_08884_, _08883_, _08879_);
  nand _59891_ (_08885_, _08884_, _08449_);
  nand _59892_ (_08886_, _08885_, _08875_);
  nand _59893_ (_08887_, _08886_, _08462_);
  nand _59894_ (_08888_, _08887_, _08865_);
  or _59895_ (_08889_, _08436_, \oc8051_golden_model_1.IRAM[1] [4]);
  or _59896_ (_08890_, _08438_, \oc8051_golden_model_1.IRAM[0] [4]);
  and _59897_ (_08891_, _08890_, _08429_);
  and _59898_ (_08892_, _08891_, _08889_);
  or _59899_ (_08893_, _08438_, \oc8051_golden_model_1.IRAM[2] [4]);
  or _59900_ (_08894_, _08436_, \oc8051_golden_model_1.IRAM[3] [4]);
  and _59901_ (_08895_, _08894_, _08443_);
  and _59902_ (_08896_, _08895_, _08893_);
  nor _59903_ (_08897_, _08896_, _08892_);
  nand _59904_ (_08898_, _08897_, _08422_);
  or _59905_ (_08899_, _08436_, \oc8051_golden_model_1.IRAM[5] [4]);
  or _59906_ (_08900_, _08438_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _59907_ (_08901_, _08900_, _08429_);
  and _59908_ (_08902_, _08901_, _08899_);
  or _59909_ (_08904_, _08438_, \oc8051_golden_model_1.IRAM[6] [4]);
  or _59910_ (_08905_, _08436_, \oc8051_golden_model_1.IRAM[7] [4]);
  and _59911_ (_08906_, _08905_, _08443_);
  and _59912_ (_08907_, _08906_, _08904_);
  nor _59913_ (_08908_, _08907_, _08902_);
  nand _59914_ (_08909_, _08908_, _08449_);
  nand _59915_ (_08910_, _08909_, _08898_);
  nand _59916_ (_08911_, _08910_, _08413_);
  or _59917_ (_08912_, _08438_, \oc8051_golden_model_1.IRAM[8] [4]);
  or _59918_ (_08913_, _08436_, \oc8051_golden_model_1.IRAM[9] [4]);
  nand _59919_ (_08915_, _08913_, _08912_);
  nand _59920_ (_08916_, _08915_, _08429_);
  or _59921_ (_08917_, _08438_, \oc8051_golden_model_1.IRAM[10] [4]);
  or _59922_ (_08918_, _08436_, \oc8051_golden_model_1.IRAM[11] [4]);
  nand _59923_ (_08919_, _08918_, _08917_);
  nand _59924_ (_08920_, _08919_, _08443_);
  nand _59925_ (_08921_, _08920_, _08916_);
  nand _59926_ (_08922_, _08921_, _08422_);
  or _59927_ (_08923_, _08438_, \oc8051_golden_model_1.IRAM[12] [4]);
  or _59928_ (_08924_, _08436_, \oc8051_golden_model_1.IRAM[13] [4]);
  nand _59929_ (_08926_, _08924_, _08923_);
  nand _59930_ (_08927_, _08926_, _08429_);
  or _59931_ (_08928_, _08438_, \oc8051_golden_model_1.IRAM[14] [4]);
  or _59932_ (_08929_, _08436_, \oc8051_golden_model_1.IRAM[15] [4]);
  nand _59933_ (_08930_, _08929_, _08928_);
  nand _59934_ (_08931_, _08930_, _08443_);
  nand _59935_ (_08932_, _08931_, _08927_);
  nand _59936_ (_08933_, _08932_, _08449_);
  nand _59937_ (_08934_, _08933_, _08922_);
  nand _59938_ (_08935_, _08934_, _08462_);
  nand _59939_ (_08937_, _08935_, _08911_);
  or _59940_ (_08938_, _08436_, \oc8051_golden_model_1.IRAM[1] [3]);
  or _59941_ (_08939_, _08438_, \oc8051_golden_model_1.IRAM[0] [3]);
  and _59942_ (_08940_, _08939_, _08429_);
  and _59943_ (_08941_, _08940_, _08938_);
  or _59944_ (_08942_, _08438_, \oc8051_golden_model_1.IRAM[2] [3]);
  or _59945_ (_08943_, _08436_, \oc8051_golden_model_1.IRAM[3] [3]);
  and _59946_ (_08944_, _08943_, _08443_);
  and _59947_ (_08945_, _08944_, _08942_);
  nor _59948_ (_08946_, _08945_, _08941_);
  nand _59949_ (_08948_, _08946_, _08422_);
  or _59950_ (_08949_, _08436_, \oc8051_golden_model_1.IRAM[5] [3]);
  or _59951_ (_08950_, _08438_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _59952_ (_08951_, _08950_, _08429_);
  and _59953_ (_08952_, _08951_, _08949_);
  or _59954_ (_08953_, _08438_, \oc8051_golden_model_1.IRAM[6] [3]);
  or _59955_ (_08954_, _08436_, \oc8051_golden_model_1.IRAM[7] [3]);
  and _59956_ (_08955_, _08954_, _08443_);
  and _59957_ (_08956_, _08955_, _08953_);
  nor _59958_ (_08957_, _08956_, _08952_);
  nand _59959_ (_08959_, _08957_, _08449_);
  nand _59960_ (_08960_, _08959_, _08948_);
  nand _59961_ (_08961_, _08960_, _08413_);
  or _59962_ (_08962_, _08438_, \oc8051_golden_model_1.IRAM[8] [3]);
  or _59963_ (_08963_, _08436_, \oc8051_golden_model_1.IRAM[9] [3]);
  nand _59964_ (_08964_, _08963_, _08962_);
  nand _59965_ (_08965_, _08964_, _08429_);
  or _59966_ (_08966_, _08438_, \oc8051_golden_model_1.IRAM[10] [3]);
  or _59967_ (_08967_, _08436_, \oc8051_golden_model_1.IRAM[11] [3]);
  nand _59968_ (_08968_, _08967_, _08966_);
  nand _59969_ (_08970_, _08968_, _08443_);
  nand _59970_ (_08971_, _08970_, _08965_);
  nand _59971_ (_08972_, _08971_, _08422_);
  or _59972_ (_08973_, _08438_, \oc8051_golden_model_1.IRAM[12] [3]);
  or _59973_ (_08974_, _08436_, \oc8051_golden_model_1.IRAM[13] [3]);
  nand _59974_ (_08975_, _08974_, _08973_);
  nand _59975_ (_08976_, _08975_, _08429_);
  or _59976_ (_08977_, _08438_, \oc8051_golden_model_1.IRAM[14] [3]);
  or _59977_ (_08978_, _08436_, \oc8051_golden_model_1.IRAM[15] [3]);
  nand _59978_ (_08979_, _08978_, _08977_);
  nand _59979_ (_08980_, _08979_, _08443_);
  nand _59980_ (_08981_, _08980_, _08976_);
  nand _59981_ (_08982_, _08981_, _08449_);
  nand _59982_ (_08983_, _08982_, _08972_);
  nand _59983_ (_08984_, _08983_, _08462_);
  nand _59984_ (_08985_, _08984_, _08961_);
  or _59985_ (_08986_, _08436_, \oc8051_golden_model_1.IRAM[1] [2]);
  or _59986_ (_08987_, _08438_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _59987_ (_08988_, _08987_, _08429_);
  and _59988_ (_08989_, _08988_, _08986_);
  or _59989_ (_08990_, _08438_, \oc8051_golden_model_1.IRAM[2] [2]);
  or _59990_ (_08991_, _08436_, \oc8051_golden_model_1.IRAM[3] [2]);
  and _59991_ (_08992_, _08991_, _08443_);
  and _59992_ (_08993_, _08992_, _08990_);
  nor _59993_ (_08994_, _08993_, _08989_);
  nand _59994_ (_08995_, _08994_, _08422_);
  or _59995_ (_08996_, _08436_, \oc8051_golden_model_1.IRAM[5] [2]);
  or _59996_ (_08997_, _08438_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _59997_ (_08998_, _08997_, _08429_);
  and _59998_ (_08999_, _08998_, _08996_);
  or _59999_ (_09000_, _08438_, \oc8051_golden_model_1.IRAM[6] [2]);
  or _60000_ (_09001_, _08436_, \oc8051_golden_model_1.IRAM[7] [2]);
  and _60001_ (_09002_, _09001_, _08443_);
  and _60002_ (_09003_, _09002_, _09000_);
  nor _60003_ (_09004_, _09003_, _08999_);
  nand _60004_ (_09005_, _09004_, _08449_);
  nand _60005_ (_09006_, _09005_, _08995_);
  nand _60006_ (_09007_, _09006_, _08413_);
  or _60007_ (_09008_, _08438_, \oc8051_golden_model_1.IRAM[8] [2]);
  or _60008_ (_09009_, _08436_, \oc8051_golden_model_1.IRAM[9] [2]);
  nand _60009_ (_09010_, _09009_, _09008_);
  nand _60010_ (_09011_, _09010_, _08429_);
  or _60011_ (_09012_, _08438_, \oc8051_golden_model_1.IRAM[10] [2]);
  or _60012_ (_09013_, _08436_, \oc8051_golden_model_1.IRAM[11] [2]);
  nand _60013_ (_09014_, _09013_, _09012_);
  nand _60014_ (_09015_, _09014_, _08443_);
  nand _60015_ (_09016_, _09015_, _09011_);
  nand _60016_ (_09017_, _09016_, _08422_);
  or _60017_ (_09018_, _08438_, \oc8051_golden_model_1.IRAM[12] [2]);
  or _60018_ (_09019_, _08436_, \oc8051_golden_model_1.IRAM[13] [2]);
  nand _60019_ (_09020_, _09019_, _09018_);
  nand _60020_ (_09021_, _09020_, _08429_);
  or _60021_ (_09022_, _08438_, \oc8051_golden_model_1.IRAM[14] [2]);
  or _60022_ (_09023_, _08436_, \oc8051_golden_model_1.IRAM[15] [2]);
  nand _60023_ (_09024_, _09023_, _09022_);
  nand _60024_ (_09025_, _09024_, _08443_);
  nand _60025_ (_09026_, _09025_, _09021_);
  nand _60026_ (_09027_, _09026_, _08449_);
  nand _60027_ (_09028_, _09027_, _09017_);
  nand _60028_ (_09029_, _09028_, _08462_);
  nand _60029_ (_09030_, _09029_, _09007_);
  or _60030_ (_09031_, _08436_, \oc8051_golden_model_1.IRAM[1] [1]);
  or _60031_ (_09032_, _08438_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _60032_ (_09033_, _09032_, _08429_);
  and _60033_ (_09034_, _09033_, _09031_);
  or _60034_ (_09035_, _08438_, \oc8051_golden_model_1.IRAM[2] [1]);
  or _60035_ (_09036_, _08436_, \oc8051_golden_model_1.IRAM[3] [1]);
  and _60036_ (_09037_, _09036_, _08443_);
  and _60037_ (_09038_, _09037_, _09035_);
  nor _60038_ (_09039_, _09038_, _09034_);
  nand _60039_ (_09040_, _09039_, _08422_);
  or _60040_ (_09041_, _08436_, \oc8051_golden_model_1.IRAM[5] [1]);
  or _60041_ (_09042_, _08438_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _60042_ (_09043_, _09042_, _08429_);
  and _60043_ (_09044_, _09043_, _09041_);
  or _60044_ (_09045_, _08438_, \oc8051_golden_model_1.IRAM[6] [1]);
  or _60045_ (_09046_, _08436_, \oc8051_golden_model_1.IRAM[7] [1]);
  and _60046_ (_09047_, _09046_, _08443_);
  and _60047_ (_09048_, _09047_, _09045_);
  nor _60048_ (_09049_, _09048_, _09044_);
  nand _60049_ (_09050_, _09049_, _08449_);
  nand _60050_ (_09051_, _09050_, _09040_);
  nand _60051_ (_09052_, _09051_, _08413_);
  or _60052_ (_09053_, _08438_, \oc8051_golden_model_1.IRAM[8] [1]);
  or _60053_ (_09054_, _08436_, \oc8051_golden_model_1.IRAM[9] [1]);
  nand _60054_ (_09055_, _09054_, _09053_);
  nand _60055_ (_09056_, _09055_, _08429_);
  or _60056_ (_09057_, _08438_, \oc8051_golden_model_1.IRAM[10] [1]);
  or _60057_ (_09058_, _08436_, \oc8051_golden_model_1.IRAM[11] [1]);
  nand _60058_ (_09059_, _09058_, _09057_);
  nand _60059_ (_09060_, _09059_, _08443_);
  nand _60060_ (_09061_, _09060_, _09056_);
  nand _60061_ (_09062_, _09061_, _08422_);
  or _60062_ (_09063_, _08438_, \oc8051_golden_model_1.IRAM[12] [1]);
  or _60063_ (_09064_, _08436_, \oc8051_golden_model_1.IRAM[13] [1]);
  nand _60064_ (_09065_, _09064_, _09063_);
  nand _60065_ (_09066_, _09065_, _08429_);
  or _60066_ (_09067_, _08438_, \oc8051_golden_model_1.IRAM[14] [1]);
  or _60067_ (_09068_, _08436_, \oc8051_golden_model_1.IRAM[15] [1]);
  nand _60068_ (_09069_, _09068_, _09067_);
  nand _60069_ (_09070_, _09069_, _08443_);
  nand _60070_ (_09071_, _09070_, _09066_);
  nand _60071_ (_09072_, _09071_, _08449_);
  nand _60072_ (_09073_, _09072_, _09062_);
  nand _60073_ (_09074_, _09073_, _08462_);
  and _60074_ (_09075_, _09074_, _09052_);
  or _60075_ (_09076_, _08436_, \oc8051_golden_model_1.IRAM[1] [0]);
  or _60076_ (_09077_, _08438_, \oc8051_golden_model_1.IRAM[0] [0]);
  and _60077_ (_09078_, _09077_, _08429_);
  and _60078_ (_09079_, _09078_, _09076_);
  or _60079_ (_09080_, _08438_, \oc8051_golden_model_1.IRAM[2] [0]);
  or _60080_ (_09081_, _08436_, \oc8051_golden_model_1.IRAM[3] [0]);
  and _60081_ (_09082_, _09081_, _08443_);
  and _60082_ (_09083_, _09082_, _09080_);
  nor _60083_ (_09084_, _09083_, _09079_);
  nand _60084_ (_09085_, _09084_, _08422_);
  or _60085_ (_09086_, _08436_, \oc8051_golden_model_1.IRAM[5] [0]);
  or _60086_ (_09087_, _08438_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _60087_ (_09088_, _09087_, _08429_);
  and _60088_ (_09089_, _09088_, _09086_);
  or _60089_ (_09090_, _08438_, \oc8051_golden_model_1.IRAM[6] [0]);
  or _60090_ (_09091_, _08436_, \oc8051_golden_model_1.IRAM[7] [0]);
  and _60091_ (_09092_, _09091_, _08443_);
  and _60092_ (_09093_, _09092_, _09090_);
  nor _60093_ (_09094_, _09093_, _09089_);
  nand _60094_ (_09095_, _09094_, _08449_);
  nand _60095_ (_09096_, _09095_, _09085_);
  nand _60096_ (_09097_, _09096_, _08413_);
  or _60097_ (_09098_, _08438_, \oc8051_golden_model_1.IRAM[8] [0]);
  or _60098_ (_09099_, _08436_, \oc8051_golden_model_1.IRAM[9] [0]);
  nand _60099_ (_09100_, _09099_, _09098_);
  nand _60100_ (_09101_, _09100_, _08429_);
  or _60101_ (_09102_, _08438_, \oc8051_golden_model_1.IRAM[10] [0]);
  or _60102_ (_09103_, _08436_, \oc8051_golden_model_1.IRAM[11] [0]);
  nand _60103_ (_09104_, _09103_, _09102_);
  nand _60104_ (_09105_, _09104_, _08443_);
  nand _60105_ (_09106_, _09105_, _09101_);
  nand _60106_ (_09107_, _09106_, _08422_);
  or _60107_ (_09108_, _08438_, \oc8051_golden_model_1.IRAM[12] [0]);
  or _60108_ (_09109_, _08436_, \oc8051_golden_model_1.IRAM[13] [0]);
  nand _60109_ (_09110_, _09109_, _09108_);
  nand _60110_ (_09111_, _09110_, _08429_);
  or _60111_ (_09112_, _08438_, \oc8051_golden_model_1.IRAM[14] [0]);
  or _60112_ (_09113_, _08436_, \oc8051_golden_model_1.IRAM[15] [0]);
  nand _60113_ (_09114_, _09113_, _09112_);
  nand _60114_ (_09115_, _09114_, _08443_);
  nand _60115_ (_09116_, _09115_, _09111_);
  nand _60116_ (_09117_, _09116_, _08449_);
  nand _60117_ (_09118_, _09117_, _09107_);
  nand _60118_ (_09119_, _09118_, _08462_);
  and _60119_ (_09120_, _09119_, _09097_);
  nor _60120_ (_09121_, _09120_, _09075_);
  and _60121_ (_09122_, _09121_, _09030_);
  and _60122_ (_09123_, _09122_, _08985_);
  and _60123_ (_09124_, _09123_, _08937_);
  and _60124_ (_09125_, _09124_, _08888_);
  and _60125_ (_09126_, _09125_, _08843_);
  nor _60126_ (_09127_, _09126_, _08798_);
  and _60127_ (_09128_, _09126_, _08798_);
  or _60128_ (_09129_, _09128_, _09127_);
  or _60129_ (_09130_, _09129_, _07052_);
  and _60130_ (_09131_, _09130_, _08797_);
  and _60131_ (_09132_, _09131_, _08796_);
  and _60132_ (_09133_, _08498_, _07050_);
  or _60133_ (_09134_, _09133_, _06127_);
  or _60134_ (_09135_, _09134_, _09132_);
  and _60135_ (_09136_, _05350_, \oc8051_golden_model_1.PC [2]);
  and _60136_ (_09137_, _09136_, \oc8051_golden_model_1.PC [3]);
  and _60137_ (_09138_, _09137_, _08387_);
  and _60138_ (_09139_, _09138_, \oc8051_golden_model_1.PC [7]);
  nor _60139_ (_09140_, _09138_, \oc8051_golden_model_1.PC [7]);
  nor _60140_ (_09141_, _09140_, _09139_);
  not _60141_ (_09142_, _09141_);
  nand _60142_ (_09143_, _09142_, _06127_);
  and _60143_ (_09144_, _09143_, _09135_);
  or _60144_ (_09145_, _09144_, _05752_);
  and _60145_ (_09146_, _08524_, _05752_);
  nor _60146_ (_09147_, _09146_, _07058_);
  and _60147_ (_09148_, _09147_, _09145_);
  and _60148_ (_09149_, _08374_, _07058_);
  and _60149_ (_09150_, _07005_, _05750_);
  or _60150_ (_09151_, _09150_, _09149_);
  or _60151_ (_09152_, _09151_, _09148_);
  nor _60152_ (_09153_, _09152_, _08281_);
  nor _60153_ (_09154_, _07609_, _06464_);
  not _60154_ (_09155_, _07223_);
  not _60155_ (_09156_, _07883_);
  not _60156_ (_09157_, _07977_);
  not _60157_ (_09158_, _08270_);
  not _60158_ (_09159_, _07353_);
  not _60159_ (_09160_, _07530_);
  not _60160_ (_09161_, _07132_);
  and _60161_ (_09162_, _09161_, _06931_);
  and _60162_ (_09163_, _09162_, _09160_);
  and _60163_ (_09164_, _09163_, _09159_);
  and _60164_ (_09165_, _09164_, _09158_);
  and _60165_ (_09166_, _09165_, _09157_);
  and _60166_ (_09167_, _09166_, _09156_);
  nor _60167_ (_09168_, _09167_, _08288_);
  and _60168_ (_09169_, _09167_, _08288_);
  nor _60169_ (_09170_, _09169_, _09168_);
  and _60170_ (_09171_, _09170_, _09155_);
  nor _60171_ (_09172_, _09171_, _09154_);
  nor _60172_ (_09173_, _09172_, _09153_);
  and _60173_ (_09174_, _09170_, _07223_);
  nor _60174_ (_09175_, _09174_, _07068_);
  not _60175_ (_09176_, _09175_);
  nor _60176_ (_09177_, _09176_, _09173_);
  and _60177_ (_09178_, _08842_, _08820_);
  and _60178_ (_09179_, _08887_, _08865_);
  and _60179_ (_09180_, _08935_, _08911_);
  and _60180_ (_09181_, _08984_, _08961_);
  and _60181_ (_09182_, _09029_, _09007_);
  and _60182_ (_09183_, _09120_, _09075_);
  and _60183_ (_09184_, _09183_, _09182_);
  and _60184_ (_09185_, _09184_, _09181_);
  and _60185_ (_09186_, _09185_, _09180_);
  and _60186_ (_09187_, _09186_, _09179_);
  and _60187_ (_09188_, _09187_, _09178_);
  nor _60188_ (_09189_, _09188_, _08798_);
  and _60189_ (_09190_, _09188_, _08798_);
  or _60190_ (_09191_, _09190_, _09189_);
  nor _60191_ (_09192_, _09191_, _07069_);
  nor _60192_ (_09193_, _09192_, _07067_);
  not _60193_ (_09194_, _09193_);
  nor _60194_ (_09195_, _09194_, _09177_);
  nor _60195_ (_09196_, _09195_, _08280_);
  nor _60196_ (_09197_, _09196_, _07305_);
  or _60197_ (_09198_, _09197_, _07634_);
  and _60198_ (_09199_, _09198_, _07633_);
  not _60199_ (_09200_, _06127_);
  and _60200_ (_09201_, \oc8051_golden_model_1.PC [9], \oc8051_golden_model_1.PC [8]);
  and _60201_ (_09202_, _09201_, \oc8051_golden_model_1.PC [10]);
  and _60202_ (_09203_, _09202_, _08389_);
  and _60203_ (_09204_, _09203_, \oc8051_golden_model_1.PC [11]);
  and _60204_ (_09205_, _09204_, \oc8051_golden_model_1.PC [12]);
  and _60205_ (_09206_, _09205_, \oc8051_golden_model_1.PC [13]);
  and _60206_ (_09207_, _09206_, \oc8051_golden_model_1.PC [14]);
  nor _60207_ (_09208_, _09207_, \oc8051_golden_model_1.PC [15]);
  and _60208_ (_09209_, _09201_, _08389_);
  and _60209_ (_09210_, _09209_, \oc8051_golden_model_1.PC [10]);
  and _60210_ (_09211_, _09210_, \oc8051_golden_model_1.PC [11]);
  and _60211_ (_09212_, _09211_, \oc8051_golden_model_1.PC [12]);
  and _60212_ (_09213_, _09212_, \oc8051_golden_model_1.PC [13]);
  and _60213_ (_09214_, _09213_, \oc8051_golden_model_1.PC [14]);
  and _60214_ (_09215_, _09214_, \oc8051_golden_model_1.PC [15]);
  nor _60215_ (_09216_, _09215_, _09208_);
  and _60216_ (_09217_, _09216_, _09200_);
  not _60217_ (_09218_, \oc8051_golden_model_1.PC [15]);
  and _60218_ (_09219_, \oc8051_golden_model_1.PC [12], \oc8051_golden_model_1.PC [13]);
  and _60219_ (_09220_, \oc8051_golden_model_1.PC [11], \oc8051_golden_model_1.PC [10]);
  and _60220_ (_09221_, _09220_, _09201_);
  and _60221_ (_09222_, _09221_, _09139_);
  and _60222_ (_09223_, _09222_, _09219_);
  and _60223_ (_09224_, _09223_, \oc8051_golden_model_1.PC [14]);
  and _60224_ (_09225_, _09224_, _09218_);
  nor _60225_ (_09226_, _09224_, _09218_);
  or _60226_ (_09227_, _09226_, _09225_);
  and _60227_ (_09228_, _09227_, _06127_);
  or _60228_ (_09229_, _09228_, _09217_);
  and _60229_ (_09230_, _09229_, _07628_);
  and _60230_ (_09231_, _09230_, _07631_);
  or _60231_ (_40751_, _09231_, _09199_);
  not _60232_ (_09232_, \oc8051_golden_model_1.B [7]);
  nor _60233_ (_09233_, _01336_, _09232_);
  nor _60234_ (_09234_, _07698_, _09232_);
  and _60235_ (_09235_, _08768_, _07698_);
  or _60236_ (_09236_, _09235_, _09234_);
  and _60237_ (_09237_, _09236_, _06284_);
  nor _60238_ (_09238_, _08361_, _09232_);
  and _60239_ (_09239_, _08374_, _08361_);
  or _60240_ (_09240_, _09239_, _09238_);
  and _60241_ (_09241_, _09240_, _06039_);
  and _60242_ (_09242_, _08498_, _07698_);
  or _60243_ (_09243_, _09242_, _09234_);
  or _60244_ (_09244_, _09243_, _06954_);
  and _60245_ (_09245_, _07698_, \oc8051_golden_model_1.ACC [7]);
  or _60246_ (_09246_, _09245_, _09234_);
  and _60247_ (_09247_, _09246_, _06938_);
  nor _60248_ (_09248_, _06938_, _09232_);
  or _60249_ (_09249_, _09248_, _06102_);
  or _60250_ (_09250_, _09249_, _09247_);
  and _60251_ (_09251_, _09250_, _06044_);
  and _60252_ (_09252_, _09251_, _09244_);
  and _60253_ (_09253_, _08503_, _08361_);
  or _60254_ (_09254_, _09253_, _09238_);
  and _60255_ (_09255_, _09254_, _06043_);
  or _60256_ (_09256_, _09255_, _06239_);
  or _60257_ (_09257_, _09256_, _09252_);
  not _60258_ (_09258_, _07698_);
  nor _60259_ (_09259_, _07785_, _09258_);
  or _60260_ (_09260_, _09259_, _09234_);
  or _60261_ (_09261_, _09260_, _06848_);
  and _60262_ (_09262_, _09261_, _09257_);
  or _60263_ (_09263_, _09262_, _06219_);
  or _60264_ (_09264_, _09246_, _06220_);
  and _60265_ (_09265_, _09264_, _06040_);
  and _60266_ (_09266_, _09265_, _09263_);
  or _60267_ (_09267_, _09266_, _09241_);
  and _60268_ (_09268_, _09267_, _06033_);
  and _60269_ (_09269_, _06114_, _06221_);
  or _60270_ (_09270_, _09238_, _08519_);
  and _60271_ (_09271_, _09254_, _06032_);
  and _60272_ (_09272_, _09271_, _09270_);
  or _60273_ (_09273_, _09272_, _09269_);
  or _60274_ (_09274_, _09273_, _09268_);
  and _60275_ (_09275_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [7]);
  and _60276_ (_09276_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [6]);
  and _60277_ (_09277_, _09276_, _09275_);
  and _60278_ (_09278_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [2]);
  and _60279_ (_09279_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  and _60280_ (_09280_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [6]);
  nor _60281_ (_09281_, _09280_, _09279_);
  nor _60282_ (_09282_, _09281_, _09277_);
  and _60283_ (_09283_, _09282_, _09278_);
  nor _60284_ (_09284_, _09283_, _09277_);
  and _60285_ (_09285_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [7]);
  and _60286_ (_09286_, _09285_, _09280_);
  and _60287_ (_09287_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [6]);
  nor _60288_ (_09288_, _09287_, _09275_);
  nor _60289_ (_09289_, _09288_, _09286_);
  not _60290_ (_09290_, _09289_);
  nor _60291_ (_09291_, _09290_, _09284_);
  and _60292_ (_09292_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [3]);
  and _60293_ (_09293_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [3]);
  and _60294_ (_09294_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [4]);
  and _60295_ (_09295_, _09294_, _09293_);
  nor _60296_ (_09296_, _09294_, _09293_);
  nor _60297_ (_09297_, _09296_, _09295_);
  and _60298_ (_09298_, _09297_, _09292_);
  nor _60299_ (_09299_, _09297_, _09292_);
  nor _60300_ (_09300_, _09299_, _09298_);
  and _60301_ (_09301_, _09290_, _09284_);
  nor _60302_ (_09302_, _09301_, _09291_);
  and _60303_ (_09303_, _09302_, _09300_);
  nor _60304_ (_09304_, _09303_, _09291_);
  not _60305_ (_09305_, _09280_);
  and _60306_ (_09306_, _09285_, _09305_);
  and _60307_ (_09307_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [5]);
  and _60308_ (_09308_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [6]);
  and _60309_ (_09309_, _09308_, _09293_);
  and _60310_ (_09310_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [4]);
  and _60311_ (_09311_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [6]);
  nor _60312_ (_09312_, _09311_, _09310_);
  nor _60313_ (_09313_, _09312_, _09309_);
  and _60314_ (_09314_, _09313_, _09307_);
  nor _60315_ (_09315_, _09313_, _09307_);
  nor _60316_ (_09316_, _09315_, _09314_);
  and _60317_ (_09317_, _09316_, _09306_);
  nor _60318_ (_09318_, _09316_, _09306_);
  nor _60319_ (_09319_, _09318_, _09317_);
  not _60320_ (_09320_, _09319_);
  nor _60321_ (_09321_, _09320_, _09304_);
  and _60322_ (_09322_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [2]);
  and _60323_ (_09323_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [7]);
  and _60324_ (_09324_, _09323_, _09322_);
  nor _60325_ (_09325_, _09298_, _09295_);
  and _60326_ (_09326_, \oc8051_golden_model_1.ACC [2], \oc8051_golden_model_1.B [7]);
  and _60327_ (_09327_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [3]);
  and _60328_ (_09328_, _09327_, _09326_);
  nor _60329_ (_09329_, _09327_, _09326_);
  nor _60330_ (_09330_, _09329_, _09328_);
  not _60331_ (_09331_, _09330_);
  nor _60332_ (_09332_, _09331_, _09325_);
  and _60333_ (_09333_, _09331_, _09325_);
  nor _60334_ (_09334_, _09333_, _09332_);
  and _60335_ (_09335_, _09334_, _09324_);
  nor _60336_ (_09336_, _09334_, _09324_);
  nor _60337_ (_09337_, _09336_, _09335_);
  and _60338_ (_09338_, _09320_, _09304_);
  nor _60339_ (_09339_, _09338_, _09321_);
  and _60340_ (_09340_, _09339_, _09337_);
  nor _60341_ (_09341_, _09340_, _09321_);
  nor _60342_ (_09342_, _09314_, _09309_);
  and _60343_ (_09343_, \oc8051_golden_model_1.ACC [3], \oc8051_golden_model_1.B [7]);
  and _60344_ (_09344_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [6]);
  and _60345_ (_09345_, _09344_, _09343_);
  nor _60346_ (_09346_, _09344_, _09343_);
  nor _60347_ (_09347_, _09346_, _09345_);
  not _60348_ (_09348_, _09347_);
  nor _60349_ (_09349_, _09348_, _09342_);
  and _60350_ (_09350_, _09348_, _09342_);
  nor _60351_ (_09351_, _09350_, _09349_);
  and _60352_ (_09352_, _09351_, _09328_);
  nor _60353_ (_09353_, _09351_, _09328_);
  nor _60354_ (_09354_, _09353_, _09352_);
  nor _60355_ (_09355_, _09317_, _09286_);
  and _60356_ (_09356_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [5]);
  and _60357_ (_09357_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [7]);
  and _60358_ (_09358_, _09357_, _09308_);
  nor _60359_ (_09359_, _09357_, _09308_);
  nor _60360_ (_09360_, _09359_, _09358_);
  and _60361_ (_09361_, _09360_, _09356_);
  nor _60362_ (_09362_, _09360_, _09356_);
  nor _60363_ (_09363_, _09362_, _09361_);
  not _60364_ (_09364_, _09363_);
  nor _60365_ (_09365_, _09364_, _09355_);
  and _60366_ (_09366_, _09364_, _09355_);
  nor _60367_ (_09367_, _09366_, _09365_);
  and _60368_ (_09368_, _09367_, _09354_);
  nor _60369_ (_09369_, _09367_, _09354_);
  nor _60370_ (_09370_, _09369_, _09368_);
  not _60371_ (_09371_, _09370_);
  nor _60372_ (_09372_, _09371_, _09341_);
  nor _60373_ (_09373_, _09335_, _09332_);
  not _60374_ (_09374_, _09373_);
  and _60375_ (_09375_, _09371_, _09341_);
  nor _60376_ (_09376_, _09375_, _09372_);
  and _60377_ (_09377_, _09376_, _09374_);
  nor _60378_ (_09378_, _09377_, _09372_);
  nor _60379_ (_09379_, _09352_, _09349_);
  not _60380_ (_09380_, _09379_);
  nor _60381_ (_09381_, _09368_, _09365_);
  not _60382_ (_09382_, _09381_);
  and _60383_ (_09383_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [7]);
  and _60384_ (_09384_, _09383_, _09308_);
  and _60385_ (_09385_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [7]);
  and _60386_ (_09386_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [6]);
  nor _60387_ (_09387_, _09386_, _09385_);
  nor _60388_ (_09388_, _09387_, _09384_);
  nor _60389_ (_09389_, _09361_, _09358_);
  and _60390_ (_09390_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [7]);
  and _60391_ (_09391_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [6]);
  and _60392_ (_09392_, _09391_, _09390_);
  nor _60393_ (_09393_, _09391_, _09390_);
  nor _60394_ (_09394_, _09393_, _09392_);
  not _60395_ (_09395_, _09394_);
  nor _60396_ (_09396_, _09395_, _09389_);
  and _60397_ (_09397_, _09395_, _09389_);
  nor _60398_ (_09398_, _09397_, _09396_);
  and _60399_ (_09399_, _09398_, _09345_);
  nor _60400_ (_09400_, _09398_, _09345_);
  nor _60401_ (_09401_, _09400_, _09399_);
  and _60402_ (_09402_, _09401_, _09388_);
  nor _60403_ (_09403_, _09401_, _09388_);
  nor _60404_ (_09404_, _09403_, _09402_);
  and _60405_ (_09405_, _09404_, _09382_);
  nor _60406_ (_09406_, _09404_, _09382_);
  nor _60407_ (_09407_, _09406_, _09405_);
  and _60408_ (_09408_, _09407_, _09380_);
  nor _60409_ (_09409_, _09407_, _09380_);
  nor _60410_ (_09410_, _09409_, _09408_);
  not _60411_ (_09411_, _09410_);
  nor _60412_ (_09412_, _09411_, _09378_);
  nor _60413_ (_09413_, _09408_, _09405_);
  nor _60414_ (_09414_, _09399_, _09396_);
  not _60415_ (_09415_, _09414_);
  and _60416_ (_09416_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [7]);
  and _60417_ (_09417_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [6]);
  and _60418_ (_09418_, _09417_, _09416_);
  nor _60419_ (_09419_, _09417_, _09416_);
  nor _60420_ (_09420_, _09419_, _09418_);
  and _60421_ (_09421_, _09420_, _09384_);
  nor _60422_ (_09422_, _09420_, _09384_);
  nor _60423_ (_09423_, _09422_, _09421_);
  and _60424_ (_09424_, _09423_, _09392_);
  nor _60425_ (_09425_, _09423_, _09392_);
  nor _60426_ (_09426_, _09425_, _09424_);
  and _60427_ (_09427_, _09426_, _09383_);
  nor _60428_ (_09428_, _09426_, _09383_);
  nor _60429_ (_09429_, _09428_, _09427_);
  and _60430_ (_09430_, _09429_, _09402_);
  nor _60431_ (_09431_, _09429_, _09402_);
  nor _60432_ (_09432_, _09431_, _09430_);
  and _60433_ (_09433_, _09432_, _09415_);
  nor _60434_ (_09434_, _09432_, _09415_);
  nor _60435_ (_09435_, _09434_, _09433_);
  not _60436_ (_09436_, _09435_);
  nor _60437_ (_09437_, _09436_, _09413_);
  and _60438_ (_09438_, _09436_, _09413_);
  nor _60439_ (_09439_, _09438_, _09437_);
  and _60440_ (_09440_, _09439_, _09412_);
  nor _60441_ (_09441_, _09433_, _09430_);
  nor _60442_ (_09442_, _09424_, _09421_);
  not _60443_ (_09443_, _09442_);
  and _60444_ (_09444_, \oc8051_golden_model_1.ACC [6], \oc8051_golden_model_1.B [7]);
  and _60445_ (_09445_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [7]);
  and _60446_ (_09446_, _09445_, _09444_);
  nor _60447_ (_09447_, _09445_, _09444_);
  nor _60448_ (_09448_, _09447_, _09446_);
  and _60449_ (_09449_, _09448_, _09418_);
  nor _60450_ (_09450_, _09448_, _09418_);
  nor _60451_ (_09451_, _09450_, _09449_);
  and _60452_ (_09452_, _09451_, _09427_);
  nor _60453_ (_09453_, _09451_, _09427_);
  nor _60454_ (_09454_, _09453_, _09452_);
  and _60455_ (_09455_, _09454_, _09443_);
  nor _60456_ (_09456_, _09454_, _09443_);
  nor _60457_ (_09457_, _09456_, _09455_);
  not _60458_ (_09458_, _09457_);
  nor _60459_ (_09459_, _09458_, _09441_);
  and _60460_ (_09460_, _09458_, _09441_);
  nor _60461_ (_09461_, _09460_, _09459_);
  and _60462_ (_09462_, _09461_, _09437_);
  nor _60463_ (_09463_, _09461_, _09437_);
  nor _60464_ (_09464_, _09463_, _09462_);
  and _60465_ (_09465_, _09464_, _09440_);
  nor _60466_ (_09466_, _09464_, _09440_);
  and _60467_ (_09467_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  and _60468_ (_09468_, _09467_, _09280_);
  and _60469_ (_09469_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [2]);
  and _60470_ (_09470_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [1]);
  nor _60471_ (_09471_, _09470_, _09276_);
  nor _60472_ (_09472_, _09471_, _09468_);
  and _60473_ (_09473_, _09472_, _09469_);
  nor _60474_ (_09474_, _09473_, _09468_);
  not _60475_ (_09475_, _09474_);
  nor _60476_ (_09476_, _09282_, _09278_);
  nor _60477_ (_09477_, _09476_, _09283_);
  and _60478_ (_09478_, _09477_, _09475_);
  and _60479_ (_09479_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [2]);
  and _60480_ (_09480_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [3]);
  and _60481_ (_09481_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [3]);
  and _60482_ (_09482_, _09481_, _09480_);
  nor _60483_ (_09483_, _09481_, _09480_);
  nor _60484_ (_09484_, _09483_, _09482_);
  and _60485_ (_09485_, _09484_, _09479_);
  nor _60486_ (_09486_, _09484_, _09479_);
  nor _60487_ (_09487_, _09486_, _09485_);
  nor _60488_ (_09488_, _09477_, _09475_);
  nor _60489_ (_09489_, _09488_, _09478_);
  and _60490_ (_09490_, _09489_, _09487_);
  nor _60491_ (_09491_, _09490_, _09478_);
  nor _60492_ (_09492_, _09302_, _09300_);
  nor _60493_ (_09493_, _09492_, _09303_);
  not _60494_ (_09494_, _09493_);
  nor _60495_ (_09495_, _09494_, _09491_);
  and _60496_ (_09496_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.ACC [0]);
  and _60497_ (_09497_, _09496_, _09323_);
  nor _60498_ (_09498_, _09485_, _09482_);
  nor _60499_ (_09499_, _09323_, _09322_);
  nor _60500_ (_09500_, _09499_, _09324_);
  not _60501_ (_09501_, _09500_);
  nor _60502_ (_09502_, _09501_, _09498_);
  and _60503_ (_09503_, _09501_, _09498_);
  nor _60504_ (_09504_, _09503_, _09502_);
  and _60505_ (_09505_, _09504_, _09497_);
  nor _60506_ (_09506_, _09504_, _09497_);
  nor _60507_ (_09507_, _09506_, _09505_);
  and _60508_ (_09508_, _09494_, _09491_);
  nor _60509_ (_09509_, _09508_, _09495_);
  and _60510_ (_09510_, _09509_, _09507_);
  nor _60511_ (_09511_, _09510_, _09495_);
  nor _60512_ (_09512_, _09339_, _09337_);
  nor _60513_ (_09513_, _09512_, _09340_);
  not _60514_ (_09514_, _09513_);
  nor _60515_ (_09515_, _09514_, _09511_);
  nor _60516_ (_09516_, _09505_, _09502_);
  not _60517_ (_09517_, _09516_);
  and _60518_ (_09518_, _09514_, _09511_);
  nor _60519_ (_09520_, _09518_, _09515_);
  and _60520_ (_09521_, _09520_, _09517_);
  nor _60521_ (_09522_, _09521_, _09515_);
  nor _60522_ (_09523_, _09376_, _09374_);
  nor _60523_ (_09524_, _09523_, _09377_);
  not _60524_ (_09525_, _09524_);
  nor _60525_ (_09526_, _09525_, _09522_);
  and _60526_ (_09527_, _09411_, _09378_);
  nor _60527_ (_09528_, _09527_, _09412_);
  and _60528_ (_09529_, _09528_, _09526_);
  nor _60529_ (_09530_, _09439_, _09412_);
  nor _60530_ (_09531_, _09530_, _09440_);
  nand _60531_ (_09532_, _09531_, _09529_);
  and _60532_ (_09533_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [1]);
  and _60533_ (_09534_, _09533_, _09467_);
  and _60534_ (_09535_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [3]);
  nor _60535_ (_09536_, _09533_, _09467_);
  nor _60536_ (_09537_, _09536_, _09534_);
  and _60537_ (_09538_, _09537_, _09535_);
  nor _60538_ (_09539_, _09538_, _09534_);
  not _60539_ (_09541_, _09539_);
  nor _60540_ (_09542_, _09472_, _09469_);
  nor _60541_ (_09543_, _09542_, _09473_);
  and _60542_ (_09544_, _09543_, _09541_);
  and _60543_ (_09545_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [5]);
  and _60544_ (_09546_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [3]);
  and _60545_ (_09547_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [2]);
  and _60546_ (_09548_, _09547_, _09546_);
  nor _60547_ (_09549_, _09547_, _09546_);
  nor _60548_ (_09550_, _09549_, _09548_);
  and _60549_ (_09551_, _09550_, _09545_);
  nor _60550_ (_09552_, _09550_, _09545_);
  nor _60551_ (_09553_, _09552_, _09551_);
  nor _60552_ (_09554_, _09543_, _09541_);
  nor _60553_ (_09555_, _09554_, _09544_);
  and _60554_ (_09556_, _09555_, _09553_);
  nor _60555_ (_09557_, _09556_, _09544_);
  not _60556_ (_09558_, _09557_);
  nor _60557_ (_09559_, _09489_, _09487_);
  nor _60558_ (_09560_, _09559_, _09490_);
  and _60559_ (_09561_, _09560_, _09558_);
  nor _60560_ (_09562_, _09551_, _09548_);
  and _60561_ (_09563_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [6]);
  and _60562_ (_09564_, \oc8051_golden_model_1.ACC [0], \oc8051_golden_model_1.B [7]);
  nor _60563_ (_09565_, _09564_, _09563_);
  nor _60564_ (_09566_, _09565_, _09497_);
  not _60565_ (_09567_, _09566_);
  nor _60566_ (_09568_, _09567_, _09562_);
  and _60567_ (_09569_, _09567_, _09562_);
  nor _60568_ (_09570_, _09569_, _09568_);
  nor _60569_ (_09571_, _09560_, _09558_);
  nor _60570_ (_09572_, _09571_, _09561_);
  and _60571_ (_09573_, _09572_, _09570_);
  nor _60572_ (_09574_, _09573_, _09561_);
  nor _60573_ (_09575_, _09509_, _09507_);
  nor _60574_ (_09576_, _09575_, _09510_);
  not _60575_ (_09577_, _09576_);
  nor _60576_ (_09578_, _09577_, _09574_);
  and _60577_ (_09579_, _09577_, _09574_);
  nor _60578_ (_09580_, _09579_, _09578_);
  and _60579_ (_09581_, _09580_, _09568_);
  nor _60580_ (_09582_, _09581_, _09578_);
  nor _60581_ (_09583_, _09520_, _09517_);
  nor _60582_ (_09584_, _09583_, _09521_);
  not _60583_ (_09585_, _09584_);
  nor _60584_ (_09586_, _09585_, _09582_);
  and _60585_ (_09587_, _09525_, _09522_);
  nor _60586_ (_09588_, _09587_, _09526_);
  and _60587_ (_09589_, _09588_, _09586_);
  nor _60588_ (_09590_, _09528_, _09526_);
  nor _60589_ (_09591_, _09590_, _09529_);
  and _60590_ (_09592_, _09591_, _09589_);
  nor _60591_ (_09593_, _09591_, _09589_);
  nor _60592_ (_09594_, _09593_, _09592_);
  and _60593_ (_09595_, \oc8051_golden_model_1.ACC [4], \oc8051_golden_model_1.B [0]);
  and _60594_ (_09596_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [3]);
  and _60595_ (_09597_, _09596_, _09595_);
  and _60596_ (_09598_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [2]);
  nor _60597_ (_09599_, _09596_, _09595_);
  nor _60598_ (_09600_, _09599_, _09597_);
  and _60599_ (_09601_, _09600_, _09598_);
  nor _60600_ (_09602_, _09601_, _09597_);
  not _60601_ (_09603_, _09602_);
  nor _60602_ (_09604_, _09537_, _09535_);
  nor _60603_ (_09605_, _09604_, _09538_);
  and _60604_ (_09606_, _09605_, _09603_);
  and _60605_ (_09607_, \oc8051_golden_model_1.B [5], \oc8051_golden_model_1.ACC [0]);
  and _60606_ (_09608_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [2]);
  and _60607_ (_09609_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [4]);
  and _60608_ (_09610_, _09609_, _09608_);
  nor _60609_ (_09611_, _09609_, _09608_);
  nor _60610_ (_09612_, _09611_, _09610_);
  and _60611_ (_09613_, _09612_, _09607_);
  nor _60612_ (_09614_, _09612_, _09607_);
  nor _60613_ (_09615_, _09614_, _09613_);
  nor _60614_ (_09616_, _09605_, _09603_);
  nor _60615_ (_09617_, _09616_, _09606_);
  and _60616_ (_09618_, _09617_, _09615_);
  nor _60617_ (_09619_, _09618_, _09606_);
  not _60618_ (_09620_, _09619_);
  nor _60619_ (_09621_, _09555_, _09553_);
  nor _60620_ (_09622_, _09621_, _09556_);
  and _60621_ (_09623_, _09622_, _09620_);
  not _60622_ (_09624_, _09496_);
  nor _60623_ (_09625_, _09613_, _09610_);
  nor _60624_ (_09626_, _09625_, _09624_);
  and _60625_ (_09627_, _09625_, _09624_);
  nor _60626_ (_09628_, _09627_, _09626_);
  nor _60627_ (_09629_, _09622_, _09620_);
  nor _60628_ (_09630_, _09629_, _09623_);
  and _60629_ (_09631_, _09630_, _09628_);
  nor _60630_ (_09632_, _09631_, _09623_);
  not _60631_ (_09633_, _09632_);
  nor _60632_ (_09634_, _09572_, _09570_);
  nor _60633_ (_09635_, _09634_, _09573_);
  and _60634_ (_09636_, _09635_, _09633_);
  nor _60635_ (_09637_, _09635_, _09633_);
  nor _60636_ (_09638_, _09637_, _09636_);
  and _60637_ (_09639_, _09638_, _09626_);
  nor _60638_ (_09640_, _09639_, _09636_);
  nor _60639_ (_09641_, _09580_, _09568_);
  nor _60640_ (_09642_, _09641_, _09581_);
  not _60641_ (_09643_, _09642_);
  nor _60642_ (_09644_, _09643_, _09640_);
  and _60643_ (_09645_, _09585_, _09582_);
  nor _60644_ (_09646_, _09645_, _09586_);
  and _60645_ (_09647_, _09646_, _09644_);
  nor _60646_ (_09648_, _09588_, _09586_);
  nor _60647_ (_09649_, _09648_, _09589_);
  nand _60648_ (_09650_, _09649_, _09647_);
  or _60649_ (_09651_, _09649_, _09647_);
  and _60650_ (_09652_, _09651_, _09650_);
  and _60651_ (_09653_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  and _60652_ (_09654_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [2]);
  and _60653_ (_09655_, _09654_, _09653_);
  and _60654_ (_09656_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [2]);
  nor _60655_ (_09657_, _09654_, _09653_);
  nor _60656_ (_09658_, _09657_, _09655_);
  and _60657_ (_09659_, _09658_, _09656_);
  nor _60658_ (_09660_, _09659_, _09655_);
  not _60659_ (_09661_, _09660_);
  nor _60660_ (_09662_, _09600_, _09598_);
  nor _60661_ (_09663_, _09662_, _09601_);
  and _60662_ (_09664_, _09663_, _09661_);
  and _60663_ (_09665_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.ACC [0]);
  and _60664_ (_09666_, _09665_, _09609_);
  and _60665_ (_09667_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [3]);
  and _60666_ (_09668_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.ACC [0]);
  nor _60667_ (_09669_, _09668_, _09667_);
  nor _60668_ (_09670_, _09669_, _09666_);
  nor _60669_ (_09671_, _09663_, _09661_);
  nor _60670_ (_09672_, _09671_, _09664_);
  and _60671_ (_09673_, _09672_, _09670_);
  nor _60672_ (_09674_, _09673_, _09664_);
  not _60673_ (_09675_, _09674_);
  nor _60674_ (_09676_, _09617_, _09615_);
  nor _60675_ (_09677_, _09676_, _09618_);
  and _60676_ (_09678_, _09677_, _09675_);
  nor _60677_ (_09679_, _09677_, _09675_);
  nor _60678_ (_09680_, _09679_, _09678_);
  and _60679_ (_09681_, _09680_, _09666_);
  nor _60680_ (_09682_, _09681_, _09678_);
  not _60681_ (_09683_, _09682_);
  nor _60682_ (_09684_, _09630_, _09628_);
  nor _60683_ (_09685_, _09684_, _09631_);
  and _60684_ (_09686_, _09685_, _09683_);
  nor _60685_ (_09687_, _09638_, _09626_);
  nor _60686_ (_09688_, _09687_, _09639_);
  and _60687_ (_09689_, _09688_, _09686_);
  and _60688_ (_09690_, _09643_, _09640_);
  nor _60689_ (_09691_, _09690_, _09644_);
  and _60690_ (_09692_, _09691_, _09689_);
  nor _60691_ (_09693_, _09646_, _09644_);
  nor _60692_ (_09694_, _09693_, _09647_);
  and _60693_ (_09696_, _09694_, _09692_);
  nor _60694_ (_09697_, _09694_, _09692_);
  nor _60695_ (_09699_, _09697_, _09696_);
  and _60696_ (_09700_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [2]);
  and _60697_ (_09702_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [1]);
  and _60698_ (_09703_, _09702_, _09700_);
  and _60699_ (_09705_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.ACC [0]);
  nor _60700_ (_09706_, _09702_, _09700_);
  nor _60701_ (_09708_, _09706_, _09703_);
  and _60702_ (_09709_, _09708_, _09705_);
  nor _60703_ (_09711_, _09709_, _09703_);
  not _60704_ (_09712_, _09711_);
  nor _60705_ (_09714_, _09658_, _09656_);
  nor _60706_ (_09715_, _09714_, _09659_);
  and _60707_ (_09717_, _09715_, _09712_);
  nor _60708_ (_09718_, _09715_, _09712_);
  nor _60709_ (_09720_, _09718_, _09717_);
  and _60710_ (_09721_, _09720_, _09665_);
  nor _60711_ (_09723_, _09721_, _09717_);
  not _60712_ (_09724_, _09723_);
  nor _60713_ (_09726_, _09672_, _09670_);
  nor _60714_ (_09727_, _09726_, _09673_);
  and _60715_ (_09729_, _09727_, _09724_);
  nor _60716_ (_09730_, _09680_, _09666_);
  nor _60717_ (_09732_, _09730_, _09681_);
  and _60718_ (_09733_, _09732_, _09729_);
  nor _60719_ (_09734_, _09685_, _09683_);
  nor _60720_ (_09735_, _09734_, _09686_);
  and _60721_ (_09736_, _09735_, _09733_);
  nor _60722_ (_09737_, _09688_, _09686_);
  nor _60723_ (_09738_, _09737_, _09689_);
  and _60724_ (_09739_, _09738_, _09736_);
  nor _60725_ (_09740_, _09691_, _09689_);
  nor _60726_ (_09741_, _09740_, _09692_);
  and _60727_ (_09742_, _09741_, _09739_);
  and _60728_ (_09743_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  and _60729_ (_09744_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.ACC [0]);
  and _60730_ (_09745_, _09744_, _09743_);
  nor _60731_ (_09746_, _09708_, _09705_);
  nor _60732_ (_09747_, _09746_, _09709_);
  and _60733_ (_09748_, _09747_, _09745_);
  nor _60734_ (_09749_, _09720_, _09665_);
  nor _60735_ (_09750_, _09749_, _09721_);
  and _60736_ (_09751_, _09750_, _09748_);
  nor _60737_ (_09752_, _09727_, _09724_);
  nor _60738_ (_09753_, _09752_, _09729_);
  and _60739_ (_09754_, _09753_, _09751_);
  nor _60740_ (_09755_, _09732_, _09729_);
  nor _60741_ (_09756_, _09755_, _09733_);
  and _60742_ (_09757_, _09756_, _09754_);
  nor _60743_ (_09758_, _09735_, _09733_);
  nor _60744_ (_09759_, _09758_, _09736_);
  and _60745_ (_09760_, _09759_, _09757_);
  nor _60746_ (_09761_, _09738_, _09736_);
  nor _60747_ (_09762_, _09761_, _09739_);
  and _60748_ (_09763_, _09762_, _09760_);
  nor _60749_ (_09764_, _09741_, _09739_);
  nor _60750_ (_09765_, _09764_, _09742_);
  and _60751_ (_09766_, _09765_, _09763_);
  nor _60752_ (_09767_, _09766_, _09742_);
  not _60753_ (_09768_, _09767_);
  and _60754_ (_09769_, _09768_, _09699_);
  or _60755_ (_09770_, _09769_, _09696_);
  nand _60756_ (_09771_, _09770_, _09652_);
  and _60757_ (_09772_, _09771_, _09650_);
  not _60758_ (_09773_, _09772_);
  and _60759_ (_09774_, _09773_, _09594_);
  or _60760_ (_09775_, _09774_, _09592_);
  or _60761_ (_09776_, _09531_, _09529_);
  and _60762_ (_09777_, _09776_, _09532_);
  nand _60763_ (_09778_, _09777_, _09775_);
  and _60764_ (_09779_, _09778_, _09532_);
  nor _60765_ (_09780_, _09779_, _09466_);
  or _60766_ (_09781_, _09780_, _09465_);
  and _60767_ (_09782_, \oc8051_golden_model_1.ACC [7], \oc8051_golden_model_1.B [7]);
  not _60768_ (_09783_, _09782_);
  nor _60769_ (_09784_, _09783_, _09417_);
  nor _60770_ (_09785_, _09784_, _09449_);
  nor _60771_ (_09786_, _09455_, _09452_);
  nor _60772_ (_09787_, _09786_, _09785_);
  and _60773_ (_09788_, _09786_, _09785_);
  nor _60774_ (_09789_, _09788_, _09787_);
  not _60775_ (_09791_, _09789_);
  nor _60776_ (_09793_, _09462_, _09459_);
  and _60777_ (_09794_, _09793_, _09791_);
  nor _60778_ (_09796_, _09793_, _09791_);
  nor _60779_ (_09797_, _09796_, _09794_);
  and _60780_ (_09799_, _09797_, _09781_);
  not _60781_ (_09800_, _09269_);
  or _60782_ (_09802_, _09787_, _09446_);
  or _60783_ (_09803_, _09802_, _09796_);
  or _60784_ (_09805_, _09803_, _09800_);
  or _60785_ (_09806_, _09805_, _09799_);
  and _60786_ (_09808_, _09806_, _06027_);
  and _60787_ (_09809_, _09808_, _09274_);
  and _60788_ (_09811_, _08376_, _08361_);
  or _60789_ (_09812_, _09811_, _09238_);
  and _60790_ (_09814_, _09812_, _06026_);
  and _60791_ (_09815_, _05659_, _05567_);
  nor _60792_ (_09817_, _09815_, _07011_);
  not _60793_ (_09818_, _09817_);
  or _60794_ (_09820_, _09818_, _09814_);
  or _60795_ (_09821_, _09820_, _09809_);
  and _60796_ (_09823_, _08485_, _07698_);
  or _60797_ (_09824_, _09234_, _07012_);
  or _60798_ (_09826_, _09824_, _09823_);
  not _60799_ (_09827_, _09815_);
  or _60800_ (_09828_, _09827_, _09260_);
  and _60801_ (_09829_, _09828_, _05669_);
  and _60802_ (_09830_, _09829_, _09826_);
  and _60803_ (_09831_, _09830_, _09821_);
  and _60804_ (_09832_, _06114_, _05659_);
  not _60805_ (_09833_, _05669_);
  and _60806_ (_09834_, _08738_, _07698_);
  or _60807_ (_09835_, _09834_, _09234_);
  and _60808_ (_09836_, _09835_, _09833_);
  or _60809_ (_09837_, _09836_, _09832_);
  or _60810_ (_09838_, _09837_, _09831_);
  not _60811_ (_09839_, _09832_);
  nor _60812_ (_09840_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [7]);
  nor _60813_ (_09841_, _09840_, _09279_);
  not _60814_ (_09842_, \oc8051_golden_model_1.B [1]);
  nor _60815_ (_09843_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [5]);
  nor _60816_ (_09844_, \oc8051_golden_model_1.B [4], \oc8051_golden_model_1.B [3]);
  and _60817_ (_09845_, _09844_, _09843_);
  and _60818_ (_09846_, _09845_, _09842_);
  nor _60819_ (_09847_, \oc8051_golden_model_1.B [2], \oc8051_golden_model_1.B [7]);
  not _60820_ (_09848_, _09847_);
  and _60821_ (_09849_, \oc8051_golden_model_1.B [0], _08393_);
  nor _60822_ (_09850_, _09849_, _09848_);
  and _60823_ (_09851_, _09850_, _09846_);
  and _60824_ (_09852_, _09851_, _09841_);
  or _60825_ (_09853_, _09851_, _08393_);
  not _60826_ (_09854_, \oc8051_golden_model_1.B [4]);
  not _60827_ (_09855_, \oc8051_golden_model_1.B [5]);
  nor _60828_ (_09856_, \oc8051_golden_model_1.B [6], \oc8051_golden_model_1.B [7]);
  and _60829_ (_09857_, _09856_, _09855_);
  and _60830_ (_09858_, _09857_, _09854_);
  nor _60831_ (_09859_, \oc8051_golden_model_1.B [3], \oc8051_golden_model_1.B [2]);
  and _60832_ (_09860_, _09859_, _09858_);
  not _60833_ (_09861_, \oc8051_golden_model_1.ACC [6]);
  and _60834_ (_09862_, \oc8051_golden_model_1.B [0], _09861_);
  nor _60835_ (_09863_, _09862_, _08393_);
  nor _60836_ (_09864_, _09863_, _09842_);
  not _60837_ (_09865_, _09864_);
  and _60838_ (_09866_, _09865_, _09860_);
  nor _60839_ (_09867_, _09866_, _09853_);
  nor _60840_ (_09868_, _09867_, _09852_);
  and _60841_ (_09869_, _09866_, \oc8051_golden_model_1.B [0]);
  nor _60842_ (_09870_, _09869_, _09861_);
  and _60843_ (_09871_, _09870_, _09842_);
  nor _60844_ (_09872_, _09870_, _09842_);
  nor _60845_ (_09873_, _09872_, _09871_);
  nor _60846_ (_09874_, \oc8051_golden_model_1.ACC [5], \oc8051_golden_model_1.B [0]);
  nor _60847_ (_09875_, _09874_, _09467_);
  nor _60848_ (_09876_, _09875_, \oc8051_golden_model_1.ACC [4]);
  not _60849_ (_09877_, \oc8051_golden_model_1.B [0]);
  and _60850_ (_09878_, \oc8051_golden_model_1.ACC [4], _09877_);
  nor _60851_ (_09879_, _09878_, \oc8051_golden_model_1.ACC [5]);
  not _60852_ (_09880_, \oc8051_golden_model_1.ACC [4]);
  and _60853_ (_09881_, _09880_, \oc8051_golden_model_1.B [0]);
  nor _60854_ (_09882_, _09881_, _09879_);
  nor _60855_ (_09883_, _09882_, _09876_);
  not _60856_ (_09884_, _09883_);
  and _60857_ (_09885_, _09884_, _09873_);
  nor _60858_ (_09886_, _09868_, \oc8051_golden_model_1.B [2]);
  nor _60859_ (_09887_, _09886_, _09871_);
  not _60860_ (_09888_, _09887_);
  nor _60861_ (_09889_, _09888_, _09885_);
  not _60862_ (_09890_, _09889_);
  and _60863_ (_09891_, \oc8051_golden_model_1.B [2], _08393_);
  nor _60864_ (_09892_, _09891_, \oc8051_golden_model_1.B [7]);
  and _60865_ (_09893_, _09892_, _09845_);
  and _60866_ (_09894_, _09893_, _09890_);
  nor _60867_ (_09895_, _09894_, _09868_);
  nor _60868_ (_09896_, _09895_, _09852_);
  nor _60869_ (_09897_, _09884_, _09873_);
  nor _60870_ (_09898_, _09897_, _09885_);
  and _60871_ (_09899_, _09898_, _09894_);
  not _60872_ (_09900_, _09870_);
  nor _60873_ (_09901_, _09894_, _09900_);
  nor _60874_ (_09902_, _09901_, _09899_);
  nor _60875_ (_09903_, _09902_, \oc8051_golden_model_1.B [2]);
  and _60876_ (_09904_, _09902_, \oc8051_golden_model_1.B [2]);
  nor _60877_ (_09905_, _09904_, _09903_);
  not _60878_ (_09906_, \oc8051_golden_model_1.ACC [5]);
  nor _60879_ (_09907_, _09894_, _09906_);
  and _60880_ (_09908_, _09894_, _09875_);
  or _60881_ (_09909_, _09908_, _09907_);
  and _60882_ (_09910_, _09909_, _09842_);
  nor _60883_ (_09911_, _09909_, _09842_);
  nor _60884_ (_09912_, _09911_, _09881_);
  nor _60885_ (_09913_, _09912_, _09910_);
  not _60886_ (_09914_, _09913_);
  and _60887_ (_09915_, _09914_, _09905_);
  nor _60888_ (_09916_, _09896_, \oc8051_golden_model_1.B [3]);
  nor _60889_ (_09917_, _09916_, _09903_);
  not _60890_ (_09918_, _09917_);
  nor _60891_ (_09919_, _09918_, _09915_);
  not _60892_ (_09920_, _09919_);
  and _60893_ (_09921_, \oc8051_golden_model_1.B [3], _08393_);
  not _60894_ (_09922_, _09921_);
  and _60895_ (_09923_, _09922_, _09858_);
  and _60896_ (_09924_, _09923_, _09920_);
  nor _60897_ (_09925_, _09924_, _09896_);
  nor _60898_ (_09926_, _09925_, _09852_);
  not _60899_ (_09927_, \oc8051_golden_model_1.B [3]);
  nor _60900_ (_09928_, _09924_, _09902_);
  nor _60901_ (_09929_, _09914_, _09905_);
  nor _60902_ (_09930_, _09929_, _09915_);
  and _60903_ (_09931_, _09930_, _09924_);
  or _60904_ (_09932_, _09931_, _09928_);
  and _60905_ (_09933_, _09932_, _09927_);
  nor _60906_ (_09934_, _09932_, _09927_);
  nor _60907_ (_09935_, _09934_, _09933_);
  not _60908_ (_09936_, _09935_);
  nor _60909_ (_09937_, _09924_, _09909_);
  nor _60910_ (_09938_, _09911_, _09910_);
  and _60911_ (_09939_, _09938_, _09881_);
  nor _60912_ (_09940_, _09938_, _09881_);
  nor _60913_ (_09941_, _09940_, _09939_);
  and _60914_ (_09942_, _09941_, _09924_);
  or _60915_ (_09943_, _09942_, _09937_);
  nor _60916_ (_09944_, _09943_, \oc8051_golden_model_1.B [2]);
  and _60917_ (_09945_, _09943_, \oc8051_golden_model_1.B [2]);
  nor _60918_ (_09946_, _09881_, _09878_);
  and _60919_ (_09947_, _09924_, _09946_);
  nor _60920_ (_09948_, _09924_, \oc8051_golden_model_1.ACC [4]);
  nor _60921_ (_09949_, _09948_, _09947_);
  and _60922_ (_09950_, _09949_, _09842_);
  nor _60923_ (_09951_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [3]);
  nor _60924_ (_09952_, _09951_, _09653_);
  nor _60925_ (_09953_, _09952_, \oc8051_golden_model_1.ACC [2]);
  and _60926_ (_09954_, _09877_, \oc8051_golden_model_1.ACC [2]);
  nor _60927_ (_09955_, _09954_, \oc8051_golden_model_1.ACC [3]);
  not _60928_ (_09956_, \oc8051_golden_model_1.ACC [2]);
  and _60929_ (_09957_, \oc8051_golden_model_1.B [0], _09956_);
  nor _60930_ (_09958_, _09957_, _09955_);
  nor _60931_ (_09959_, _09958_, _09953_);
  not _60932_ (_09960_, _09959_);
  nor _60933_ (_09961_, _09949_, _09842_);
  nor _60934_ (_09962_, _09961_, _09950_);
  and _60935_ (_09963_, _09962_, _09960_);
  nor _60936_ (_09964_, _09963_, _09950_);
  nor _60937_ (_09965_, _09964_, _09945_);
  nor _60938_ (_09966_, _09965_, _09944_);
  nor _60939_ (_09967_, _09966_, _09936_);
  nor _60940_ (_09968_, _09926_, \oc8051_golden_model_1.B [4]);
  nor _60941_ (_09969_, _09968_, _09933_);
  not _60942_ (_09970_, _09969_);
  nor _60943_ (_09971_, _09970_, _09967_);
  not _60944_ (_09972_, _09857_);
  and _60945_ (_09973_, \oc8051_golden_model_1.B [4], _08393_);
  nor _60946_ (_09974_, _09973_, _09972_);
  not _60947_ (_09975_, _09974_);
  nor _60948_ (_09976_, _09975_, _09971_);
  nor _60949_ (_09977_, _09976_, _09926_);
  nor _60950_ (_09978_, _09977_, _09852_);
  and _60951_ (_09979_, _09856_, \oc8051_golden_model_1.ACC [7]);
  nor _60952_ (_09980_, _09979_, _09857_);
  nor _60953_ (_09981_, _09978_, \oc8051_golden_model_1.B [5]);
  and _60954_ (_09982_, _09966_, _09936_);
  nor _60955_ (_09983_, _09982_, _09967_);
  not _60956_ (_09984_, _09983_);
  and _60957_ (_09985_, _09984_, _09976_);
  nor _60958_ (_09986_, _09976_, _09932_);
  nor _60959_ (_09987_, _09986_, _09985_);
  and _60960_ (_09988_, _09987_, _09854_);
  nor _60961_ (_09989_, _09987_, _09854_);
  nor _60962_ (_09990_, _09989_, _09988_);
  not _60963_ (_09991_, _09990_);
  nor _60964_ (_09992_, _09976_, _09943_);
  nor _60965_ (_09993_, _09945_, _09944_);
  and _60966_ (_09994_, _09993_, _09964_);
  nor _60967_ (_09995_, _09993_, _09964_);
  nor _60968_ (_09996_, _09995_, _09994_);
  not _60969_ (_09997_, _09996_);
  and _60970_ (_09998_, _09997_, _09976_);
  nor _60971_ (_09999_, _09998_, _09992_);
  nor _60972_ (_10000_, _09999_, \oc8051_golden_model_1.B [3]);
  and _60973_ (_10001_, _09999_, \oc8051_golden_model_1.B [3]);
  not _60974_ (_10002_, \oc8051_golden_model_1.B [2]);
  nor _60975_ (_10003_, _09962_, _09960_);
  nor _60976_ (_10004_, _10003_, _09963_);
  not _60977_ (_10005_, _10004_);
  and _60978_ (_10006_, _10005_, _09976_);
  nor _60979_ (_10007_, _09976_, _09949_);
  nor _60980_ (_10008_, _10007_, _10006_);
  and _60981_ (_10009_, _10008_, _10002_);
  not _60982_ (_10010_, \oc8051_golden_model_1.ACC [3]);
  nor _60983_ (_10011_, _09976_, _10010_);
  and _60984_ (_10012_, _09976_, _09952_);
  or _60985_ (_10013_, _10012_, _10011_);
  and _60986_ (_10014_, _10013_, _09842_);
  nor _60987_ (_10015_, _10013_, _09842_);
  nor _60988_ (_10016_, _10015_, _09957_);
  nor _60989_ (_10017_, _10016_, _10014_);
  nor _60990_ (_10018_, _10008_, _10002_);
  nor _60991_ (_10019_, _10018_, _10009_);
  not _60992_ (_10020_, _10019_);
  nor _60993_ (_10021_, _10020_, _10017_);
  nor _60994_ (_10022_, _10021_, _10009_);
  nor _60995_ (_10023_, _10022_, _10001_);
  nor _60996_ (_10024_, _10023_, _10000_);
  nor _60997_ (_10025_, _10024_, _09991_);
  or _60998_ (_10026_, _10025_, _09988_);
  nor _60999_ (_10027_, _10026_, _09981_);
  nor _61000_ (_10028_, _10027_, _09980_);
  nor _61001_ (_10029_, _10028_, _09978_);
  nor _61002_ (_10030_, _10029_, _09852_);
  not _61003_ (_10031_, _10028_);
  and _61004_ (_10032_, _10024_, _09991_);
  nor _61005_ (_10033_, _10032_, _10025_);
  nor _61006_ (_10034_, _10033_, _10031_);
  nor _61007_ (_10035_, _10028_, _09987_);
  nor _61008_ (_10036_, _10035_, _10034_);
  and _61009_ (_10037_, _10036_, _09855_);
  nor _61010_ (_10038_, _10036_, _09855_);
  nor _61011_ (_10039_, _10038_, _10037_);
  nor _61012_ (_10040_, _10028_, _09999_);
  nor _61013_ (_10041_, _10001_, _10000_);
  nor _61014_ (_10042_, _10041_, _10022_);
  and _61015_ (_10043_, _10041_, _10022_);
  or _61016_ (_10044_, _10043_, _10042_);
  and _61017_ (_10045_, _10044_, _10028_);
  or _61018_ (_10046_, _10045_, _10040_);
  and _61019_ (_10047_, _10046_, _09854_);
  nor _61020_ (_10048_, _10046_, _09854_);
  and _61021_ (_10049_, _10020_, _10017_);
  nor _61022_ (_10050_, _10049_, _10021_);
  nor _61023_ (_10051_, _10050_, _10031_);
  nor _61024_ (_10052_, _10028_, _10008_);
  nor _61025_ (_10053_, _10052_, _10051_);
  and _61026_ (_10054_, _10053_, _09927_);
  nor _61027_ (_10055_, _10015_, _10014_);
  nor _61028_ (_10056_, _10055_, _09957_);
  and _61029_ (_10057_, _10055_, _09957_);
  or _61030_ (_10058_, _10057_, _10056_);
  nor _61031_ (_10059_, _10058_, _10031_);
  nor _61032_ (_10060_, _10028_, _10013_);
  nor _61033_ (_10061_, _10060_, _10059_);
  and _61034_ (_10062_, _10061_, _10002_);
  nor _61035_ (_10063_, _10061_, _10002_);
  nor _61036_ (_10064_, _10028_, \oc8051_golden_model_1.ACC [2]);
  nor _61037_ (_10065_, _09957_, _09954_);
  and _61038_ (_10066_, _10028_, _10065_);
  nor _61039_ (_10067_, _10066_, _10064_);
  and _61040_ (_10068_, _10067_, _09842_);
  and _61041_ (_10069_, _05784_, \oc8051_golden_model_1.B [0]);
  not _61042_ (_10070_, _10069_);
  nor _61043_ (_10071_, _10067_, _09842_);
  nor _61044_ (_10072_, _10071_, _10068_);
  and _61045_ (_10073_, _10072_, _10070_);
  nor _61046_ (_10074_, _10073_, _10068_);
  nor _61047_ (_10075_, _10074_, _10063_);
  nor _61048_ (_10076_, _10075_, _10062_);
  not _61049_ (_10077_, _10076_);
  nor _61050_ (_10078_, _10053_, _09927_);
  nor _61051_ (_10079_, _10078_, _10054_);
  and _61052_ (_10080_, _10079_, _10077_);
  nor _61053_ (_10081_, _10080_, _10054_);
  nor _61054_ (_10082_, _10081_, _10048_);
  nor _61055_ (_10083_, _10082_, _10047_);
  not _61056_ (_10084_, _10083_);
  and _61057_ (_10085_, _10084_, _10039_);
  nor _61058_ (_10086_, _10030_, \oc8051_golden_model_1.B [6]);
  or _61059_ (_10087_, _10086_, _10037_);
  or _61060_ (_10088_, _10087_, _10085_);
  not _61061_ (_10089_, \oc8051_golden_model_1.B [6]);
  or _61062_ (_10090_, _10089_, \oc8051_golden_model_1.ACC [7]);
  and _61063_ (_10091_, _10090_, _09232_);
  and _61064_ (_10092_, _10091_, _10088_);
  nor _61065_ (_10093_, _10092_, _10030_);
  or _61066_ (_10094_, _10093_, _09852_);
  nor _61067_ (_10095_, _10094_, \oc8051_golden_model_1.B [7]);
  nor _61068_ (_10096_, _10095_, _09782_);
  nor _61069_ (_10097_, _10084_, _10039_);
  nor _61070_ (_10098_, _10097_, _10085_);
  and _61071_ (_10099_, _10098_, _10092_);
  not _61072_ (_10100_, _10036_);
  nor _61073_ (_10101_, _10092_, _10100_);
  nor _61074_ (_10102_, _10101_, _10099_);
  and _61075_ (_10103_, _10102_, \oc8051_golden_model_1.B [6]);
  not _61076_ (_10104_, _10103_);
  nor _61077_ (_10105_, _10104_, _10096_);
  nor _61078_ (_10106_, _10063_, _10062_);
  or _61079_ (_10107_, _10106_, _10074_);
  nand _61080_ (_10108_, _10106_, _10074_);
  and _61081_ (_10109_, _10108_, _10107_);
  and _61082_ (_10110_, _10109_, _10092_);
  nor _61083_ (_10111_, _10092_, _10061_);
  nor _61084_ (_10112_, _10111_, _10110_);
  and _61085_ (_10113_, _10112_, _09927_);
  nor _61086_ (_10114_, _10112_, _09927_);
  nor _61087_ (_10115_, _10114_, _10113_);
  nor _61088_ (_10116_, _10072_, _10070_);
  nor _61089_ (_10117_, _10116_, _10073_);
  and _61090_ (_10118_, _10117_, _10092_);
  not _61091_ (_10119_, _10067_);
  nor _61092_ (_10120_, _10092_, _10119_);
  nor _61093_ (_10121_, _10120_, _10118_);
  and _61094_ (_10122_, _10121_, \oc8051_golden_model_1.B [2]);
  nor _61095_ (_10123_, _10121_, \oc8051_golden_model_1.B [2]);
  nor _61096_ (_10124_, _10123_, _10122_);
  and _61097_ (_10125_, _10124_, _10115_);
  or _61098_ (_10126_, _10092_, \oc8051_golden_model_1.ACC [1]);
  nor _61099_ (_10127_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.B [0]);
  or _61100_ (_10128_, _10127_, _09743_);
  nand _61101_ (_10129_, _10092_, _10128_);
  and _61102_ (_10130_, _10129_, _10126_);
  and _61103_ (_10131_, _10130_, _09842_);
  nor _61104_ (_10132_, _10130_, _09842_);
  and _61105_ (_10133_, _09877_, \oc8051_golden_model_1.ACC [0]);
  not _61106_ (_10134_, _10133_);
  nor _61107_ (_10135_, _10134_, _10132_);
  nor _61108_ (_10136_, _10135_, _10131_);
  and _61109_ (_10137_, _10136_, _10125_);
  not _61110_ (_10138_, _10137_);
  and _61111_ (_10139_, _10122_, _10115_);
  nor _61112_ (_10140_, _10139_, _10114_);
  and _61113_ (_10141_, _10140_, _10138_);
  nor _61114_ (_10142_, _10079_, _10077_);
  nor _61115_ (_10143_, _10142_, _10080_);
  and _61116_ (_10144_, _10143_, _10092_);
  not _61117_ (_10145_, _10053_);
  nor _61118_ (_10146_, _10092_, _10145_);
  nor _61119_ (_10147_, _10146_, _10144_);
  and _61120_ (_10148_, _10147_, \oc8051_golden_model_1.B [4]);
  nor _61121_ (_10149_, _10147_, \oc8051_golden_model_1.B [4]);
  nor _61122_ (_10150_, _10149_, _10148_);
  nor _61123_ (_10151_, _10048_, _10047_);
  or _61124_ (_10152_, _10151_, _10081_);
  nand _61125_ (_10153_, _10151_, _10081_);
  and _61126_ (_10154_, _10153_, _10152_);
  and _61127_ (_10155_, _10154_, _10092_);
  nor _61128_ (_10156_, _10092_, _10046_);
  nor _61129_ (_10157_, _10156_, _10155_);
  nor _61130_ (_10158_, _10157_, _09855_);
  and _61131_ (_10159_, _10157_, _09855_);
  nor _61132_ (_10160_, _10159_, _10158_);
  and _61133_ (_10161_, _10160_, _10150_);
  nor _61134_ (_10162_, _10102_, \oc8051_golden_model_1.B [6]);
  nor _61135_ (_10163_, _10162_, _10103_);
  not _61136_ (_10164_, _10163_);
  nor _61137_ (_10165_, _10164_, _10096_);
  and _61138_ (_10166_, _10165_, _10161_);
  not _61139_ (_10167_, _10166_);
  nor _61140_ (_10168_, _10167_, _10141_);
  and _61141_ (_10169_, _10030_, \oc8051_golden_model_1.B [7]);
  and _61142_ (_10170_, _10160_, _10148_);
  nor _61143_ (_10171_, _10170_, _10158_);
  not _61144_ (_10172_, _10171_);
  and _61145_ (_10173_, _10172_, _10165_);
  or _61146_ (_10174_, _10173_, _10169_);
  or _61147_ (_10175_, _10174_, _10168_);
  nor _61148_ (_10176_, _10175_, _10105_);
  nor _61149_ (_10177_, _10132_, _10131_);
  and _61150_ (_10178_, \oc8051_golden_model_1.B [0], _05758_);
  not _61151_ (_10179_, _10178_);
  and _61152_ (_10180_, _10179_, _10177_);
  and _61153_ (_10181_, _10180_, _10134_);
  and _61154_ (_10182_, _10181_, _10125_);
  and _61155_ (_10183_, _10182_, _10166_);
  nor _61156_ (_10184_, _10183_, _10176_);
  and _61157_ (_10185_, _10184_, _10094_);
  or _61158_ (_10186_, _10185_, _09852_);
  or _61159_ (_10187_, _10186_, _09839_);
  and _61160_ (_10188_, _10187_, _06020_);
  and _61161_ (_10189_, _10188_, _09838_);
  and _61162_ (_10190_, _08549_, _07698_);
  or _61163_ (_10191_, _10190_, _09234_);
  and _61164_ (_10192_, _10191_, _06019_);
  or _61165_ (_10193_, _10192_, _06112_);
  or _61166_ (_10194_, _10193_, _10189_);
  and _61167_ (_10195_, _08760_, _07698_);
  or _61168_ (_10196_, _10195_, _09234_);
  or _61169_ (_10197_, _10196_, _08751_);
  and _61170_ (_10198_, _10197_, _08756_);
  and _61171_ (_10199_, _10198_, _10194_);
  or _61172_ (_10200_, _10199_, _09237_);
  and _61173_ (_10201_, _10200_, _07032_);
  or _61174_ (_10202_, _09234_, _07788_);
  and _61175_ (_10203_, _10191_, _06108_);
  and _61176_ (_10204_, _10203_, _10202_);
  or _61177_ (_10205_, _10204_, _10201_);
  and _61178_ (_10206_, _10205_, _06278_);
  and _61179_ (_10207_, _09246_, _06277_);
  and _61180_ (_10208_, _10207_, _10202_);
  or _61181_ (_10209_, _10208_, _06130_);
  or _61182_ (_10210_, _10209_, _10206_);
  and _61183_ (_10211_, _08759_, _07698_);
  or _61184_ (_10212_, _09234_, _08777_);
  or _61185_ (_10213_, _10212_, _10211_);
  and _61186_ (_10214_, _10213_, _08782_);
  and _61187_ (_10215_, _10214_, _10210_);
  nor _61188_ (_10216_, _08767_, _09258_);
  or _61189_ (_10217_, _10216_, _09234_);
  and _61190_ (_10218_, _10217_, _06292_);
  or _61191_ (_10219_, _10218_, _06316_);
  or _61192_ (_10220_, _10219_, _10215_);
  or _61193_ (_10221_, _09243_, _06718_);
  and _61194_ (_10222_, _10221_, _05653_);
  and _61195_ (_10223_, _10222_, _10220_);
  and _61196_ (_10224_, _09240_, _05652_);
  or _61197_ (_10225_, _10224_, _06047_);
  or _61198_ (_10226_, _10225_, _10223_);
  and _61199_ (_10227_, _08279_, _07698_);
  or _61200_ (_10228_, _09234_, _06048_);
  or _61201_ (_10229_, _10228_, _10227_);
  and _61202_ (_10230_, _10229_, _01336_);
  and _61203_ (_10231_, _10230_, _10226_);
  or _61204_ (_10232_, _10231_, _09233_);
  and _61205_ (_40752_, _10232_, _42882_);
  nor _61206_ (_10233_, _01336_, _08393_);
  and _61207_ (_10234_, _06931_, \oc8051_golden_model_1.PSW [7]);
  and _61208_ (_10235_, _10234_, _09161_);
  and _61209_ (_10236_, _10235_, _09160_);
  and _61210_ (_10237_, _10236_, _09159_);
  and _61211_ (_10238_, _10237_, _09158_);
  and _61212_ (_10239_, _10238_, _09157_);
  and _61213_ (_10240_, _10239_, _09156_);
  and _61214_ (_10241_, _10240_, _08288_);
  nor _61215_ (_10242_, _10240_, _08288_);
  or _61216_ (_10243_, _10242_, _10241_);
  and _61217_ (_10244_, _10243_, \oc8051_golden_model_1.ACC [7]);
  nor _61218_ (_10245_, _10243_, \oc8051_golden_model_1.ACC [7]);
  nor _61219_ (_10246_, _10245_, _10244_);
  nor _61220_ (_10247_, _10239_, _09156_);
  nor _61221_ (_10248_, _10247_, _10240_);
  and _61222_ (_10249_, _10248_, \oc8051_golden_model_1.ACC [6]);
  nor _61223_ (_10250_, _10248_, _09861_);
  and _61224_ (_10251_, _10248_, _09861_);
  nor _61225_ (_10252_, _10251_, _10250_);
  not _61226_ (_10253_, _10252_);
  nor _61227_ (_10254_, _10238_, _09157_);
  nor _61228_ (_10255_, _10254_, _10239_);
  and _61229_ (_10256_, _10255_, \oc8051_golden_model_1.ACC [5]);
  nor _61230_ (_10257_, _10255_, _09906_);
  and _61231_ (_10258_, _10255_, _09906_);
  nor _61232_ (_10259_, _10258_, _10257_);
  nor _61233_ (_10260_, _10237_, _09158_);
  nor _61234_ (_10261_, _10260_, _10238_);
  nand _61235_ (_10262_, _10261_, \oc8051_golden_model_1.ACC [4]);
  nor _61236_ (_10263_, _10261_, _09880_);
  and _61237_ (_10264_, _10261_, _09880_);
  or _61238_ (_10265_, _10264_, _10263_);
  nor _61239_ (_10266_, _10236_, _09159_);
  nor _61240_ (_10267_, _10266_, _10237_);
  and _61241_ (_10268_, _10267_, \oc8051_golden_model_1.ACC [3]);
  nor _61242_ (_10269_, _10267_, _10010_);
  and _61243_ (_10270_, _10267_, _10010_);
  nor _61244_ (_10271_, _10270_, _10269_);
  nor _61245_ (_10272_, _10235_, _09160_);
  nor _61246_ (_10273_, _10272_, _10236_);
  and _61247_ (_10274_, _10273_, \oc8051_golden_model_1.ACC [2]);
  nor _61248_ (_10275_, _10273_, _09956_);
  and _61249_ (_10276_, _10273_, _09956_);
  nor _61250_ (_10277_, _10276_, _10275_);
  nor _61251_ (_10278_, _10234_, _09161_);
  nor _61252_ (_10279_, _10278_, _10235_);
  and _61253_ (_10280_, _10279_, \oc8051_golden_model_1.ACC [1]);
  and _61254_ (_10281_, _10279_, _05784_);
  nor _61255_ (_10282_, _10279_, _05784_);
  nor _61256_ (_10283_, _10282_, _10281_);
  nor _61257_ (_10284_, _06931_, \oc8051_golden_model_1.PSW [7]);
  nor _61258_ (_10285_, _10284_, _10234_);
  and _61259_ (_10286_, _10285_, \oc8051_golden_model_1.ACC [0]);
  not _61260_ (_10287_, _10286_);
  nor _61261_ (_10288_, _10287_, _10283_);
  nor _61262_ (_10289_, _10288_, _10280_);
  nor _61263_ (_10290_, _10289_, _10277_);
  nor _61264_ (_10291_, _10290_, _10274_);
  nor _61265_ (_10292_, _10291_, _10271_);
  or _61266_ (_10293_, _10292_, _10268_);
  nand _61267_ (_10294_, _10293_, _10265_);
  and _61268_ (_10295_, _10294_, _10262_);
  nor _61269_ (_10296_, _10295_, _10259_);
  or _61270_ (_10297_, _10296_, _10256_);
  and _61271_ (_10298_, _10297_, _10253_);
  nor _61272_ (_10299_, _10298_, _10249_);
  nor _61273_ (_10300_, _10299_, _10246_);
  and _61274_ (_10301_, _10299_, _10246_);
  nor _61275_ (_10302_, _10301_, _10300_);
  and _61276_ (_10303_, _05731_, _05567_);
  not _61277_ (_10304_, _10303_);
  or _61278_ (_10305_, _10304_, _10302_);
  and _61279_ (_10306_, _06114_, _05671_);
  not _61280_ (_10307_, _10306_);
  and _61281_ (_10308_, _08127_, \oc8051_golden_model_1.PSW [7]);
  and _61282_ (_10309_, _10308_, _08078_);
  and _61283_ (_10310_, _10309_, _08177_);
  and _61284_ (_10311_, _10310_, _08029_);
  and _61285_ (_10312_, _10311_, _08273_);
  and _61286_ (_10313_, _10312_, _07980_);
  and _61287_ (_10314_, _10313_, _07886_);
  nor _61288_ (_10315_, _10314_, _07787_);
  and _61289_ (_10316_, _10314_, _07787_);
  nor _61290_ (_10317_, _10316_, _10315_);
  and _61291_ (_10318_, _10317_, \oc8051_golden_model_1.ACC [7]);
  nor _61292_ (_10319_, _10317_, \oc8051_golden_model_1.ACC [7]);
  nor _61293_ (_10320_, _10319_, _10318_);
  not _61294_ (_10321_, _10320_);
  nor _61295_ (_10322_, _10313_, _07886_);
  nor _61296_ (_10323_, _10322_, _10314_);
  nor _61297_ (_10324_, _10323_, _09861_);
  nor _61298_ (_10325_, _10312_, _07980_);
  nor _61299_ (_10326_, _10325_, _10313_);
  and _61300_ (_10327_, _10326_, _09906_);
  nor _61301_ (_10328_, _10326_, _09906_);
  nor _61302_ (_10329_, _10328_, _10327_);
  not _61303_ (_10330_, _10329_);
  nor _61304_ (_10331_, _10311_, _08273_);
  nor _61305_ (_10332_, _10331_, _10312_);
  nor _61306_ (_10333_, _10332_, _09880_);
  and _61307_ (_10334_, _10332_, _09880_);
  or _61308_ (_10335_, _10334_, _10333_);
  or _61309_ (_10336_, _10335_, _10330_);
  nor _61310_ (_10337_, _10310_, _08029_);
  nor _61311_ (_10338_, _10337_, _10311_);
  nor _61312_ (_10339_, _10338_, _10010_);
  and _61313_ (_10340_, _10338_, _10010_);
  nor _61314_ (_10341_, _10340_, _10339_);
  nor _61315_ (_10342_, _10309_, _08177_);
  nor _61316_ (_10343_, _10342_, _10310_);
  nor _61317_ (_10344_, _10343_, _09956_);
  and _61318_ (_10345_, _10343_, _09956_);
  nor _61319_ (_10346_, _10345_, _10344_);
  and _61320_ (_10347_, _10346_, _10341_);
  nor _61321_ (_10348_, _10308_, _08078_);
  nor _61322_ (_10349_, _10348_, _10309_);
  nor _61323_ (_10350_, _10349_, _05784_);
  and _61324_ (_10351_, _10349_, _05784_);
  nor _61325_ (_10352_, _08127_, \oc8051_golden_model_1.PSW [7]);
  nor _61326_ (_10353_, _10352_, _10308_);
  and _61327_ (_10354_, _10353_, _05758_);
  nor _61328_ (_10355_, _10354_, _10351_);
  or _61329_ (_10356_, _10355_, _10350_);
  nand _61330_ (_10357_, _10356_, _10347_);
  and _61331_ (_10358_, _10344_, _10341_);
  nor _61332_ (_10359_, _10358_, _10339_);
  and _61333_ (_10360_, _10359_, _10357_);
  nor _61334_ (_10361_, _10360_, _10336_);
  and _61335_ (_10362_, _10333_, _10329_);
  nor _61336_ (_10363_, _10362_, _10328_);
  not _61337_ (_10364_, _10363_);
  nor _61338_ (_10365_, _10364_, _10361_);
  and _61339_ (_10366_, _10323_, _09861_);
  nor _61340_ (_10367_, _10324_, _10366_);
  not _61341_ (_10368_, _10367_);
  nor _61342_ (_10369_, _10368_, _10365_);
  or _61343_ (_10370_, _10369_, _10324_);
  and _61344_ (_10371_, _10370_, _10321_);
  nor _61345_ (_10372_, _10370_, _10321_);
  or _61346_ (_10373_, _10372_, _10371_);
  or _61347_ (_10374_, _10373_, _06267_);
  and _61348_ (_10375_, _10374_, _10307_);
  and _61349_ (_10376_, _06114_, _06037_);
  nand _61350_ (_10377_, _10376_, _10010_);
  nor _61351_ (_10378_, _05693_, _08382_);
  nand _61352_ (_10379_, _10378_, _07785_);
  nor _61353_ (_10380_, _08359_, _08393_);
  and _61354_ (_10381_, _08503_, _08359_);
  or _61355_ (_10382_, _10381_, _10380_);
  or _61356_ (_10383_, _10382_, _06044_);
  and _61357_ (_10384_, _10383_, _06848_);
  nor _61358_ (_10385_, _07701_, _08393_);
  and _61359_ (_10386_, _08498_, _07701_);
  or _61360_ (_10387_, _10386_, _10385_);
  and _61361_ (_10388_, _10387_, _06102_);
  and _61362_ (_10389_, _06114_, _06523_);
  not _61363_ (_10390_, _10389_);
  or _61364_ (_10391_, _10390_, _08485_);
  nor _61365_ (_10392_, _06137_, _05697_);
  not _61366_ (_10393_, _10392_);
  nor _61367_ (_10394_, _05667_, _05661_);
  and _61368_ (_10395_, _10394_, _06523_);
  nor _61369_ (_10396_, _10395_, _06528_);
  and _61370_ (_10397_, _06133_, _06523_);
  nor _61371_ (_10398_, _10397_, _06525_);
  and _61372_ (_10399_, _10398_, _10396_);
  and _61373_ (_10400_, _10399_, _10393_);
  nor _61374_ (_10401_, _10400_, _07785_);
  or _61375_ (_10402_, _06530_, \oc8051_golden_model_1.ACC [7]);
  nand _61376_ (_10403_, _06530_, \oc8051_golden_model_1.ACC [7]);
  and _61377_ (_10404_, _10403_, _10402_);
  and _61378_ (_10405_, _10404_, _10400_);
  or _61379_ (_10406_, _10405_, _10389_);
  or _61380_ (_10407_, _10406_, _10401_);
  and _61381_ (_10408_, _06954_, _05698_);
  and _61382_ (_10409_, _10408_, _10407_);
  and _61383_ (_10410_, _10409_, _10391_);
  or _61384_ (_10411_, _10410_, _10388_);
  and _61385_ (_10412_, _06114_, _06042_);
  not _61386_ (_10413_, _10412_);
  and _61387_ (_10414_, _10413_, _10411_);
  nor _61388_ (_10415_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [2]);
  nor _61389_ (_10416_, _10415_, _10010_);
  and _61390_ (_10417_, _10416_, \oc8051_golden_model_1.ACC [4]);
  and _61391_ (_10418_, _10417_, \oc8051_golden_model_1.ACC [5]);
  and _61392_ (_10419_, _10418_, \oc8051_golden_model_1.ACC [6]);
  and _61393_ (_10420_, _10419_, \oc8051_golden_model_1.ACC [7]);
  nor _61394_ (_10421_, _10419_, \oc8051_golden_model_1.ACC [7]);
  nor _61395_ (_10422_, _10421_, _10420_);
  nor _61396_ (_10423_, _10417_, \oc8051_golden_model_1.ACC [5]);
  nor _61397_ (_10424_, _10423_, _10418_);
  nor _61398_ (_10425_, _10418_, \oc8051_golden_model_1.ACC [6]);
  nor _61399_ (_10426_, _10425_, _10419_);
  nor _61400_ (_10427_, _10426_, _10424_);
  not _61401_ (_10428_, _10427_);
  nand _61402_ (_10429_, _10428_, _10422_);
  nor _61403_ (_10430_, _10420_, \oc8051_golden_model_1.PSW [7]);
  and _61404_ (_10431_, _10430_, _10429_);
  nor _61405_ (_10432_, _10431_, _10427_);
  or _61406_ (_10433_, _10432_, _10422_);
  and _61407_ (_10434_, _10429_, _10412_);
  and _61408_ (_10435_, _10434_, _10433_);
  or _61409_ (_10436_, _10435_, _06043_);
  or _61410_ (_10437_, _10436_, _10414_);
  and _61411_ (_10438_, _10437_, _10384_);
  not _61412_ (_10439_, _07701_);
  nor _61413_ (_10440_, _07785_, _10439_);
  or _61414_ (_10441_, _10440_, _10385_);
  and _61415_ (_10442_, _10441_, _06239_);
  or _61416_ (_10443_, _10442_, _10378_);
  or _61417_ (_10444_, _10443_, _10438_);
  and _61418_ (_10445_, _10444_, _10379_);
  or _61419_ (_10446_, _10445_, _06970_);
  or _61420_ (_10447_, _08485_, _06971_);
  and _61421_ (_10448_, _10447_, _06220_);
  and _61422_ (_10449_, _10448_, _10446_);
  nor _61423_ (_10450_, _07787_, _06220_);
  or _61424_ (_10451_, _10450_, _10376_);
  or _61425_ (_10452_, _10451_, _10449_);
  and _61426_ (_10453_, _10452_, _10377_);
  or _61427_ (_10454_, _10453_, _06039_);
  and _61428_ (_10455_, _08374_, _08359_);
  or _61429_ (_10456_, _10455_, _10380_);
  or _61430_ (_10457_, _10456_, _06040_);
  and _61431_ (_10458_, _10457_, _06033_);
  and _61432_ (_10459_, _10458_, _10454_);
  or _61433_ (_10460_, _10380_, _08519_);
  and _61434_ (_10461_, _10382_, _06032_);
  and _61435_ (_10462_, _10461_, _10460_);
  or _61436_ (_10463_, _10462_, _09269_);
  or _61437_ (_10464_, _10463_, _10459_);
  nor _61438_ (_10465_, _09762_, _09760_);
  nor _61439_ (_10466_, _10465_, _09763_);
  or _61440_ (_10467_, _10466_, _09800_);
  and _61441_ (_10468_, _05671_, _05567_);
  not _61442_ (_10469_, _10468_);
  and _61443_ (_10470_, _10469_, _10467_);
  and _61444_ (_10471_, _10470_, _10464_);
  nor _61445_ (_10472_, _10263_, _10257_);
  nor _61446_ (_10473_, _10472_, _10258_);
  not _61447_ (_10474_, _10259_);
  or _61448_ (_10475_, _10265_, _10474_);
  and _61449_ (_10476_, _10277_, _10271_);
  and _61450_ (_10477_, _10285_, _05758_);
  nor _61451_ (_10478_, _10477_, _10281_);
  or _61452_ (_10479_, _10478_, _10282_);
  nand _61453_ (_10480_, _10479_, _10476_);
  and _61454_ (_10481_, _10275_, _10271_);
  nor _61455_ (_10482_, _10481_, _10269_);
  and _61456_ (_10483_, _10482_, _10480_);
  nor _61457_ (_10484_, _10483_, _10475_);
  nor _61458_ (_10485_, _10484_, _10473_);
  nor _61459_ (_10486_, _10485_, _10253_);
  or _61460_ (_10487_, _10486_, _10250_);
  nor _61461_ (_10488_, _10487_, _10246_);
  and _61462_ (_10489_, _10487_, _10246_);
  or _61463_ (_10490_, _10489_, _10488_);
  nor _61464_ (_10491_, _10490_, _10469_);
  nor _61465_ (_10492_, _10491_, _10471_);
  and _61466_ (_10493_, _10394_, _05671_);
  nor _61467_ (_10494_, _10493_, _10492_);
  and _61468_ (_10495_, _09188_, \oc8051_golden_model_1.PSW [7]);
  nor _61469_ (_10496_, _10495_, _08798_);
  and _61470_ (_10497_, _10495_, _08798_);
  nor _61471_ (_10498_, _10497_, _10496_);
  and _61472_ (_10499_, _10498_, \oc8051_golden_model_1.ACC [7]);
  nor _61473_ (_10500_, _10498_, \oc8051_golden_model_1.ACC [7]);
  nor _61474_ (_10501_, _10500_, _10499_);
  not _61475_ (_10502_, _10501_);
  and _61476_ (_10503_, _09187_, \oc8051_golden_model_1.PSW [7]);
  nor _61477_ (_10504_, _10503_, _09178_);
  nor _61478_ (_10505_, _10504_, _10495_);
  nor _61479_ (_10506_, _10505_, _09861_);
  and _61480_ (_10507_, _09186_, \oc8051_golden_model_1.PSW [7]);
  nor _61481_ (_10508_, _10507_, _09179_);
  nor _61482_ (_10509_, _10508_, _10503_);
  and _61483_ (_10510_, _10509_, _09906_);
  nor _61484_ (_10511_, _10509_, _09906_);
  and _61485_ (_10512_, _09185_, \oc8051_golden_model_1.PSW [7]);
  nor _61486_ (_10513_, _10512_, _09180_);
  nor _61487_ (_10514_, _10513_, _10507_);
  nor _61488_ (_10515_, _10514_, _09880_);
  nor _61489_ (_10516_, _10515_, _10511_);
  nor _61490_ (_10517_, _10516_, _10510_);
  nor _61491_ (_10518_, _10511_, _10510_);
  not _61492_ (_10519_, _10518_);
  and _61493_ (_10520_, _10514_, _09880_);
  or _61494_ (_10521_, _10520_, _10515_);
  or _61495_ (_10522_, _10521_, _10519_);
  and _61496_ (_10523_, _09184_, \oc8051_golden_model_1.PSW [7]);
  nor _61497_ (_10524_, _10523_, _09181_);
  nor _61498_ (_10525_, _10524_, _10512_);
  nor _61499_ (_10526_, _10525_, _10010_);
  and _61500_ (_10527_, _10525_, _10010_);
  nor _61501_ (_10528_, _10527_, _10526_);
  and _61502_ (_10529_, _09183_, \oc8051_golden_model_1.PSW [7]);
  nor _61503_ (_10530_, _10529_, _09182_);
  nor _61504_ (_10531_, _10530_, _10523_);
  nor _61505_ (_10532_, _10531_, _09956_);
  and _61506_ (_10533_, _10531_, _09956_);
  nor _61507_ (_10534_, _10533_, _10532_);
  and _61508_ (_10535_, _10534_, _10528_);
  and _61509_ (_10536_, _09120_, \oc8051_golden_model_1.PSW [7]);
  nor _61510_ (_10537_, _10536_, _09075_);
  nor _61511_ (_10538_, _10537_, _10529_);
  nor _61512_ (_10539_, _10538_, _05784_);
  and _61513_ (_10540_, _10538_, _05784_);
  nor _61514_ (_10541_, _09120_, \oc8051_golden_model_1.PSW [7]);
  nor _61515_ (_10542_, _10541_, _10536_);
  and _61516_ (_10543_, _10542_, _05758_);
  nor _61517_ (_10544_, _10543_, _10540_);
  or _61518_ (_10545_, _10544_, _10539_);
  nand _61519_ (_10546_, _10545_, _10535_);
  and _61520_ (_10547_, _10532_, _10528_);
  nor _61521_ (_10548_, _10547_, _10526_);
  and _61522_ (_10549_, _10548_, _10546_);
  nor _61523_ (_10550_, _10549_, _10522_);
  nor _61524_ (_10551_, _10550_, _10517_);
  and _61525_ (_10552_, _10505_, _09861_);
  nor _61526_ (_10553_, _10506_, _10552_);
  not _61527_ (_10554_, _10553_);
  nor _61528_ (_10555_, _10554_, _10551_);
  or _61529_ (_10556_, _10555_, _10506_);
  and _61530_ (_10557_, _10556_, _10502_);
  nor _61531_ (_10558_, _10556_, _10502_);
  or _61532_ (_10559_, _10558_, _10557_);
  and _61533_ (_10560_, _10559_, _10493_);
  nor _61534_ (_10561_, _10560_, _10494_);
  nor _61535_ (_10562_, _10561_, _06591_);
  and _61536_ (_10563_, _10559_, _06591_);
  or _61537_ (_10564_, _10563_, _10562_);
  or _61538_ (_10565_, _10564_, _06261_);
  and _61539_ (_10566_, _10565_, _10375_);
  and _61540_ (_10567_, _08375_, _06299_);
  and _61541_ (_10568_, _10567_, _07697_);
  and _61542_ (_10569_, _10567_, _07690_);
  and _61543_ (_10570_, _10569_, _07414_);
  nor _61544_ (_10571_, _10570_, _05952_);
  nor _61545_ (_10572_, _10571_, _10568_);
  nor _61546_ (_10573_, _10572_, _08393_);
  and _61547_ (_10574_, _10572_, _08393_);
  nor _61548_ (_10575_, _10574_, _10573_);
  nor _61549_ (_10576_, _10569_, _07414_);
  nor _61550_ (_10577_, _10576_, _10570_);
  nor _61551_ (_10578_, _10577_, _09861_);
  and _61552_ (_10579_, _10567_, _07674_);
  nor _61553_ (_10580_, _10579_, _07683_);
  nor _61554_ (_10581_, _10580_, _10569_);
  and _61555_ (_10582_, _10581_, _09906_);
  nor _61556_ (_10583_, _10581_, _09906_);
  nor _61557_ (_10584_, _10567_, _07674_);
  nor _61558_ (_10585_, _10584_, _10579_);
  nor _61559_ (_10586_, _10585_, _09880_);
  nor _61560_ (_10587_, _10586_, _10583_);
  nor _61561_ (_10588_, _10587_, _10582_);
  nor _61562_ (_10589_, _10583_, _10582_);
  not _61563_ (_10590_, _10589_);
  and _61564_ (_10591_, _10585_, _09880_);
  or _61565_ (_10592_, _10591_, _10586_);
  or _61566_ (_10593_, _10592_, _10590_);
  nor _61567_ (_10594_, _08375_, _06299_);
  nor _61568_ (_10595_, _10594_, _10567_);
  nor _61569_ (_10596_, _10595_, _10010_);
  and _61570_ (_10597_, _10595_, _10010_);
  nor _61571_ (_10598_, _10597_, _10596_);
  and _61572_ (_10599_, _07639_, \oc8051_golden_model_1.PSW [7]);
  nor _61573_ (_10600_, _10599_, _07477_);
  or _61574_ (_10601_, _10600_, _08375_);
  and _61575_ (_10602_, _10601_, \oc8051_golden_model_1.ACC [2]);
  nor _61576_ (_10603_, _10601_, \oc8051_golden_model_1.ACC [2]);
  nor _61577_ (_10604_, _10603_, _10602_);
  and _61578_ (_10605_, _10604_, _10598_);
  not _61579_ (_10606_, \oc8051_golden_model_1.PSW [7]);
  nor _61580_ (_10607_, _06016_, _10606_);
  nor _61581_ (_10608_, _10607_, _07076_);
  nor _61582_ (_10609_, _10608_, _10599_);
  nor _61583_ (_10610_, _10609_, _05784_);
  and _61584_ (_10611_, _10609_, _05784_);
  nor _61585_ (_10612_, _06016_, \oc8051_golden_model_1.PSW [7]);
  and _61586_ (_10613_, _06016_, \oc8051_golden_model_1.PSW [7]);
  nor _61587_ (_10614_, _10613_, _10612_);
  nor _61588_ (_10615_, _10614_, \oc8051_golden_model_1.ACC [0]);
  nor _61589_ (_10616_, _10615_, _10611_);
  or _61590_ (_10617_, _10616_, _10610_);
  nand _61591_ (_10618_, _10617_, _10605_);
  and _61592_ (_10619_, _10602_, _10598_);
  nor _61593_ (_10620_, _10619_, _10596_);
  and _61594_ (_10621_, _10620_, _10618_);
  nor _61595_ (_10622_, _10621_, _10593_);
  nor _61596_ (_10623_, _10622_, _10588_);
  and _61597_ (_10624_, _10577_, _09861_);
  nor _61598_ (_10625_, _10578_, _10624_);
  not _61599_ (_10626_, _10625_);
  nor _61600_ (_10627_, _10626_, _10623_);
  or _61601_ (_10628_, _10627_, _10578_);
  nor _61602_ (_10629_, _10628_, _10575_);
  and _61603_ (_10630_, _10628_, _10575_);
  or _61604_ (_10631_, _10630_, _10629_);
  nor _61605_ (_10632_, _10631_, _10307_);
  or _61606_ (_10633_, _10632_, _05676_);
  or _61607_ (_10634_, _10633_, _10566_);
  or _61608_ (_10635_, _05952_, _05675_);
  and _61609_ (_10636_, _10635_, _06027_);
  and _61610_ (_10637_, _10636_, _10634_);
  and _61611_ (_10638_, _08376_, _08359_);
  or _61612_ (_10639_, _10638_, _10380_);
  and _61613_ (_10640_, _10639_, _06026_);
  or _61614_ (_10641_, _10640_, _09818_);
  or _61615_ (_10642_, _10641_, _10637_);
  and _61616_ (_10643_, _08485_, _07701_);
  or _61617_ (_10644_, _10385_, _07012_);
  or _61618_ (_10645_, _10644_, _10643_);
  or _61619_ (_10646_, _10441_, _09827_);
  and _61620_ (_10647_, _10646_, _05669_);
  and _61621_ (_10648_, _10647_, _10645_);
  and _61622_ (_10649_, _10648_, _10642_);
  and _61623_ (_10650_, _08738_, _07701_);
  or _61624_ (_10651_, _10650_, _10385_);
  and _61625_ (_10652_, _10651_, _09833_);
  or _61626_ (_10653_, _10652_, _09832_);
  or _61627_ (_10654_, _10653_, _10649_);
  or _61628_ (_10655_, _09851_, _09839_);
  and _61629_ (_10656_, _10655_, _05664_);
  and _61630_ (_10657_, _10656_, _10654_);
  and _61631_ (_10658_, _05952_, _05663_);
  or _61632_ (_10659_, _10658_, _06019_);
  or _61633_ (_10660_, _10659_, _10657_);
  and _61634_ (_10661_, _06114_, _05723_);
  not _61635_ (_10662_, _10661_);
  and _61636_ (_10663_, _08549_, _07701_);
  or _61637_ (_10664_, _10663_, _10385_);
  or _61638_ (_10665_, _10664_, _06020_);
  and _61639_ (_10666_, _10665_, _10662_);
  and _61640_ (_10667_, _10666_, _10660_);
  and _61641_ (_10668_, _10661_, _05952_);
  and _61642_ (_10669_, _07005_, _05726_);
  or _61643_ (_10670_, _10669_, _10668_);
  or _61644_ (_10671_, _10670_, _10667_);
  and _61645_ (_10672_, _07785_, _08393_);
  nor _61646_ (_10673_, _07785_, _08393_);
  nor _61647_ (_10674_, _10673_, _10672_);
  not _61648_ (_10675_, _10669_);
  or _61649_ (_10676_, _10675_, _10674_);
  nor _61650_ (_10677_, _06137_, _06644_);
  not _61651_ (_10678_, _10677_);
  and _61652_ (_10679_, _10678_, _10676_);
  and _61653_ (_10680_, _10679_, _10671_);
  and _61654_ (_10681_, _07002_, _05726_);
  and _61655_ (_10682_, _10677_, _10674_);
  or _61656_ (_10683_, _10682_, _10681_);
  or _61657_ (_10684_, _10683_, _10680_);
  and _61658_ (_10685_, _06103_, _05726_);
  not _61659_ (_10686_, _10685_);
  not _61660_ (_10687_, _10681_);
  or _61661_ (_10688_, _10687_, _10674_);
  and _61662_ (_10689_, _10688_, _10686_);
  and _61663_ (_10690_, _10689_, _10684_);
  and _61664_ (_10691_, _08798_, _08393_);
  and _61665_ (_10692_, _08485_, \oc8051_golden_model_1.ACC [7]);
  nor _61666_ (_10693_, _10692_, _10691_);
  and _61667_ (_10694_, _10685_, _10693_);
  or _61668_ (_10695_, _10694_, _06282_);
  or _61669_ (_10697_, _10695_, _10690_);
  and _61670_ (_10698_, _06114_, _05726_);
  not _61671_ (_10699_, _10698_);
  or _61672_ (_10700_, _08768_, _06283_);
  and _61673_ (_10701_, _10700_, _10699_);
  and _61674_ (_10702_, _10701_, _10697_);
  nor _61675_ (_10703_, _05952_, \oc8051_golden_model_1.ACC [7]);
  and _61676_ (_10704_, _05952_, \oc8051_golden_model_1.ACC [7]);
  nor _61677_ (_10705_, _10704_, _10703_);
  and _61678_ (_10706_, _10698_, _10705_);
  or _61679_ (_10708_, _10706_, _06112_);
  or _61680_ (_10709_, _10708_, _10702_);
  and _61681_ (_10710_, _08760_, _07701_);
  or _61682_ (_10711_, _10710_, _10385_);
  or _61683_ (_10712_, _10711_, _08751_);
  and _61684_ (_10713_, _10712_, _08756_);
  and _61685_ (_10714_, _10713_, _10709_);
  and _61686_ (_10715_, _10385_, _06284_);
  or _61687_ (_10716_, _10715_, _06482_);
  or _61688_ (_10717_, _10716_, _10714_);
  not _61689_ (_10719_, _10673_);
  nand _61690_ (_10720_, _10719_, _06482_);
  and _61691_ (_10721_, _06096_, _05735_);
  not _61692_ (_10722_, _10721_);
  not _61693_ (_10723_, _06490_);
  and _61694_ (_10724_, _06133_, _05735_);
  nor _61695_ (_10725_, _10724_, _06835_);
  and _61696_ (_10726_, _10725_, _10723_);
  and _61697_ (_10727_, _10726_, _10722_);
  and _61698_ (_10728_, _10727_, _10720_);
  and _61699_ (_10730_, _10728_, _10717_);
  and _61700_ (_10731_, _06103_, _05735_);
  nor _61701_ (_10732_, _10727_, _10719_);
  or _61702_ (_10733_, _10732_, _10731_);
  or _61703_ (_10734_, _10733_, _10730_);
  not _61704_ (_10735_, _06279_);
  not _61705_ (_10736_, _10731_);
  or _61706_ (_10737_, _10736_, _10692_);
  and _61707_ (_10738_, _10737_, _10735_);
  and _61708_ (_10739_, _10738_, _10734_);
  and _61709_ (_10741_, _06114_, _05735_);
  nor _61710_ (_10742_, _10741_, _06279_);
  not _61711_ (_10743_, _10742_);
  or _61712_ (_10744_, _10741_, _08766_);
  and _61713_ (_10745_, _10744_, _10743_);
  or _61714_ (_10746_, _10745_, _10739_);
  not _61715_ (_10747_, _10741_);
  or _61716_ (_10748_, _10747_, _10704_);
  and _61717_ (_10749_, _10748_, _07032_);
  and _61718_ (_10750_, _10749_, _10746_);
  and _61719_ (_10752_, _06450_, _05739_);
  nand _61720_ (_10753_, _10664_, _06108_);
  nor _61721_ (_10754_, _10753_, _08767_);
  or _61722_ (_10755_, _10754_, _10752_);
  or _61723_ (_10756_, _10755_, _10750_);
  not _61724_ (_10757_, _05739_);
  nor _61725_ (_10758_, _06460_, _06229_);
  nor _61726_ (_10759_, _10758_, _10757_);
  not _61727_ (_10760_, _10759_);
  nand _61728_ (_10761_, _10672_, _10752_);
  and _61729_ (_10763_, _10761_, _10760_);
  and _61730_ (_10764_, _10763_, _10756_);
  and _61731_ (_10765_, _06133_, _05739_);
  nor _61732_ (_10766_, _10765_, _06665_);
  not _61733_ (_10767_, _10766_);
  nor _61734_ (_10768_, _10760_, _10672_);
  or _61735_ (_10769_, _10768_, _10767_);
  or _61736_ (_10770_, _10769_, _10764_);
  nand _61737_ (_10771_, _10767_, _10672_);
  and _61738_ (_10772_, _10771_, _06668_);
  and _61739_ (_10773_, _10772_, _10770_);
  nor _61740_ (_10774_, _10672_, _06668_);
  and _61741_ (_10775_, _06103_, _05739_);
  or _61742_ (_10776_, _10775_, _10774_);
  or _61743_ (_10777_, _10776_, _10773_);
  nand _61744_ (_10778_, _10775_, _10691_);
  and _61745_ (_10779_, _10778_, _06291_);
  and _61746_ (_10780_, _10779_, _10777_);
  and _61747_ (_10781_, _06114_, _05739_);
  nor _61748_ (_10782_, _08767_, _06291_);
  or _61749_ (_10783_, _10782_, _10781_);
  or _61750_ (_10784_, _10783_, _10780_);
  nand _61751_ (_10785_, _10781_, _10703_);
  and _61752_ (_10786_, _10785_, _08777_);
  and _61753_ (_10787_, _10786_, _10784_);
  and _61754_ (_10788_, _08759_, _07701_);
  or _61755_ (_10789_, _10788_, _10385_);
  and _61756_ (_10790_, _10789_, _06130_);
  or _61757_ (_10791_, _10790_, _10303_);
  or _61758_ (_10792_, _10791_, _10787_);
  and _61759_ (_10793_, _10792_, _10305_);
  and _61760_ (_10794_, _06103_, _05731_);
  or _61761_ (_10795_, _10794_, _10793_);
  not _61762_ (_10796_, _10794_);
  nand _61763_ (_10797_, _10505_, \oc8051_golden_model_1.ACC [6]);
  and _61764_ (_10798_, _10509_, \oc8051_golden_model_1.ACC [5]);
  nand _61765_ (_10799_, _10514_, \oc8051_golden_model_1.ACC [4]);
  and _61766_ (_10800_, _10525_, \oc8051_golden_model_1.ACC [3]);
  and _61767_ (_10801_, _10531_, \oc8051_golden_model_1.ACC [2]);
  and _61768_ (_10802_, _10538_, \oc8051_golden_model_1.ACC [1]);
  nor _61769_ (_10803_, _10540_, _10539_);
  and _61770_ (_10804_, _10542_, \oc8051_golden_model_1.ACC [0]);
  not _61771_ (_10805_, _10804_);
  nor _61772_ (_10806_, _10805_, _10803_);
  nor _61773_ (_10807_, _10806_, _10802_);
  nor _61774_ (_10808_, _10807_, _10534_);
  nor _61775_ (_10809_, _10808_, _10801_);
  nor _61776_ (_10810_, _10809_, _10528_);
  or _61777_ (_10811_, _10810_, _10800_);
  nand _61778_ (_10812_, _10811_, _10521_);
  and _61779_ (_10813_, _10812_, _10799_);
  nor _61780_ (_10814_, _10813_, _10518_);
  or _61781_ (_10815_, _10814_, _10798_);
  nand _61782_ (_10816_, _10815_, _10554_);
  and _61783_ (_10817_, _10816_, _10797_);
  nor _61784_ (_10818_, _10817_, _10501_);
  and _61785_ (_10819_, _10817_, _10501_);
  nor _61786_ (_10820_, _10819_, _10818_);
  or _61787_ (_10821_, _10820_, _10796_);
  and _61788_ (_10822_, _10821_, _06289_);
  and _61789_ (_10823_, _10822_, _10795_);
  and _61790_ (_10824_, _06114_, _05731_);
  nor _61791_ (_10825_, _10824_, _06288_);
  not _61792_ (_10826_, _10825_);
  and _61793_ (_10827_, _10323_, \oc8051_golden_model_1.ACC [6]);
  and _61794_ (_10828_, _10326_, \oc8051_golden_model_1.ACC [5]);
  nand _61795_ (_10829_, _10332_, \oc8051_golden_model_1.ACC [4]);
  and _61796_ (_10830_, _10338_, \oc8051_golden_model_1.ACC [3]);
  and _61797_ (_10831_, _10343_, \oc8051_golden_model_1.ACC [2]);
  and _61798_ (_10832_, _10349_, \oc8051_golden_model_1.ACC [1]);
  nor _61799_ (_10833_, _10351_, _10350_);
  not _61800_ (_10834_, _10833_);
  and _61801_ (_10835_, _10353_, \oc8051_golden_model_1.ACC [0]);
  and _61802_ (_10836_, _10835_, _10834_);
  nor _61803_ (_10837_, _10836_, _10832_);
  nor _61804_ (_10838_, _10837_, _10346_);
  nor _61805_ (_10839_, _10838_, _10831_);
  nor _61806_ (_10840_, _10839_, _10341_);
  or _61807_ (_10841_, _10840_, _10830_);
  nand _61808_ (_10842_, _10841_, _10335_);
  and _61809_ (_10843_, _10842_, _10829_);
  nor _61810_ (_10844_, _10843_, _10329_);
  or _61811_ (_10845_, _10844_, _10828_);
  and _61812_ (_10846_, _10845_, _10368_);
  nor _61813_ (_10847_, _10846_, _10827_);
  nor _61814_ (_10848_, _10847_, _10320_);
  and _61815_ (_10849_, _10847_, _10320_);
  nor _61816_ (_10850_, _10849_, _10848_);
  or _61817_ (_10851_, _10850_, _10824_);
  and _61818_ (_10852_, _10851_, _10826_);
  or _61819_ (_10853_, _10852_, _10823_);
  and _61820_ (_10854_, _05731_, _06107_);
  not _61821_ (_10855_, _10854_);
  not _61822_ (_10856_, _10824_);
  nand _61823_ (_10857_, _10577_, \oc8051_golden_model_1.ACC [6]);
  and _61824_ (_10858_, _10581_, \oc8051_golden_model_1.ACC [5]);
  nand _61825_ (_10859_, _10585_, \oc8051_golden_model_1.ACC [4]);
  and _61826_ (_10860_, _10595_, \oc8051_golden_model_1.ACC [3]);
  nor _61827_ (_10861_, _10601_, _09956_);
  and _61828_ (_10862_, _10609_, \oc8051_golden_model_1.ACC [1]);
  nor _61829_ (_10863_, _10611_, _10610_);
  not _61830_ (_10864_, _10863_);
  nor _61831_ (_10865_, _10614_, _05758_);
  and _61832_ (_10866_, _10865_, _10864_);
  nor _61833_ (_10867_, _10866_, _10862_);
  nor _61834_ (_10868_, _10867_, _10604_);
  nor _61835_ (_10869_, _10868_, _10861_);
  nor _61836_ (_10870_, _10869_, _10598_);
  or _61837_ (_10871_, _10870_, _10860_);
  nand _61838_ (_10872_, _10871_, _10592_);
  and _61839_ (_10873_, _10872_, _10859_);
  nor _61840_ (_10874_, _10873_, _10589_);
  or _61841_ (_10875_, _10874_, _10858_);
  nand _61842_ (_10876_, _10875_, _10626_);
  and _61843_ (_10877_, _10876_, _10857_);
  nor _61844_ (_10878_, _10877_, _10575_);
  and _61845_ (_10879_, _10877_, _10575_);
  nor _61846_ (_10880_, _10879_, _10878_);
  or _61847_ (_10881_, _10880_, _10856_);
  and _61848_ (_10882_, _10881_, _10855_);
  and _61849_ (_10883_, _10882_, _10853_);
  nand _61850_ (_10884_, _10854_, \oc8051_golden_model_1.ACC [6]);
  and _61851_ (_10885_, _07002_, _05746_);
  not _61852_ (_10886_, _10885_);
  and _61853_ (_10887_, _07005_, _05746_);
  nor _61854_ (_10888_, _06137_, _06841_);
  nor _61855_ (_10889_, _10888_, _10887_);
  and _61856_ (_10890_, _10889_, _10886_);
  nand _61857_ (_10891_, _10890_, _10884_);
  or _61858_ (_10892_, _10891_, _10883_);
  nor _61859_ (_10893_, _07883_, _09861_);
  not _61860_ (_10894_, _10893_);
  nand _61861_ (_10895_, _07883_, _09861_);
  and _61862_ (_10896_, _10894_, _10895_);
  nor _61863_ (_10897_, _07977_, _09906_);
  and _61864_ (_10898_, _07977_, _09906_);
  nor _61865_ (_10899_, _10898_, _10897_);
  not _61866_ (_10900_, _10899_);
  nor _61867_ (_10901_, _08270_, _09880_);
  nand _61868_ (_10902_, _08270_, _09880_);
  not _61869_ (_10903_, _10901_);
  and _61870_ (_10904_, _10903_, _10902_);
  nor _61871_ (_10905_, _07353_, _10010_);
  and _61872_ (_10906_, _07353_, _10010_);
  nor _61873_ (_10907_, _07530_, _09956_);
  and _61874_ (_10908_, _07530_, _09956_);
  nor _61875_ (_10909_, _10907_, _10908_);
  nor _61876_ (_10910_, _07132_, _05784_);
  and _61877_ (_10911_, _07132_, _05784_);
  nor _61878_ (_10912_, _10910_, _10911_);
  and _61879_ (_10913_, _06931_, \oc8051_golden_model_1.ACC [0]);
  and _61880_ (_10914_, _10913_, _10912_);
  nor _61881_ (_10915_, _10914_, _10910_);
  not _61882_ (_10916_, _10915_);
  and _61883_ (_10917_, _10916_, _10909_);
  nor _61884_ (_10918_, _10917_, _10907_);
  nor _61885_ (_10919_, _10918_, _10906_);
  or _61886_ (_10920_, _10919_, _10905_);
  and _61887_ (_10921_, _10920_, _10904_);
  nor _61888_ (_10922_, _10921_, _10901_);
  nor _61889_ (_10923_, _10922_, _10900_);
  or _61890_ (_10924_, _10923_, _10897_);
  nand _61891_ (_10925_, _10924_, _10896_);
  and _61892_ (_10926_, _10925_, _10894_);
  nor _61893_ (_10927_, _10926_, _10674_);
  and _61894_ (_10928_, _10926_, _10674_);
  or _61895_ (_10929_, _10928_, _10927_);
  or _61896_ (_10930_, _10929_, _10890_);
  and _61897_ (_10931_, _10930_, _10892_);
  and _61898_ (_10932_, _06103_, _05746_);
  or _61899_ (_10933_, _10932_, _10931_);
  not _61900_ (_10934_, _10932_);
  and _61901_ (_10935_, _09178_, \oc8051_golden_model_1.ACC [6]);
  or _61902_ (_10936_, _09178_, \oc8051_golden_model_1.ACC [6]);
  not _61903_ (_10937_, _10935_);
  and _61904_ (_10938_, _10937_, _10936_);
  and _61905_ (_10939_, _09179_, \oc8051_golden_model_1.ACC [5]);
  and _61906_ (_10940_, _08888_, _09906_);
  or _61907_ (_10941_, _10940_, _10939_);
  or _61908_ (_10942_, _08937_, _09880_);
  or _61909_ (_10943_, _09180_, \oc8051_golden_model_1.ACC [4]);
  and _61910_ (_10944_, _10942_, _10943_);
  and _61911_ (_10945_, _09181_, \oc8051_golden_model_1.ACC [3]);
  and _61912_ (_10946_, _08985_, _10010_);
  and _61913_ (_10947_, _09182_, \oc8051_golden_model_1.ACC [2]);
  and _61914_ (_10948_, _09030_, _09956_);
  nor _61915_ (_10949_, _10947_, _10948_);
  not _61916_ (_10950_, _10949_);
  and _61917_ (_10951_, _09075_, \oc8051_golden_model_1.ACC [1]);
  or _61918_ (_10952_, _09075_, \oc8051_golden_model_1.ACC [1]);
  not _61919_ (_10953_, _10951_);
  and _61920_ (_10954_, _10953_, _10952_);
  and _61921_ (_10955_, _09120_, \oc8051_golden_model_1.ACC [0]);
  and _61922_ (_10956_, _10955_, _10954_);
  nor _61923_ (_10957_, _10956_, _10951_);
  nor _61924_ (_10958_, _10957_, _10950_);
  nor _61925_ (_10959_, _10958_, _10947_);
  nor _61926_ (_10960_, _10959_, _10946_);
  or _61927_ (_10961_, _10960_, _10945_);
  nand _61928_ (_10962_, _10961_, _10944_);
  and _61929_ (_10963_, _10962_, _10942_);
  nor _61930_ (_10964_, _10963_, _10941_);
  or _61931_ (_10965_, _10964_, _10939_);
  and _61932_ (_10966_, _10965_, _10938_);
  nor _61933_ (_10967_, _10966_, _10935_);
  and _61934_ (_10968_, _10967_, _10693_);
  nor _61935_ (_10969_, _10967_, _10693_);
  or _61936_ (_10970_, _10969_, _10968_);
  or _61937_ (_10971_, _10970_, _10934_);
  and _61938_ (_10972_, _10971_, _06052_);
  and _61939_ (_10973_, _10972_, _10933_);
  and _61940_ (_10974_, _06114_, _05746_);
  nor _61941_ (_10975_, _10974_, _06051_);
  not _61942_ (_10976_, _10975_);
  nor _61943_ (_10977_, _07885_, _09861_);
  not _61944_ (_10978_, _10977_);
  and _61945_ (_10979_, _07885_, _09861_);
  nor _61946_ (_10980_, _10979_, _10977_);
  nor _61947_ (_10981_, _07979_, _09906_);
  and _61948_ (_10982_, _07979_, _09906_);
  nor _61949_ (_10983_, _08272_, _09880_);
  not _61950_ (_10984_, _10983_);
  and _61951_ (_10985_, _08272_, _09880_);
  nor _61952_ (_10986_, _10985_, _10983_);
  nor _61953_ (_10987_, _08028_, _10010_);
  and _61954_ (_10988_, _08028_, _10010_);
  nor _61955_ (_10989_, _08176_, _09956_);
  and _61956_ (_10990_, _08176_, _09956_);
  nor _61957_ (_10991_, _10990_, _10989_);
  nor _61958_ (_10992_, _08077_, _05784_);
  and _61959_ (_10993_, _08077_, _05784_);
  nor _61960_ (_10994_, _10993_, _10992_);
  and _61961_ (_10995_, _08127_, \oc8051_golden_model_1.ACC [0]);
  and _61962_ (_10996_, _10995_, _10994_);
  nor _61963_ (_10997_, _10996_, _10992_);
  not _61964_ (_10998_, _10997_);
  and _61965_ (_10999_, _10998_, _10991_);
  nor _61966_ (_11000_, _10999_, _10989_);
  nor _61967_ (_11001_, _11000_, _10988_);
  or _61968_ (_11002_, _11001_, _10987_);
  nand _61969_ (_11003_, _11002_, _10986_);
  and _61970_ (_11004_, _11003_, _10984_);
  nor _61971_ (_11005_, _11004_, _10982_);
  or _61972_ (_11006_, _11005_, _10981_);
  nand _61973_ (_11007_, _11006_, _10980_);
  and _61974_ (_11008_, _11007_, _10978_);
  and _61975_ (_11009_, _11008_, _08768_);
  nor _61976_ (_11010_, _11008_, _08768_);
  or _61977_ (_11011_, _11010_, _10974_);
  or _61978_ (_11012_, _11011_, _11009_);
  and _61979_ (_11013_, _11012_, _10976_);
  or _61980_ (_11014_, _11013_, _10973_);
  and _61981_ (_11015_, _05746_, _06107_);
  not _61982_ (_11016_, _11015_);
  nor _61983_ (_11017_, _06084_, _09861_);
  not _61984_ (_11018_, _11017_);
  and _61985_ (_11019_, _06084_, _09861_);
  nor _61986_ (_11020_, _11017_, _11019_);
  nor _61987_ (_11021_, _06359_, _09906_);
  and _61988_ (_11022_, _06359_, _09906_);
  nor _61989_ (_11023_, _06758_, _09880_);
  not _61990_ (_11024_, _11023_);
  and _61991_ (_11025_, _06758_, _09880_);
  or _61992_ (_11026_, _11025_, _11023_);
  not _61993_ (_11027_, _11026_);
  nor _61994_ (_11028_, _05983_, _10010_);
  and _61995_ (_11029_, _05983_, _10010_);
  nor _61996_ (_11030_, _06403_, _09956_);
  and _61997_ (_11031_, _06403_, _09956_);
  or _61998_ (_11032_, _11031_, _11030_);
  nor _61999_ (_11033_, _06799_, _05784_);
  and _62000_ (_11034_, _06799_, _05784_);
  nor _62001_ (_11035_, _11033_, _11034_);
  nor _62002_ (_11036_, _06016_, _05758_);
  and _62003_ (_11037_, _11036_, _11035_);
  nor _62004_ (_11038_, _11037_, _11033_);
  nor _62005_ (_11039_, _11038_, _11032_);
  nor _62006_ (_11040_, _11039_, _11030_);
  nor _62007_ (_11041_, _11040_, _11029_);
  or _62008_ (_11042_, _11041_, _11028_);
  nand _62009_ (_11043_, _11042_, _11027_);
  and _62010_ (_11044_, _11043_, _11024_);
  nor _62011_ (_11045_, _11044_, _11022_);
  or _62012_ (_11046_, _11045_, _11021_);
  nand _62013_ (_11047_, _11046_, _11020_);
  and _62014_ (_11048_, _11047_, _11018_);
  and _62015_ (_11049_, _11048_, _10705_);
  not _62016_ (_11050_, _10974_);
  nor _62017_ (_11051_, _11048_, _10705_);
  or _62018_ (_11052_, _11051_, _11050_);
  or _62019_ (_11053_, _11052_, _11049_);
  and _62020_ (_11054_, _11053_, _11016_);
  and _62021_ (_11055_, _11054_, _11014_);
  and _62022_ (_11056_, _11015_, \oc8051_golden_model_1.ACC [6]);
  or _62023_ (_11057_, _11056_, _06316_);
  or _62024_ (_11058_, _11057_, _11055_);
  and _62025_ (_11059_, _06114_, _05495_);
  not _62026_ (_11060_, _11059_);
  or _62027_ (_11061_, _10387_, _06718_);
  and _62028_ (_11062_, _11061_, _11060_);
  and _62029_ (_11063_, _11062_, _11058_);
  and _62030_ (_11064_, _06107_, _05495_);
  and _62031_ (_11065_, _10415_, _05758_);
  and _62032_ (_11066_, _11065_, _10010_);
  and _62033_ (_11067_, _11066_, _09880_);
  and _62034_ (_11068_, _11067_, _09906_);
  and _62035_ (_11069_, _11068_, _09861_);
  nor _62036_ (_11070_, _11069_, _08393_);
  and _62037_ (_11071_, _11069_, _08393_);
  or _62038_ (_11072_, _11071_, _11070_);
  and _62039_ (_11073_, _11072_, _11059_);
  or _62040_ (_11074_, _11073_, _11064_);
  or _62041_ (_11075_, _11074_, _11063_);
  nand _62042_ (_11076_, _11064_, _10606_);
  and _62043_ (_11077_, _11076_, _05653_);
  and _62044_ (_11078_, _11077_, _11075_);
  and _62045_ (_11079_, _10456_, _05652_);
  or _62046_ (_11080_, _11079_, _06047_);
  or _62047_ (_11081_, _11080_, _11078_);
  and _62048_ (_11082_, _06114_, _05750_);
  not _62049_ (_11083_, _11082_);
  and _62050_ (_11084_, _08279_, _07701_);
  or _62051_ (_11085_, _10385_, _06048_);
  or _62052_ (_11086_, _11085_, _11084_);
  and _62053_ (_11087_, _11086_, _11083_);
  and _62054_ (_11088_, _11087_, _11081_);
  and _62055_ (_11089_, _05750_, _06107_);
  and _62056_ (_11090_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  and _62057_ (_11091_, _11090_, \oc8051_golden_model_1.ACC [2]);
  and _62058_ (_11092_, _11091_, \oc8051_golden_model_1.ACC [3]);
  and _62059_ (_11093_, _11092_, \oc8051_golden_model_1.ACC [4]);
  and _62060_ (_11094_, _11093_, \oc8051_golden_model_1.ACC [5]);
  and _62061_ (_11095_, _11094_, \oc8051_golden_model_1.ACC [6]);
  or _62062_ (_11096_, _11095_, \oc8051_golden_model_1.ACC [7]);
  nand _62063_ (_11097_, _11095_, \oc8051_golden_model_1.ACC [7]);
  and _62064_ (_11098_, _11097_, _11096_);
  and _62065_ (_11099_, _11098_, _11082_);
  or _62066_ (_11100_, _11099_, _11089_);
  or _62067_ (_11101_, _11100_, _11088_);
  nand _62068_ (_11102_, _11089_, _05758_);
  and _62069_ (_11103_, _11102_, _01336_);
  and _62070_ (_11104_, _11103_, _11101_);
  or _62071_ (_11105_, _11104_, _10233_);
  and _62072_ (_40753_, _11105_, _42882_);
  not _62073_ (_11106_, \oc8051_golden_model_1.PCON [7]);
  nor _62074_ (_11107_, _01336_, _11106_);
  nor _62075_ (_11108_, _07641_, _11106_);
  not _62076_ (_11109_, _07641_);
  nor _62077_ (_11110_, _08767_, _11109_);
  or _62078_ (_11111_, _11110_, _11108_);
  and _62079_ (_11112_, _11111_, _06292_);
  or _62080_ (_11113_, _11108_, _07788_);
  and _62081_ (_11114_, _08549_, _07641_);
  or _62082_ (_11115_, _11114_, _11108_);
  and _62083_ (_11116_, _11115_, _06108_);
  and _62084_ (_11117_, _11116_, _11113_);
  and _62085_ (_11118_, _08768_, _07641_);
  or _62086_ (_11119_, _11118_, _11108_);
  and _62087_ (_11120_, _11119_, _06284_);
  or _62088_ (_11121_, _11115_, _06020_);
  and _62089_ (_11122_, _08498_, _07641_);
  or _62090_ (_11123_, _11122_, _11108_);
  or _62091_ (_11124_, _11123_, _06954_);
  and _62092_ (_11125_, _07641_, \oc8051_golden_model_1.ACC [7]);
  or _62093_ (_11126_, _11125_, _11108_);
  and _62094_ (_11127_, _11126_, _06938_);
  nor _62095_ (_11128_, _06938_, _11106_);
  or _62096_ (_11129_, _11128_, _06102_);
  or _62097_ (_11130_, _11129_, _11127_);
  and _62098_ (_11131_, _11130_, _06848_);
  and _62099_ (_11132_, _11131_, _11124_);
  nor _62100_ (_11133_, _07785_, _11109_);
  or _62101_ (_11134_, _11133_, _11108_);
  and _62102_ (_11135_, _11134_, _06239_);
  or _62103_ (_11136_, _11135_, _11132_);
  and _62104_ (_11137_, _11136_, _06220_);
  and _62105_ (_11138_, _11126_, _06219_);
  or _62106_ (_11139_, _11138_, _09818_);
  or _62107_ (_11140_, _11139_, _11137_);
  and _62108_ (_11141_, _08485_, _07641_);
  or _62109_ (_11142_, _11108_, _07012_);
  or _62110_ (_11143_, _11142_, _11141_);
  or _62111_ (_11144_, _11134_, _09827_);
  and _62112_ (_11145_, _11144_, _05669_);
  and _62113_ (_11146_, _11145_, _11143_);
  and _62114_ (_11147_, _11146_, _11140_);
  and _62115_ (_11148_, _08738_, _07641_);
  or _62116_ (_11149_, _11148_, _11108_);
  and _62117_ (_11150_, _11149_, _09833_);
  or _62118_ (_11151_, _11150_, _06019_);
  or _62119_ (_11152_, _11151_, _11147_);
  and _62120_ (_11153_, _11152_, _11121_);
  or _62121_ (_11154_, _11153_, _06112_);
  and _62122_ (_11155_, _08760_, _07641_);
  or _62123_ (_11156_, _11155_, _11108_);
  or _62124_ (_11157_, _11156_, _08751_);
  and _62125_ (_11158_, _11157_, _08756_);
  and _62126_ (_11159_, _11158_, _11154_);
  or _62127_ (_11160_, _11159_, _11120_);
  and _62128_ (_11161_, _11160_, _07032_);
  or _62129_ (_11162_, _11161_, _11117_);
  and _62130_ (_11163_, _11162_, _06278_);
  and _62131_ (_11164_, _11126_, _06277_);
  and _62132_ (_11165_, _11164_, _11113_);
  or _62133_ (_11166_, _11165_, _06130_);
  or _62134_ (_11167_, _11166_, _11163_);
  and _62135_ (_11168_, _08759_, _07641_);
  or _62136_ (_11169_, _11108_, _08777_);
  or _62137_ (_11170_, _11169_, _11168_);
  and _62138_ (_11171_, _11170_, _08782_);
  and _62139_ (_11172_, _11171_, _11167_);
  or _62140_ (_11173_, _11172_, _11112_);
  and _62141_ (_11174_, _11173_, _06718_);
  and _62142_ (_11175_, _11123_, _06316_);
  or _62143_ (_11176_, _11175_, _06047_);
  or _62144_ (_11177_, _11176_, _11174_);
  and _62145_ (_11178_, _08279_, _07641_);
  or _62146_ (_11179_, _11108_, _06048_);
  or _62147_ (_11180_, _11179_, _11178_);
  and _62148_ (_11181_, _11180_, _01336_);
  and _62149_ (_11182_, _11181_, _11177_);
  or _62150_ (_11183_, _11182_, _11107_);
  and _62151_ (_40756_, _11183_, _42882_);
  and _62152_ (_11184_, _01340_, \oc8051_golden_model_1.TMOD [7]);
  not _62153_ (_11185_, _07653_);
  and _62154_ (_11186_, _11185_, \oc8051_golden_model_1.TMOD [7]);
  nor _62155_ (_11187_, _08767_, _11185_);
  or _62156_ (_11188_, _11187_, _11186_);
  and _62157_ (_11189_, _11188_, _06292_);
  and _62158_ (_11190_, _08768_, _07653_);
  or _62159_ (_11191_, _11190_, _11186_);
  and _62160_ (_11192_, _11191_, _06284_);
  and _62161_ (_11193_, _08549_, _07653_);
  or _62162_ (_11194_, _11193_, _11186_);
  or _62163_ (_11195_, _11194_, _06020_);
  and _62164_ (_11196_, _08498_, _07653_);
  or _62165_ (_11197_, _11196_, _11186_);
  or _62166_ (_11198_, _11197_, _06954_);
  and _62167_ (_11199_, _07653_, \oc8051_golden_model_1.ACC [7]);
  or _62168_ (_11200_, _11199_, _11186_);
  and _62169_ (_11201_, _11200_, _06938_);
  and _62170_ (_11202_, _06939_, \oc8051_golden_model_1.TMOD [7]);
  or _62171_ (_11203_, _11202_, _06102_);
  or _62172_ (_11204_, _11203_, _11201_);
  and _62173_ (_11205_, _11204_, _06848_);
  and _62174_ (_11206_, _11205_, _11198_);
  nor _62175_ (_11207_, _07785_, _11185_);
  or _62176_ (_11208_, _11207_, _11186_);
  and _62177_ (_11209_, _11208_, _06239_);
  or _62178_ (_11210_, _11209_, _11206_);
  and _62179_ (_11211_, _11210_, _06220_);
  and _62180_ (_11212_, _11200_, _06219_);
  or _62181_ (_11213_, _11212_, _09818_);
  or _62182_ (_11214_, _11213_, _11211_);
  and _62183_ (_11215_, _08485_, _07653_);
  or _62184_ (_11216_, _11186_, _07012_);
  or _62185_ (_11217_, _11216_, _11215_);
  or _62186_ (_11218_, _11208_, _09827_);
  and _62187_ (_11219_, _11218_, _05669_);
  and _62188_ (_11220_, _11219_, _11217_);
  and _62189_ (_11221_, _11220_, _11214_);
  and _62190_ (_11222_, _08738_, _07653_);
  or _62191_ (_11223_, _11222_, _11186_);
  and _62192_ (_11224_, _11223_, _09833_);
  or _62193_ (_11225_, _11224_, _06019_);
  or _62194_ (_11226_, _11225_, _11221_);
  and _62195_ (_11227_, _11226_, _11195_);
  or _62196_ (_11228_, _11227_, _06112_);
  and _62197_ (_11229_, _08760_, _07653_);
  or _62198_ (_11230_, _11186_, _08751_);
  or _62199_ (_11231_, _11230_, _11229_);
  and _62200_ (_11232_, _11231_, _08756_);
  and _62201_ (_11233_, _11232_, _11228_);
  or _62202_ (_11234_, _11233_, _11192_);
  and _62203_ (_11235_, _11234_, _07032_);
  or _62204_ (_11236_, _11186_, _07788_);
  and _62205_ (_11237_, _11194_, _06108_);
  and _62206_ (_11238_, _11237_, _11236_);
  or _62207_ (_11239_, _11238_, _11235_);
  and _62208_ (_11240_, _11239_, _06278_);
  and _62209_ (_11241_, _11200_, _06277_);
  and _62210_ (_11242_, _11241_, _11236_);
  or _62211_ (_11243_, _11242_, _06130_);
  or _62212_ (_11244_, _11243_, _11240_);
  and _62213_ (_11245_, _08759_, _07653_);
  or _62214_ (_11246_, _11186_, _08777_);
  or _62215_ (_11247_, _11246_, _11245_);
  and _62216_ (_11248_, _11247_, _08782_);
  and _62217_ (_11249_, _11248_, _11244_);
  or _62218_ (_11250_, _11249_, _11189_);
  and _62219_ (_11251_, _11250_, _06718_);
  and _62220_ (_11252_, _11197_, _06316_);
  or _62221_ (_11253_, _11252_, _06047_);
  or _62222_ (_11254_, _11253_, _11251_);
  and _62223_ (_11255_, _08279_, _07653_);
  or _62224_ (_11256_, _11186_, _06048_);
  or _62225_ (_11257_, _11256_, _11255_);
  and _62226_ (_11258_, _11257_, _01336_);
  and _62227_ (_11259_, _11258_, _11254_);
  or _62228_ (_11260_, _11259_, _11184_);
  and _62229_ (_40757_, _11260_, _42882_);
  not _62230_ (_11261_, \oc8051_golden_model_1.DPL [7]);
  nor _62231_ (_11262_, _01336_, _11261_);
  nor _62232_ (_11263_, _07733_, _11261_);
  not _62233_ (_11264_, _07733_);
  nor _62234_ (_11265_, _08767_, _11264_);
  or _62235_ (_11266_, _11265_, _11263_);
  and _62236_ (_11267_, _11266_, _06292_);
  and _62237_ (_11268_, _08768_, _07733_);
  or _62238_ (_11269_, _11268_, _11263_);
  and _62239_ (_11270_, _11269_, _06284_);
  and _62240_ (_11271_, _08549_, _07733_);
  or _62241_ (_11272_, _11271_, _11263_);
  or _62242_ (_11273_, _11272_, _06020_);
  and _62243_ (_11274_, _08498_, _07733_);
  or _62244_ (_11275_, _11274_, _11263_);
  or _62245_ (_11276_, _11275_, _06954_);
  and _62246_ (_11277_, _07733_, \oc8051_golden_model_1.ACC [7]);
  or _62247_ (_11278_, _11277_, _11263_);
  and _62248_ (_11279_, _11278_, _06938_);
  nor _62249_ (_11280_, _06938_, _11261_);
  or _62250_ (_11281_, _11280_, _06102_);
  or _62251_ (_11282_, _11281_, _11279_);
  and _62252_ (_11283_, _11282_, _06848_);
  and _62253_ (_11284_, _11283_, _11276_);
  nor _62254_ (_11285_, _07785_, _11264_);
  or _62255_ (_11286_, _11285_, _11263_);
  and _62256_ (_11287_, _11286_, _06239_);
  or _62257_ (_11288_, _11287_, _06219_);
  or _62258_ (_11289_, _11288_, _11284_);
  nor _62259_ (_11290_, _05701_, _05662_);
  not _62260_ (_11291_, _11290_);
  or _62261_ (_11292_, _11278_, _06220_);
  and _62262_ (_11293_, _11292_, _11291_);
  and _62263_ (_11294_, _11293_, _11289_);
  and _62264_ (_11295_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  and _62265_ (_11296_, _11295_, \oc8051_golden_model_1.DPL [2]);
  and _62266_ (_11297_, _11296_, \oc8051_golden_model_1.DPL [3]);
  and _62267_ (_11298_, _11297_, \oc8051_golden_model_1.DPL [4]);
  and _62268_ (_11299_, _11298_, \oc8051_golden_model_1.DPL [5]);
  and _62269_ (_11300_, _11299_, \oc8051_golden_model_1.DPL [6]);
  nor _62270_ (_11301_, _11300_, \oc8051_golden_model_1.DPL [7]);
  and _62271_ (_11302_, _11300_, \oc8051_golden_model_1.DPL [7]);
  nor _62272_ (_11303_, _11302_, _11301_);
  and _62273_ (_11304_, _11303_, _11290_);
  or _62274_ (_11305_, _11304_, _11294_);
  and _62275_ (_11306_, _11305_, _06111_);
  nor _62276_ (_11307_, _08332_, _06111_);
  or _62277_ (_11308_, _11307_, _09818_);
  or _62278_ (_11309_, _11308_, _11306_);
  and _62279_ (_11310_, _08485_, _07733_);
  or _62280_ (_11311_, _11263_, _07012_);
  or _62281_ (_11312_, _11311_, _11310_);
  or _62282_ (_11313_, _11286_, _09827_);
  and _62283_ (_11314_, _11313_, _05669_);
  and _62284_ (_11315_, _11314_, _11312_);
  and _62285_ (_11316_, _11315_, _11309_);
  and _62286_ (_11317_, _08738_, _07733_);
  or _62287_ (_11318_, _11317_, _11263_);
  and _62288_ (_11319_, _11318_, _09833_);
  or _62289_ (_11320_, _11319_, _06019_);
  or _62290_ (_11321_, _11320_, _11316_);
  and _62291_ (_11322_, _11321_, _11273_);
  or _62292_ (_11323_, _11322_, _06112_);
  and _62293_ (_11324_, _08760_, _07733_);
  or _62294_ (_11325_, _11263_, _08751_);
  or _62295_ (_11326_, _11325_, _11324_);
  and _62296_ (_11327_, _11326_, _08756_);
  and _62297_ (_11328_, _11327_, _11323_);
  or _62298_ (_11329_, _11328_, _11270_);
  and _62299_ (_11330_, _11329_, _07032_);
  or _62300_ (_11331_, _11263_, _07788_);
  and _62301_ (_11332_, _11272_, _06108_);
  and _62302_ (_11333_, _11332_, _11331_);
  or _62303_ (_11334_, _11333_, _11330_);
  and _62304_ (_11335_, _11334_, _06278_);
  and _62305_ (_11336_, _11278_, _06277_);
  and _62306_ (_11337_, _11336_, _11331_);
  or _62307_ (_11338_, _11337_, _06130_);
  or _62308_ (_11339_, _11338_, _11335_);
  and _62309_ (_11340_, _08759_, _07733_);
  or _62310_ (_11341_, _11263_, _08777_);
  or _62311_ (_11342_, _11341_, _11340_);
  and _62312_ (_11343_, _11342_, _08782_);
  and _62313_ (_11344_, _11343_, _11339_);
  or _62314_ (_11345_, _11344_, _11267_);
  and _62315_ (_11346_, _11345_, _06718_);
  and _62316_ (_11347_, _11275_, _06316_);
  or _62317_ (_11348_, _11347_, _06047_);
  or _62318_ (_11349_, _11348_, _11346_);
  and _62319_ (_11350_, _08279_, _07733_);
  or _62320_ (_11351_, _11263_, _06048_);
  or _62321_ (_11352_, _11351_, _11350_);
  and _62322_ (_11353_, _11352_, _01336_);
  and _62323_ (_11354_, _11353_, _11349_);
  or _62324_ (_11355_, _11354_, _11262_);
  and _62325_ (_40758_, _11355_, _42882_);
  not _62326_ (_11356_, \oc8051_golden_model_1.DPH [7]);
  nor _62327_ (_11357_, _01336_, _11356_);
  nor _62328_ (_11358_, _07802_, _11356_);
  not _62329_ (_11359_, _07724_);
  nor _62330_ (_11360_, _08767_, _11359_);
  or _62331_ (_11361_, _11360_, _11358_);
  and _62332_ (_11362_, _11361_, _06292_);
  and _62333_ (_11363_, _08768_, _07724_);
  or _62334_ (_11364_, _11363_, _11358_);
  and _62335_ (_11365_, _11364_, _06284_);
  and _62336_ (_11366_, _08549_, _07802_);
  or _62337_ (_11367_, _11366_, _11358_);
  or _62338_ (_11368_, _11367_, _06020_);
  and _62339_ (_11369_, _08498_, _07724_);
  or _62340_ (_11370_, _11369_, _11358_);
  or _62341_ (_11371_, _11370_, _06954_);
  and _62342_ (_11372_, _07802_, \oc8051_golden_model_1.ACC [7]);
  or _62343_ (_11373_, _11372_, _11358_);
  and _62344_ (_11374_, _11373_, _06938_);
  nor _62345_ (_11375_, _06938_, _11356_);
  or _62346_ (_11376_, _11375_, _06102_);
  or _62347_ (_11377_, _11376_, _11374_);
  and _62348_ (_11378_, _11377_, _06848_);
  and _62349_ (_11379_, _11378_, _11371_);
  nor _62350_ (_11380_, _07785_, _11359_);
  or _62351_ (_11381_, _11380_, _11358_);
  and _62352_ (_11382_, _11381_, _06239_);
  or _62353_ (_11383_, _11382_, _06219_);
  or _62354_ (_11384_, _11383_, _11379_);
  or _62355_ (_11385_, _11373_, _06220_);
  and _62356_ (_11386_, _11385_, _11291_);
  and _62357_ (_11387_, _11386_, _11384_);
  and _62358_ (_11388_, _11302_, \oc8051_golden_model_1.DPH [0]);
  and _62359_ (_11389_, _11388_, \oc8051_golden_model_1.DPH [1]);
  and _62360_ (_11390_, _11389_, \oc8051_golden_model_1.DPH [2]);
  and _62361_ (_11391_, _11390_, \oc8051_golden_model_1.DPH [3]);
  and _62362_ (_11392_, _11391_, \oc8051_golden_model_1.DPH [4]);
  and _62363_ (_11393_, _11392_, \oc8051_golden_model_1.DPH [5]);
  and _62364_ (_11394_, _11393_, \oc8051_golden_model_1.DPH [6]);
  nand _62365_ (_11395_, _11394_, \oc8051_golden_model_1.DPH [7]);
  or _62366_ (_11396_, _11394_, \oc8051_golden_model_1.DPH [7]);
  and _62367_ (_11397_, _11396_, _11290_);
  and _62368_ (_11398_, _11397_, _11395_);
  or _62369_ (_11399_, _11398_, _11387_);
  and _62370_ (_11400_, _11399_, _06111_);
  and _62371_ (_11401_, _06110_, _05952_);
  or _62372_ (_11402_, _11401_, _09818_);
  or _62373_ (_11403_, _11402_, _11400_);
  or _62374_ (_11404_, _11358_, _07012_);
  and _62375_ (_11405_, _08485_, _07802_);
  or _62376_ (_11406_, _11405_, _11404_);
  or _62377_ (_11407_, _11381_, _09827_);
  and _62378_ (_11408_, _11407_, _05669_);
  and _62379_ (_11409_, _11408_, _11406_);
  and _62380_ (_11410_, _11409_, _11403_);
  and _62381_ (_11411_, _08738_, _07724_);
  or _62382_ (_11412_, _11411_, _11358_);
  and _62383_ (_11413_, _11412_, _09833_);
  or _62384_ (_11414_, _11413_, _06019_);
  or _62385_ (_11415_, _11414_, _11410_);
  and _62386_ (_11416_, _11415_, _11368_);
  or _62387_ (_11417_, _11416_, _06112_);
  and _62388_ (_11418_, _08760_, _07724_);
  or _62389_ (_11419_, _11358_, _08751_);
  or _62390_ (_11420_, _11419_, _11418_);
  and _62391_ (_11421_, _11420_, _08756_);
  and _62392_ (_11422_, _11421_, _11417_);
  or _62393_ (_11423_, _11422_, _11365_);
  and _62394_ (_11424_, _11423_, _07032_);
  or _62395_ (_11425_, _11358_, _07788_);
  and _62396_ (_11426_, _11367_, _06108_);
  and _62397_ (_11427_, _11426_, _11425_);
  or _62398_ (_11428_, _11427_, _11424_);
  and _62399_ (_11429_, _11428_, _06278_);
  and _62400_ (_11430_, _11373_, _06277_);
  and _62401_ (_11431_, _11430_, _11425_);
  or _62402_ (_11432_, _11431_, _06130_);
  or _62403_ (_11433_, _11432_, _11429_);
  and _62404_ (_11434_, _08759_, _07724_);
  or _62405_ (_11435_, _11358_, _08777_);
  or _62406_ (_11436_, _11435_, _11434_);
  and _62407_ (_11437_, _11436_, _08782_);
  and _62408_ (_11438_, _11437_, _11433_);
  or _62409_ (_11439_, _11438_, _11362_);
  and _62410_ (_11440_, _11439_, _06718_);
  and _62411_ (_11441_, _11370_, _06316_);
  or _62412_ (_11442_, _11441_, _06047_);
  or _62413_ (_11443_, _11442_, _11440_);
  and _62414_ (_11444_, _08279_, _07724_);
  or _62415_ (_11445_, _11358_, _06048_);
  or _62416_ (_11446_, _11445_, _11444_);
  and _62417_ (_11447_, _11446_, _01336_);
  and _62418_ (_11448_, _11447_, _11443_);
  or _62419_ (_11449_, _11448_, _11357_);
  and _62420_ (_40759_, _11449_, _42882_);
  and _62421_ (_11450_, _01340_, \oc8051_golden_model_1.TL1 [7]);
  not _62422_ (_11451_, _07667_);
  and _62423_ (_11452_, _11451_, \oc8051_golden_model_1.TL1 [7]);
  nor _62424_ (_11453_, _08767_, _11451_);
  or _62425_ (_11454_, _11453_, _11452_);
  and _62426_ (_11455_, _11454_, _06292_);
  and _62427_ (_11456_, _08768_, _07667_);
  or _62428_ (_11457_, _11456_, _11452_);
  and _62429_ (_11458_, _11457_, _06284_);
  and _62430_ (_11459_, _08549_, _07667_);
  or _62431_ (_11460_, _11459_, _11452_);
  or _62432_ (_11461_, _11460_, _06020_);
  and _62433_ (_11462_, _08498_, _07667_);
  or _62434_ (_11463_, _11462_, _11452_);
  or _62435_ (_11464_, _11463_, _06954_);
  and _62436_ (_11465_, _07667_, \oc8051_golden_model_1.ACC [7]);
  or _62437_ (_11466_, _11465_, _11452_);
  and _62438_ (_11467_, _11466_, _06938_);
  and _62439_ (_11468_, _06939_, \oc8051_golden_model_1.TL1 [7]);
  or _62440_ (_11469_, _11468_, _06102_);
  or _62441_ (_11470_, _11469_, _11467_);
  and _62442_ (_11471_, _11470_, _06848_);
  and _62443_ (_11472_, _11471_, _11464_);
  nor _62444_ (_11473_, _07785_, _11451_);
  or _62445_ (_11474_, _11473_, _11452_);
  and _62446_ (_11475_, _11474_, _06239_);
  or _62447_ (_11476_, _11475_, _11472_);
  and _62448_ (_11477_, _11476_, _06220_);
  and _62449_ (_11478_, _11466_, _06219_);
  or _62450_ (_11479_, _11478_, _09818_);
  or _62451_ (_11480_, _11479_, _11477_);
  and _62452_ (_11481_, _08485_, _07667_);
  or _62453_ (_11482_, _11452_, _07012_);
  or _62454_ (_11483_, _11482_, _11481_);
  or _62455_ (_11484_, _11474_, _09827_);
  and _62456_ (_11485_, _11484_, _05669_);
  and _62457_ (_11486_, _11485_, _11483_);
  and _62458_ (_11487_, _11486_, _11480_);
  and _62459_ (_11488_, _08738_, _07667_);
  or _62460_ (_11489_, _11488_, _11452_);
  and _62461_ (_11490_, _11489_, _09833_);
  or _62462_ (_11491_, _11490_, _06019_);
  or _62463_ (_11492_, _11491_, _11487_);
  and _62464_ (_11493_, _11492_, _11461_);
  or _62465_ (_11494_, _11493_, _06112_);
  and _62466_ (_11495_, _08760_, _07667_);
  or _62467_ (_11496_, _11495_, _11452_);
  or _62468_ (_11497_, _11496_, _08751_);
  and _62469_ (_11498_, _11497_, _08756_);
  and _62470_ (_11499_, _11498_, _11494_);
  or _62471_ (_11500_, _11499_, _11458_);
  and _62472_ (_11501_, _11500_, _07032_);
  or _62473_ (_11502_, _11452_, _07788_);
  and _62474_ (_11503_, _11460_, _06108_);
  and _62475_ (_11504_, _11503_, _11502_);
  or _62476_ (_11505_, _11504_, _11501_);
  and _62477_ (_11506_, _11505_, _06278_);
  and _62478_ (_11507_, _11466_, _06277_);
  and _62479_ (_11508_, _11507_, _11502_);
  or _62480_ (_11509_, _11508_, _06130_);
  or _62481_ (_11510_, _11509_, _11506_);
  and _62482_ (_11511_, _08759_, _07667_);
  or _62483_ (_11512_, _11452_, _08777_);
  or _62484_ (_11513_, _11512_, _11511_);
  and _62485_ (_11514_, _11513_, _08782_);
  and _62486_ (_11515_, _11514_, _11510_);
  or _62487_ (_11516_, _11515_, _11455_);
  and _62488_ (_11517_, _11516_, _06718_);
  and _62489_ (_11518_, _11463_, _06316_);
  or _62490_ (_11519_, _11518_, _06047_);
  or _62491_ (_11520_, _11519_, _11517_);
  and _62492_ (_11521_, _08279_, _07667_);
  or _62493_ (_11522_, _11452_, _06048_);
  or _62494_ (_11523_, _11522_, _11521_);
  and _62495_ (_11524_, _11523_, _01336_);
  and _62496_ (_11525_, _11524_, _11520_);
  or _62497_ (_11526_, _11525_, _11450_);
  and _62498_ (_40760_, _11526_, _42882_);
  and _62499_ (_11527_, _01340_, \oc8051_golden_model_1.TL0 [7]);
  not _62500_ (_11528_, _07659_);
  and _62501_ (_11529_, _11528_, \oc8051_golden_model_1.TL0 [7]);
  nor _62502_ (_11530_, _08767_, _11528_);
  or _62503_ (_11531_, _11530_, _11529_);
  and _62504_ (_11532_, _11531_, _06292_);
  and _62505_ (_11533_, _08768_, _07659_);
  or _62506_ (_11534_, _11533_, _11529_);
  and _62507_ (_11535_, _11534_, _06284_);
  and _62508_ (_11536_, _08549_, _07659_);
  or _62509_ (_11537_, _11536_, _11529_);
  or _62510_ (_11538_, _11537_, _06020_);
  and _62511_ (_11539_, _08498_, _07659_);
  or _62512_ (_11540_, _11539_, _11529_);
  or _62513_ (_11541_, _11540_, _06954_);
  and _62514_ (_11542_, _07659_, \oc8051_golden_model_1.ACC [7]);
  or _62515_ (_11543_, _11542_, _11529_);
  and _62516_ (_11544_, _11543_, _06938_);
  and _62517_ (_11545_, _06939_, \oc8051_golden_model_1.TL0 [7]);
  or _62518_ (_11546_, _11545_, _06102_);
  or _62519_ (_11547_, _11546_, _11544_);
  and _62520_ (_11548_, _11547_, _06848_);
  and _62521_ (_11549_, _11548_, _11541_);
  nor _62522_ (_11550_, _07785_, _11528_);
  or _62523_ (_11551_, _11550_, _11529_);
  and _62524_ (_11552_, _11551_, _06239_);
  or _62525_ (_11553_, _11552_, _11549_);
  and _62526_ (_11554_, _11553_, _06220_);
  and _62527_ (_11555_, _11543_, _06219_);
  or _62528_ (_11556_, _11555_, _09818_);
  or _62529_ (_11557_, _11556_, _11554_);
  and _62530_ (_11558_, _08485_, _07659_);
  or _62531_ (_11559_, _11529_, _07012_);
  or _62532_ (_11560_, _11559_, _11558_);
  or _62533_ (_11561_, _11551_, _09827_);
  and _62534_ (_11562_, _11561_, _05669_);
  and _62535_ (_11563_, _11562_, _11560_);
  and _62536_ (_11564_, _11563_, _11557_);
  and _62537_ (_11565_, _08738_, _07659_);
  or _62538_ (_11566_, _11565_, _11529_);
  and _62539_ (_11567_, _11566_, _09833_);
  or _62540_ (_11568_, _11567_, _06019_);
  or _62541_ (_11569_, _11568_, _11564_);
  and _62542_ (_11570_, _11569_, _11538_);
  or _62543_ (_11571_, _11570_, _06112_);
  and _62544_ (_11572_, _08760_, _07659_);
  or _62545_ (_11573_, _11529_, _08751_);
  or _62546_ (_11574_, _11573_, _11572_);
  and _62547_ (_11575_, _11574_, _08756_);
  and _62548_ (_11576_, _11575_, _11571_);
  or _62549_ (_11577_, _11576_, _11535_);
  and _62550_ (_11578_, _11577_, _07032_);
  or _62551_ (_11579_, _11529_, _07788_);
  and _62552_ (_11580_, _11537_, _06108_);
  and _62553_ (_11581_, _11580_, _11579_);
  or _62554_ (_11582_, _11581_, _11578_);
  and _62555_ (_11583_, _11582_, _06278_);
  and _62556_ (_11584_, _11543_, _06277_);
  and _62557_ (_11585_, _11584_, _11579_);
  or _62558_ (_11586_, _11585_, _06130_);
  or _62559_ (_11587_, _11586_, _11583_);
  and _62560_ (_11588_, _08759_, _07659_);
  or _62561_ (_11589_, _11529_, _08777_);
  or _62562_ (_11590_, _11589_, _11588_);
  and _62563_ (_11591_, _11590_, _08782_);
  and _62564_ (_11592_, _11591_, _11587_);
  or _62565_ (_11593_, _11592_, _11532_);
  and _62566_ (_11594_, _11593_, _06718_);
  and _62567_ (_11595_, _11540_, _06316_);
  or _62568_ (_11596_, _11595_, _06047_);
  or _62569_ (_11597_, _11596_, _11594_);
  and _62570_ (_11598_, _08279_, _07659_);
  or _62571_ (_11599_, _11529_, _06048_);
  or _62572_ (_11600_, _11599_, _11598_);
  and _62573_ (_11601_, _11600_, _01336_);
  and _62574_ (_11602_, _11601_, _11597_);
  or _62575_ (_11603_, _11602_, _11527_);
  and _62576_ (_40762_, _11603_, _42882_);
  and _62577_ (_11604_, _01340_, \oc8051_golden_model_1.TCON [7]);
  not _62578_ (_11605_, _07648_);
  and _62579_ (_11606_, _11605_, \oc8051_golden_model_1.TCON [7]);
  and _62580_ (_11607_, _08768_, _07648_);
  or _62581_ (_11608_, _11607_, _11606_);
  and _62582_ (_11609_, _11608_, _06284_);
  and _62583_ (_11610_, _08549_, _07648_);
  or _62584_ (_11611_, _11610_, _11606_);
  or _62585_ (_11612_, _11611_, _06020_);
  and _62586_ (_11613_, _08498_, _07648_);
  or _62587_ (_11614_, _11613_, _11606_);
  or _62588_ (_11615_, _11614_, _06954_);
  and _62589_ (_11616_, _07648_, \oc8051_golden_model_1.ACC [7]);
  or _62590_ (_11617_, _11616_, _11606_);
  and _62591_ (_11618_, _11617_, _06938_);
  and _62592_ (_11619_, _06939_, \oc8051_golden_model_1.TCON [7]);
  or _62593_ (_11620_, _11619_, _06102_);
  or _62594_ (_11621_, _11620_, _11618_);
  and _62595_ (_11622_, _11621_, _06044_);
  and _62596_ (_11623_, _11622_, _11615_);
  not _62597_ (_11624_, _08341_);
  and _62598_ (_11625_, _11624_, \oc8051_golden_model_1.TCON [7]);
  and _62599_ (_11626_, _08503_, _08341_);
  or _62600_ (_11627_, _11626_, _11625_);
  and _62601_ (_11628_, _11627_, _06043_);
  or _62602_ (_11629_, _11628_, _06239_);
  or _62603_ (_11630_, _11629_, _11623_);
  nor _62604_ (_11631_, _07785_, _11605_);
  or _62605_ (_11632_, _11631_, _11606_);
  or _62606_ (_11633_, _11632_, _06848_);
  and _62607_ (_11634_, _11633_, _11630_);
  or _62608_ (_11635_, _11634_, _06219_);
  or _62609_ (_11636_, _11617_, _06220_);
  and _62610_ (_11637_, _11636_, _06040_);
  and _62611_ (_11638_, _11637_, _11635_);
  and _62612_ (_11639_, _08374_, _08341_);
  or _62613_ (_11640_, _11639_, _11625_);
  and _62614_ (_11641_, _11640_, _06039_);
  or _62615_ (_11642_, _11641_, _06032_);
  or _62616_ (_11643_, _11642_, _11638_);
  or _62617_ (_11644_, _11625_, _08519_);
  and _62618_ (_11645_, _11644_, _11627_);
  or _62619_ (_11646_, _11645_, _06033_);
  and _62620_ (_11647_, _11646_, _06027_);
  and _62621_ (_11648_, _11647_, _11643_);
  and _62622_ (_11649_, _08376_, _08341_);
  or _62623_ (_11650_, _11649_, _11625_);
  and _62624_ (_11651_, _11650_, _06026_);
  or _62625_ (_11652_, _11651_, _09818_);
  or _62626_ (_11653_, _11652_, _11648_);
  and _62627_ (_11654_, _08485_, _07648_);
  or _62628_ (_11655_, _11606_, _07012_);
  or _62629_ (_11656_, _11655_, _11654_);
  or _62630_ (_11657_, _11632_, _09827_);
  and _62631_ (_11658_, _11657_, _05669_);
  and _62632_ (_11659_, _11658_, _11656_);
  and _62633_ (_11660_, _11659_, _11653_);
  and _62634_ (_11661_, _08738_, _07648_);
  or _62635_ (_11662_, _11661_, _11606_);
  and _62636_ (_11663_, _11662_, _09833_);
  or _62637_ (_11664_, _11663_, _06019_);
  or _62638_ (_11665_, _11664_, _11660_);
  and _62639_ (_11666_, _11665_, _11612_);
  or _62640_ (_11667_, _11666_, _06112_);
  and _62641_ (_11668_, _08760_, _07648_);
  or _62642_ (_11669_, _11606_, _08751_);
  or _62643_ (_11670_, _11669_, _11668_);
  and _62644_ (_11671_, _11670_, _08756_);
  and _62645_ (_11672_, _11671_, _11667_);
  or _62646_ (_11673_, _11672_, _11609_);
  and _62647_ (_11674_, _11673_, _07032_);
  or _62648_ (_11675_, _11606_, _07788_);
  and _62649_ (_11676_, _11611_, _06108_);
  and _62650_ (_11677_, _11676_, _11675_);
  or _62651_ (_11678_, _11677_, _11674_);
  and _62652_ (_11679_, _11678_, _06278_);
  and _62653_ (_11680_, _11617_, _06277_);
  and _62654_ (_11681_, _11680_, _11675_);
  or _62655_ (_11682_, _11681_, _06130_);
  or _62656_ (_11683_, _11682_, _11679_);
  and _62657_ (_11684_, _08759_, _07648_);
  or _62658_ (_11685_, _11606_, _08777_);
  or _62659_ (_11686_, _11685_, _11684_);
  and _62660_ (_11687_, _11686_, _08782_);
  and _62661_ (_11688_, _11687_, _11683_);
  nor _62662_ (_11689_, _08767_, _11605_);
  or _62663_ (_11690_, _11689_, _11606_);
  and _62664_ (_11691_, _11690_, _06292_);
  or _62665_ (_11692_, _11691_, _06316_);
  or _62666_ (_11693_, _11692_, _11688_);
  or _62667_ (_11694_, _11614_, _06718_);
  and _62668_ (_11695_, _11694_, _05653_);
  and _62669_ (_11696_, _11695_, _11693_);
  and _62670_ (_11697_, _11640_, _05652_);
  or _62671_ (_11698_, _11697_, _06047_);
  or _62672_ (_11699_, _11698_, _11696_);
  and _62673_ (_11700_, _08279_, _07648_);
  or _62674_ (_11701_, _11606_, _06048_);
  or _62675_ (_11702_, _11701_, _11700_);
  and _62676_ (_11703_, _11702_, _01336_);
  and _62677_ (_11704_, _11703_, _11699_);
  or _62678_ (_11705_, _11704_, _11604_);
  and _62679_ (_40763_, _11705_, _42882_);
  and _62680_ (_11706_, _01340_, \oc8051_golden_model_1.TH1 [7]);
  not _62681_ (_11707_, _07670_);
  and _62682_ (_11708_, _11707_, \oc8051_golden_model_1.TH1 [7]);
  nor _62683_ (_11709_, _08767_, _11707_);
  or _62684_ (_11710_, _11709_, _11708_);
  and _62685_ (_11711_, _11710_, _06292_);
  or _62686_ (_11712_, _11708_, _07788_);
  and _62687_ (_11713_, _08549_, _07670_);
  or _62688_ (_11714_, _11713_, _11708_);
  and _62689_ (_11715_, _11714_, _06108_);
  and _62690_ (_11716_, _11715_, _11712_);
  and _62691_ (_11717_, _08768_, _07670_);
  or _62692_ (_11718_, _11717_, _11708_);
  and _62693_ (_11719_, _11718_, _06284_);
  or _62694_ (_11720_, _11714_, _06020_);
  and _62695_ (_11721_, _08498_, _07670_);
  or _62696_ (_11722_, _11721_, _11708_);
  or _62697_ (_11723_, _11722_, _06954_);
  and _62698_ (_11724_, _07670_, \oc8051_golden_model_1.ACC [7]);
  or _62699_ (_11725_, _11724_, _11708_);
  and _62700_ (_11726_, _11725_, _06938_);
  and _62701_ (_11727_, _06939_, \oc8051_golden_model_1.TH1 [7]);
  or _62702_ (_11728_, _11727_, _06102_);
  or _62703_ (_11729_, _11728_, _11726_);
  and _62704_ (_11730_, _11729_, _06848_);
  and _62705_ (_11731_, _11730_, _11723_);
  nor _62706_ (_11732_, _07785_, _11707_);
  or _62707_ (_11733_, _11732_, _11708_);
  and _62708_ (_11734_, _11733_, _06239_);
  or _62709_ (_11735_, _11734_, _11731_);
  and _62710_ (_11736_, _11735_, _06220_);
  and _62711_ (_11737_, _11725_, _06219_);
  or _62712_ (_11738_, _11737_, _09818_);
  or _62713_ (_11739_, _11738_, _11736_);
  and _62714_ (_11740_, _08485_, _07670_);
  or _62715_ (_11741_, _11708_, _07012_);
  or _62716_ (_11742_, _11741_, _11740_);
  or _62717_ (_11743_, _11733_, _09827_);
  and _62718_ (_11744_, _11743_, _05669_);
  and _62719_ (_11745_, _11744_, _11742_);
  and _62720_ (_11746_, _11745_, _11739_);
  and _62721_ (_11747_, _08738_, _07670_);
  or _62722_ (_11748_, _11747_, _11708_);
  and _62723_ (_11749_, _11748_, _09833_);
  or _62724_ (_11750_, _11749_, _06019_);
  or _62725_ (_11751_, _11750_, _11746_);
  and _62726_ (_11752_, _11751_, _11720_);
  or _62727_ (_11753_, _11752_, _06112_);
  and _62728_ (_11754_, _08760_, _07670_);
  or _62729_ (_11755_, _11754_, _11708_);
  or _62730_ (_11756_, _11755_, _08751_);
  and _62731_ (_11757_, _11756_, _08756_);
  and _62732_ (_11758_, _11757_, _11753_);
  or _62733_ (_11759_, _11758_, _11719_);
  and _62734_ (_11760_, _11759_, _07032_);
  or _62735_ (_11761_, _11760_, _11716_);
  and _62736_ (_11762_, _11761_, _06278_);
  and _62737_ (_11763_, _11725_, _06277_);
  and _62738_ (_11764_, _11763_, _11712_);
  or _62739_ (_11765_, _11764_, _06130_);
  or _62740_ (_11766_, _11765_, _11762_);
  and _62741_ (_11767_, _08759_, _07670_);
  or _62742_ (_11768_, _11708_, _08777_);
  or _62743_ (_11769_, _11768_, _11767_);
  and _62744_ (_11770_, _11769_, _08782_);
  and _62745_ (_11771_, _11770_, _11766_);
  or _62746_ (_11772_, _11771_, _11711_);
  and _62747_ (_11773_, _11772_, _06718_);
  and _62748_ (_11774_, _11722_, _06316_);
  or _62749_ (_11775_, _11774_, _06047_);
  or _62750_ (_11776_, _11775_, _11773_);
  and _62751_ (_11777_, _08279_, _07670_);
  or _62752_ (_11778_, _11708_, _06048_);
  or _62753_ (_11779_, _11778_, _11777_);
  and _62754_ (_11780_, _11779_, _01336_);
  and _62755_ (_11781_, _11780_, _11776_);
  or _62756_ (_11782_, _11781_, _11706_);
  and _62757_ (_40764_, _11782_, _42882_);
  and _62758_ (_11783_, _01340_, \oc8051_golden_model_1.TH0 [7]);
  not _62759_ (_11784_, _07663_);
  and _62760_ (_11785_, _11784_, \oc8051_golden_model_1.TH0 [7]);
  nor _62761_ (_11786_, _08767_, _11784_);
  or _62762_ (_11787_, _11786_, _11785_);
  and _62763_ (_11788_, _11787_, _06292_);
  and _62764_ (_11789_, _08768_, _07663_);
  or _62765_ (_11790_, _11789_, _11785_);
  and _62766_ (_11791_, _11790_, _06284_);
  and _62767_ (_11792_, _08549_, _07663_);
  or _62768_ (_11793_, _11792_, _11785_);
  or _62769_ (_11794_, _11793_, _06020_);
  and _62770_ (_11795_, _08498_, _07663_);
  or _62771_ (_11796_, _11795_, _11785_);
  or _62772_ (_11797_, _11796_, _06954_);
  and _62773_ (_11798_, _07663_, \oc8051_golden_model_1.ACC [7]);
  or _62774_ (_11799_, _11798_, _11785_);
  and _62775_ (_11800_, _11799_, _06938_);
  and _62776_ (_11801_, _06939_, \oc8051_golden_model_1.TH0 [7]);
  or _62777_ (_11802_, _11801_, _06102_);
  or _62778_ (_11803_, _11802_, _11800_);
  and _62779_ (_11804_, _11803_, _06848_);
  and _62780_ (_11805_, _11804_, _11797_);
  nor _62781_ (_11806_, _07785_, _11784_);
  or _62782_ (_11807_, _11806_, _11785_);
  and _62783_ (_11808_, _11807_, _06239_);
  or _62784_ (_11809_, _11808_, _11805_);
  and _62785_ (_11810_, _11809_, _06220_);
  and _62786_ (_11811_, _11799_, _06219_);
  or _62787_ (_11812_, _11811_, _09818_);
  or _62788_ (_11813_, _11812_, _11810_);
  and _62789_ (_11814_, _08485_, _07663_);
  or _62790_ (_11815_, _11785_, _07012_);
  or _62791_ (_11816_, _11815_, _11814_);
  or _62792_ (_11817_, _11807_, _09827_);
  and _62793_ (_11818_, _11817_, _05669_);
  and _62794_ (_11819_, _11818_, _11816_);
  and _62795_ (_11820_, _11819_, _11813_);
  and _62796_ (_11821_, _08738_, _07663_);
  or _62797_ (_11822_, _11821_, _11785_);
  and _62798_ (_11823_, _11822_, _09833_);
  or _62799_ (_11824_, _11823_, _06019_);
  or _62800_ (_11825_, _11824_, _11820_);
  and _62801_ (_11826_, _11825_, _11794_);
  or _62802_ (_11827_, _11826_, _06112_);
  and _62803_ (_11828_, _08760_, _07663_);
  or _62804_ (_11829_, _11785_, _08751_);
  or _62805_ (_11830_, _11829_, _11828_);
  and _62806_ (_11831_, _11830_, _08756_);
  and _62807_ (_11832_, _11831_, _11827_);
  or _62808_ (_11833_, _11832_, _11791_);
  and _62809_ (_11834_, _11833_, _07032_);
  or _62810_ (_11835_, _11785_, _07788_);
  and _62811_ (_11836_, _11793_, _06108_);
  and _62812_ (_11837_, _11836_, _11835_);
  or _62813_ (_11838_, _11837_, _11834_);
  and _62814_ (_11839_, _11838_, _06278_);
  and _62815_ (_11840_, _11799_, _06277_);
  and _62816_ (_11841_, _11840_, _11835_);
  or _62817_ (_11842_, _11841_, _06130_);
  or _62818_ (_11843_, _11842_, _11839_);
  and _62819_ (_11844_, _08759_, _07663_);
  or _62820_ (_11845_, _11785_, _08777_);
  or _62821_ (_11846_, _11845_, _11844_);
  and _62822_ (_11847_, _11846_, _08782_);
  and _62823_ (_11848_, _11847_, _11843_);
  or _62824_ (_11849_, _11848_, _11788_);
  and _62825_ (_11850_, _11849_, _06718_);
  and _62826_ (_11851_, _11796_, _06316_);
  or _62827_ (_11852_, _11851_, _06047_);
  or _62828_ (_11853_, _11852_, _11850_);
  and _62829_ (_11854_, _08279_, _07663_);
  or _62830_ (_11855_, _11785_, _06048_);
  or _62831_ (_11856_, _11855_, _11854_);
  and _62832_ (_11857_, _11856_, _01336_);
  and _62833_ (_11858_, _11857_, _11853_);
  or _62834_ (_11859_, _11858_, _11783_);
  and _62835_ (_40765_, _11859_, _42882_);
  not _62836_ (_11860_, _05331_);
  and _62837_ (_11861_, _08387_, _11860_);
  and _62838_ (_11862_, _11861_, \oc8051_golden_model_1.PC [7]);
  and _62839_ (_11863_, _11862_, _09201_);
  and _62840_ (_11864_, _11863_, \oc8051_golden_model_1.PC [10]);
  and _62841_ (_11865_, _11864_, \oc8051_golden_model_1.PC [11]);
  and _62842_ (_11866_, _11865_, \oc8051_golden_model_1.PC [12]);
  and _62843_ (_11867_, _11866_, \oc8051_golden_model_1.PC [13]);
  and _62844_ (_11868_, _11867_, \oc8051_golden_model_1.PC [14]);
  or _62845_ (_11869_, _11868_, \oc8051_golden_model_1.PC [15]);
  nand _62846_ (_11870_, _11868_, \oc8051_golden_model_1.PC [15]);
  and _62847_ (_11871_, _11870_, _11869_);
  and _62848_ (_11872_, _10934_, _10890_);
  or _62849_ (_11873_, _11872_, _11871_);
  nor _62850_ (_11874_, _09206_, \oc8051_golden_model_1.PC [14]);
  nor _62851_ (_11875_, _11874_, _09207_);
  and _62852_ (_11876_, _11875_, _05952_);
  nor _62853_ (_11877_, _11875_, _05952_);
  nor _62854_ (_11878_, _11877_, _11876_);
  nor _62855_ (_11879_, _09205_, \oc8051_golden_model_1.PC [13]);
  nor _62856_ (_11880_, _11879_, _09206_);
  and _62857_ (_11881_, _11880_, _05952_);
  nor _62858_ (_11882_, _11880_, _05952_);
  nor _62859_ (_11883_, _09204_, \oc8051_golden_model_1.PC [12]);
  nor _62860_ (_11884_, _11883_, _09205_);
  and _62861_ (_11885_, _11884_, _05952_);
  nor _62862_ (_11886_, _09209_, \oc8051_golden_model_1.PC [10]);
  nor _62863_ (_11887_, _11886_, _09210_);
  and _62864_ (_11888_, _11887_, _05952_);
  not _62865_ (_11889_, _11888_);
  nor _62866_ (_11890_, _09210_, \oc8051_golden_model_1.PC [11]);
  nor _62867_ (_11891_, _11890_, _09211_);
  and _62868_ (_11892_, _11891_, _05952_);
  nor _62869_ (_11893_, _11891_, _05952_);
  nor _62870_ (_11894_, _11893_, _11892_);
  nor _62871_ (_11895_, _11887_, _05952_);
  nor _62872_ (_11896_, _11895_, _11888_);
  and _62873_ (_11897_, _11896_, _11894_);
  and _62874_ (_11898_, _08389_, \oc8051_golden_model_1.PC [8]);
  nor _62875_ (_11899_, _11898_, \oc8051_golden_model_1.PC [9]);
  nor _62876_ (_11900_, _11899_, _09209_);
  and _62877_ (_11901_, _11900_, _05952_);
  nor _62878_ (_11902_, _11900_, _05952_);
  nor _62879_ (_11903_, _11902_, _11901_);
  and _62880_ (_11904_, _08391_, _05952_);
  nor _62881_ (_11905_, _08391_, _05952_);
  and _62882_ (_11906_, _08386_, _05850_);
  nor _62883_ (_11907_, _11906_, \oc8051_golden_model_1.PC [6]);
  nor _62884_ (_11908_, _11907_, _08388_);
  not _62885_ (_11909_, _11908_);
  nor _62886_ (_11910_, _11909_, _06084_);
  and _62887_ (_11911_, _11909_, _06084_);
  nor _62888_ (_11912_, _11911_, _11910_);
  not _62889_ (_11913_, _11912_);
  and _62890_ (_11914_, _05850_, \oc8051_golden_model_1.PC [4]);
  nor _62891_ (_11915_, _11914_, \oc8051_golden_model_1.PC [5]);
  nor _62892_ (_11916_, _11915_, _11906_);
  not _62893_ (_11917_, _11916_);
  nor _62894_ (_11918_, _11917_, _06359_);
  and _62895_ (_11919_, _11917_, _06359_);
  nor _62896_ (_11920_, _05850_, \oc8051_golden_model_1.PC [4]);
  nor _62897_ (_11921_, _11920_, _11914_);
  not _62898_ (_11922_, _11921_);
  nor _62899_ (_11923_, _11922_, _06758_);
  nor _62900_ (_11924_, _05983_, _06148_);
  and _62901_ (_11925_, _05983_, _06148_);
  nor _62902_ (_11926_, _06403_, _05804_);
  nor _62903_ (_11927_, _06799_, \oc8051_golden_model_1.PC [1]);
  nor _62904_ (_11928_, _06016_, _05346_);
  and _62905_ (_11929_, _06799_, \oc8051_golden_model_1.PC [1]);
  nor _62906_ (_11930_, _11929_, _11927_);
  and _62907_ (_11931_, _11930_, _11928_);
  nor _62908_ (_11932_, _11931_, _11927_);
  and _62909_ (_11933_, _06403_, _05804_);
  nor _62910_ (_11934_, _11933_, _11926_);
  not _62911_ (_11935_, _11934_);
  nor _62912_ (_11936_, _11935_, _11932_);
  nor _62913_ (_11937_, _11936_, _11926_);
  nor _62914_ (_11938_, _11937_, _11925_);
  nor _62915_ (_11939_, _11938_, _11924_);
  and _62916_ (_11940_, _11922_, _06758_);
  nor _62917_ (_11941_, _11940_, _11923_);
  not _62918_ (_11942_, _11941_);
  nor _62919_ (_11943_, _11942_, _11939_);
  nor _62920_ (_11944_, _11943_, _11923_);
  nor _62921_ (_11945_, _11944_, _11919_);
  nor _62922_ (_11946_, _11945_, _11918_);
  nor _62923_ (_11947_, _11946_, _11913_);
  nor _62924_ (_11948_, _11947_, _11910_);
  nor _62925_ (_11949_, _11948_, _11905_);
  or _62926_ (_11950_, _11949_, _11904_);
  nor _62927_ (_11951_, _08389_, \oc8051_golden_model_1.PC [8]);
  nor _62928_ (_11952_, _11951_, _11898_);
  and _62929_ (_11953_, _11952_, _05952_);
  nor _62930_ (_11954_, _11952_, _05952_);
  nor _62931_ (_11955_, _11954_, _11953_);
  and _62932_ (_11956_, _11955_, _11950_);
  and _62933_ (_11957_, _11956_, _11903_);
  and _62934_ (_11958_, _11957_, _11897_);
  nor _62935_ (_11959_, _11953_, _11901_);
  not _62936_ (_11960_, _11959_);
  and _62937_ (_11961_, _11960_, _11897_);
  or _62938_ (_11962_, _11961_, _11892_);
  nor _62939_ (_11963_, _11962_, _11958_);
  and _62940_ (_11964_, _11963_, _11889_);
  nor _62941_ (_11965_, _11884_, _05952_);
  nor _62942_ (_11966_, _11965_, _11885_);
  not _62943_ (_11967_, _11966_);
  nor _62944_ (_11968_, _11967_, _11964_);
  nor _62945_ (_11969_, _11968_, _11885_);
  nor _62946_ (_11970_, _11969_, _11882_);
  nor _62947_ (_11971_, _11970_, _11881_);
  not _62948_ (_11972_, _11971_);
  and _62949_ (_11973_, _11972_, _11878_);
  nor _62950_ (_11974_, _11973_, _11876_);
  nor _62951_ (_11975_, _09216_, _05952_);
  and _62952_ (_11976_, _09216_, _05952_);
  nor _62953_ (_11977_, _11976_, _11975_);
  and _62954_ (_11978_, _11977_, _11974_);
  nor _62955_ (_11979_, _11977_, _11974_);
  or _62956_ (_11980_, _11979_, _11978_);
  or _62957_ (_11981_, _11980_, _10606_);
  and _62958_ (_11982_, _05739_, _05650_);
  or _62959_ (_11983_, _09216_, \oc8051_golden_model_1.PSW [7]);
  and _62960_ (_11984_, _11983_, _11982_);
  and _62961_ (_11985_, _11984_, _11981_);
  nor _62962_ (_11986_, _10781_, _06290_);
  not _62963_ (_11987_, _11986_);
  or _62964_ (_11988_, _06093_, _06135_);
  and _62965_ (_11989_, _11988_, _05739_);
  not _62966_ (_11990_, _11989_);
  and _62967_ (_11991_, _07002_, _05739_);
  nor _62968_ (_11992_, _10775_, _11991_);
  and _62969_ (_11993_, _11992_, _11990_);
  or _62970_ (_11994_, _11993_, _11871_);
  nor _62971_ (_11995_, _06093_, _06229_);
  nor _62972_ (_11996_, _11995_, _06656_);
  not _62973_ (_11997_, _11996_);
  and _62974_ (_11998_, _06227_, _05735_);
  and _62975_ (_11999_, _07002_, _05735_);
  or _62976_ (_12000_, _11999_, _10731_);
  nor _62977_ (_12001_, _12000_, _11998_);
  and _62978_ (_12002_, _12001_, _11997_);
  or _62979_ (_12003_, _12002_, _11871_);
  not _62980_ (_12004_, _07248_);
  nor _62981_ (_12005_, _11988_, _12004_);
  nor _62982_ (_12006_, _12005_, _06644_);
  not _62983_ (_12007_, _12006_);
  or _62984_ (_12008_, _12007_, _11871_);
  or _62985_ (_12009_, _09216_, _08742_);
  not _62986_ (_12010_, _09227_);
  nor _62987_ (_12011_, _12010_, _05669_);
  nor _62988_ (_12012_, _05685_, _05662_);
  not _62989_ (_12013_, _12012_);
  and _62990_ (_12014_, _09202_, _09139_);
  and _62991_ (_12015_, _12014_, \oc8051_golden_model_1.PC [11]);
  and _62992_ (_12016_, _12015_, \oc8051_golden_model_1.PC [12]);
  and _62993_ (_12017_, _12016_, \oc8051_golden_model_1.PC [13]);
  and _62994_ (_12018_, _12017_, \oc8051_golden_model_1.PC [14]);
  nor _62995_ (_12019_, _12017_, \oc8051_golden_model_1.PC [14]);
  nor _62996_ (_12020_, _12019_, _12018_);
  not _62997_ (_12021_, _12020_);
  nor _62998_ (_12022_, _12021_, _08332_);
  and _62999_ (_12023_, _12021_, _08332_);
  nor _63000_ (_12024_, _12023_, _12022_);
  not _63001_ (_12025_, _12024_);
  nor _63002_ (_12026_, _12016_, \oc8051_golden_model_1.PC [13]);
  nor _63003_ (_12027_, _12026_, _12017_);
  not _63004_ (_12028_, _12027_);
  nor _63005_ (_12029_, _12028_, _08332_);
  and _63006_ (_12030_, _12028_, _08332_);
  nor _63007_ (_12031_, _12015_, \oc8051_golden_model_1.PC [12]);
  nor _63008_ (_12032_, _12031_, _12016_);
  not _63009_ (_12033_, _12032_);
  nor _63010_ (_12034_, _12033_, _08332_);
  nor _63011_ (_12035_, _12014_, \oc8051_golden_model_1.PC [11]);
  nor _63012_ (_12036_, _12035_, _12015_);
  not _63013_ (_12037_, _12036_);
  nor _63014_ (_12038_, _12037_, _08332_);
  and _63015_ (_12039_, _12037_, _08332_);
  nor _63016_ (_12040_, _12039_, _12038_);
  and _63017_ (_12041_, _09201_, _09139_);
  nor _63018_ (_12042_, _12041_, \oc8051_golden_model_1.PC [10]);
  nor _63019_ (_12043_, _12042_, _12014_);
  not _63020_ (_12044_, _12043_);
  nor _63021_ (_12045_, _12044_, _08332_);
  and _63022_ (_12046_, _12044_, _08332_);
  nor _63023_ (_12047_, _12046_, _12045_);
  and _63024_ (_12048_, _12047_, _12040_);
  and _63025_ (_12049_, _09139_, \oc8051_golden_model_1.PC [8]);
  nor _63026_ (_12050_, _12049_, \oc8051_golden_model_1.PC [9]);
  nor _63027_ (_12051_, _12050_, _12041_);
  not _63028_ (_12052_, _12051_);
  nor _63029_ (_12053_, _12052_, _08332_);
  and _63030_ (_12054_, _12052_, _08332_);
  nor _63031_ (_12055_, _12054_, _12053_);
  nor _63032_ (_12056_, _09142_, _08332_);
  and _63033_ (_12057_, _09142_, _08332_);
  nor _63034_ (_12058_, _12057_, _12056_);
  not _63035_ (_12059_, _12058_);
  and _63036_ (_12060_, _09137_, _08386_);
  nor _63037_ (_12061_, _12060_, \oc8051_golden_model_1.PC [6]);
  nor _63038_ (_12062_, _12061_, _09138_);
  not _63039_ (_12063_, _12062_);
  nor _63040_ (_12064_, _12063_, _08647_);
  and _63041_ (_12065_, _12063_, _08647_);
  nor _63042_ (_12066_, _12065_, _12064_);
  and _63043_ (_12067_, _09137_, \oc8051_golden_model_1.PC [4]);
  nor _63044_ (_12068_, _12067_, \oc8051_golden_model_1.PC [5]);
  nor _63045_ (_12069_, _12068_, _12060_);
  not _63046_ (_12070_, _12069_);
  nor _63047_ (_12071_, _12070_, _08612_);
  and _63048_ (_12072_, _12070_, _08612_);
  nor _63049_ (_12073_, _09137_, \oc8051_golden_model_1.PC [4]);
  nor _63050_ (_12074_, _12073_, _12067_);
  not _63051_ (_12075_, _12074_);
  nor _63052_ (_12076_, _12075_, _08581_);
  nor _63053_ (_12077_, _09136_, \oc8051_golden_model_1.PC [3]);
  nor _63054_ (_12078_, _12077_, _09137_);
  not _63055_ (_12079_, _12078_);
  nor _63056_ (_12080_, _12079_, _06215_);
  and _63057_ (_12081_, _12079_, _06215_);
  nor _63058_ (_12082_, _05350_, \oc8051_golden_model_1.PC [2]);
  nor _63059_ (_12083_, _12082_, _09136_);
  not _63060_ (_12084_, _12083_);
  nor _63061_ (_12085_, _12084_, _06445_);
  not _63062_ (_12086_, _05777_);
  nor _63063_ (_12087_, _06832_, _12086_);
  nor _63064_ (_12088_, _06633_, \oc8051_golden_model_1.PC [0]);
  and _63065_ (_12089_, _06832_, _12086_);
  nor _63066_ (_12090_, _12089_, _12087_);
  and _63067_ (_12091_, _12090_, _12088_);
  nor _63068_ (_12092_, _12091_, _12087_);
  and _63069_ (_12093_, _12084_, _06445_);
  nor _63070_ (_12094_, _12093_, _12085_);
  not _63071_ (_12095_, _12094_);
  nor _63072_ (_12096_, _12095_, _12092_);
  nor _63073_ (_12097_, _12096_, _12085_);
  nor _63074_ (_12098_, _12097_, _12081_);
  nor _63075_ (_12099_, _12098_, _12080_);
  and _63076_ (_12100_, _12075_, _08581_);
  nor _63077_ (_12101_, _12100_, _12076_);
  not _63078_ (_12102_, _12101_);
  nor _63079_ (_12103_, _12102_, _12099_);
  nor _63080_ (_12104_, _12103_, _12076_);
  nor _63081_ (_12105_, _12104_, _12072_);
  or _63082_ (_12106_, _12105_, _12071_);
  and _63083_ (_12107_, _12106_, _12066_);
  nor _63084_ (_12108_, _12107_, _12064_);
  nor _63085_ (_12109_, _12108_, _12059_);
  nor _63086_ (_12110_, _12109_, _12056_);
  nor _63087_ (_12111_, _09139_, \oc8051_golden_model_1.PC [8]);
  nor _63088_ (_12112_, _12111_, _12049_);
  not _63089_ (_12113_, _12112_);
  nor _63090_ (_12114_, _12113_, _08332_);
  and _63091_ (_12115_, _12113_, _08332_);
  nor _63092_ (_12116_, _12115_, _12114_);
  not _63093_ (_12117_, _12116_);
  nor _63094_ (_12118_, _12117_, _12110_);
  and _63095_ (_12119_, _12118_, _12055_);
  and _63096_ (_12120_, _12119_, _12048_);
  nor _63097_ (_12121_, _12114_, _12053_);
  not _63098_ (_12122_, _12121_);
  and _63099_ (_12123_, _12122_, _12048_);
  or _63100_ (_12124_, _12123_, _12045_);
  or _63101_ (_12125_, _12124_, _12120_);
  nor _63102_ (_12126_, _12125_, _12038_);
  and _63103_ (_12127_, _12033_, _08332_);
  nor _63104_ (_12128_, _12127_, _12034_);
  not _63105_ (_12129_, _12128_);
  nor _63106_ (_12130_, _12129_, _12126_);
  nor _63107_ (_12131_, _12130_, _12034_);
  nor _63108_ (_12132_, _12131_, _12030_);
  nor _63109_ (_12133_, _12132_, _12029_);
  nor _63110_ (_12134_, _12133_, _12025_);
  nor _63111_ (_12135_, _12134_, _12022_);
  and _63112_ (_12136_, _12010_, _08332_);
  nor _63113_ (_12137_, _12010_, _08332_);
  nor _63114_ (_12138_, _12137_, _12136_);
  and _63115_ (_12139_, _12138_, _12135_);
  nor _63116_ (_12140_, _12138_, _12135_);
  or _63117_ (_12141_, _12140_, _12139_);
  or _63118_ (_12142_, _09181_, _05983_);
  or _63119_ (_12143_, _08985_, _06299_);
  and _63120_ (_12144_, _12143_, _12142_);
  or _63121_ (_12145_, _09182_, _06403_);
  or _63122_ (_12146_, _09030_, _07477_);
  and _63123_ (_12147_, _12146_, _12145_);
  and _63124_ (_12148_, _12147_, _12144_);
  nand _63125_ (_12149_, _09120_, _06016_);
  nand _63126_ (_12150_, _09074_, _09052_);
  or _63127_ (_12151_, _12150_, _07076_);
  or _63128_ (_12152_, _09075_, _06799_);
  and _63129_ (_12153_, _12152_, _12151_);
  and _63130_ (_12154_, _12153_, _12149_);
  and _63131_ (_12155_, _12154_, _12148_);
  or _63132_ (_12156_, _09120_, _06016_);
  and _63133_ (_12157_, _08798_, _05952_);
  nor _63134_ (_12158_, _12157_, _08531_);
  or _63135_ (_12159_, _09178_, _06084_);
  or _63136_ (_12160_, _08843_, _07414_);
  and _63137_ (_12161_, _12160_, _12159_);
  and _63138_ (_12162_, _12161_, _12158_);
  or _63139_ (_12163_, _09179_, _06359_);
  or _63140_ (_12164_, _08888_, _07683_);
  and _63141_ (_12165_, _12164_, _12163_);
  or _63142_ (_12166_, _09180_, _06758_);
  or _63143_ (_12167_, _08937_, _07674_);
  and _63144_ (_12168_, _12167_, _12166_);
  and _63145_ (_12169_, _12168_, _12165_);
  and _63146_ (_12170_, _12169_, _12162_);
  and _63147_ (_12171_, _12170_, _12156_);
  and _63148_ (_12172_, _12171_, _12155_);
  or _63149_ (_12173_, _12172_, _12141_);
  nand _63150_ (_12174_, _12171_, _12155_);
  or _63151_ (_12175_, _12174_, _09227_);
  and _63152_ (_12176_, _12175_, _06104_);
  and _63153_ (_12177_, _12176_, _12173_);
  and _63154_ (_12178_, _09216_, _06219_);
  and _63155_ (_12179_, _06244_, _05690_);
  or _63156_ (_12180_, _12179_, _09216_);
  nor _63157_ (_12181_, _05689_, _05662_);
  nor _63158_ (_12182_, _12181_, _10412_);
  and _63159_ (_12183_, _07885_, _07787_);
  and _63160_ (_12184_, _12183_, _08489_);
  and _63161_ (_12185_, _08127_, _08077_);
  and _63162_ (_12186_, _08492_, _12185_);
  nand _63163_ (_12187_, _12186_, _12184_);
  or _63164_ (_12188_, _12187_, _09227_);
  and _63165_ (_12189_, _12186_, _12184_);
  or _63166_ (_12190_, _12189_, _12141_);
  and _63167_ (_12191_, _12190_, _06102_);
  and _63168_ (_12192_, _12191_, _12188_);
  and _63169_ (_12193_, _07132_, _06931_);
  and _63170_ (_12194_, _07883_, _07785_);
  and _63171_ (_12195_, _12194_, _12193_);
  and _63172_ (_12196_, _08290_, _08289_);
  and _63173_ (_12197_, _12196_, _12195_);
  and _63174_ (_12198_, _12197_, _09216_);
  nand _63175_ (_12199_, _12196_, _12195_);
  and _63176_ (_12200_, _12199_, _11980_);
  or _63177_ (_12201_, _12200_, _08383_);
  or _63178_ (_12202_, _12201_, _12198_);
  nor _63179_ (_12203_, _06933_, _05697_);
  not _63180_ (_12204_, _12203_);
  and _63181_ (_12205_, _12204_, _10400_);
  nor _63182_ (_12206_, _06938_, _06943_);
  or _63183_ (_12207_, _12206_, _09216_);
  or _63184_ (_12208_, _06530_, _06943_);
  or _63185_ (_12209_, _06938_, \oc8051_golden_model_1.PC [15]);
  or _63186_ (_12210_, _12209_, _12208_);
  or _63187_ (_12211_, _12210_, _07250_);
  nand _63188_ (_12212_, _12211_, _12207_);
  nand _63189_ (_12213_, _12212_, _12205_);
  nor _63190_ (_12214_, _07250_, _06530_);
  and _63191_ (_12215_, _12214_, _12205_);
  or _63192_ (_12216_, _12215_, _11871_);
  and _63193_ (_12217_, _12216_, _12213_);
  or _63194_ (_12218_, _12217_, _08384_);
  nor _63195_ (_12219_, _06948_, _06102_);
  and _63196_ (_12220_, _12219_, _12218_);
  and _63197_ (_12221_, _12220_, _12202_);
  or _63198_ (_12222_, _12221_, _12192_);
  and _63199_ (_12223_, _12222_, _12182_);
  not _63200_ (_12224_, _12179_);
  and _63201_ (_12225_, _12182_, _06949_);
  not _63202_ (_12226_, _12225_);
  and _63203_ (_12227_, _12226_, _11871_);
  or _63204_ (_12228_, _12227_, _12224_);
  or _63205_ (_12229_, _12228_, _12223_);
  and _63206_ (_12230_, _12229_, _12180_);
  nor _63207_ (_12231_, _10378_, _06970_);
  not _63208_ (_12232_, _12231_);
  or _63209_ (_12233_, _12232_, _12230_);
  or _63210_ (_12234_, _12231_, _11871_);
  and _63211_ (_12235_, _12234_, _06220_);
  and _63212_ (_12236_, _12235_, _12233_);
  or _63213_ (_12237_, _12236_, _12178_);
  nor _63214_ (_12238_, _05693_, _05662_);
  nor _63215_ (_12239_, _12238_, _10376_);
  and _63216_ (_12240_, _12239_, _12237_);
  not _63217_ (_12241_, _12239_);
  and _63218_ (_12242_, _12241_, _11871_);
  not _63219_ (_12243_, _05694_);
  nor _63220_ (_12244_, _06038_, _12243_);
  and _63221_ (_12245_, _12244_, _06040_);
  not _63222_ (_12246_, _12245_);
  or _63223_ (_12247_, _12246_, _12242_);
  or _63224_ (_12248_, _12247_, _12240_);
  or _63225_ (_12249_, _12245_, _09216_);
  and _63226_ (_12250_, _12249_, _12248_);
  not _63227_ (_12251_, _06138_);
  and _63228_ (_12252_, _07002_, _06031_);
  and _63229_ (_12253_, _07005_, _06031_);
  nor _63230_ (_12254_, _12253_, _12252_);
  and _63231_ (_12255_, _12254_, _12251_);
  not _63232_ (_12256_, _12255_);
  or _63233_ (_12257_, _12256_, _12250_);
  not _63234_ (_12258_, _06104_);
  not _63235_ (_12259_, _07786_);
  and _63236_ (_12260_, _07785_, _05952_);
  nor _63237_ (_12261_, _12260_, _12259_);
  nor _63238_ (_12262_, _07883_, _07414_);
  and _63239_ (_12263_, _07883_, _07414_);
  nor _63240_ (_12264_, _12263_, _12262_);
  and _63241_ (_12265_, _12264_, _12261_);
  nor _63242_ (_12266_, _07977_, _07683_);
  and _63243_ (_12267_, _07977_, _07683_);
  nor _63244_ (_12268_, _12267_, _12266_);
  and _63245_ (_12269_, _08270_, _07674_);
  nor _63246_ (_12270_, _08270_, _07674_);
  nor _63247_ (_12271_, _12270_, _12269_);
  and _63248_ (_12272_, _12271_, _12268_);
  and _63249_ (_12273_, _12272_, _12265_);
  and _63250_ (_12274_, _07353_, _06299_);
  nor _63251_ (_12275_, _07353_, _06299_);
  nor _63252_ (_12276_, _12275_, _12274_);
  and _63253_ (_12277_, _07530_, _07477_);
  nor _63254_ (_12278_, _07530_, _07477_);
  nor _63255_ (_12279_, _12278_, _12277_);
  and _63256_ (_12280_, _12279_, _12276_);
  nor _63257_ (_12281_, _07132_, _07076_);
  and _63258_ (_12282_, _07132_, _07076_);
  nor _63259_ (_12283_, _12282_, _12281_);
  and _63260_ (_12284_, _06931_, _06016_);
  nor _63261_ (_12285_, _06931_, _06016_);
  nor _63262_ (_12286_, _12285_, _12284_);
  and _63263_ (_12287_, _12286_, _12283_);
  and _63264_ (_12288_, _12287_, _12280_);
  and _63265_ (_12289_, _12288_, _12273_);
  or _63266_ (_12290_, _12289_, _12141_);
  nand _63267_ (_12291_, _12289_, _12010_);
  and _63268_ (_12292_, _12291_, _12290_);
  or _63269_ (_12293_, _12292_, _12255_);
  and _63270_ (_12294_, _12293_, _12258_);
  and _63271_ (_12295_, _12294_, _12257_);
  or _63272_ (_12296_, _12295_, _06121_);
  or _63273_ (_12297_, _12296_, _12177_);
  not _63274_ (_12298_, _06115_);
  nor _63275_ (_12299_, _10988_, _10987_);
  nor _63276_ (_12300_, _12299_, _10991_);
  not _63277_ (_12301_, _10994_);
  nor _63278_ (_12302_, _08127_, \oc8051_golden_model_1.ACC [0]);
  or _63279_ (_12303_, _12302_, _10995_);
  and _63280_ (_12304_, _12303_, _12301_);
  and _63281_ (_12305_, _12304_, _12300_);
  nor _63282_ (_12306_, _10981_, _10982_);
  nor _63283_ (_12307_, _12306_, _10986_);
  nor _63284_ (_12308_, _10980_, _08768_);
  and _63285_ (_12309_, _12308_, _12307_);
  and _63286_ (_12310_, _12309_, _12305_);
  and _63287_ (_12311_, _12310_, _09227_);
  not _63288_ (_12312_, _12310_);
  and _63289_ (_12313_, _12312_, _12141_);
  or _63290_ (_12314_, _12313_, _06509_);
  or _63291_ (_12315_, _12314_, _12311_);
  and _63292_ (_12316_, _12315_, _12298_);
  and _63293_ (_12317_, _12316_, _12297_);
  not _63294_ (_12318_, _11032_);
  nor _63295_ (_12319_, _11028_, _11029_);
  nor _63296_ (_12320_, _12319_, _12318_);
  and _63297_ (_12321_, _06016_, _05758_);
  nor _63298_ (_12322_, _12321_, _11036_);
  nor _63299_ (_12323_, _12322_, _11035_);
  and _63300_ (_12324_, _12323_, _12320_);
  nor _63301_ (_12325_, _11021_, _11022_);
  nor _63302_ (_12326_, _12325_, _11027_);
  nor _63303_ (_12327_, _11020_, _10705_);
  and _63304_ (_12328_, _12327_, _12326_);
  and _63305_ (_12329_, _12328_, _12324_);
  or _63306_ (_12330_, _12329_, _12141_);
  nand _63307_ (_12331_, _12329_, _12010_);
  and _63308_ (_12332_, _12331_, _06115_);
  and _63309_ (_12333_, _12332_, _12330_);
  or _63310_ (_12334_, _12333_, _12317_);
  and _63311_ (_12335_, _12334_, _12013_);
  nand _63312_ (_12336_, _12012_, _11871_);
  nor _63313_ (_12337_, _06032_, _07355_);
  and _63314_ (_12338_, _06222_, _05609_);
  nor _63315_ (_12339_, _12338_, _06253_);
  and _63316_ (_12340_, _12339_, _06231_);
  and _63317_ (_12341_, _06460_, _06221_);
  nor _63318_ (_12342_, _07248_, _05701_);
  nor _63319_ (_12343_, _12342_, _12341_);
  and _63320_ (_12344_, _12343_, _12340_);
  and _63321_ (_12345_, _12344_, _12337_);
  nand _63322_ (_12346_, _12345_, _12336_);
  or _63323_ (_12347_, _12346_, _12335_);
  nor _63324_ (_12348_, _05701_, _05668_);
  not _63325_ (_12349_, _12348_);
  nor _63326_ (_12350_, _11290_, _09269_);
  and _63327_ (_12351_, _12350_, _12349_);
  or _63328_ (_12352_, _12345_, _09216_);
  and _63329_ (_12353_, _12352_, _12351_);
  and _63330_ (_12354_, _12353_, _12347_);
  not _63331_ (_12355_, _12351_);
  and _63332_ (_12356_, _12355_, _11871_);
  and _63333_ (_12357_, _06252_, _05702_);
  not _63334_ (_12358_, _12357_);
  or _63335_ (_12359_, _12358_, _12356_);
  or _63336_ (_12360_, _12359_, _12354_);
  and _63337_ (_12361_, _06103_, _05671_);
  nor _63338_ (_12362_, _10468_, _12361_);
  or _63339_ (_12363_, _12357_, _09216_);
  and _63340_ (_12364_, _12363_, _12362_);
  and _63341_ (_12365_, _12364_, _12360_);
  nor _63342_ (_12366_, _10306_, _06261_);
  not _63343_ (_12367_, _12366_);
  not _63344_ (_12368_, _12362_);
  and _63345_ (_12369_, _12368_, _11871_);
  or _63346_ (_12370_, _12369_, _12367_);
  or _63347_ (_12371_, _12370_, _12365_);
  or _63348_ (_12372_, _12366_, _09216_);
  and _63349_ (_12373_, _12372_, _05675_);
  and _63350_ (_12374_, _12373_, _12371_);
  nand _63351_ (_12375_, _11871_, _05676_);
  nor _63352_ (_12376_, _06026_, _06023_);
  nand _63353_ (_12377_, _12376_, _12375_);
  or _63354_ (_12378_, _12377_, _12374_);
  or _63355_ (_12379_, _12376_, _09216_);
  and _63356_ (_12380_, _12379_, _06111_);
  and _63357_ (_12381_, _12380_, _12378_);
  nand _63358_ (_12382_, _09227_, _06110_);
  nand _63359_ (_12383_, _12382_, _09817_);
  or _63360_ (_12384_, _12383_, _12381_);
  or _63361_ (_12385_, _09817_, _09216_);
  and _63362_ (_12386_, _12385_, _05669_);
  and _63363_ (_12387_, _12386_, _12384_);
  or _63364_ (_12388_, _12387_, _12011_);
  nor _63365_ (_12389_, _09832_, _05663_);
  and _63366_ (_12390_, _12389_, _12388_);
  nor _63367_ (_12391_, _06089_, _05719_);
  not _63368_ (_12392_, _12391_);
  not _63369_ (_12393_, _12389_);
  and _63370_ (_12394_, _12393_, _11871_);
  or _63371_ (_12395_, _12394_, _12392_);
  or _63372_ (_12396_, _12395_, _12390_);
  and _63373_ (_12397_, _05659_, _05650_);
  not _63374_ (_12398_, _12397_);
  or _63375_ (_12399_, _12391_, _09216_);
  and _63376_ (_12400_, _12399_, _12398_);
  and _63377_ (_12401_, _12400_, _12396_);
  and _63378_ (_12402_, _12397_, _11980_);
  or _63379_ (_12403_, _12402_, _08743_);
  or _63380_ (_12404_, _12403_, _12401_);
  and _63381_ (_12405_, _12404_, _12009_);
  or _63382_ (_12406_, _12405_, _06019_);
  nand _63383_ (_12407_, _12010_, _06019_);
  and _63384_ (_12408_, _12407_, _10662_);
  and _63385_ (_12409_, _12408_, _12406_);
  and _63386_ (_12410_, _10661_, _09216_);
  or _63387_ (_12411_, _12410_, _12409_);
  and _63388_ (_12412_, _05723_, _06107_);
  not _63389_ (_12413_, _12412_);
  and _63390_ (_12414_, _12413_, _12411_);
  nor _63391_ (_12415_, _06088_, _05724_);
  not _63392_ (_12416_, _12415_);
  and _63393_ (_12417_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  nor _63394_ (_12418_, \oc8051_golden_model_1.DPL [7], \oc8051_golden_model_1.ACC [7]);
  and _63395_ (_12419_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _63396_ (_12420_, \oc8051_golden_model_1.DPL [6], \oc8051_golden_model_1.ACC [6]);
  nor _63397_ (_12421_, _12420_, _12419_);
  not _63398_ (_12422_, _12421_);
  and _63399_ (_12423_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _63400_ (_12424_, \oc8051_golden_model_1.DPL [5], \oc8051_golden_model_1.ACC [5]);
  nor _63401_ (_12425_, _12424_, _12423_);
  not _63402_ (_12426_, _12425_);
  and _63403_ (_12427_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _63404_ (_12428_, _05862_, _05857_);
  nor _63405_ (_12429_, \oc8051_golden_model_1.DPL [4], \oc8051_golden_model_1.ACC [4]);
  nor _63406_ (_12430_, _12429_, _12427_);
  not _63407_ (_12431_, _12430_);
  nor _63408_ (_12432_, _12431_, _12428_);
  nor _63409_ (_12433_, _12432_, _12427_);
  nor _63410_ (_12434_, _12433_, _12426_);
  nor _63411_ (_12435_, _12434_, _12423_);
  nor _63412_ (_12436_, _12435_, _12422_);
  nor _63413_ (_12437_, _12436_, _12419_);
  nor _63414_ (_12438_, _12437_, _12418_);
  or _63415_ (_12439_, _12438_, _12417_);
  and _63416_ (_12440_, _12439_, \oc8051_golden_model_1.DPH [0]);
  and _63417_ (_12441_, _12440_, \oc8051_golden_model_1.DPH [1]);
  and _63418_ (_12442_, _12441_, \oc8051_golden_model_1.DPH [2]);
  and _63419_ (_12443_, _12442_, \oc8051_golden_model_1.DPH [3]);
  and _63420_ (_12444_, _12443_, \oc8051_golden_model_1.DPH [4]);
  and _63421_ (_12445_, _12444_, \oc8051_golden_model_1.DPH [5]);
  and _63422_ (_12446_, _12445_, \oc8051_golden_model_1.DPH [6]);
  nand _63423_ (_12447_, _12446_, \oc8051_golden_model_1.DPH [7]);
  or _63424_ (_12448_, _12446_, \oc8051_golden_model_1.DPH [7]);
  and _63425_ (_12449_, _12448_, _12412_);
  and _63426_ (_12450_, _12449_, _12447_);
  or _63427_ (_12451_, _12450_, _12416_);
  or _63428_ (_12452_, _12451_, _12414_);
  and _63429_ (_12453_, _05723_, _05650_);
  not _63430_ (_12454_, _12453_);
  or _63431_ (_12455_, _12415_, _09216_);
  and _63432_ (_12456_, _12455_, _12454_);
  and _63433_ (_12457_, _12456_, _12452_);
  or _63434_ (_12458_, _11980_, _11071_);
  not _63435_ (_12459_, _11071_);
  or _63436_ (_12460_, _12459_, _09216_);
  and _63437_ (_12461_, _12460_, _12453_);
  and _63438_ (_12462_, _12461_, _12458_);
  or _63439_ (_12463_, _12462_, _12006_);
  or _63440_ (_12464_, _12463_, _12457_);
  and _63441_ (_12465_, _12464_, _12008_);
  nor _63442_ (_12466_, _10698_, _06282_);
  not _63443_ (_12467_, _12466_);
  or _63444_ (_12468_, _12467_, _12465_);
  or _63445_ (_12469_, _12466_, _09216_);
  and _63446_ (_12470_, _12469_, _08751_);
  and _63447_ (_12471_, _12470_, _12468_);
  nand _63448_ (_12472_, _09227_, _06112_);
  nor _63449_ (_12473_, _06284_, _05727_);
  nand _63450_ (_12474_, _12473_, _12472_);
  or _63451_ (_12475_, _12474_, _12471_);
  and _63452_ (_12476_, _05726_, _05650_);
  not _63453_ (_12477_, _12476_);
  or _63454_ (_12478_, _12473_, _09216_);
  and _63455_ (_12479_, _12478_, _12477_);
  and _63456_ (_12480_, _12479_, _12475_);
  not _63457_ (_12481_, _12002_);
  or _63458_ (_12482_, _11980_, _12459_);
  or _63459_ (_12483_, _11071_, _09216_);
  and _63460_ (_12484_, _12483_, _12476_);
  and _63461_ (_12485_, _12484_, _12482_);
  or _63462_ (_12486_, _12485_, _12481_);
  or _63463_ (_12487_, _12486_, _12480_);
  and _63464_ (_12488_, _12487_, _12003_);
  or _63465_ (_12489_, _12488_, _10743_);
  or _63466_ (_12490_, _10742_, _09216_);
  and _63467_ (_12491_, _12490_, _07032_);
  and _63468_ (_12492_, _12491_, _12489_);
  nand _63469_ (_12493_, _09227_, _06108_);
  nor _63470_ (_12494_, _06277_, _05736_);
  nand _63471_ (_12495_, _12494_, _12493_);
  or _63472_ (_12496_, _12495_, _12492_);
  and _63473_ (_12497_, _05735_, _05650_);
  not _63474_ (_12498_, _12497_);
  or _63475_ (_12499_, _12494_, _09216_);
  and _63476_ (_12500_, _12499_, _12498_);
  and _63477_ (_12501_, _12500_, _12496_);
  not _63478_ (_12502_, _11993_);
  or _63479_ (_12503_, _11980_, \oc8051_golden_model_1.PSW [7]);
  or _63480_ (_12504_, _09216_, _10606_);
  and _63481_ (_12505_, _12504_, _12497_);
  and _63482_ (_12506_, _12505_, _12503_);
  or _63483_ (_12507_, _12506_, _12502_);
  or _63484_ (_12508_, _12507_, _12501_);
  and _63485_ (_12509_, _12508_, _11994_);
  or _63486_ (_12510_, _12509_, _11987_);
  or _63487_ (_12511_, _11986_, _09216_);
  and _63488_ (_12512_, _12511_, _08777_);
  and _63489_ (_12513_, _12512_, _12510_);
  nand _63490_ (_12514_, _09227_, _06130_);
  nor _63491_ (_12515_, _06292_, _05740_);
  nand _63492_ (_12516_, _12515_, _12514_);
  or _63493_ (_12517_, _12516_, _12513_);
  not _63494_ (_12518_, _11982_);
  or _63495_ (_12519_, _12515_, _09216_);
  and _63496_ (_12520_, _12519_, _12518_);
  and _63497_ (_12521_, _12520_, _12517_);
  or _63498_ (_12522_, _12521_, _11985_);
  nor _63499_ (_12523_, _10794_, _10303_);
  and _63500_ (_12524_, _12523_, _12522_);
  not _63501_ (_12525_, _12523_);
  and _63502_ (_12526_, _12525_, _11871_);
  or _63503_ (_12527_, _12526_, _10826_);
  or _63504_ (_12528_, _12527_, _12524_);
  or _63505_ (_12529_, _10825_, _09216_);
  and _63506_ (_12530_, _12529_, _10855_);
  and _63507_ (_12531_, _12530_, _12528_);
  and _63508_ (_12532_, _11871_, _10854_);
  or _63509_ (_12533_, _12532_, _06298_);
  or _63510_ (_12534_, _12533_, _12531_);
  nand _63511_ (_12535_, _07785_, _06298_);
  and _63512_ (_12536_, _12535_, _12534_);
  or _63513_ (_12537_, _12536_, _05732_);
  or _63514_ (_12538_, _09216_, _05734_);
  and _63515_ (_12539_, _12538_, _06306_);
  and _63516_ (_12540_, _12539_, _12537_);
  not _63517_ (_12541_, _11872_);
  not _63518_ (_12542_, _07732_);
  and _63519_ (_12543_, _07638_, \oc8051_golden_model_1.P0 [2]);
  and _63520_ (_12544_, _08341_, \oc8051_golden_model_1.TCON [2]);
  and _63521_ (_12545_, _08345_, \oc8051_golden_model_1.P1 [2]);
  and _63522_ (_12546_, _08347_, \oc8051_golden_model_1.SCON [2]);
  and _63523_ (_12547_, _08349_, \oc8051_golden_model_1.P2 [2]);
  and _63524_ (_12548_, _08351_, \oc8051_golden_model_1.IE [2]);
  and _63525_ (_12549_, _08353_, \oc8051_golden_model_1.P3 [2]);
  and _63526_ (_12550_, _08357_, \oc8051_golden_model_1.IP [2]);
  and _63527_ (_12551_, _08355_, \oc8051_golden_model_1.PSW [2]);
  and _63528_ (_12552_, _08359_, \oc8051_golden_model_1.ACC [2]);
  and _63529_ (_12553_, _08361_, \oc8051_golden_model_1.B [2]);
  or _63530_ (_12554_, _12553_, _12552_);
  or _63531_ (_12555_, _12554_, _12551_);
  or _63532_ (_12556_, _12555_, _12550_);
  or _63533_ (_12557_, _12556_, _12549_);
  or _63534_ (_12558_, _12557_, _12548_);
  or _63535_ (_12559_, _12558_, _12547_);
  or _63536_ (_12560_, _12559_, _12546_);
  or _63537_ (_12561_, _12560_, _12545_);
  or _63538_ (_12562_, _12561_, _12544_);
  nor _63539_ (_12563_, _12562_, _12543_);
  and _63540_ (_12564_, _12563_, _08175_);
  nor _63541_ (_12565_, _12564_, _12542_);
  not _63542_ (_12566_, _07726_);
  and _63543_ (_12567_, _08357_, \oc8051_golden_model_1.IP [1]);
  and _63544_ (_12568_, _08355_, \oc8051_golden_model_1.PSW [1]);
  and _63545_ (_12569_, _08359_, \oc8051_golden_model_1.ACC [1]);
  and _63546_ (_12570_, _08361_, \oc8051_golden_model_1.B [1]);
  or _63547_ (_12571_, _12570_, _12569_);
  or _63548_ (_12572_, _12571_, _12568_);
  and _63549_ (_12573_, _08341_, \oc8051_golden_model_1.TCON [1]);
  and _63550_ (_12574_, _07638_, \oc8051_golden_model_1.P0 [1]);
  and _63551_ (_12575_, _08345_, \oc8051_golden_model_1.P1 [1]);
  or _63552_ (_12576_, _12575_, _12574_);
  or _63553_ (_12577_, _12576_, _12573_);
  and _63554_ (_12578_, _08353_, \oc8051_golden_model_1.P3 [1]);
  and _63555_ (_12579_, _08351_, \oc8051_golden_model_1.IE [1]);
  or _63556_ (_12580_, _12579_, _12578_);
  and _63557_ (_12581_, _08347_, \oc8051_golden_model_1.SCON [1]);
  and _63558_ (_12582_, _08349_, \oc8051_golden_model_1.P2 [1]);
  or _63559_ (_12583_, _12582_, _12581_);
  or _63560_ (_12584_, _12583_, _12580_);
  or _63561_ (_12585_, _12584_, _12577_);
  or _63562_ (_12586_, _12585_, _12572_);
  nor _63563_ (_12587_, _12586_, _12567_);
  and _63564_ (_12588_, _12587_, _08076_);
  nor _63565_ (_12589_, _12588_, _12566_);
  nor _63566_ (_12590_, _12589_, _12565_);
  and _63567_ (_12591_, _07644_, _06403_);
  not _63568_ (_12592_, _12591_);
  and _63569_ (_12593_, _07638_, \oc8051_golden_model_1.P0 [0]);
  and _63570_ (_12594_, _08341_, \oc8051_golden_model_1.TCON [0]);
  and _63571_ (_12595_, _08345_, \oc8051_golden_model_1.P1 [0]);
  and _63572_ (_12596_, _08347_, \oc8051_golden_model_1.SCON [0]);
  and _63573_ (_12597_, _08349_, \oc8051_golden_model_1.P2 [0]);
  and _63574_ (_12598_, _08351_, \oc8051_golden_model_1.IE [0]);
  and _63575_ (_12599_, _08353_, \oc8051_golden_model_1.P3 [0]);
  and _63576_ (_12600_, _08357_, \oc8051_golden_model_1.IP [0]);
  and _63577_ (_12601_, _08355_, \oc8051_golden_model_1.PSW [0]);
  and _63578_ (_12602_, _08359_, \oc8051_golden_model_1.ACC [0]);
  and _63579_ (_12603_, _08361_, \oc8051_golden_model_1.B [0]);
  or _63580_ (_12604_, _12603_, _12602_);
  or _63581_ (_12605_, _12604_, _12601_);
  or _63582_ (_12606_, _12605_, _12600_);
  or _63583_ (_12607_, _12606_, _12599_);
  or _63584_ (_12608_, _12607_, _12598_);
  or _63585_ (_12609_, _12608_, _12597_);
  or _63586_ (_12610_, _12609_, _12596_);
  or _63587_ (_12611_, _12610_, _12595_);
  or _63588_ (_12612_, _12611_, _12594_);
  nor _63589_ (_12613_, _12612_, _12593_);
  not _63590_ (_12614_, _12613_);
  nor _63591_ (_12615_, _12614_, _08126_);
  nor _63592_ (_12616_, _12615_, _12592_);
  and _63593_ (_12617_, _07638_, \oc8051_golden_model_1.P0 [5]);
  and _63594_ (_12618_, _08341_, \oc8051_golden_model_1.TCON [5]);
  and _63595_ (_12619_, _08345_, \oc8051_golden_model_1.P1 [5]);
  and _63596_ (_12620_, _08347_, \oc8051_golden_model_1.SCON [5]);
  and _63597_ (_12621_, _08349_, \oc8051_golden_model_1.P2 [5]);
  and _63598_ (_12622_, _08351_, \oc8051_golden_model_1.IE [5]);
  and _63599_ (_12623_, _08353_, \oc8051_golden_model_1.P3 [5]);
  and _63600_ (_12624_, _08357_, \oc8051_golden_model_1.IP [5]);
  and _63601_ (_12625_, _08355_, \oc8051_golden_model_1.PSW [5]);
  and _63602_ (_12626_, _08359_, \oc8051_golden_model_1.ACC [5]);
  and _63603_ (_12627_, _08361_, \oc8051_golden_model_1.B [5]);
  or _63604_ (_12628_, _12627_, _12626_);
  or _63605_ (_12629_, _12628_, _12625_);
  or _63606_ (_12630_, _12629_, _12624_);
  or _63607_ (_12631_, _12630_, _12623_);
  or _63608_ (_12632_, _12631_, _12622_);
  or _63609_ (_12633_, _12632_, _12621_);
  or _63610_ (_12634_, _12633_, _12620_);
  or _63611_ (_12635_, _12634_, _12619_);
  or _63612_ (_12636_, _12635_, _12618_);
  nor _63613_ (_12637_, _12636_, _12617_);
  and _63614_ (_12638_, _12637_, _07978_);
  and _63615_ (_12639_, _07650_, _07477_);
  not _63616_ (_12640_, _12639_);
  nor _63617_ (_12641_, _12640_, _12638_);
  nor _63618_ (_12642_, _12641_, _12616_);
  and _63619_ (_12643_, _12642_, _12590_);
  not _63620_ (_12644_, _07723_);
  and _63621_ (_12645_, _08357_, \oc8051_golden_model_1.IP [3]);
  and _63622_ (_12646_, _08355_, \oc8051_golden_model_1.PSW [3]);
  and _63623_ (_12647_, _08361_, \oc8051_golden_model_1.B [3]);
  and _63624_ (_12648_, _08359_, \oc8051_golden_model_1.ACC [3]);
  or _63625_ (_12649_, _12648_, _12647_);
  or _63626_ (_12650_, _12649_, _12646_);
  and _63627_ (_12651_, _08341_, \oc8051_golden_model_1.TCON [3]);
  and _63628_ (_12652_, _07638_, \oc8051_golden_model_1.P0 [3]);
  and _63629_ (_12653_, _08345_, \oc8051_golden_model_1.P1 [3]);
  or _63630_ (_12654_, _12653_, _12652_);
  or _63631_ (_12655_, _12654_, _12651_);
  and _63632_ (_12656_, _08353_, \oc8051_golden_model_1.P3 [3]);
  and _63633_ (_12657_, _08351_, \oc8051_golden_model_1.IE [3]);
  or _63634_ (_12658_, _12657_, _12656_);
  and _63635_ (_12659_, _08347_, \oc8051_golden_model_1.SCON [3]);
  and _63636_ (_12660_, _08349_, \oc8051_golden_model_1.P2 [3]);
  or _63637_ (_12661_, _12660_, _12659_);
  or _63638_ (_12662_, _12661_, _12658_);
  or _63639_ (_12663_, _12662_, _12655_);
  or _63640_ (_12664_, _12663_, _12650_);
  nor _63641_ (_12665_, _12664_, _12645_);
  and _63642_ (_12666_, _12665_, _08027_);
  nor _63643_ (_12667_, _12666_, _12644_);
  nor _63644_ (_12668_, _12667_, _08518_);
  and _63645_ (_12669_, _07638_, \oc8051_golden_model_1.P0 [6]);
  and _63646_ (_12670_, _08341_, \oc8051_golden_model_1.TCON [6]);
  and _63647_ (_12671_, _08345_, \oc8051_golden_model_1.P1 [6]);
  and _63648_ (_12672_, _08347_, \oc8051_golden_model_1.SCON [6]);
  and _63649_ (_12673_, _08349_, \oc8051_golden_model_1.P2 [6]);
  and _63650_ (_12674_, _08351_, \oc8051_golden_model_1.IE [6]);
  and _63651_ (_12675_, _08353_, \oc8051_golden_model_1.P3 [6]);
  and _63652_ (_12676_, _08357_, \oc8051_golden_model_1.IP [6]);
  and _63653_ (_12677_, _08355_, \oc8051_golden_model_1.PSW [6]);
  and _63654_ (_12678_, _08359_, \oc8051_golden_model_1.ACC [6]);
  and _63655_ (_12679_, _08361_, \oc8051_golden_model_1.B [6]);
  or _63656_ (_12680_, _12679_, _12678_);
  or _63657_ (_12681_, _12680_, _12677_);
  or _63658_ (_12682_, _12681_, _12676_);
  or _63659_ (_12683_, _12682_, _12675_);
  or _63660_ (_12684_, _12683_, _12674_);
  or _63661_ (_12685_, _12684_, _12673_);
  or _63662_ (_12686_, _12685_, _12672_);
  or _63663_ (_12687_, _12686_, _12671_);
  or _63664_ (_12688_, _12687_, _12670_);
  nor _63665_ (_12689_, _12688_, _12669_);
  and _63666_ (_12690_, _12689_, _07884_);
  and _63667_ (_12691_, _07656_, _07477_);
  not _63668_ (_12692_, _12691_);
  nor _63669_ (_12693_, _12692_, _12690_);
  and _63670_ (_12694_, _08349_, \oc8051_golden_model_1.P2 [4]);
  and _63671_ (_12695_, _08351_, \oc8051_golden_model_1.IE [4]);
  and _63672_ (_12696_, _08353_, \oc8051_golden_model_1.P3 [4]);
  or _63673_ (_12697_, _12696_, _12695_);
  nor _63674_ (_12698_, _12697_, _12694_);
  and _63675_ (_12699_, _08341_, \oc8051_golden_model_1.TCON [4]);
  and _63676_ (_12700_, _08345_, \oc8051_golden_model_1.P1 [4]);
  and _63677_ (_12701_, _07638_, \oc8051_golden_model_1.P0 [4]);
  or _63678_ (_12702_, _12701_, _12700_);
  nor _63679_ (_12703_, _12702_, _12699_);
  and _63680_ (_12704_, _08357_, \oc8051_golden_model_1.IP [4]);
  and _63681_ (_12705_, _08361_, \oc8051_golden_model_1.B [4]);
  and _63682_ (_12706_, _08359_, \oc8051_golden_model_1.ACC [4]);
  or _63683_ (_12707_, _12706_, _12705_);
  nor _63684_ (_12708_, _12707_, _12704_);
  and _63685_ (_12709_, _08347_, \oc8051_golden_model_1.SCON [4]);
  and _63686_ (_12710_, _08355_, \oc8051_golden_model_1.PSW [4]);
  nor _63687_ (_12711_, _12710_, _12709_);
  and _63688_ (_12712_, _12711_, _12708_);
  and _63689_ (_12714_, _12712_, _12703_);
  and _63690_ (_12715_, _12714_, _12698_);
  and _63691_ (_12716_, _12715_, _08271_);
  and _63692_ (_12717_, _07644_, _07477_);
  not _63693_ (_12718_, _12717_);
  nor _63694_ (_12719_, _12718_, _12716_);
  nor _63695_ (_12720_, _12719_, _12693_);
  and _63696_ (_12721_, _12720_, _12668_);
  and _63697_ (_12722_, _12721_, _12643_);
  not _63698_ (_12723_, _12722_);
  or _63699_ (_12724_, _12141_, _12723_);
  or _63700_ (_12725_, _09227_, _12722_);
  and _63701_ (_12726_, _12725_, _06129_);
  and _63702_ (_12727_, _12726_, _12724_);
  or _63703_ (_12728_, _12727_, _12541_);
  or _63704_ (_12729_, _12728_, _12540_);
  and _63705_ (_12730_, _12729_, _11873_);
  or _63706_ (_12731_, _12730_, _10976_);
  or _63707_ (_12732_, _10975_, _09216_);
  and _63708_ (_12733_, _12732_, _11016_);
  and _63709_ (_12735_, _12733_, _12731_);
  and _63710_ (_12736_, _11871_, _11015_);
  or _63711_ (_12737_, _12736_, _06049_);
  or _63712_ (_12738_, _12737_, _12735_);
  nand _63713_ (_12739_, _07785_, _06049_);
  and _63714_ (_12740_, _12739_, _12738_);
  or _63715_ (_12741_, _12740_, _05747_);
  or _63716_ (_12742_, _09216_, _05748_);
  and _63717_ (_12743_, _12742_, _06704_);
  and _63718_ (_12744_, _12743_, _12741_);
  or _63719_ (_12745_, _12141_, _12722_);
  nand _63720_ (_12746_, _12010_, _12722_);
  and _63721_ (_12747_, _12746_, _12745_);
  and _63722_ (_12748_, _12747_, _06126_);
  and _63723_ (_12749_, _08287_, _07052_);
  not _63724_ (_12750_, _12749_);
  or _63725_ (_12751_, _12750_, _12748_);
  or _63726_ (_12752_, _12751_, _12744_);
  or _63727_ (_12753_, _12749_, _11871_);
  and _63728_ (_12754_, _12753_, _06718_);
  and _63729_ (_12755_, _12754_, _12752_);
  nor _63730_ (_12756_, _11064_, _11059_);
  nand _63731_ (_12757_, _09216_, _06316_);
  nand _63732_ (_12758_, _12757_, _12756_);
  or _63733_ (_12759_, _12758_, _12755_);
  or _63734_ (_12760_, _11871_, _12756_);
  and _63735_ (_12761_, _12760_, _09200_);
  and _63736_ (_12762_, _12761_, _12759_);
  and _63737_ (_12763_, _06127_, _05952_);
  or _63738_ (_12764_, _12763_, _05752_);
  or _63739_ (_12765_, _12764_, _12762_);
  not _63740_ (_12766_, _05752_);
  or _63741_ (_12767_, _09216_, _12766_);
  and _63742_ (_12768_, _12767_, _05653_);
  and _63743_ (_12769_, _12768_, _12765_);
  and _63744_ (_12770_, _12747_, _05652_);
  and _63745_ (_12771_, _09154_, _07069_);
  not _63746_ (_12772_, _12771_);
  or _63747_ (_12773_, _12772_, _12770_);
  or _63748_ (_12774_, _12773_, _12769_);
  or _63749_ (_12775_, _12771_, _11871_);
  and _63750_ (_12776_, _12775_, _06048_);
  and _63751_ (_12777_, _12776_, _12774_);
  nand _63752_ (_12778_, _09216_, _06047_);
  nor _63753_ (_12779_, _11089_, _11082_);
  nand _63754_ (_12780_, _12779_, _12778_);
  or _63755_ (_12781_, _12780_, _12777_);
  not _63756_ (_12782_, _06119_);
  or _63757_ (_12783_, _12779_, _11871_);
  and _63758_ (_12784_, _12783_, _12782_);
  and _63759_ (_12785_, _12784_, _12781_);
  and _63760_ (_12786_, _06119_, _05952_);
  or _63761_ (_12787_, _12786_, _05751_);
  or _63762_ (_12788_, _12787_, _12785_);
  and _63763_ (_12789_, _05750_, _05650_);
  not _63764_ (_12790_, _12789_);
  not _63765_ (_12791_, _05751_);
  or _63766_ (_12792_, _09216_, _12791_);
  and _63767_ (_12793_, _12792_, _12790_);
  and _63768_ (_12794_, _12793_, _12788_);
  and _63769_ (_12795_, _12789_, _11871_);
  or _63770_ (_12796_, _12795_, _12794_);
  or _63771_ (_12797_, _12796_, _01340_);
  or _63772_ (_12798_, _01336_, \oc8051_golden_model_1.PC [15]);
  and _63773_ (_12799_, _12798_, _42882_);
  and _63774_ (_40766_, _12799_, _12797_);
  not _63775_ (_12800_, _07686_);
  and _63776_ (_12801_, _12800_, \oc8051_golden_model_1.P2 [7]);
  and _63777_ (_12802_, _08768_, _07686_);
  or _63778_ (_12803_, _12802_, _12801_);
  and _63779_ (_12804_, _12803_, _06284_);
  and _63780_ (_12805_, _08549_, _07686_);
  or _63781_ (_12806_, _12805_, _12801_);
  or _63782_ (_12807_, _12806_, _06020_);
  and _63783_ (_12808_, _08498_, _07686_);
  or _63784_ (_12809_, _12808_, _12801_);
  or _63785_ (_12810_, _12809_, _06954_);
  and _63786_ (_12811_, _07686_, \oc8051_golden_model_1.ACC [7]);
  or _63787_ (_12812_, _12811_, _12801_);
  and _63788_ (_12813_, _12812_, _06938_);
  and _63789_ (_12814_, _06939_, \oc8051_golden_model_1.P2 [7]);
  or _63790_ (_12815_, _12814_, _06102_);
  or _63791_ (_12816_, _12815_, _12813_);
  and _63792_ (_12817_, _12816_, _06044_);
  and _63793_ (_12818_, _12817_, _12810_);
  not _63794_ (_12819_, _08349_);
  and _63795_ (_12820_, _12819_, \oc8051_golden_model_1.P2 [7]);
  and _63796_ (_12821_, _08503_, _08349_);
  or _63797_ (_12822_, _12821_, _12820_);
  and _63798_ (_12823_, _12822_, _06043_);
  or _63799_ (_12824_, _12823_, _06239_);
  or _63800_ (_12825_, _12824_, _12818_);
  nor _63801_ (_12826_, _07785_, _12800_);
  or _63802_ (_12827_, _12826_, _12801_);
  or _63803_ (_12828_, _12827_, _06848_);
  and _63804_ (_12829_, _12828_, _12825_);
  or _63805_ (_12830_, _12829_, _06219_);
  or _63806_ (_12831_, _12812_, _06220_);
  and _63807_ (_12832_, _12831_, _06040_);
  and _63808_ (_12833_, _12832_, _12830_);
  and _63809_ (_12834_, _08374_, _08349_);
  or _63810_ (_12835_, _12834_, _12820_);
  and _63811_ (_12836_, _12835_, _06039_);
  or _63812_ (_12837_, _12836_, _06032_);
  or _63813_ (_12838_, _12837_, _12833_);
  or _63814_ (_12839_, _12820_, _08519_);
  and _63815_ (_12840_, _12839_, _12822_);
  or _63816_ (_12841_, _12840_, _06033_);
  and _63817_ (_12842_, _12841_, _06027_);
  and _63818_ (_12843_, _12842_, _12838_);
  and _63819_ (_12844_, _08376_, _08349_);
  or _63820_ (_12845_, _12844_, _12820_);
  and _63821_ (_12846_, _12845_, _06026_);
  or _63822_ (_12847_, _12846_, _09818_);
  or _63823_ (_12848_, _12847_, _12843_);
  and _63824_ (_12849_, _08485_, _07686_);
  or _63825_ (_12850_, _12801_, _07012_);
  or _63826_ (_12851_, _12850_, _12849_);
  or _63827_ (_12852_, _12827_, _09827_);
  and _63828_ (_12853_, _12852_, _05669_);
  and _63829_ (_12854_, _12853_, _12851_);
  and _63830_ (_12855_, _12854_, _12848_);
  and _63831_ (_12856_, _08738_, _07686_);
  or _63832_ (_12857_, _12856_, _12801_);
  and _63833_ (_12858_, _12857_, _09833_);
  or _63834_ (_12859_, _12858_, _06019_);
  or _63835_ (_12860_, _12859_, _12855_);
  and _63836_ (_12861_, _12860_, _12807_);
  or _63837_ (_12862_, _12861_, _06112_);
  and _63838_ (_12863_, _08760_, _07686_);
  or _63839_ (_12864_, _12801_, _08751_);
  or _63840_ (_12865_, _12864_, _12863_);
  and _63841_ (_12866_, _12865_, _08756_);
  and _63842_ (_12867_, _12866_, _12862_);
  or _63843_ (_12868_, _12867_, _12804_);
  and _63844_ (_12869_, _12868_, _07032_);
  or _63845_ (_12870_, _12801_, _07788_);
  and _63846_ (_12871_, _12806_, _06108_);
  and _63847_ (_12872_, _12871_, _12870_);
  or _63848_ (_12873_, _12872_, _12869_);
  and _63849_ (_12874_, _12873_, _06278_);
  and _63850_ (_12875_, _12812_, _06277_);
  and _63851_ (_12876_, _12875_, _12870_);
  or _63852_ (_12877_, _12876_, _06130_);
  or _63853_ (_12878_, _12877_, _12874_);
  and _63854_ (_12879_, _08759_, _07686_);
  or _63855_ (_12880_, _12801_, _08777_);
  or _63856_ (_12881_, _12880_, _12879_);
  and _63857_ (_12882_, _12881_, _08782_);
  and _63858_ (_12883_, _12882_, _12878_);
  nor _63859_ (_12884_, _08767_, _12800_);
  or _63860_ (_12885_, _12884_, _12801_);
  and _63861_ (_12886_, _12885_, _06292_);
  or _63862_ (_12887_, _12886_, _06316_);
  or _63863_ (_12888_, _12887_, _12883_);
  or _63864_ (_12889_, _12809_, _06718_);
  and _63865_ (_12890_, _12889_, _05653_);
  and _63866_ (_12891_, _12890_, _12888_);
  and _63867_ (_12892_, _12835_, _05652_);
  or _63868_ (_12893_, _12892_, _06047_);
  or _63869_ (_12894_, _12893_, _12891_);
  and _63870_ (_12895_, _08279_, _07686_);
  or _63871_ (_12896_, _12801_, _06048_);
  or _63872_ (_12897_, _12896_, _12895_);
  and _63873_ (_12898_, _12897_, _01336_);
  and _63874_ (_12899_, _12898_, _12894_);
  nor _63875_ (_12900_, \oc8051_golden_model_1.P2 [7], rst);
  nor _63876_ (_12901_, _12900_, _00000_);
  or _63877_ (_40768_, _12901_, _12899_);
  not _63878_ (_12902_, _07692_);
  and _63879_ (_12903_, _12902_, \oc8051_golden_model_1.P3 [7]);
  and _63880_ (_12904_, _08768_, _07692_);
  or _63881_ (_12905_, _12904_, _12903_);
  and _63882_ (_12906_, _12905_, _06284_);
  and _63883_ (_12907_, _08549_, _07692_);
  or _63884_ (_12908_, _12907_, _12903_);
  or _63885_ (_12909_, _12908_, _06020_);
  and _63886_ (_12910_, _08498_, _07692_);
  or _63887_ (_12911_, _12910_, _12903_);
  or _63888_ (_12912_, _12911_, _06954_);
  and _63889_ (_12913_, _07692_, \oc8051_golden_model_1.ACC [7]);
  or _63890_ (_12914_, _12913_, _12903_);
  and _63891_ (_12915_, _12914_, _06938_);
  and _63892_ (_12916_, _06939_, \oc8051_golden_model_1.P3 [7]);
  or _63893_ (_12917_, _12916_, _06102_);
  or _63894_ (_12918_, _12917_, _12915_);
  and _63895_ (_12919_, _12918_, _06044_);
  and _63896_ (_12920_, _12919_, _12912_);
  not _63897_ (_12921_, _08353_);
  and _63898_ (_12922_, _12921_, \oc8051_golden_model_1.P3 [7]);
  and _63899_ (_12923_, _08503_, _08353_);
  or _63900_ (_12924_, _12923_, _12922_);
  and _63901_ (_12925_, _12924_, _06043_);
  or _63902_ (_12926_, _12925_, _06239_);
  or _63903_ (_12927_, _12926_, _12920_);
  nor _63904_ (_12928_, _07785_, _12902_);
  or _63905_ (_12929_, _12928_, _12903_);
  or _63906_ (_12930_, _12929_, _06848_);
  and _63907_ (_12931_, _12930_, _12927_);
  or _63908_ (_12932_, _12931_, _06219_);
  or _63909_ (_12933_, _12914_, _06220_);
  and _63910_ (_12934_, _12933_, _06040_);
  and _63911_ (_12935_, _12934_, _12932_);
  and _63912_ (_12936_, _08374_, _08353_);
  or _63913_ (_12937_, _12936_, _12922_);
  and _63914_ (_12938_, _12937_, _06039_);
  or _63915_ (_12939_, _12938_, _06032_);
  or _63916_ (_12940_, _12939_, _12935_);
  or _63917_ (_12941_, _12922_, _08519_);
  and _63918_ (_12942_, _12941_, _12924_);
  or _63919_ (_12943_, _12942_, _06033_);
  and _63920_ (_12944_, _12943_, _06027_);
  and _63921_ (_12945_, _12944_, _12940_);
  and _63922_ (_12946_, _08376_, _08353_);
  or _63923_ (_12947_, _12946_, _12922_);
  and _63924_ (_12948_, _12947_, _06026_);
  or _63925_ (_12949_, _12948_, _09818_);
  or _63926_ (_12950_, _12949_, _12945_);
  and _63927_ (_12951_, _08485_, _07692_);
  or _63928_ (_12952_, _12903_, _07012_);
  or _63929_ (_12953_, _12952_, _12951_);
  or _63930_ (_12954_, _12929_, _09827_);
  and _63931_ (_12955_, _12954_, _05669_);
  and _63932_ (_12956_, _12955_, _12953_);
  and _63933_ (_12957_, _12956_, _12950_);
  and _63934_ (_12958_, _08738_, _07692_);
  or _63935_ (_12959_, _12958_, _12903_);
  and _63936_ (_12960_, _12959_, _09833_);
  or _63937_ (_12961_, _12960_, _06019_);
  or _63938_ (_12962_, _12961_, _12957_);
  and _63939_ (_12963_, _12962_, _12909_);
  or _63940_ (_12964_, _12963_, _06112_);
  and _63941_ (_12965_, _08760_, _07692_);
  or _63942_ (_12966_, _12965_, _12903_);
  or _63943_ (_12967_, _12966_, _08751_);
  and _63944_ (_12968_, _12967_, _08756_);
  and _63945_ (_12969_, _12968_, _12964_);
  or _63946_ (_12970_, _12969_, _12906_);
  and _63947_ (_12971_, _12970_, _07032_);
  or _63948_ (_12972_, _12903_, _07788_);
  and _63949_ (_12973_, _12908_, _06108_);
  and _63950_ (_12974_, _12973_, _12972_);
  or _63951_ (_12975_, _12974_, _12971_);
  and _63952_ (_12976_, _12975_, _06278_);
  and _63953_ (_12977_, _12914_, _06277_);
  and _63954_ (_12978_, _12977_, _12972_);
  or _63955_ (_12979_, _12978_, _06130_);
  or _63956_ (_12980_, _12979_, _12976_);
  and _63957_ (_12981_, _08759_, _07692_);
  or _63958_ (_12982_, _12903_, _08777_);
  or _63959_ (_12983_, _12982_, _12981_);
  and _63960_ (_12984_, _12983_, _08782_);
  and _63961_ (_12985_, _12984_, _12980_);
  nor _63962_ (_12986_, _08767_, _12902_);
  or _63963_ (_12987_, _12986_, _12903_);
  and _63964_ (_12988_, _12987_, _06292_);
  or _63965_ (_12989_, _12988_, _06316_);
  or _63966_ (_12990_, _12989_, _12985_);
  or _63967_ (_12991_, _12911_, _06718_);
  and _63968_ (_12992_, _12991_, _05653_);
  and _63969_ (_12993_, _12992_, _12990_);
  and _63970_ (_12994_, _12937_, _05652_);
  or _63971_ (_12995_, _12994_, _06047_);
  or _63972_ (_12996_, _12995_, _12993_);
  and _63973_ (_12997_, _08279_, _07692_);
  or _63974_ (_12998_, _12903_, _06048_);
  or _63975_ (_12999_, _12998_, _12997_);
  and _63976_ (_13000_, _12999_, _01336_);
  and _63977_ (_13001_, _13000_, _12996_);
  nor _63978_ (_13002_, \oc8051_golden_model_1.P3 [7], rst);
  nor _63979_ (_13003_, _13002_, _00000_);
  or _63980_ (_40769_, _13003_, _13001_);
  nor _63981_ (_13004_, \oc8051_golden_model_1.P0 [7], rst);
  nor _63982_ (_13005_, _13004_, _00000_);
  not _63983_ (_13006_, _07730_);
  and _63984_ (_13007_, _13006_, \oc8051_golden_model_1.P0 [7]);
  and _63985_ (_13008_, _08768_, _07730_);
  or _63986_ (_13009_, _13008_, _13007_);
  and _63987_ (_13010_, _13009_, _06284_);
  and _63988_ (_13011_, _08549_, _07730_);
  or _63989_ (_13012_, _13011_, _13007_);
  or _63990_ (_13013_, _13012_, _06020_);
  and _63991_ (_13014_, _08498_, _07730_);
  or _63992_ (_13015_, _13014_, _13007_);
  or _63993_ (_13016_, _13015_, _06954_);
  and _63994_ (_13017_, _07730_, \oc8051_golden_model_1.ACC [7]);
  or _63995_ (_13018_, _13017_, _13007_);
  and _63996_ (_13019_, _13018_, _06938_);
  and _63997_ (_13020_, _06939_, \oc8051_golden_model_1.P0 [7]);
  or _63998_ (_13021_, _13020_, _06102_);
  or _63999_ (_13022_, _13021_, _13019_);
  and _64000_ (_13023_, _13022_, _06044_);
  and _64001_ (_13024_, _13023_, _13016_);
  not _64002_ (_13025_, _07638_);
  and _64003_ (_13026_, _13025_, \oc8051_golden_model_1.P0 [7]);
  and _64004_ (_13027_, _08503_, _07638_);
  or _64005_ (_13028_, _13027_, _13026_);
  and _64006_ (_13029_, _13028_, _06043_);
  or _64007_ (_13030_, _13029_, _06239_);
  or _64008_ (_13031_, _13030_, _13024_);
  nor _64009_ (_13032_, _07785_, _13006_);
  or _64010_ (_13033_, _13032_, _13007_);
  or _64011_ (_13034_, _13033_, _06848_);
  and _64012_ (_13035_, _13034_, _13031_);
  or _64013_ (_13036_, _13035_, _06219_);
  or _64014_ (_13037_, _13018_, _06220_);
  and _64015_ (_13038_, _13037_, _06040_);
  and _64016_ (_13039_, _13038_, _13036_);
  and _64017_ (_13040_, _08374_, _07638_);
  or _64018_ (_13041_, _13040_, _13026_);
  and _64019_ (_13042_, _13041_, _06039_);
  or _64020_ (_13043_, _13042_, _06032_);
  or _64021_ (_13044_, _13043_, _13039_);
  or _64022_ (_13045_, _13026_, _08519_);
  and _64023_ (_13046_, _13045_, _13028_);
  or _64024_ (_13047_, _13046_, _06033_);
  and _64025_ (_13048_, _13047_, _06027_);
  and _64026_ (_13049_, _13048_, _13044_);
  and _64027_ (_13050_, _08376_, _07638_);
  or _64028_ (_13051_, _13050_, _13026_);
  and _64029_ (_13052_, _13051_, _06026_);
  or _64030_ (_13053_, _13052_, _09818_);
  or _64031_ (_13054_, _13053_, _13049_);
  and _64032_ (_13055_, _08485_, _07730_);
  or _64033_ (_13056_, _13007_, _07012_);
  or _64034_ (_13057_, _13056_, _13055_);
  or _64035_ (_13058_, _13033_, _09827_);
  and _64036_ (_13059_, _13058_, _05669_);
  and _64037_ (_13060_, _13059_, _13057_);
  and _64038_ (_13061_, _13060_, _13054_);
  and _64039_ (_13062_, _08738_, _07730_);
  or _64040_ (_13063_, _13062_, _13007_);
  and _64041_ (_13064_, _13063_, _09833_);
  or _64042_ (_13065_, _13064_, _06019_);
  or _64043_ (_13066_, _13065_, _13061_);
  and _64044_ (_13067_, _13066_, _13013_);
  or _64045_ (_13068_, _13067_, _06112_);
  and _64046_ (_13069_, _08760_, _07730_);
  or _64047_ (_13070_, _13007_, _08751_);
  or _64048_ (_13071_, _13070_, _13069_);
  and _64049_ (_13072_, _13071_, _08756_);
  and _64050_ (_13073_, _13072_, _13068_);
  or _64051_ (_13074_, _13073_, _13010_);
  and _64052_ (_13075_, _13074_, _07032_);
  or _64053_ (_13076_, _13007_, _07788_);
  and _64054_ (_13077_, _13012_, _06108_);
  and _64055_ (_13078_, _13077_, _13076_);
  or _64056_ (_13079_, _13078_, _13075_);
  and _64057_ (_13080_, _13079_, _06278_);
  and _64058_ (_13081_, _13018_, _06277_);
  and _64059_ (_13082_, _13081_, _13076_);
  or _64060_ (_13083_, _13082_, _06130_);
  or _64061_ (_13084_, _13083_, _13080_);
  and _64062_ (_13085_, _08759_, _07730_);
  or _64063_ (_13086_, _13007_, _08777_);
  or _64064_ (_13087_, _13086_, _13085_);
  and _64065_ (_13088_, _13087_, _08782_);
  and _64066_ (_13089_, _13088_, _13084_);
  nor _64067_ (_13090_, _08767_, _13006_);
  or _64068_ (_13091_, _13090_, _13007_);
  and _64069_ (_13092_, _13091_, _06292_);
  or _64070_ (_13093_, _13092_, _06316_);
  or _64071_ (_13094_, _13093_, _13089_);
  or _64072_ (_13095_, _13015_, _06718_);
  and _64073_ (_13096_, _13095_, _05653_);
  and _64074_ (_13097_, _13096_, _13094_);
  and _64075_ (_13098_, _13041_, _05652_);
  or _64076_ (_13099_, _13098_, _06047_);
  or _64077_ (_13100_, _13099_, _13097_);
  and _64078_ (_13101_, _08279_, _07730_);
  or _64079_ (_13102_, _13007_, _06048_);
  or _64080_ (_13103_, _13102_, _13101_);
  and _64081_ (_13104_, _13103_, _01336_);
  and _64082_ (_13105_, _13104_, _13100_);
  or _64083_ (_40770_, _13105_, _13005_);
  nor _64084_ (_13106_, \oc8051_golden_model_1.P1 [7], rst);
  nor _64085_ (_13107_, _13106_, _00000_);
  not _64086_ (_13108_, _07677_);
  and _64087_ (_13109_, _13108_, \oc8051_golden_model_1.P1 [7]);
  and _64088_ (_13110_, _08768_, _07677_);
  or _64089_ (_13111_, _13110_, _13109_);
  and _64090_ (_13112_, _13111_, _06284_);
  and _64091_ (_13113_, _08549_, _07677_);
  or _64092_ (_13114_, _13113_, _13109_);
  or _64093_ (_13115_, _13114_, _06020_);
  and _64094_ (_13116_, _08498_, _07677_);
  or _64095_ (_13117_, _13116_, _13109_);
  or _64096_ (_13118_, _13117_, _06954_);
  and _64097_ (_13119_, _07677_, \oc8051_golden_model_1.ACC [7]);
  or _64098_ (_13120_, _13119_, _13109_);
  and _64099_ (_13121_, _13120_, _06938_);
  and _64100_ (_13122_, _06939_, \oc8051_golden_model_1.P1 [7]);
  or _64101_ (_13123_, _13122_, _06102_);
  or _64102_ (_13124_, _13123_, _13121_);
  and _64103_ (_13125_, _13124_, _06044_);
  and _64104_ (_13126_, _13125_, _13118_);
  not _64105_ (_13127_, _08345_);
  and _64106_ (_13128_, _13127_, \oc8051_golden_model_1.P1 [7]);
  and _64107_ (_13129_, _08503_, _08345_);
  or _64108_ (_13130_, _13129_, _13128_);
  and _64109_ (_13131_, _13130_, _06043_);
  or _64110_ (_13132_, _13131_, _06239_);
  or _64111_ (_13133_, _13132_, _13126_);
  nor _64112_ (_13134_, _07785_, _13108_);
  or _64113_ (_13135_, _13134_, _13109_);
  or _64114_ (_13136_, _13135_, _06848_);
  and _64115_ (_13137_, _13136_, _13133_);
  or _64116_ (_13138_, _13137_, _06219_);
  or _64117_ (_13139_, _13120_, _06220_);
  and _64118_ (_13140_, _13139_, _06040_);
  and _64119_ (_13141_, _13140_, _13138_);
  and _64120_ (_13142_, _08374_, _08345_);
  or _64121_ (_13143_, _13142_, _13128_);
  and _64122_ (_13144_, _13143_, _06039_);
  or _64123_ (_13145_, _13144_, _06032_);
  or _64124_ (_13146_, _13145_, _13141_);
  or _64125_ (_13147_, _13128_, _08519_);
  and _64126_ (_13148_, _13147_, _13130_);
  or _64127_ (_13149_, _13148_, _06033_);
  and _64128_ (_13150_, _13149_, _06027_);
  and _64129_ (_13151_, _13150_, _13146_);
  and _64130_ (_13152_, _08376_, _08345_);
  or _64131_ (_13153_, _13152_, _13128_);
  and _64132_ (_13154_, _13153_, _06026_);
  or _64133_ (_13155_, _13154_, _09818_);
  or _64134_ (_13156_, _13155_, _13151_);
  and _64135_ (_13157_, _08485_, _07677_);
  or _64136_ (_13158_, _13109_, _07012_);
  or _64137_ (_13159_, _13158_, _13157_);
  or _64138_ (_13160_, _13135_, _09827_);
  and _64139_ (_13161_, _13160_, _05669_);
  and _64140_ (_13162_, _13161_, _13159_);
  and _64141_ (_13163_, _13162_, _13156_);
  and _64142_ (_13164_, _08738_, _07677_);
  or _64143_ (_13165_, _13164_, _13109_);
  and _64144_ (_13166_, _13165_, _09833_);
  or _64145_ (_13167_, _13166_, _06019_);
  or _64146_ (_13168_, _13167_, _13163_);
  and _64147_ (_13169_, _13168_, _13115_);
  or _64148_ (_13170_, _13169_, _06112_);
  and _64149_ (_13171_, _08760_, _07677_);
  or _64150_ (_13172_, _13171_, _13109_);
  or _64151_ (_13173_, _13172_, _08751_);
  and _64152_ (_13174_, _13173_, _08756_);
  and _64153_ (_13175_, _13174_, _13170_);
  or _64154_ (_13176_, _13175_, _13112_);
  and _64155_ (_13177_, _13176_, _07032_);
  or _64156_ (_13178_, _13109_, _07788_);
  and _64157_ (_13179_, _13114_, _06108_);
  and _64158_ (_13180_, _13179_, _13178_);
  or _64159_ (_13181_, _13180_, _13177_);
  and _64160_ (_13182_, _13181_, _06278_);
  and _64161_ (_13183_, _13120_, _06277_);
  and _64162_ (_13184_, _13183_, _13178_);
  or _64163_ (_13185_, _13184_, _06130_);
  or _64164_ (_13186_, _13185_, _13182_);
  and _64165_ (_13187_, _08759_, _07677_);
  or _64166_ (_13188_, _13109_, _08777_);
  or _64167_ (_13189_, _13188_, _13187_);
  and _64168_ (_13190_, _13189_, _08782_);
  and _64169_ (_13191_, _13190_, _13186_);
  nor _64170_ (_13192_, _08767_, _13108_);
  or _64171_ (_13193_, _13192_, _13109_);
  and _64172_ (_13194_, _13193_, _06292_);
  or _64173_ (_13195_, _13194_, _06316_);
  or _64174_ (_13196_, _13195_, _13191_);
  or _64175_ (_13197_, _13117_, _06718_);
  and _64176_ (_13198_, _13197_, _05653_);
  and _64177_ (_13199_, _13198_, _13196_);
  and _64178_ (_13200_, _13143_, _05652_);
  or _64179_ (_13201_, _13200_, _06047_);
  or _64180_ (_13202_, _13201_, _13199_);
  and _64181_ (_13203_, _08279_, _07677_);
  or _64182_ (_13204_, _13109_, _06048_);
  or _64183_ (_13205_, _13204_, _13203_);
  and _64184_ (_13206_, _13205_, _01336_);
  and _64185_ (_13207_, _13206_, _13202_);
  or _64186_ (_40771_, _13207_, _13107_);
  and _64187_ (_13208_, _01340_, \oc8051_golden_model_1.IP [7]);
  not _64188_ (_13209_, _07694_);
  and _64189_ (_13210_, _13209_, \oc8051_golden_model_1.IP [7]);
  and _64190_ (_13211_, _08768_, _07694_);
  or _64191_ (_13212_, _13211_, _13210_);
  and _64192_ (_13213_, _13212_, _06284_);
  and _64193_ (_13214_, _08549_, _07694_);
  or _64194_ (_13215_, _13214_, _13210_);
  or _64195_ (_13216_, _13215_, _06020_);
  and _64196_ (_13217_, _08498_, _07694_);
  or _64197_ (_13218_, _13217_, _13210_);
  or _64198_ (_13219_, _13218_, _06954_);
  and _64199_ (_13220_, _07694_, \oc8051_golden_model_1.ACC [7]);
  or _64200_ (_13221_, _13220_, _13210_);
  and _64201_ (_13222_, _13221_, _06938_);
  and _64202_ (_13223_, _06939_, \oc8051_golden_model_1.IP [7]);
  or _64203_ (_13224_, _13223_, _06102_);
  or _64204_ (_13225_, _13224_, _13222_);
  and _64205_ (_13226_, _13225_, _06044_);
  and _64206_ (_13227_, _13226_, _13219_);
  not _64207_ (_13228_, _08357_);
  and _64208_ (_13229_, _13228_, \oc8051_golden_model_1.IP [7]);
  and _64209_ (_13230_, _08503_, _08357_);
  or _64210_ (_13231_, _13230_, _13229_);
  and _64211_ (_13232_, _13231_, _06043_);
  or _64212_ (_13233_, _13232_, _06239_);
  or _64213_ (_13234_, _13233_, _13227_);
  nor _64214_ (_13235_, _07785_, _13209_);
  or _64215_ (_13236_, _13235_, _13210_);
  or _64216_ (_13237_, _13236_, _06848_);
  and _64217_ (_13238_, _13237_, _13234_);
  or _64218_ (_13239_, _13238_, _06219_);
  or _64219_ (_13240_, _13221_, _06220_);
  and _64220_ (_13241_, _13240_, _06040_);
  and _64221_ (_13242_, _13241_, _13239_);
  and _64222_ (_13243_, _08374_, _08357_);
  or _64223_ (_13244_, _13243_, _13229_);
  and _64224_ (_13245_, _13244_, _06039_);
  or _64225_ (_13246_, _13245_, _06032_);
  or _64226_ (_13247_, _13246_, _13242_);
  or _64227_ (_13248_, _13229_, _08519_);
  and _64228_ (_13249_, _13248_, _13231_);
  or _64229_ (_13250_, _13249_, _06033_);
  and _64230_ (_13251_, _13250_, _06027_);
  and _64231_ (_13252_, _13251_, _13247_);
  and _64232_ (_13253_, _08376_, _08357_);
  or _64233_ (_13254_, _13253_, _13229_);
  and _64234_ (_13255_, _13254_, _06026_);
  or _64235_ (_13256_, _13255_, _09818_);
  or _64236_ (_13257_, _13256_, _13252_);
  and _64237_ (_13258_, _08485_, _07694_);
  or _64238_ (_13259_, _13210_, _07012_);
  or _64239_ (_13260_, _13259_, _13258_);
  or _64240_ (_13261_, _13236_, _09827_);
  and _64241_ (_13262_, _13261_, _05669_);
  and _64242_ (_13263_, _13262_, _13260_);
  and _64243_ (_13264_, _13263_, _13257_);
  and _64244_ (_13265_, _08738_, _07694_);
  or _64245_ (_13266_, _13265_, _13210_);
  and _64246_ (_13267_, _13266_, _09833_);
  or _64247_ (_13268_, _13267_, _06019_);
  or _64248_ (_13269_, _13268_, _13264_);
  and _64249_ (_13270_, _13269_, _13216_);
  or _64250_ (_13271_, _13270_, _06112_);
  and _64251_ (_13272_, _08760_, _07694_);
  or _64252_ (_13273_, _13210_, _08751_);
  or _64253_ (_13274_, _13273_, _13272_);
  and _64254_ (_13275_, _13274_, _08756_);
  and _64255_ (_13276_, _13275_, _13271_);
  or _64256_ (_13277_, _13276_, _13213_);
  and _64257_ (_13278_, _13277_, _07032_);
  or _64258_ (_13279_, _13210_, _07788_);
  and _64259_ (_13280_, _13215_, _06108_);
  and _64260_ (_13281_, _13280_, _13279_);
  or _64261_ (_13282_, _13281_, _13278_);
  and _64262_ (_13283_, _13282_, _06278_);
  and _64263_ (_13284_, _13221_, _06277_);
  and _64264_ (_13285_, _13284_, _13279_);
  or _64265_ (_13286_, _13285_, _06130_);
  or _64266_ (_13287_, _13286_, _13283_);
  and _64267_ (_13288_, _08759_, _07694_);
  or _64268_ (_13289_, _13210_, _08777_);
  or _64269_ (_13290_, _13289_, _13288_);
  and _64270_ (_13291_, _13290_, _08782_);
  and _64271_ (_13292_, _13291_, _13287_);
  nor _64272_ (_13293_, _08767_, _13209_);
  or _64273_ (_13294_, _13293_, _13210_);
  and _64274_ (_13295_, _13294_, _06292_);
  or _64275_ (_13296_, _13295_, _06316_);
  or _64276_ (_13297_, _13296_, _13292_);
  or _64277_ (_13298_, _13218_, _06718_);
  and _64278_ (_13299_, _13298_, _05653_);
  and _64279_ (_13300_, _13299_, _13297_);
  and _64280_ (_13301_, _13244_, _05652_);
  or _64281_ (_13302_, _13301_, _06047_);
  or _64282_ (_13303_, _13302_, _13300_);
  and _64283_ (_13304_, _08279_, _07694_);
  or _64284_ (_13305_, _13210_, _06048_);
  or _64285_ (_13306_, _13305_, _13304_);
  and _64286_ (_13307_, _13306_, _01336_);
  and _64287_ (_13308_, _13307_, _13303_);
  or _64288_ (_13309_, _13308_, _13208_);
  and _64289_ (_40772_, _13309_, _42882_);
  and _64290_ (_13310_, _01340_, \oc8051_golden_model_1.IE [7]);
  not _64291_ (_13311_, _07688_);
  and _64292_ (_13312_, _13311_, \oc8051_golden_model_1.IE [7]);
  and _64293_ (_13313_, _08768_, _07688_);
  or _64294_ (_13314_, _13313_, _13312_);
  and _64295_ (_13315_, _13314_, _06284_);
  and _64296_ (_13316_, _08549_, _07688_);
  or _64297_ (_13317_, _13316_, _13312_);
  or _64298_ (_13318_, _13317_, _06020_);
  and _64299_ (_13319_, _08498_, _07688_);
  or _64300_ (_13320_, _13319_, _13312_);
  or _64301_ (_13321_, _13320_, _06954_);
  and _64302_ (_13322_, _07688_, \oc8051_golden_model_1.ACC [7]);
  or _64303_ (_13323_, _13322_, _13312_);
  and _64304_ (_13324_, _13323_, _06938_);
  and _64305_ (_13325_, _06939_, \oc8051_golden_model_1.IE [7]);
  or _64306_ (_13326_, _13325_, _06102_);
  or _64307_ (_13327_, _13326_, _13324_);
  and _64308_ (_13328_, _13327_, _06044_);
  and _64309_ (_13329_, _13328_, _13321_);
  not _64310_ (_13330_, _08351_);
  and _64311_ (_13331_, _13330_, \oc8051_golden_model_1.IE [7]);
  and _64312_ (_13332_, _08503_, _08351_);
  or _64313_ (_13333_, _13332_, _13331_);
  and _64314_ (_13334_, _13333_, _06043_);
  or _64315_ (_13335_, _13334_, _06239_);
  or _64316_ (_13336_, _13335_, _13329_);
  nor _64317_ (_13337_, _07785_, _13311_);
  or _64318_ (_13338_, _13337_, _13312_);
  or _64319_ (_13339_, _13338_, _06848_);
  and _64320_ (_13340_, _13339_, _13336_);
  or _64321_ (_13341_, _13340_, _06219_);
  or _64322_ (_13342_, _13323_, _06220_);
  and _64323_ (_13343_, _13342_, _06040_);
  and _64324_ (_13344_, _13343_, _13341_);
  and _64325_ (_13345_, _08374_, _08351_);
  or _64326_ (_13346_, _13345_, _13331_);
  and _64327_ (_13347_, _13346_, _06039_);
  or _64328_ (_13348_, _13347_, _06032_);
  or _64329_ (_13349_, _13348_, _13344_);
  or _64330_ (_13350_, _13331_, _08519_);
  and _64331_ (_13351_, _13350_, _13333_);
  or _64332_ (_13352_, _13351_, _06033_);
  and _64333_ (_13353_, _13352_, _06027_);
  and _64334_ (_13354_, _13353_, _13349_);
  and _64335_ (_13355_, _08376_, _08351_);
  or _64336_ (_13356_, _13355_, _13331_);
  and _64337_ (_13357_, _13356_, _06026_);
  or _64338_ (_13358_, _13357_, _09818_);
  or _64339_ (_13359_, _13358_, _13354_);
  and _64340_ (_13360_, _08485_, _07688_);
  or _64341_ (_13361_, _13312_, _07012_);
  or _64342_ (_13362_, _13361_, _13360_);
  or _64343_ (_13363_, _13338_, _09827_);
  and _64344_ (_13364_, _13363_, _05669_);
  and _64345_ (_13365_, _13364_, _13362_);
  and _64346_ (_13366_, _13365_, _13359_);
  and _64347_ (_13367_, _08738_, _07688_);
  or _64348_ (_13368_, _13367_, _13312_);
  and _64349_ (_13369_, _13368_, _09833_);
  or _64350_ (_13370_, _13369_, _06019_);
  or _64351_ (_13371_, _13370_, _13366_);
  and _64352_ (_13372_, _13371_, _13318_);
  or _64353_ (_13373_, _13372_, _06112_);
  and _64354_ (_13374_, _08760_, _07688_);
  or _64355_ (_13375_, _13374_, _13312_);
  or _64356_ (_13376_, _13375_, _08751_);
  and _64357_ (_13377_, _13376_, _08756_);
  and _64358_ (_13378_, _13377_, _13373_);
  or _64359_ (_13379_, _13378_, _13315_);
  and _64360_ (_13380_, _13379_, _07032_);
  or _64361_ (_13381_, _13312_, _07788_);
  and _64362_ (_13382_, _13317_, _06108_);
  and _64363_ (_13383_, _13382_, _13381_);
  or _64364_ (_13384_, _13383_, _13380_);
  and _64365_ (_13385_, _13384_, _06278_);
  and _64366_ (_13386_, _13323_, _06277_);
  and _64367_ (_13387_, _13386_, _13381_);
  or _64368_ (_13388_, _13387_, _06130_);
  or _64369_ (_13389_, _13388_, _13385_);
  and _64370_ (_13390_, _08759_, _07688_);
  or _64371_ (_13391_, _13312_, _08777_);
  or _64372_ (_13392_, _13391_, _13390_);
  and _64373_ (_13393_, _13392_, _08782_);
  and _64374_ (_13394_, _13393_, _13389_);
  nor _64375_ (_13395_, _08767_, _13311_);
  or _64376_ (_13396_, _13395_, _13312_);
  and _64377_ (_13397_, _13396_, _06292_);
  or _64378_ (_13398_, _13397_, _06316_);
  or _64379_ (_13399_, _13398_, _13394_);
  or _64380_ (_13400_, _13320_, _06718_);
  and _64381_ (_13401_, _13400_, _05653_);
  and _64382_ (_13402_, _13401_, _13399_);
  and _64383_ (_13403_, _13346_, _05652_);
  or _64384_ (_13404_, _13403_, _06047_);
  or _64385_ (_13405_, _13404_, _13402_);
  and _64386_ (_13406_, _08279_, _07688_);
  or _64387_ (_13407_, _13312_, _06048_);
  or _64388_ (_13408_, _13407_, _13406_);
  and _64389_ (_13409_, _13408_, _01336_);
  and _64390_ (_13410_, _13409_, _13405_);
  or _64391_ (_13411_, _13410_, _13310_);
  and _64392_ (_40774_, _13411_, _42882_);
  and _64393_ (_13412_, _01340_, \oc8051_golden_model_1.SCON [7]);
  not _64394_ (_13413_, _07679_);
  and _64395_ (_13414_, _13413_, \oc8051_golden_model_1.SCON [7]);
  and _64396_ (_13415_, _08768_, _07679_);
  or _64397_ (_13416_, _13415_, _13414_);
  and _64398_ (_13417_, _13416_, _06284_);
  and _64399_ (_13418_, _08549_, _07679_);
  or _64400_ (_13419_, _13418_, _13414_);
  or _64401_ (_13420_, _13419_, _06020_);
  and _64402_ (_13421_, _08498_, _07679_);
  or _64403_ (_13422_, _13421_, _13414_);
  or _64404_ (_13423_, _13422_, _06954_);
  and _64405_ (_13424_, _07679_, \oc8051_golden_model_1.ACC [7]);
  or _64406_ (_13425_, _13424_, _13414_);
  and _64407_ (_13426_, _13425_, _06938_);
  and _64408_ (_13427_, _06939_, \oc8051_golden_model_1.SCON [7]);
  or _64409_ (_13428_, _13427_, _06102_);
  or _64410_ (_13429_, _13428_, _13426_);
  and _64411_ (_13430_, _13429_, _06044_);
  and _64412_ (_13431_, _13430_, _13423_);
  not _64413_ (_13432_, _08347_);
  and _64414_ (_13433_, _13432_, \oc8051_golden_model_1.SCON [7]);
  and _64415_ (_13434_, _08503_, _08347_);
  or _64416_ (_13435_, _13434_, _13433_);
  and _64417_ (_13436_, _13435_, _06043_);
  or _64418_ (_13437_, _13436_, _06239_);
  or _64419_ (_13438_, _13437_, _13431_);
  nor _64420_ (_13439_, _07785_, _13413_);
  or _64421_ (_13440_, _13439_, _13414_);
  or _64422_ (_13441_, _13440_, _06848_);
  and _64423_ (_13442_, _13441_, _13438_);
  or _64424_ (_13443_, _13442_, _06219_);
  or _64425_ (_13444_, _13425_, _06220_);
  and _64426_ (_13445_, _13444_, _06040_);
  and _64427_ (_13446_, _13445_, _13443_);
  and _64428_ (_13447_, _08374_, _08347_);
  or _64429_ (_13448_, _13447_, _13433_);
  and _64430_ (_13449_, _13448_, _06039_);
  or _64431_ (_13450_, _13449_, _06032_);
  or _64432_ (_13451_, _13450_, _13446_);
  or _64433_ (_13452_, _13433_, _08519_);
  and _64434_ (_13453_, _13452_, _13435_);
  or _64435_ (_13454_, _13453_, _06033_);
  and _64436_ (_13455_, _13454_, _06027_);
  and _64437_ (_13456_, _13455_, _13451_);
  and _64438_ (_13457_, _08376_, _08347_);
  or _64439_ (_13458_, _13457_, _13433_);
  and _64440_ (_13459_, _13458_, _06026_);
  or _64441_ (_13460_, _13459_, _09818_);
  or _64442_ (_13461_, _13460_, _13456_);
  and _64443_ (_13462_, _08485_, _07679_);
  or _64444_ (_13463_, _13414_, _07012_);
  or _64445_ (_13464_, _13463_, _13462_);
  or _64446_ (_13465_, _13440_, _09827_);
  and _64447_ (_13466_, _13465_, _05669_);
  and _64448_ (_13467_, _13466_, _13464_);
  and _64449_ (_13468_, _13467_, _13461_);
  and _64450_ (_13469_, _08738_, _07679_);
  or _64451_ (_13470_, _13469_, _13414_);
  and _64452_ (_13471_, _13470_, _09833_);
  or _64453_ (_13472_, _13471_, _06019_);
  or _64454_ (_13473_, _13472_, _13468_);
  and _64455_ (_13474_, _13473_, _13420_);
  or _64456_ (_13475_, _13474_, _06112_);
  and _64457_ (_13476_, _08760_, _07679_);
  or _64458_ (_13477_, _13476_, _13414_);
  or _64459_ (_13478_, _13477_, _08751_);
  and _64460_ (_13479_, _13478_, _08756_);
  and _64461_ (_13480_, _13479_, _13475_);
  or _64462_ (_13481_, _13480_, _13417_);
  and _64463_ (_13482_, _13481_, _07032_);
  or _64464_ (_13483_, _13414_, _07788_);
  and _64465_ (_13484_, _13419_, _06108_);
  and _64466_ (_13485_, _13484_, _13483_);
  or _64467_ (_13486_, _13485_, _13482_);
  and _64468_ (_13487_, _13486_, _06278_);
  and _64469_ (_13488_, _13425_, _06277_);
  and _64470_ (_13489_, _13488_, _13483_);
  or _64471_ (_13490_, _13489_, _06130_);
  or _64472_ (_13491_, _13490_, _13487_);
  and _64473_ (_13492_, _08759_, _07679_);
  or _64474_ (_13493_, _13414_, _08777_);
  or _64475_ (_13494_, _13493_, _13492_);
  and _64476_ (_13495_, _13494_, _08782_);
  and _64477_ (_13496_, _13495_, _13491_);
  nor _64478_ (_13497_, _08767_, _13413_);
  or _64479_ (_13498_, _13497_, _13414_);
  and _64480_ (_13499_, _13498_, _06292_);
  or _64481_ (_13500_, _13499_, _06316_);
  or _64482_ (_13501_, _13500_, _13496_);
  or _64483_ (_13502_, _13422_, _06718_);
  and _64484_ (_13503_, _13502_, _05653_);
  and _64485_ (_13504_, _13503_, _13501_);
  and _64486_ (_13505_, _13448_, _05652_);
  or _64487_ (_13506_, _13505_, _06047_);
  or _64488_ (_13507_, _13506_, _13504_);
  and _64489_ (_13508_, _08279_, _07679_);
  or _64490_ (_13509_, _13414_, _06048_);
  or _64491_ (_13510_, _13509_, _13508_);
  and _64492_ (_13511_, _13510_, _01336_);
  and _64493_ (_13512_, _13511_, _13507_);
  or _64494_ (_13513_, _13512_, _13412_);
  and _64495_ (_40775_, _13513_, _42882_);
  not _64496_ (_13514_, \oc8051_golden_model_1.SP [7]);
  nor _64497_ (_13515_, _01336_, _13514_);
  and _64498_ (_13516_, _07360_, \oc8051_golden_model_1.SP [4]);
  and _64499_ (_13517_, _13516_, \oc8051_golden_model_1.SP [5]);
  and _64500_ (_13518_, _13517_, \oc8051_golden_model_1.SP [6]);
  or _64501_ (_13519_, _13518_, \oc8051_golden_model_1.SP [7]);
  nand _64502_ (_13520_, _13518_, \oc8051_golden_model_1.SP [7]);
  and _64503_ (_13521_, _13520_, _13519_);
  or _64504_ (_13522_, _13521_, _07059_);
  nor _64505_ (_13523_, _07727_, _13514_);
  and _64506_ (_13524_, _08768_, _07727_);
  or _64507_ (_13525_, _13524_, _13523_);
  and _64508_ (_13526_, _13525_, _06284_);
  and _64509_ (_13527_, _13517_, \oc8051_golden_model_1.SP [0]);
  and _64510_ (_13528_, _13527_, \oc8051_golden_model_1.SP [6]);
  nor _64511_ (_13529_, _13528_, _13514_);
  and _64512_ (_13530_, _13528_, _13514_);
  or _64513_ (_13531_, _13530_, _13529_);
  and _64514_ (_13532_, _13531_, _06038_);
  and _64515_ (_13533_, _08498_, _07727_);
  or _64516_ (_13534_, _13533_, _13523_);
  or _64517_ (_13535_, _13534_, _06954_);
  and _64518_ (_13536_, _07833_, \oc8051_golden_model_1.ACC [7]);
  or _64519_ (_13537_, _13536_, _13523_);
  or _64520_ (_13538_, _13537_, _06939_);
  or _64521_ (_13539_, _06938_, \oc8051_golden_model_1.SP [7]);
  and _64522_ (_13540_, _13539_, _07233_);
  and _64523_ (_13541_, _13540_, _13538_);
  and _64524_ (_13542_, _13521_, _06943_);
  or _64525_ (_13543_, _13542_, _06102_);
  or _64526_ (_13544_, _13543_, _13541_);
  and _64527_ (_13545_, _13544_, _05690_);
  and _64528_ (_13546_, _13545_, _13535_);
  and _64529_ (_13547_, _13521_, _07272_);
  or _64530_ (_13548_, _13547_, _06239_);
  or _64531_ (_13549_, _13548_, _13546_);
  not _64532_ (_13550_, \oc8051_golden_model_1.SP [6]);
  not _64533_ (_13551_, \oc8051_golden_model_1.SP [5]);
  not _64534_ (_13552_, \oc8051_golden_model_1.SP [4]);
  and _64535_ (_13553_, _08403_, _13552_);
  and _64536_ (_13554_, _13553_, _13551_);
  and _64537_ (_13555_, _13554_, _13550_);
  and _64538_ (_13556_, _13555_, _06029_);
  nor _64539_ (_13557_, _13556_, _13514_);
  and _64540_ (_13558_, _13556_, _13514_);
  nor _64541_ (_13559_, _13558_, _13557_);
  nand _64542_ (_13560_, _13559_, _06239_);
  and _64543_ (_13561_, _13560_, _13549_);
  or _64544_ (_13562_, _13561_, _06219_);
  or _64545_ (_13563_, _13537_, _06220_);
  and _64546_ (_13564_, _13563_, _07364_);
  and _64547_ (_13565_, _13564_, _13562_);
  or _64548_ (_13566_, _13565_, _13532_);
  and _64549_ (_13567_, _13566_, _07271_);
  not _64550_ (_13568_, _07271_);
  and _64551_ (_13569_, _13521_, _13568_);
  or _64552_ (_13570_, _13569_, _09818_);
  or _64553_ (_13571_, _13570_, _13567_);
  or _64554_ (_13572_, _13523_, _07012_);
  and _64555_ (_13573_, _08485_, _07833_);
  or _64556_ (_13574_, _13573_, _13572_);
  not _64557_ (_13575_, _07727_);
  nor _64558_ (_13576_, _07785_, _13575_);
  or _64559_ (_13577_, _13523_, _09827_);
  or _64560_ (_13578_, _13577_, _13576_);
  and _64561_ (_13579_, _13578_, _05669_);
  and _64562_ (_13580_, _13579_, _13574_);
  and _64563_ (_13581_, _13580_, _13571_);
  and _64564_ (_13582_, _08738_, _07727_);
  or _64565_ (_13583_, _13582_, _13523_);
  and _64566_ (_13584_, _13583_, _09833_);
  or _64567_ (_13585_, _13584_, _06019_);
  or _64568_ (_13586_, _13585_, _13581_);
  not _64569_ (_13587_, _05724_);
  and _64570_ (_13588_, _08549_, _07833_);
  or _64571_ (_13589_, _13588_, _13523_);
  or _64572_ (_13590_, _13589_, _06020_);
  and _64573_ (_13591_, _13590_, _13587_);
  and _64574_ (_13592_, _13591_, _13586_);
  and _64575_ (_13593_, _13521_, _05724_);
  or _64576_ (_13594_, _13593_, _06112_);
  or _64577_ (_13595_, _13594_, _13592_);
  and _64578_ (_13596_, _08760_, _07833_);
  or _64579_ (_13597_, _13596_, _13523_);
  or _64580_ (_13598_, _13597_, _08751_);
  and _64581_ (_13599_, _13598_, _08756_);
  and _64582_ (_13600_, _13599_, _13595_);
  or _64583_ (_13601_, _13600_, _13526_);
  and _64584_ (_13602_, _13601_, _07032_);
  or _64585_ (_13603_, _13523_, _07788_);
  and _64586_ (_13604_, _13589_, _06108_);
  and _64587_ (_13605_, _13604_, _13603_);
  or _64588_ (_13606_, _13605_, _13602_);
  and _64589_ (_13607_, _13606_, _12494_);
  and _64590_ (_13608_, _13521_, _05736_);
  or _64591_ (_13609_, _13608_, _06130_);
  and _64592_ (_13610_, _13537_, _06277_);
  and _64593_ (_13611_, _13610_, _13603_);
  or _64594_ (_13612_, _13611_, _13609_);
  or _64595_ (_13613_, _13612_, _13607_);
  and _64596_ (_13614_, _08759_, _07727_);
  or _64597_ (_13615_, _13523_, _08777_);
  or _64598_ (_13616_, _13615_, _13614_);
  and _64599_ (_13617_, _13616_, _13613_);
  or _64600_ (_13618_, _13617_, _06292_);
  not _64601_ (_13619_, _06298_);
  nor _64602_ (_13620_, _08767_, _13575_);
  or _64603_ (_13621_, _13523_, _08782_);
  or _64604_ (_13622_, _13621_, _13620_);
  and _64605_ (_13623_, _13622_, _13619_);
  and _64606_ (_13624_, _13623_, _13618_);
  or _64607_ (_13625_, _13555_, \oc8051_golden_model_1.SP [7]);
  nand _64608_ (_13626_, _13555_, \oc8051_golden_model_1.SP [7]);
  and _64609_ (_13627_, _13626_, _13625_);
  and _64610_ (_13628_, _13627_, _06298_);
  or _64611_ (_13629_, _13628_, _05732_);
  or _64612_ (_13630_, _13629_, _13624_);
  or _64613_ (_13631_, _13521_, _05734_);
  and _64614_ (_13632_, _13631_, _13630_);
  or _64615_ (_13633_, _13632_, _06049_);
  or _64616_ (_13634_, _13627_, _06050_);
  and _64617_ (_13635_, _13634_, _06718_);
  and _64618_ (_13636_, _13635_, _13633_);
  and _64619_ (_13637_, _13534_, _06316_);
  or _64620_ (_13638_, _13637_, _07458_);
  or _64621_ (_13639_, _13638_, _13636_);
  and _64622_ (_13640_, _13639_, _13522_);
  or _64623_ (_13641_, _13640_, _06047_);
  and _64624_ (_13642_, _08279_, _07727_);
  or _64625_ (_13643_, _13523_, _06048_);
  or _64626_ (_13644_, _13643_, _13642_);
  and _64627_ (_13645_, _13644_, _01336_);
  and _64628_ (_13646_, _13645_, _13641_);
  or _64629_ (_13648_, _13646_, _13515_);
  and _64630_ (_40776_, _13648_, _42882_);
  and _64631_ (_13649_, _01340_, \oc8051_golden_model_1.SBUF [7]);
  not _64632_ (_13650_, _07681_);
  and _64633_ (_13651_, _13650_, \oc8051_golden_model_1.SBUF [7]);
  nor _64634_ (_13652_, _08767_, _13650_);
  or _64635_ (_13653_, _13652_, _13651_);
  and _64636_ (_13654_, _13653_, _06292_);
  or _64637_ (_13655_, _13651_, _07788_);
  and _64638_ (_13656_, _08549_, _07681_);
  or _64639_ (_13658_, _13656_, _13651_);
  and _64640_ (_13659_, _13658_, _06108_);
  and _64641_ (_13660_, _13659_, _13655_);
  and _64642_ (_13661_, _08768_, _07681_);
  or _64643_ (_13662_, _13661_, _13651_);
  and _64644_ (_13663_, _13662_, _06284_);
  or _64645_ (_13664_, _13658_, _06020_);
  and _64646_ (_13665_, _08498_, _07681_);
  or _64647_ (_13666_, _13665_, _13651_);
  or _64648_ (_13667_, _13666_, _06954_);
  and _64649_ (_13669_, _07681_, \oc8051_golden_model_1.ACC [7]);
  or _64650_ (_13670_, _13669_, _13651_);
  and _64651_ (_13671_, _13670_, _06938_);
  and _64652_ (_13672_, _06939_, \oc8051_golden_model_1.SBUF [7]);
  or _64653_ (_13673_, _13672_, _06102_);
  or _64654_ (_13674_, _13673_, _13671_);
  and _64655_ (_13675_, _13674_, _06848_);
  and _64656_ (_13676_, _13675_, _13667_);
  nor _64657_ (_13677_, _07785_, _13650_);
  or _64658_ (_13678_, _13677_, _13651_);
  and _64659_ (_13680_, _13678_, _06239_);
  or _64660_ (_13681_, _13680_, _13676_);
  and _64661_ (_13682_, _13681_, _06220_);
  and _64662_ (_13683_, _13670_, _06219_);
  or _64663_ (_13684_, _13683_, _09818_);
  or _64664_ (_13685_, _13684_, _13682_);
  and _64665_ (_13686_, _08485_, _07681_);
  or _64666_ (_13687_, _13651_, _07012_);
  or _64667_ (_13688_, _13687_, _13686_);
  or _64668_ (_13689_, _13678_, _09827_);
  and _64669_ (_13691_, _13689_, _05669_);
  and _64670_ (_13692_, _13691_, _13688_);
  and _64671_ (_13693_, _13692_, _13685_);
  and _64672_ (_13694_, _08738_, _07681_);
  or _64673_ (_13695_, _13694_, _13651_);
  and _64674_ (_13696_, _13695_, _09833_);
  or _64675_ (_13697_, _13696_, _06019_);
  or _64676_ (_13698_, _13697_, _13693_);
  and _64677_ (_13699_, _13698_, _13664_);
  or _64678_ (_13700_, _13699_, _06112_);
  and _64679_ (_13702_, _08760_, _07681_);
  or _64680_ (_13703_, _13651_, _08751_);
  or _64681_ (_13704_, _13703_, _13702_);
  and _64682_ (_13705_, _13704_, _08756_);
  and _64683_ (_13706_, _13705_, _13700_);
  or _64684_ (_13707_, _13706_, _13663_);
  and _64685_ (_13708_, _13707_, _07032_);
  or _64686_ (_13709_, _13708_, _13660_);
  and _64687_ (_13710_, _13709_, _06278_);
  and _64688_ (_13711_, _13670_, _06277_);
  and _64689_ (_13713_, _13711_, _13655_);
  or _64690_ (_13714_, _13713_, _06130_);
  or _64691_ (_13715_, _13714_, _13710_);
  and _64692_ (_13716_, _08759_, _07681_);
  or _64693_ (_13717_, _13651_, _08777_);
  or _64694_ (_13718_, _13717_, _13716_);
  and _64695_ (_13719_, _13718_, _08782_);
  and _64696_ (_13720_, _13719_, _13715_);
  or _64697_ (_13721_, _13720_, _13654_);
  and _64698_ (_13722_, _13721_, _06718_);
  and _64699_ (_13724_, _13666_, _06316_);
  or _64700_ (_13725_, _13724_, _06047_);
  or _64701_ (_13726_, _13725_, _13722_);
  and _64702_ (_13727_, _08279_, _07681_);
  or _64703_ (_13728_, _13651_, _06048_);
  or _64704_ (_13729_, _13728_, _13727_);
  and _64705_ (_13730_, _13729_, _01336_);
  and _64706_ (_13731_, _13730_, _13726_);
  or _64707_ (_13732_, _13731_, _13649_);
  and _64708_ (_40777_, _13732_, _42882_);
  nor _64709_ (_13734_, _01336_, _10606_);
  nor _64710_ (_13735_, _08355_, _10606_);
  and _64711_ (_13736_, _08374_, _08355_);
  or _64712_ (_13737_, _13736_, _13735_);
  or _64713_ (_13738_, _13737_, _05653_);
  not _64714_ (_13739_, _10704_);
  or _64715_ (_13740_, _11048_, _10703_);
  and _64716_ (_13741_, _13740_, _10974_);
  nand _64717_ (_13742_, _13741_, _13739_);
  nor _64718_ (_13743_, _07705_, _10606_);
  not _64719_ (_13745_, _07705_);
  nor _64720_ (_13746_, _08767_, _13745_);
  or _64721_ (_13747_, _13746_, _13743_);
  and _64722_ (_13748_, _13747_, _06292_);
  and _64723_ (_13749_, _08768_, _07705_);
  or _64724_ (_13750_, _13749_, _13743_);
  and _64725_ (_13751_, _13750_, _06284_);
  and _64726_ (_13752_, _08738_, _07705_);
  or _64727_ (_13753_, _13752_, _13743_);
  and _64728_ (_13754_, _13753_, _09833_);
  and _64729_ (_13756_, _10314_, _07788_);
  and _64730_ (_13757_, _10324_, _10320_);
  nor _64731_ (_13758_, _13757_, _10318_);
  nand _64732_ (_13759_, _10367_, _10320_);
  or _64733_ (_13760_, _13759_, _10365_);
  and _64734_ (_13761_, _13760_, _13758_);
  or _64735_ (_13762_, _13761_, _13756_);
  and _64736_ (_13763_, _13762_, _06261_);
  not _64737_ (_13764_, _06250_);
  not _64738_ (_13765_, _06251_);
  nor _64739_ (_13767_, _12722_, _13765_);
  nand _64740_ (_13768_, _07979_, \oc8051_golden_model_1.ACC [5]);
  nor _64741_ (_13769_, _07979_, \oc8051_golden_model_1.ACC [5]);
  nor _64742_ (_13770_, _08272_, \oc8051_golden_model_1.ACC [4]);
  or _64743_ (_13771_, _13770_, _13769_);
  and _64744_ (_13772_, _13771_, _13768_);
  and _64745_ (_13773_, _13772_, _12308_);
  nor _64746_ (_13774_, _07787_, \oc8051_golden_model_1.ACC [7]);
  or _64747_ (_13775_, _07885_, \oc8051_golden_model_1.ACC [6]);
  nor _64748_ (_13776_, _13775_, _08768_);
  or _64749_ (_13778_, _13776_, _13774_);
  or _64750_ (_13779_, _13778_, _13773_);
  nand _64751_ (_13780_, _08028_, \oc8051_golden_model_1.ACC [3]);
  nor _64752_ (_13781_, _08028_, \oc8051_golden_model_1.ACC [3]);
  nor _64753_ (_13782_, _08176_, \oc8051_golden_model_1.ACC [2]);
  or _64754_ (_13783_, _13782_, _13781_);
  and _64755_ (_13784_, _13783_, _13780_);
  nor _64756_ (_13785_, _08077_, \oc8051_golden_model_1.ACC [1]);
  nor _64757_ (_13786_, _08127_, _05758_);
  nor _64758_ (_13787_, _13786_, _10994_);
  or _64759_ (_13789_, _13787_, _13785_);
  and _64760_ (_13790_, _13789_, _12300_);
  or _64761_ (_13791_, _13790_, _13784_);
  and _64762_ (_13792_, _13791_, _12309_);
  or _64763_ (_13793_, _13792_, _13779_);
  nor _64764_ (_13794_, _12310_, _06509_);
  and _64765_ (_13795_, _13794_, _13793_);
  and _64766_ (_13796_, _08498_, _07705_);
  or _64767_ (_13797_, _13796_, _13743_);
  or _64768_ (_13798_, _13797_, _06954_);
  and _64769_ (_13799_, _07705_, \oc8051_golden_model_1.ACC [7]);
  or _64770_ (_13800_, _13799_, _13743_);
  and _64771_ (_13801_, _13800_, _06938_);
  nor _64772_ (_13802_, _06938_, _10606_);
  or _64773_ (_13803_, _13802_, _06102_);
  or _64774_ (_13804_, _13803_, _13801_);
  and _64775_ (_13805_, _13804_, _10413_);
  and _64776_ (_13806_, _13805_, _13798_);
  nor _64777_ (_13807_, _10431_, _10413_);
  not _64778_ (_13808_, _12181_);
  nand _64779_ (_13809_, _13808_, _06244_);
  or _64780_ (_13810_, _13809_, _13807_);
  or _64781_ (_13811_, _13810_, _13806_);
  and _64782_ (_13812_, _08503_, _08355_);
  or _64783_ (_13813_, _13812_, _13735_);
  or _64784_ (_13814_, _13813_, _06044_);
  nor _64785_ (_13815_, _07785_, _13745_);
  or _64786_ (_13816_, _13815_, _13743_);
  or _64787_ (_13817_, _13816_, _06848_);
  and _64788_ (_13818_, _13817_, _13814_);
  and _64789_ (_13819_, _13818_, _13811_);
  or _64790_ (_13820_, _13819_, _06219_);
  or _64791_ (_13821_, _13800_, _06220_);
  nor _64792_ (_13822_, _12238_, _06039_);
  and _64793_ (_13823_, _13822_, _13821_);
  and _64794_ (_13824_, _13823_, _13820_);
  and _64795_ (_13825_, _13737_, _06039_);
  or _64796_ (_13826_, _13825_, _12256_);
  or _64797_ (_13827_, _13826_, _13824_);
  not _64798_ (_13828_, _12289_);
  nor _64799_ (_13829_, _12284_, _12281_);
  or _64800_ (_13830_, _12282_, _13829_);
  and _64801_ (_13831_, _13830_, _12280_);
  nor _64802_ (_13832_, _12277_, _12274_);
  nor _64803_ (_13833_, _12275_, _13832_);
  or _64804_ (_13834_, _13833_, _13831_);
  and _64805_ (_13835_, _13834_, _12273_);
  and _64806_ (_13836_, _12268_, _12269_);
  or _64807_ (_13837_, _13836_, _12267_);
  and _64808_ (_13838_, _13837_, _12265_);
  and _64809_ (_13839_, _12263_, _07786_);
  or _64810_ (_13840_, _13839_, _12260_);
  or _64811_ (_13841_, _13840_, _13838_);
  or _64812_ (_13842_, _13841_, _13835_);
  and _64813_ (_13843_, _13842_, _13828_);
  or _64814_ (_13844_, _13843_, _12255_);
  and _64815_ (_13845_, _13844_, _12258_);
  and _64816_ (_13846_, _13845_, _13827_);
  and _64817_ (_13847_, _06513_, _06031_);
  and _64818_ (_13848_, _10394_, _06031_);
  nor _64819_ (_13849_, _13848_, _13847_);
  not _64820_ (_13850_, _13849_);
  not _64821_ (_13851_, _12145_);
  nand _64822_ (_13852_, _12143_, _13851_);
  nand _64823_ (_13853_, _13852_, _12142_);
  not _64824_ (_13854_, _12152_);
  or _64825_ (_13855_, _12154_, _13854_);
  and _64826_ (_13856_, _13855_, _12148_);
  or _64827_ (_13857_, _13856_, _13853_);
  and _64828_ (_13858_, _13857_, _12170_);
  nand _64829_ (_13859_, _12166_, _12163_);
  and _64830_ (_13860_, _12164_, _13859_);
  and _64831_ (_13861_, _13860_, _12162_);
  not _64832_ (_13862_, _12157_);
  and _64833_ (_13863_, _12159_, _13862_);
  nor _64834_ (_13864_, _13863_, _08531_);
  or _64835_ (_13865_, _13864_, _13861_);
  or _64836_ (_13866_, _13865_, _13858_);
  and _64837_ (_13867_, _13866_, _12174_);
  and _64838_ (_13868_, _13867_, _13850_);
  or _64839_ (_13869_, _13868_, _13846_);
  and _64840_ (_13870_, _13869_, _06509_);
  or _64841_ (_13871_, _13870_, _13795_);
  and _64842_ (_13872_, _13871_, _12298_);
  nor _64843_ (_13873_, _06799_, \oc8051_golden_model_1.ACC [1]);
  and _64844_ (_13874_, _06799_, \oc8051_golden_model_1.ACC [1]);
  and _64845_ (_13875_, _06016_, \oc8051_golden_model_1.ACC [0]);
  nor _64846_ (_13876_, _13875_, _13874_);
  or _64847_ (_13877_, _13876_, _13873_);
  and _64848_ (_13878_, _13877_, _12320_);
  nand _64849_ (_13879_, _05983_, \oc8051_golden_model_1.ACC [3]);
  nor _64850_ (_13880_, _05983_, \oc8051_golden_model_1.ACC [3]);
  nor _64851_ (_13881_, _06403_, \oc8051_golden_model_1.ACC [2]);
  or _64852_ (_13882_, _13881_, _13880_);
  and _64853_ (_13883_, _13882_, _13879_);
  or _64854_ (_13884_, _13883_, _13878_);
  and _64855_ (_13885_, _13884_, _12328_);
  nand _64856_ (_13886_, _06359_, \oc8051_golden_model_1.ACC [5]);
  nor _64857_ (_13887_, _06359_, \oc8051_golden_model_1.ACC [5]);
  nor _64858_ (_13888_, _06758_, \oc8051_golden_model_1.ACC [4]);
  or _64859_ (_13889_, _13888_, _13887_);
  and _64860_ (_13890_, _13889_, _13886_);
  and _64861_ (_13891_, _13890_, _12327_);
  and _64862_ (_13892_, _05952_, _08393_);
  or _64863_ (_13893_, _06084_, \oc8051_golden_model_1.ACC [6]);
  nor _64864_ (_13894_, _13893_, _10705_);
  or _64865_ (_13895_, _13894_, _13892_);
  or _64866_ (_13896_, _13895_, _13891_);
  or _64867_ (_13897_, _13896_, _13885_);
  nor _64868_ (_13898_, _12329_, _12298_);
  and _64869_ (_13899_, _13898_, _13897_);
  or _64870_ (_13900_, _13899_, _12012_);
  or _64871_ (_13901_, _13900_, _13872_);
  nand _64872_ (_13902_, _12012_, \oc8051_golden_model_1.PSW [7]);
  and _64873_ (_13903_, _13902_, _06033_);
  and _64874_ (_13904_, _13903_, _13901_);
  and _64875_ (_13905_, _08520_, _08355_);
  or _64876_ (_13906_, _13905_, _13735_);
  and _64877_ (_13907_, _13906_, _06032_);
  nor _64878_ (_13908_, _13907_, _13904_);
  nor _64879_ (_13909_, _13908_, _06253_);
  and _64880_ (_13910_, _06253_, \oc8051_golden_model_1.PSW [7]);
  and _64881_ (_13911_, _13910_, _12722_);
  or _64882_ (_13912_, _13911_, _13909_);
  nor _64883_ (_13913_, _09269_, _06251_);
  and _64884_ (_13914_, _13913_, _13912_);
  or _64885_ (_13915_, _13914_, _13767_);
  and _64886_ (_13916_, _13915_, _13764_);
  or _64887_ (_13917_, _12722_, \oc8051_golden_model_1.PSW [7]);
  and _64888_ (_13918_, _13917_, _06250_);
  or _64889_ (_13919_, _13918_, _10468_);
  or _64890_ (_13920_, _13919_, _13916_);
  and _64891_ (_13921_, _10250_, _10246_);
  nor _64892_ (_13922_, _13921_, _10244_);
  nand _64893_ (_13923_, _10252_, _10246_);
  or _64894_ (_13924_, _13923_, _10485_);
  and _64895_ (_13925_, _13924_, _13922_);
  or _64896_ (_13926_, _10469_, _10241_);
  or _64897_ (_13927_, _13926_, _13925_);
  and _64898_ (_13928_, _13927_, _13920_);
  or _64899_ (_13929_, _13928_, _12361_);
  and _64900_ (_13930_, _10506_, _10501_);
  nor _64901_ (_13931_, _13930_, _10499_);
  nand _64902_ (_13932_, _10553_, _10501_);
  or _64903_ (_13933_, _13932_, _10551_);
  and _64904_ (_13934_, _13933_, _13931_);
  not _64905_ (_13935_, _12361_);
  and _64906_ (_13936_, _10495_, _08485_);
  or _64907_ (_13937_, _13936_, _13935_);
  or _64908_ (_13938_, _13937_, _13934_);
  and _64909_ (_13939_, _13938_, _06267_);
  and _64910_ (_13940_, _13939_, _13929_);
  or _64911_ (_13941_, _13940_, _13763_);
  and _64912_ (_13942_, _13941_, _10307_);
  and _64913_ (_13943_, _10578_, _10575_);
  nor _64914_ (_13944_, _13943_, _10573_);
  nand _64915_ (_13945_, _10625_, _10575_);
  or _64916_ (_13946_, _13945_, _10623_);
  and _64917_ (_13947_, _13946_, _13944_);
  or _64918_ (_13948_, _13947_, _10568_);
  and _64919_ (_13949_, _13948_, _10306_);
  or _64920_ (_13950_, _13949_, _09818_);
  or _64921_ (_13951_, _13950_, _13942_);
  and _64922_ (_13952_, _08485_, _07705_);
  or _64923_ (_13953_, _13743_, _07012_);
  or _64924_ (_13954_, _13953_, _13952_);
  or _64925_ (_13955_, _13816_, _09827_);
  and _64926_ (_13956_, _13955_, _05669_);
  and _64927_ (_13957_, _13956_, _13954_);
  and _64928_ (_13958_, _13957_, _13951_);
  or _64929_ (_13959_, _13958_, _13754_);
  nor _64930_ (_13960_, _09832_, _06089_);
  and _64931_ (_13961_, _13960_, _13959_);
  nor _64932_ (_13962_, _12722_, _10606_);
  and _64933_ (_13963_, _13962_, _06089_);
  or _64934_ (_13964_, _13963_, _06019_);
  or _64935_ (_13965_, _13964_, _13961_);
  and _64936_ (_13966_, _08549_, _07705_);
  or _64937_ (_13967_, _13966_, _13743_);
  or _64938_ (_13968_, _13967_, _06020_);
  and _64939_ (_13969_, _13968_, _13965_);
  or _64940_ (_13970_, _13969_, _06088_);
  nand _64941_ (_13971_, _12722_, _10606_);
  or _64942_ (_13972_, _13971_, _06636_);
  and _64943_ (_13973_, _13972_, _13970_);
  or _64944_ (_13974_, _13973_, _06112_);
  and _64945_ (_13975_, _08760_, _07705_);
  or _64946_ (_13976_, _13975_, _13743_);
  or _64947_ (_13977_, _13976_, _08751_);
  and _64948_ (_13978_, _13977_, _08756_);
  and _64949_ (_13979_, _13978_, _13974_);
  or _64950_ (_13980_, _13979_, _13751_);
  and _64951_ (_13981_, _13980_, _07032_);
  or _64952_ (_13982_, _13743_, _07788_);
  and _64953_ (_13983_, _13967_, _06108_);
  and _64954_ (_13984_, _13983_, _13982_);
  or _64955_ (_13985_, _13984_, _13981_);
  and _64956_ (_13986_, _13985_, _06278_);
  and _64957_ (_13987_, _13800_, _06277_);
  and _64958_ (_13988_, _13987_, _13982_);
  or _64959_ (_13989_, _13988_, _06130_);
  or _64960_ (_13990_, _13989_, _13986_);
  and _64961_ (_13991_, _08759_, _07705_);
  or _64962_ (_13992_, _13743_, _08777_);
  or _64963_ (_13993_, _13992_, _13991_);
  and _64964_ (_13994_, _13993_, _08782_);
  and _64965_ (_13995_, _13994_, _13990_);
  or _64966_ (_13996_, _13995_, _13748_);
  and _64967_ (_13997_, _13996_, _10304_);
  nor _64968_ (_13998_, _10243_, _08393_);
  or _64969_ (_13999_, _13998_, _10300_);
  or _64970_ (_14000_, _13999_, _10241_);
  and _64971_ (_14001_, _14000_, _10303_);
  or _64972_ (_14002_, _14001_, _10794_);
  or _64973_ (_14003_, _14002_, _13997_);
  or _64974_ (_14004_, _10796_, _13936_);
  nor _64975_ (_14005_, _10498_, _08393_);
  or _64976_ (_14006_, _14005_, _10818_);
  or _64977_ (_14007_, _14006_, _14004_);
  and _64978_ (_14008_, _14007_, _06289_);
  and _64979_ (_14009_, _14008_, _14003_);
  nor _64980_ (_14010_, _10317_, _08393_);
  or _64981_ (_14011_, _14010_, _10848_);
  or _64982_ (_14012_, _10824_, _13756_);
  or _64983_ (_14013_, _14012_, _14011_);
  and _64984_ (_14014_, _14013_, _10826_);
  or _64985_ (_14015_, _14014_, _14009_);
  and _64986_ (_14016_, _10572_, \oc8051_golden_model_1.ACC [7]);
  or _64987_ (_14017_, _14016_, _10878_);
  or _64988_ (_14018_, _10856_, _10568_);
  or _64989_ (_14019_, _14018_, _14017_);
  and _64990_ (_14020_, _14019_, _10855_);
  and _64991_ (_14021_, _14020_, _14015_);
  nand _64992_ (_14022_, _10885_, _06545_);
  and _64993_ (_14023_, _14022_, _10889_);
  nand _64994_ (_14024_, _10854_, \oc8051_golden_model_1.ACC [7]);
  nand _64995_ (_14025_, _14024_, _14023_);
  or _64996_ (_14026_, _14025_, _14021_);
  or _64997_ (_14027_, _10926_, _10672_);
  nand _64998_ (_14028_, _14027_, _10719_);
  nor _64999_ (_14029_, _14028_, _14023_);
  nor _65000_ (_14030_, _14029_, _06693_);
  and _65001_ (_14031_, _14030_, _14026_);
  and _65002_ (_14032_, _14028_, _06693_);
  or _65003_ (_14033_, _14032_, _10932_);
  or _65004_ (_14034_, _14033_, _14031_);
  and _65005_ (_14035_, _10966_, _10693_);
  nor _65006_ (_14036_, _10935_, _10692_);
  nor _65007_ (_14037_, _14036_, _10691_);
  or _65008_ (_14038_, _14037_, _10934_);
  or _65009_ (_14039_, _14038_, _14035_);
  and _65010_ (_14040_, _14039_, _06052_);
  and _65011_ (_14041_, _14040_, _14034_);
  not _65012_ (_14042_, _08767_);
  not _65013_ (_14043_, _08766_);
  nand _65014_ (_14044_, _11008_, _14043_);
  and _65015_ (_14045_, _14044_, _06051_);
  and _65016_ (_14046_, _14045_, _14042_);
  or _65017_ (_14047_, _14046_, _10974_);
  or _65018_ (_14048_, _14047_, _14041_);
  and _65019_ (_14049_, _14048_, _13742_);
  or _65020_ (_14050_, _14049_, _06316_);
  nor _65021_ (_14051_, _13797_, _06718_);
  nor _65022_ (_14052_, _14051_, _11064_);
  and _65023_ (_14053_, _14052_, _14050_);
  and _65024_ (_14054_, _11064_, \oc8051_golden_model_1.ACC [0]);
  or _65025_ (_14055_, _14054_, _05652_);
  or _65026_ (_14056_, _14055_, _14053_);
  and _65027_ (_14057_, _14056_, _13738_);
  or _65028_ (_14058_, _14057_, _06047_);
  and _65029_ (_14059_, _08279_, _07705_);
  or _65030_ (_14060_, _13743_, _06048_);
  or _65031_ (_14061_, _14060_, _14059_);
  and _65032_ (_14062_, _14061_, _01336_);
  and _65033_ (_14063_, _14062_, _14058_);
  or _65034_ (_14064_, _14063_, _13734_);
  and _65035_ (_40778_, _14064_, _42882_);
  and _65036_ (_14065_, _12112_, _06127_);
  not _65037_ (_14066_, _11952_);
  nor _65038_ (_14067_, _14066_, _06127_);
  or _65039_ (_14068_, _14067_, _14065_);
  nor _65040_ (_14069_, _08403_, _07360_);
  not _65041_ (_14070_, _14069_);
  and _65042_ (_14071_, _14070_, _07628_);
  and _65043_ (_14072_, _14071_, _07081_);
  not _65044_ (_14073_, _14072_);
  or _65045_ (_14074_, _14073_, _14068_);
  nor _65046_ (_14075_, _07476_, _07305_);
  nor _65047_ (_14076_, _14075_, _07615_);
  nor _65048_ (_14077_, _07305_, _07074_);
  nor _65049_ (_14078_, _14077_, _07306_);
  and _65050_ (_14079_, _14078_, _07304_);
  and _65051_ (_14080_, _14079_, _14076_);
  nand _65052_ (_14081_, _06127_, \oc8051_golden_model_1.PC [0]);
  nand _65053_ (_14082_, _12302_, _08783_);
  or _65054_ (_14083_, _08127_, _08672_);
  and _65055_ (_14084_, _08127_, _08672_);
  not _65056_ (_14085_, _14084_);
  and _65057_ (_14086_, _14085_, _14083_);
  and _65058_ (_14087_, _14086_, _08752_);
  or _65059_ (_14088_, _07009_, _06931_);
  or _65060_ (_14089_, _08127_, _06233_);
  nor _65061_ (_14090_, _12615_, _12591_);
  or _65062_ (_14091_, _14090_, _08378_);
  nor _65063_ (_14092_, _08127_, _08381_);
  nand _65064_ (_14093_, _08384_, _06931_);
  nand _65065_ (_14094_, _06943_, _05346_);
  or _65066_ (_14095_, _06943_, \oc8051_golden_model_1.ACC [0]);
  and _65067_ (_14096_, _14095_, _14094_);
  nor _65068_ (_14097_, _14096_, _08384_);
  nor _65069_ (_14098_, _14097_, _06955_);
  and _65070_ (_14099_, _14098_, _14093_);
  or _65071_ (_14100_, _14099_, _14092_);
  and _65072_ (_14101_, _14100_, _08380_);
  nand _65073_ (_14102_, _12615_, _12592_);
  and _65074_ (_14103_, _14102_, _06953_);
  or _65075_ (_14104_, _14103_, _07272_);
  or _65076_ (_14105_, _14104_, _14101_);
  nor _65077_ (_14106_, _05690_, \oc8051_golden_model_1.PC [0]);
  nor _65078_ (_14107_, _14106_, _06963_);
  and _65079_ (_14108_, _14107_, _14105_);
  and _65080_ (_14109_, _06963_, _06931_);
  or _65081_ (_14110_, _14109_, _06975_);
  or _65082_ (_14111_, _14110_, _14108_);
  and _65083_ (_14112_, _14111_, _14091_);
  or _65084_ (_14113_, _14112_, _06038_);
  or _65085_ (_14114_, _08127_, _07364_);
  and _65086_ (_14115_, _14114_, _06036_);
  and _65087_ (_14116_, _14115_, _14113_);
  nor _65088_ (_14117_, _12616_, _06036_);
  and _65089_ (_14118_, _14117_, _14102_);
  or _65090_ (_14119_, _14118_, _14116_);
  and _65091_ (_14120_, _14119_, _05686_);
  or _65092_ (_14121_, _05686_, _05346_);
  nand _65093_ (_14122_, _06233_, _14121_);
  or _65094_ (_14123_, _14122_, _14120_);
  and _65095_ (_14124_, _14123_, _14089_);
  or _65096_ (_14125_, _14124_, _06992_);
  and _65097_ (_14126_, _09120_, _06053_);
  nand _65098_ (_14127_, _08124_, _06992_);
  or _65099_ (_14128_, _14127_, _14126_);
  and _65100_ (_14129_, _14128_, _14125_);
  or _65101_ (_14130_, _14129_, _06991_);
  nand _65102_ (_14131_, _12591_, _10606_);
  and _65103_ (_14132_, _14131_, _14102_);
  or _65104_ (_14133_, _14132_, _07308_);
  and _65105_ (_14134_, _14133_, _05673_);
  and _65106_ (_14135_, _14134_, _14130_);
  or _65107_ (_14136_, _05673_, _05346_);
  nand _65108_ (_14137_, _07009_, _14136_);
  or _65109_ (_14138_, _14137_, _14135_);
  and _65110_ (_14139_, _14138_, _14088_);
  or _65111_ (_14140_, _14139_, _07013_);
  or _65112_ (_14141_, _09120_, _07231_);
  and _65113_ (_14142_, _14141_, _08545_);
  and _65114_ (_14143_, _14142_, _14140_);
  and _65115_ (_14144_, _08332_, _06931_);
  and _65116_ (_14145_, _08668_, \oc8051_golden_model_1.SCON [0]);
  and _65117_ (_14146_, _08677_, \oc8051_golden_model_1.SBUF [0]);
  or _65118_ (_14147_, _14146_, _14145_);
  and _65119_ (_14148_, _08660_, \oc8051_golden_model_1.P0 [0]);
  and _65120_ (_14149_, _08682_, \oc8051_golden_model_1.P1 [0]);
  or _65121_ (_14150_, _14149_, _14148_);
  or _65122_ (_14151_, _14150_, _14147_);
  and _65123_ (_14152_, _08680_, \oc8051_golden_model_1.TCON [0]);
  and _65124_ (_14153_, _08654_, \oc8051_golden_model_1.ACC [0]);
  or _65125_ (_14154_, _14153_, _14152_);
  and _65126_ (_14155_, _08675_, \oc8051_golden_model_1.TMOD [0]);
  and _65127_ (_14156_, _08702_, \oc8051_golden_model_1.TL0 [0]);
  or _65128_ (_14157_, _14156_, _14155_);
  or _65129_ (_14158_, _14157_, _14154_);
  and _65130_ (_14159_, _08693_, \oc8051_golden_model_1.IE [0]);
  and _65131_ (_14160_, _08695_, \oc8051_golden_model_1.P3 [0]);
  or _65132_ (_14161_, _14160_, _14159_);
  and _65133_ (_14162_, _08687_, \oc8051_golden_model_1.P2 [0]);
  and _65134_ (_14163_, _08690_, \oc8051_golden_model_1.IP [0]);
  or _65135_ (_14164_, _14163_, _14162_);
  or _65136_ (_14165_, _14164_, _14161_);
  and _65137_ (_14166_, _08650_, \oc8051_golden_model_1.B [0]);
  and _65138_ (_14167_, _08704_, \oc8051_golden_model_1.PSW [0]);
  or _65139_ (_14168_, _14167_, _14166_);
  or _65140_ (_14169_, _14168_, _14165_);
  or _65141_ (_14170_, _14169_, _14158_);
  or _65142_ (_14171_, _14170_, _14151_);
  and _65143_ (_14172_, _08732_, \oc8051_golden_model_1.PCON [0]);
  and _65144_ (_14173_, _08725_, \oc8051_golden_model_1.TH1 [0]);
  and _65145_ (_14174_, _08712_, \oc8051_golden_model_1.TH0 [0]);
  or _65146_ (_14175_, _14174_, _14173_);
  or _65147_ (_14176_, _14175_, _14172_);
  and _65148_ (_14177_, _08716_, \oc8051_golden_model_1.TL1 [0]);
  and _65149_ (_14178_, _08723_, \oc8051_golden_model_1.DPH [0]);
  or _65150_ (_14179_, _14178_, _14177_);
  and _65151_ (_14180_, _08728_, \oc8051_golden_model_1.DPL [0]);
  and _65152_ (_14181_, _08719_, \oc8051_golden_model_1.SP [0]);
  or _65153_ (_14182_, _14181_, _14180_);
  or _65154_ (_14183_, _14182_, _14179_);
  or _65155_ (_14184_, _14183_, _14176_);
  or _65156_ (_14185_, _14184_, _14171_);
  or _65157_ (_14186_, _14185_, _14144_);
  and _65158_ (_14187_, _14186_, _07010_);
  or _65159_ (_14188_, _14187_, _08743_);
  or _65160_ (_14189_, _14188_, _14143_);
  and _65161_ (_14190_, _08743_, _06016_);
  nor _65162_ (_14191_, _14190_, _06021_);
  and _65163_ (_14192_, _14191_, _14189_);
  and _65164_ (_14193_, _08672_, _06021_);
  or _65165_ (_14194_, _14193_, _05724_);
  or _65166_ (_14195_, _14194_, _14192_);
  and _65167_ (_14196_, _05724_, _05346_);
  nor _65168_ (_14197_, _14196_, _08752_);
  and _65169_ (_14198_, _14197_, _14195_);
  or _65170_ (_14199_, _14198_, _14087_);
  and _65171_ (_14200_, _14199_, _08765_);
  nor _65172_ (_14201_, _12303_, _08765_);
  or _65173_ (_14202_, _14201_, _14200_);
  and _65174_ (_14203_, _14202_, _08764_);
  and _65175_ (_14204_, _14084_, _08301_);
  or _65176_ (_14205_, _14204_, _14203_);
  and _65177_ (_14206_, _14205_, _08300_);
  and _65178_ (_14207_, _10995_, _07031_);
  or _65179_ (_14208_, _14207_, _05736_);
  or _65180_ (_14209_, _14208_, _14206_);
  and _65181_ (_14210_, _05736_, _05346_);
  nor _65182_ (_14211_, _14210_, _08778_);
  and _65183_ (_14212_, _14211_, _14209_);
  and _65184_ (_14213_, _14083_, _08778_);
  or _65185_ (_14214_, _14213_, _08783_);
  or _65186_ (_14215_, _14214_, _14212_);
  and _65187_ (_14216_, _14215_, _14082_);
  or _65188_ (_14217_, _14216_, _05732_);
  nand _65189_ (_14218_, _05732_, _05346_);
  and _65190_ (_14219_, _14218_, _08287_);
  and _65191_ (_14220_, _14219_, _14217_);
  nand _65192_ (_14221_, _07052_, _06931_);
  and _65193_ (_14222_, _14221_, _12750_);
  or _65194_ (_14223_, _14222_, _14220_);
  nand _65195_ (_14224_, _09120_, _07051_);
  and _65196_ (_14225_, _14224_, _08797_);
  and _65197_ (_14226_, _14225_, _14223_);
  nor _65198_ (_14227_, _08127_, _08797_);
  or _65199_ (_14228_, _14227_, _06127_);
  or _65200_ (_14229_, _14228_, _14226_);
  and _65201_ (_14230_, _14229_, _14081_);
  or _65202_ (_14231_, _14230_, _05752_);
  and _65203_ (_14232_, _05752_, _05346_);
  nor _65204_ (_14233_, _14232_, _07058_);
  and _65205_ (_14234_, _14233_, _14231_);
  not _65206_ (_14235_, _09154_);
  and _65207_ (_14236_, _14090_, _07058_);
  or _65208_ (_14237_, _14236_, _14235_);
  or _65209_ (_14238_, _14237_, _14234_);
  nand _65210_ (_14239_, _14235_, _06931_);
  and _65211_ (_14240_, _14239_, _07069_);
  and _65212_ (_14241_, _14240_, _14238_);
  nor _65213_ (_14242_, _09120_, _07069_);
  or _65214_ (_14243_, _14242_, _07067_);
  or _65215_ (_14244_, _14243_, _14241_);
  nand _65216_ (_14245_, _08127_, _07067_);
  and _65217_ (_14246_, _14245_, _07304_);
  and _65218_ (_14247_, _14246_, _14244_);
  and _65219_ (_14248_, _14247_, _14080_);
  or _65220_ (_14249_, _14080_, _06505_);
  nand _65221_ (_14250_, _14249_, _14073_);
  or _65222_ (_14251_, _14250_, _14248_);
  and _65223_ (_40792_, _14251_, _14074_);
  or _65224_ (_14252_, _14080_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _65225_ (_14253_, _14252_, _14073_);
  not _65226_ (_14254_, _14080_);
  nor _65227_ (_14255_, _09162_, _08291_);
  and _65228_ (_14256_, _14255_, _14235_);
  nor _65229_ (_14257_, _14255_, _06866_);
  or _65230_ (_14258_, _14257_, _07210_);
  and _65231_ (_14259_, _05732_, _05312_);
  nand _65232_ (_14260_, _08077_, _06832_);
  nor _65233_ (_14261_, _08077_, _06832_);
  not _65234_ (_14262_, _14261_);
  and _65235_ (_14263_, _14262_, _14260_);
  and _65236_ (_14264_, _14263_, _08752_);
  nand _65237_ (_14265_, _07132_, _08541_);
  nand _65238_ (_14266_, _12588_, _12566_);
  nand _65239_ (_14267_, _07726_, _10606_);
  and _65240_ (_14268_, _14267_, _06991_);
  and _65241_ (_14269_, _14268_, _14266_);
  or _65242_ (_14270_, _12150_, _05952_);
  nand _65243_ (_14271_, _14270_, _08075_);
  and _65244_ (_14272_, _14271_, _06992_);
  nor _65245_ (_14273_, _12588_, _07726_);
  or _65246_ (_14274_, _14273_, _08378_);
  nand _65247_ (_14275_, _14255_, _08384_);
  and _65248_ (_14276_, _06943_, _05312_);
  and _65249_ (_14277_, _11988_, _06042_);
  nor _65250_ (_14278_, _06943_, _05784_);
  or _65251_ (_14279_, _14278_, _14277_);
  or _65252_ (_14280_, _14279_, _07139_);
  or _65253_ (_14281_, _14280_, _14276_);
  and _65254_ (_14282_, _14281_, _14275_);
  and _65255_ (_14283_, _14282_, _08381_);
  nor _65256_ (_14284_, _08491_, _08128_);
  nor _65257_ (_14285_, _14284_, _08381_);
  or _65258_ (_14286_, _14285_, _14283_);
  or _65259_ (_14287_, _14286_, _06953_);
  or _65260_ (_14288_, _14266_, _08380_);
  and _65261_ (_14289_, _14288_, _14287_);
  or _65262_ (_14290_, _14289_, _07272_);
  nor _65263_ (_14291_, _05690_, _05312_);
  nor _65264_ (_14292_, _14291_, _06963_);
  and _65265_ (_14293_, _14292_, _14290_);
  and _65266_ (_14294_, _09161_, _06963_);
  or _65267_ (_14295_, _14294_, _06975_);
  or _65268_ (_14296_, _14295_, _14293_);
  and _65269_ (_14297_, _14296_, _14274_);
  or _65270_ (_14298_, _14297_, _06038_);
  nand _65271_ (_14299_, _08077_, _06038_);
  and _65272_ (_14300_, _14299_, _06036_);
  and _65273_ (_14301_, _14300_, _14298_);
  not _65274_ (_14302_, _12589_);
  and _65275_ (_14303_, _14266_, _14302_);
  and _65276_ (_14304_, _14303_, _06035_);
  or _65277_ (_14305_, _14304_, _14301_);
  and _65278_ (_14306_, _14305_, _05686_);
  or _65279_ (_14307_, _05686_, \oc8051_golden_model_1.PC [1]);
  nand _65280_ (_14308_, _06233_, _14307_);
  or _65281_ (_14309_, _14308_, _14306_);
  nand _65282_ (_14310_, _08077_, _06573_);
  and _65283_ (_14311_, _14310_, _06993_);
  and _65284_ (_14312_, _14311_, _14309_);
  or _65285_ (_14313_, _14312_, _14272_);
  and _65286_ (_14314_, _14313_, _07308_);
  or _65287_ (_14315_, _14314_, _14269_);
  and _65288_ (_14316_, _14315_, _05673_);
  or _65289_ (_14317_, _05673_, \oc8051_golden_model_1.PC [1]);
  nand _65290_ (_14318_, _07009_, _14317_);
  or _65291_ (_14319_, _14318_, _14316_);
  and _65292_ (_14320_, _14319_, _14265_);
  or _65293_ (_14321_, _14320_, _07013_);
  or _65294_ (_14322_, _09075_, _07231_);
  and _65295_ (_14323_, _14322_, _08545_);
  and _65296_ (_14324_, _14323_, _14321_);
  nor _65297_ (_14325_, _08549_, _07132_);
  and _65298_ (_14326_, _08675_, \oc8051_golden_model_1.TMOD [1]);
  and _65299_ (_14327_, _08682_, \oc8051_golden_model_1.P1 [1]);
  or _65300_ (_14328_, _14327_, _14326_);
  and _65301_ (_14329_, _08702_, \oc8051_golden_model_1.TL0 [1]);
  and _65302_ (_14330_, _08650_, \oc8051_golden_model_1.B [1]);
  or _65303_ (_14331_, _14330_, _14329_);
  or _65304_ (_14332_, _14331_, _14328_);
  and _65305_ (_14333_, _08660_, \oc8051_golden_model_1.P0 [1]);
  and _65306_ (_14334_, _08680_, \oc8051_golden_model_1.TCON [1]);
  or _65307_ (_14335_, _14334_, _14333_);
  and _65308_ (_14336_, _08668_, \oc8051_golden_model_1.SCON [1]);
  and _65309_ (_14337_, _08704_, \oc8051_golden_model_1.PSW [1]);
  or _65310_ (_14338_, _14337_, _14336_);
  or _65311_ (_14339_, _14338_, _14335_);
  and _65312_ (_14340_, _08693_, \oc8051_golden_model_1.IE [1]);
  and _65313_ (_14341_, _08690_, \oc8051_golden_model_1.IP [1]);
  or _65314_ (_14342_, _14341_, _14340_);
  and _65315_ (_14343_, _08687_, \oc8051_golden_model_1.P2 [1]);
  and _65316_ (_14344_, _08695_, \oc8051_golden_model_1.P3 [1]);
  or _65317_ (_14345_, _14344_, _14343_);
  or _65318_ (_14346_, _14345_, _14342_);
  and _65319_ (_14347_, _08677_, \oc8051_golden_model_1.SBUF [1]);
  and _65320_ (_14348_, _08654_, \oc8051_golden_model_1.ACC [1]);
  or _65321_ (_14349_, _14348_, _14347_);
  or _65322_ (_14350_, _14349_, _14346_);
  or _65323_ (_14351_, _14350_, _14339_);
  or _65324_ (_14352_, _14351_, _14332_);
  and _65325_ (_14353_, _08716_, \oc8051_golden_model_1.TL1 [1]);
  and _65326_ (_14354_, _08732_, \oc8051_golden_model_1.PCON [1]);
  and _65327_ (_14355_, _08725_, \oc8051_golden_model_1.TH1 [1]);
  or _65328_ (_14356_, _14355_, _14354_);
  or _65329_ (_14357_, _14356_, _14353_);
  and _65330_ (_14358_, _08712_, \oc8051_golden_model_1.TH0 [1]);
  and _65331_ (_14359_, _08719_, \oc8051_golden_model_1.SP [1]);
  or _65332_ (_14360_, _14359_, _14358_);
  and _65333_ (_14361_, _08728_, \oc8051_golden_model_1.DPL [1]);
  and _65334_ (_14362_, _08723_, \oc8051_golden_model_1.DPH [1]);
  or _65335_ (_14363_, _14362_, _14361_);
  or _65336_ (_14364_, _14363_, _14360_);
  or _65337_ (_14365_, _14364_, _14357_);
  or _65338_ (_14366_, _14365_, _14352_);
  or _65339_ (_14367_, _14366_, _14325_);
  and _65340_ (_14368_, _14367_, _07010_);
  or _65341_ (_14369_, _14368_, _08743_);
  or _65342_ (_14370_, _14369_, _14324_);
  and _65343_ (_14371_, _08743_, _06799_);
  nor _65344_ (_14372_, _14371_, _06021_);
  and _65345_ (_14373_, _14372_, _14370_);
  and _65346_ (_14374_, _08699_, _06021_);
  or _65347_ (_14375_, _14374_, _05724_);
  or _65348_ (_14376_, _14375_, _14373_);
  and _65349_ (_14377_, _05724_, \oc8051_golden_model_1.PC [1]);
  nor _65350_ (_14378_, _14377_, _08752_);
  and _65351_ (_14379_, _14378_, _14376_);
  or _65352_ (_14380_, _14379_, _14264_);
  and _65353_ (_14381_, _14380_, _08765_);
  and _65354_ (_14382_, _10994_, _08757_);
  or _65355_ (_14383_, _14382_, _08301_);
  or _65356_ (_14384_, _14383_, _14381_);
  or _65357_ (_14385_, _14261_, _08764_);
  and _65358_ (_14386_, _14385_, _08300_);
  and _65359_ (_14387_, _14386_, _14384_);
  and _65360_ (_14388_, _10992_, _07031_);
  or _65361_ (_14389_, _14388_, _05736_);
  or _65362_ (_14390_, _14389_, _14387_);
  and _65363_ (_14391_, _05736_, \oc8051_golden_model_1.PC [1]);
  nor _65364_ (_14392_, _14391_, _08778_);
  and _65365_ (_14393_, _14392_, _14390_);
  and _65366_ (_14394_, _14260_, _08778_);
  or _65367_ (_14395_, _14394_, _08783_);
  or _65368_ (_14396_, _14395_, _14393_);
  nand _65369_ (_14397_, _10993_, _08783_);
  and _65370_ (_14398_, _14397_, _05734_);
  and _65371_ (_14399_, _14398_, _14396_);
  nor _65372_ (_14400_, _14399_, _14259_);
  nor _65373_ (_14401_, _14400_, _07278_);
  not _65374_ (_14402_, _14255_);
  nand _65375_ (_14403_, _14402_, _07278_);
  nand _65376_ (_14404_, _14403_, _06459_);
  or _65377_ (_14405_, _14404_, _14401_);
  or _65378_ (_14406_, _14402_, _06459_);
  and _65379_ (_14407_, _14406_, _06866_);
  and _65380_ (_14408_, _14407_, _14405_);
  or _65381_ (_14409_, _14408_, _14258_);
  nand _65382_ (_14410_, _14255_, _07210_);
  and _65383_ (_14411_, _14410_, _07052_);
  and _65384_ (_14412_, _14411_, _14409_);
  nor _65385_ (_14413_, _09183_, _09121_);
  nor _65386_ (_14414_, _14413_, _07052_);
  or _65387_ (_14415_, _14414_, _14412_);
  and _65388_ (_14416_, _14415_, _08797_);
  nor _65389_ (_14417_, _14284_, _08797_);
  or _65390_ (_14418_, _14417_, _06127_);
  or _65391_ (_14419_, _14418_, _14416_);
  nand _65392_ (_14420_, _06127_, _12086_);
  and _65393_ (_14421_, _14420_, _12766_);
  and _65394_ (_14422_, _14421_, _14419_);
  and _65395_ (_14423_, _05752_, _05312_);
  or _65396_ (_14424_, _07058_, _14423_);
  or _65397_ (_14425_, _14424_, _14422_);
  or _65398_ (_14426_, _14273_, _07295_);
  and _65399_ (_14427_, _14426_, _09154_);
  and _65400_ (_14428_, _14427_, _14425_);
  or _65401_ (_14429_, _14428_, _14256_);
  and _65402_ (_14430_, _14429_, _07069_);
  and _65403_ (_14431_, _14413_, _07068_);
  or _65404_ (_14432_, _14431_, _07067_);
  or _65405_ (_14433_, _14432_, _14430_);
  or _65406_ (_14434_, _14284_, _07232_);
  and _65407_ (_14435_, _14434_, _07304_);
  and _65408_ (_14436_, _14435_, _14433_);
  or _65409_ (_14437_, _14436_, _14254_);
  and _65410_ (_14438_, _14437_, _14253_);
  nor _65411_ (_14439_, _07627_, _01340_);
  and _65412_ (_14440_, _14439_, _42882_);
  nor _65413_ (_14441_, _07627_, _06029_);
  and _65414_ (_14442_, _14441_, _01336_);
  and _65415_ (_14443_, _14442_, _42882_);
  not _65416_ (_14444_, _14443_);
  or _65417_ (_14445_, _07627_, \oc8051_golden_model_1.SP [1]);
  or _65418_ (_14446_, _14445_, _01340_);
  or _65419_ (_14447_, _14446_, rst);
  and _65420_ (_14448_, _14447_, _14444_);
  not _65421_ (_14449_, _07622_);
  or _65422_ (_14450_, _07627_, _14449_);
  or _65423_ (_14451_, _14450_, _01340_);
  or _65424_ (_14452_, _14451_, rst);
  not _65425_ (_14453_, _07625_);
  or _65426_ (_14454_, _07627_, _14453_);
  or _65427_ (_14455_, _14454_, _01340_);
  or _65428_ (_14456_, _14455_, rst);
  and _65429_ (_14457_, _14456_, _14452_);
  and _65430_ (_14458_, _14457_, _14448_);
  and _65431_ (_14459_, _14458_, _14440_);
  not _65432_ (_14460_, _07627_);
  not _65433_ (_14461_, _11900_);
  nor _65434_ (_14462_, _14461_, _06127_);
  and _65435_ (_14463_, _12051_, _06127_);
  or _65436_ (_14464_, _14463_, _14462_);
  and _65437_ (_14465_, _14464_, _14460_);
  and _65438_ (_14466_, _14465_, _01336_);
  and _65439_ (_14467_, _14466_, _42882_);
  and _65440_ (_14468_, _14467_, _14459_);
  or _65441_ (_40793_, _14468_, _14438_);
  or _65442_ (_14469_, _14080_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _65443_ (_14470_, _14469_, _14073_);
  nor _65444_ (_14471_, _09162_, _09160_);
  nor _65445_ (_14472_, _14471_, _09163_);
  and _65446_ (_14473_, _14472_, _14235_);
  and _65447_ (_14474_, _05803_, _05732_);
  nand _65448_ (_14475_, _07530_, _08541_);
  or _65449_ (_14476_, _09030_, _05952_);
  nand _65450_ (_14477_, _14476_, _08174_);
  and _65451_ (_14478_, _14477_, _06992_);
  nor _65452_ (_14479_, _12564_, _07732_);
  or _65453_ (_14480_, _14479_, _08378_);
  and _65454_ (_14481_, _08291_, _07530_);
  nor _65455_ (_14482_, _08291_, _07530_);
  or _65456_ (_14483_, _14482_, _14481_);
  or _65457_ (_14484_, _14483_, _08383_);
  nor _65458_ (_14485_, _06943_, _09956_);
  and _65459_ (_14486_, _06943_, _05803_);
  or _65460_ (_14487_, _14486_, _08384_);
  or _65461_ (_14488_, _14487_, _14485_);
  and _65462_ (_14489_, _14488_, _14484_);
  and _65463_ (_14490_, _14489_, _08381_);
  nand _65464_ (_14491_, _08491_, _08176_);
  or _65465_ (_14492_, _08491_, _08176_);
  nand _65466_ (_14493_, _14492_, _14491_);
  and _65467_ (_14494_, _14493_, _06955_);
  or _65468_ (_14495_, _14494_, _14490_);
  and _65469_ (_14496_, _14495_, _08380_);
  nand _65470_ (_14497_, _12564_, _12542_);
  and _65471_ (_14498_, _14497_, _06953_);
  or _65472_ (_14499_, _14498_, _07272_);
  or _65473_ (_14500_, _14499_, _14496_);
  nor _65474_ (_14501_, _05803_, _05690_);
  nor _65475_ (_14502_, _14501_, _06963_);
  and _65476_ (_14503_, _14502_, _14500_);
  and _65477_ (_14504_, _09160_, _06963_);
  or _65478_ (_14505_, _14504_, _06975_);
  or _65479_ (_14506_, _14505_, _14503_);
  and _65480_ (_14507_, _14506_, _14480_);
  or _65481_ (_14508_, _14507_, _06038_);
  nand _65482_ (_14509_, _08176_, _06038_);
  and _65483_ (_14510_, _14509_, _06036_);
  and _65484_ (_14511_, _14510_, _14508_);
  not _65485_ (_14512_, _12565_);
  and _65486_ (_14513_, _14497_, _14512_);
  and _65487_ (_14514_, _14513_, _06035_);
  or _65488_ (_14515_, _14514_, _14511_);
  and _65489_ (_14516_, _14515_, _05686_);
  or _65490_ (_14517_, _05804_, _05686_);
  nand _65491_ (_14518_, _06233_, _14517_);
  or _65492_ (_14519_, _14518_, _14516_);
  nand _65493_ (_14520_, _08176_, _06573_);
  and _65494_ (_14521_, _14520_, _06993_);
  and _65495_ (_14522_, _14521_, _14519_);
  or _65496_ (_14523_, _14522_, _14478_);
  and _65497_ (_14524_, _14523_, _07308_);
  nand _65498_ (_14525_, _07732_, _10606_);
  and _65499_ (_14526_, _14525_, _06991_);
  and _65500_ (_14527_, _14526_, _14497_);
  or _65501_ (_14528_, _14527_, _14524_);
  and _65502_ (_14529_, _14528_, _05673_);
  or _65503_ (_14530_, _05804_, _05673_);
  nand _65504_ (_14531_, _07009_, _14530_);
  or _65505_ (_14532_, _14531_, _14529_);
  and _65506_ (_14533_, _14532_, _14475_);
  or _65507_ (_14534_, _14533_, _07013_);
  or _65508_ (_14535_, _09182_, _07231_);
  and _65509_ (_14536_, _14535_, _08545_);
  and _65510_ (_14537_, _14536_, _14534_);
  nor _65511_ (_14538_, _08549_, _07530_);
  and _65512_ (_14539_, _08668_, \oc8051_golden_model_1.SCON [2]);
  and _65513_ (_14540_, _08650_, \oc8051_golden_model_1.B [2]);
  or _65514_ (_14541_, _14540_, _14539_);
  and _65515_ (_14542_, _08702_, \oc8051_golden_model_1.TL0 [2]);
  and _65516_ (_14543_, _08704_, \oc8051_golden_model_1.PSW [2]);
  or _65517_ (_14544_, _14543_, _14542_);
  or _65518_ (_14545_, _14544_, _14541_);
  and _65519_ (_14546_, _08675_, \oc8051_golden_model_1.TMOD [2]);
  and _65520_ (_14547_, _08682_, \oc8051_golden_model_1.P1 [2]);
  or _65521_ (_14548_, _14547_, _14546_);
  and _65522_ (_14549_, _08680_, \oc8051_golden_model_1.TCON [2]);
  and _65523_ (_14550_, _08677_, \oc8051_golden_model_1.SBUF [2]);
  or _65524_ (_14551_, _14550_, _14549_);
  or _65525_ (_14552_, _14551_, _14548_);
  and _65526_ (_14553_, _08687_, \oc8051_golden_model_1.P2 [2]);
  and _65527_ (_14554_, _08690_, \oc8051_golden_model_1.IP [2]);
  or _65528_ (_14555_, _14554_, _14553_);
  and _65529_ (_14556_, _08693_, \oc8051_golden_model_1.IE [2]);
  and _65530_ (_14557_, _08695_, \oc8051_golden_model_1.P3 [2]);
  or _65531_ (_14558_, _14557_, _14556_);
  or _65532_ (_14559_, _14558_, _14555_);
  and _65533_ (_14560_, _08660_, \oc8051_golden_model_1.P0 [2]);
  and _65534_ (_14561_, _08654_, \oc8051_golden_model_1.ACC [2]);
  or _65535_ (_14562_, _14561_, _14560_);
  or _65536_ (_14563_, _14562_, _14559_);
  or _65537_ (_14564_, _14563_, _14552_);
  or _65538_ (_14565_, _14564_, _14545_);
  and _65539_ (_14566_, _08725_, \oc8051_golden_model_1.TH1 [2]);
  and _65540_ (_14567_, _08716_, \oc8051_golden_model_1.TL1 [2]);
  and _65541_ (_14568_, _08719_, \oc8051_golden_model_1.SP [2]);
  or _65542_ (_14569_, _14568_, _14567_);
  or _65543_ (_14570_, _14569_, _14566_);
  and _65544_ (_14571_, _08728_, \oc8051_golden_model_1.DPL [2]);
  and _65545_ (_14572_, _08732_, \oc8051_golden_model_1.PCON [2]);
  or _65546_ (_14573_, _14572_, _14571_);
  and _65547_ (_14574_, _08723_, \oc8051_golden_model_1.DPH [2]);
  and _65548_ (_14575_, _08712_, \oc8051_golden_model_1.TH0 [2]);
  or _65549_ (_14576_, _14575_, _14574_);
  or _65550_ (_14577_, _14576_, _14573_);
  or _65551_ (_14578_, _14577_, _14570_);
  or _65552_ (_14579_, _14578_, _14565_);
  or _65553_ (_14580_, _14579_, _14538_);
  and _65554_ (_14581_, _14580_, _07010_);
  or _65555_ (_14582_, _14581_, _08743_);
  or _65556_ (_14583_, _14582_, _14537_);
  and _65557_ (_14584_, _08743_, _06403_);
  nor _65558_ (_14585_, _14584_, _06021_);
  and _65559_ (_14586_, _14585_, _14583_);
  and _65560_ (_14587_, _08730_, _06021_);
  or _65561_ (_14588_, _14587_, _05724_);
  or _65562_ (_14589_, _14588_, _14586_);
  and _65563_ (_14590_, _05804_, _05724_);
  nor _65564_ (_14591_, _14590_, _08752_);
  and _65565_ (_14592_, _14591_, _14589_);
  nand _65566_ (_14593_, _08176_, _06445_);
  nor _65567_ (_14594_, _08176_, _06445_);
  not _65568_ (_14595_, _14594_);
  and _65569_ (_14596_, _14595_, _14593_);
  and _65570_ (_14597_, _14596_, _08752_);
  or _65571_ (_14598_, _14597_, _14592_);
  and _65572_ (_14599_, _14598_, _08765_);
  and _65573_ (_14600_, _10991_, _08757_);
  or _65574_ (_14601_, _14600_, _14599_);
  and _65575_ (_14602_, _14601_, _08764_);
  and _65576_ (_14603_, _14594_, _08301_);
  or _65577_ (_14604_, _14603_, _14602_);
  and _65578_ (_14605_, _14604_, _08300_);
  and _65579_ (_14606_, _10989_, _07031_);
  or _65580_ (_14607_, _14606_, _05736_);
  or _65581_ (_14608_, _14607_, _14605_);
  and _65582_ (_14609_, _05804_, _05736_);
  nor _65583_ (_14610_, _14609_, _08778_);
  and _65584_ (_14611_, _14610_, _14608_);
  and _65585_ (_14612_, _14593_, _08778_);
  or _65586_ (_14613_, _14612_, _08783_);
  or _65587_ (_14614_, _14613_, _14611_);
  nand _65588_ (_14615_, _10990_, _08783_);
  and _65589_ (_14616_, _14615_, _05734_);
  and _65590_ (_14617_, _14616_, _14614_);
  or _65591_ (_14618_, _14617_, _14474_);
  and _65592_ (_14619_, _14618_, _08283_);
  and _65593_ (_14620_, _06133_, _05495_);
  not _65594_ (_14621_, _14620_);
  and _65595_ (_14622_, _08285_, _14621_);
  not _65596_ (_14623_, _14622_);
  or _65597_ (_14624_, _14623_, _06708_);
  and _65598_ (_14625_, _14483_, _08282_);
  or _65599_ (_14626_, _14625_, _14624_);
  or _65600_ (_14627_, _14626_, _14619_);
  not _65601_ (_14628_, _14624_);
  or _65602_ (_14629_, _14628_, _14483_);
  and _65603_ (_14630_, _14629_, _07052_);
  and _65604_ (_14631_, _14630_, _14627_);
  nor _65605_ (_14632_, _09121_, _09030_);
  or _65606_ (_14633_, _14632_, _09122_);
  and _65607_ (_14634_, _14633_, _07051_);
  or _65608_ (_14635_, _14634_, _14631_);
  and _65609_ (_14636_, _14635_, _08797_);
  and _65610_ (_14637_, _14493_, _07050_);
  or _65611_ (_14638_, _14637_, _06127_);
  or _65612_ (_14639_, _14638_, _14636_);
  nand _65613_ (_14640_, _12084_, _06127_);
  and _65614_ (_14641_, _14640_, _12766_);
  and _65615_ (_14642_, _14641_, _14639_);
  and _65616_ (_14643_, _05803_, _05752_);
  or _65617_ (_14644_, _07058_, _14643_);
  or _65618_ (_14645_, _14644_, _14642_);
  or _65619_ (_14646_, _14479_, _07295_);
  and _65620_ (_14647_, _14646_, _09154_);
  and _65621_ (_14648_, _14647_, _14645_);
  or _65622_ (_14649_, _14648_, _14473_);
  and _65623_ (_14650_, _14649_, _07069_);
  or _65624_ (_14651_, _09183_, _09182_);
  nor _65625_ (_14652_, _09184_, _07069_);
  and _65626_ (_14653_, _14652_, _14651_);
  or _65627_ (_14654_, _14653_, _07067_);
  or _65628_ (_14655_, _14654_, _14650_);
  nor _65629_ (_14656_, _08177_, _08128_);
  nor _65630_ (_14657_, _14656_, _08178_);
  or _65631_ (_14658_, _14657_, _07232_);
  and _65632_ (_14659_, _14658_, _07304_);
  and _65633_ (_14660_, _14659_, _14655_);
  or _65634_ (_14661_, _14660_, _14254_);
  and _65635_ (_14662_, _14661_, _14470_);
  and _65636_ (_14663_, _12043_, _06127_);
  not _65637_ (_14664_, _11887_);
  nor _65638_ (_14665_, _14664_, _06127_);
  or _65639_ (_14666_, _14665_, _14663_);
  and _65640_ (_14667_, _14666_, _14460_);
  and _65641_ (_14668_, _14667_, _01336_);
  and _65642_ (_14669_, _14668_, _42882_);
  and _65643_ (_14670_, _14669_, _14459_);
  or _65644_ (_40794_, _14670_, _14662_);
  and _65645_ (_14671_, _14491_, _08029_);
  or _65646_ (_14672_, _14671_, _08493_);
  or _65647_ (_14673_, _14672_, _08797_);
  nor _65648_ (_14674_, _14481_, _07353_);
  or _65649_ (_14675_, _14674_, _08292_);
  or _65650_ (_14676_, _14675_, _08286_);
  nor _65651_ (_14677_, _08028_, _06215_);
  and _65652_ (_14678_, _14677_, _08301_);
  nor _65653_ (_14679_, _06148_, _05673_);
  nand _65654_ (_14680_, _08028_, _06573_);
  nor _65655_ (_14681_, _12666_, _07723_);
  or _65656_ (_14682_, _14681_, _08378_);
  nand _65657_ (_14683_, _12666_, _12644_);
  or _65658_ (_14684_, _14683_, _08380_);
  and _65659_ (_14685_, _14672_, _06955_);
  or _65660_ (_14686_, _14675_, _08383_);
  and _65661_ (_14687_, _06943_, _05853_);
  nor _65662_ (_14688_, _06943_, _10010_);
  or _65663_ (_14689_, _14688_, _14687_);
  nor _65664_ (_14690_, _14689_, _08384_);
  nor _65665_ (_14691_, _14690_, _06955_);
  and _65666_ (_14692_, _14691_, _14686_);
  or _65667_ (_14693_, _14692_, _06953_);
  or _65668_ (_14694_, _14693_, _14685_);
  and _65669_ (_14695_, _14694_, _14684_);
  or _65670_ (_14696_, _14695_, _07272_);
  nor _65671_ (_14697_, _05853_, _05690_);
  nor _65672_ (_14698_, _14697_, _06963_);
  and _65673_ (_14699_, _14698_, _14696_);
  and _65674_ (_14700_, _09159_, _06963_);
  or _65675_ (_14701_, _14700_, _06975_);
  or _65676_ (_14702_, _14701_, _14699_);
  and _65677_ (_14703_, _14702_, _14682_);
  or _65678_ (_14704_, _14703_, _06038_);
  nand _65679_ (_14705_, _08028_, _06038_);
  and _65680_ (_14706_, _14705_, _06036_);
  and _65681_ (_14707_, _14706_, _14704_);
  not _65682_ (_14708_, _12667_);
  and _65683_ (_14709_, _14683_, _14708_);
  and _65684_ (_14710_, _14709_, _06035_);
  or _65685_ (_14711_, _14710_, _14707_);
  and _65686_ (_14712_, _14711_, _05686_);
  or _65687_ (_14713_, _06148_, _05686_);
  nand _65688_ (_14714_, _06233_, _14713_);
  or _65689_ (_14715_, _14714_, _14712_);
  and _65690_ (_14716_, _14715_, _14680_);
  or _65691_ (_14717_, _14716_, _06992_);
  and _65692_ (_14718_, _09181_, _06053_);
  nand _65693_ (_14719_, _08026_, _06992_);
  or _65694_ (_14720_, _14719_, _14718_);
  and _65695_ (_14721_, _14720_, _14717_);
  or _65696_ (_14722_, _14721_, _06991_);
  and _65697_ (_14723_, _07723_, \oc8051_golden_model_1.PSW [7]);
  or _65698_ (_14724_, _14681_, _14723_);
  or _65699_ (_14725_, _14724_, _07308_);
  and _65700_ (_14726_, _14725_, _05673_);
  and _65701_ (_14727_, _14726_, _14722_);
  or _65702_ (_14728_, _14727_, _14679_);
  and _65703_ (_14729_, _14728_, _07009_);
  nor _65704_ (_14730_, _07353_, _07009_);
  or _65705_ (_14731_, _14730_, _07013_);
  or _65706_ (_14732_, _14731_, _14729_);
  or _65707_ (_14733_, _09181_, _07231_);
  and _65708_ (_14734_, _14733_, _08545_);
  and _65709_ (_14735_, _14734_, _14732_);
  nor _65710_ (_14736_, _08549_, _07353_);
  and _65711_ (_14737_, _08654_, \oc8051_golden_model_1.ACC [3]);
  and _65712_ (_14738_, _08650_, \oc8051_golden_model_1.B [3]);
  or _65713_ (_14739_, _14738_, _14737_);
  and _65714_ (_14740_, _08660_, \oc8051_golden_model_1.P0 [3]);
  and _65715_ (_14741_, _08704_, \oc8051_golden_model_1.PSW [3]);
  or _65716_ (_14742_, _14741_, _14740_);
  or _65717_ (_14743_, _14742_, _14739_);
  and _65718_ (_14744_, _08680_, \oc8051_golden_model_1.TCON [3]);
  and _65719_ (_14745_, _08682_, \oc8051_golden_model_1.P1 [3]);
  or _65720_ (_14746_, _14745_, _14744_);
  and _65721_ (_14747_, _08668_, \oc8051_golden_model_1.SCON [3]);
  and _65722_ (_14748_, _08677_, \oc8051_golden_model_1.SBUF [3]);
  or _65723_ (_14749_, _14748_, _14747_);
  or _65724_ (_14750_, _14749_, _14746_);
  and _65725_ (_14751_, _08687_, \oc8051_golden_model_1.P2 [3]);
  and _65726_ (_14752_, _08690_, \oc8051_golden_model_1.IP [3]);
  or _65727_ (_14753_, _14752_, _14751_);
  and _65728_ (_14754_, _08693_, \oc8051_golden_model_1.IE [3]);
  and _65729_ (_14755_, _08695_, \oc8051_golden_model_1.P3 [3]);
  or _65730_ (_14756_, _14755_, _14754_);
  or _65731_ (_14757_, _14756_, _14753_);
  and _65732_ (_14758_, _08675_, \oc8051_golden_model_1.TMOD [3]);
  and _65733_ (_14759_, _08702_, \oc8051_golden_model_1.TL0 [3]);
  or _65734_ (_14760_, _14759_, _14758_);
  or _65735_ (_14761_, _14760_, _14757_);
  or _65736_ (_14762_, _14761_, _14750_);
  or _65737_ (_14763_, _14762_, _14743_);
  and _65738_ (_14764_, _08728_, \oc8051_golden_model_1.DPL [3]);
  and _65739_ (_14765_, _08732_, \oc8051_golden_model_1.PCON [3]);
  and _65740_ (_14766_, _08716_, \oc8051_golden_model_1.TL1 [3]);
  or _65741_ (_14767_, _14766_, _14765_);
  or _65742_ (_14768_, _14767_, _14764_);
  and _65743_ (_14769_, _08725_, \oc8051_golden_model_1.TH1 [3]);
  and _65744_ (_14770_, _08712_, \oc8051_golden_model_1.TH0 [3]);
  or _65745_ (_14771_, _14770_, _14769_);
  and _65746_ (_14772_, _08723_, \oc8051_golden_model_1.DPH [3]);
  and _65747_ (_14773_, _08719_, \oc8051_golden_model_1.SP [3]);
  or _65748_ (_14774_, _14773_, _14772_);
  or _65749_ (_14775_, _14774_, _14771_);
  or _65750_ (_14776_, _14775_, _14768_);
  or _65751_ (_14777_, _14776_, _14763_);
  or _65752_ (_14778_, _14777_, _14736_);
  and _65753_ (_14779_, _14778_, _07010_);
  or _65754_ (_14780_, _14779_, _08743_);
  or _65755_ (_14781_, _14780_, _14735_);
  and _65756_ (_14782_, _08743_, _05983_);
  nor _65757_ (_14783_, _14782_, _06021_);
  and _65758_ (_14784_, _14783_, _14781_);
  and _65759_ (_14785_, _08662_, _06021_);
  or _65760_ (_14786_, _14785_, _05724_);
  or _65761_ (_14787_, _14786_, _14784_);
  and _65762_ (_14788_, _06148_, _05724_);
  nor _65763_ (_14789_, _14788_, _08752_);
  and _65764_ (_14790_, _14789_, _14787_);
  not _65765_ (_14791_, _14677_);
  nand _65766_ (_14792_, _08028_, _06215_);
  and _65767_ (_14793_, _14792_, _14791_);
  and _65768_ (_14794_, _14793_, _08752_);
  or _65769_ (_14795_, _14794_, _08757_);
  or _65770_ (_14796_, _14795_, _14790_);
  or _65771_ (_14797_, _12299_, _08765_);
  and _65772_ (_14798_, _14797_, _08764_);
  and _65773_ (_14799_, _14798_, _14796_);
  or _65774_ (_14800_, _14799_, _14678_);
  and _65775_ (_14801_, _14800_, _08300_);
  and _65776_ (_14802_, _10987_, _07031_);
  or _65777_ (_14803_, _14802_, _05736_);
  or _65778_ (_14804_, _14803_, _14801_);
  and _65779_ (_14805_, _06148_, _05736_);
  nor _65780_ (_14806_, _14805_, _08778_);
  and _65781_ (_14807_, _14806_, _14804_);
  and _65782_ (_14808_, _14792_, _08778_);
  or _65783_ (_14809_, _14808_, _08783_);
  or _65784_ (_14810_, _14809_, _14807_);
  nand _65785_ (_14811_, _10988_, _08783_);
  and _65786_ (_14812_, _14811_, _05734_);
  and _65787_ (_14813_, _14812_, _14810_);
  nand _65788_ (_14814_, _05853_, _05732_);
  nand _65789_ (_14815_, _08286_, _14814_);
  or _65790_ (_14816_, _14815_, _14813_);
  and _65791_ (_14817_, _14816_, _14676_);
  or _65792_ (_14818_, _14817_, _07210_);
  or _65793_ (_14819_, _14675_, _07211_);
  and _65794_ (_14820_, _14819_, _07052_);
  and _65795_ (_14821_, _14820_, _14818_);
  nor _65796_ (_14822_, _09122_, _08985_);
  or _65797_ (_14823_, _14822_, _09123_);
  and _65798_ (_14824_, _14823_, _07051_);
  or _65799_ (_14825_, _14824_, _07050_);
  or _65800_ (_14826_, _14825_, _14821_);
  and _65801_ (_14827_, _14826_, _14673_);
  or _65802_ (_14828_, _14827_, _06127_);
  nand _65803_ (_14829_, _12079_, _06127_);
  and _65804_ (_14830_, _14829_, _12766_);
  and _65805_ (_14831_, _14830_, _14828_);
  and _65806_ (_14832_, _05853_, _05752_);
  or _65807_ (_14833_, _07058_, _14832_);
  or _65808_ (_14834_, _14833_, _14831_);
  or _65809_ (_14835_, _14681_, _07295_);
  and _65810_ (_14836_, _14835_, _09154_);
  and _65811_ (_14837_, _14836_, _14834_);
  nor _65812_ (_14838_, _09163_, _09159_);
  nor _65813_ (_14839_, _14838_, _09164_);
  and _65814_ (_14840_, _14839_, _14235_);
  or _65815_ (_14841_, _14840_, _14837_);
  and _65816_ (_14842_, _14841_, _07069_);
  or _65817_ (_14843_, _09184_, _09181_);
  nor _65818_ (_14844_, _09185_, _07069_);
  and _65819_ (_14845_, _14844_, _14843_);
  or _65820_ (_14846_, _14845_, _07067_);
  or _65821_ (_14847_, _14846_, _14842_);
  nor _65822_ (_14848_, _08178_, _08029_);
  nor _65823_ (_14849_, _14848_, _08179_);
  or _65824_ (_14850_, _14849_, _07232_);
  and _65825_ (_14851_, _14850_, _07304_);
  and _65826_ (_14852_, _14851_, _14847_);
  or _65827_ (_14853_, _14852_, _14254_);
  or _65828_ (_14854_, _14080_, \oc8051_golden_model_1.IRAM[0] [3]);
  and _65829_ (_14855_, _14854_, _14073_);
  and _65830_ (_14856_, _14855_, _14853_);
  and _65831_ (_14857_, _11891_, _09200_);
  and _65832_ (_14858_, _12036_, _06127_);
  or _65833_ (_14859_, _14858_, _14857_);
  and _65834_ (_14860_, _14859_, _14460_);
  and _65835_ (_14861_, _14860_, _01336_);
  and _65836_ (_14862_, _14861_, _42882_);
  and _65837_ (_14863_, _14862_, _14459_);
  or _65838_ (_40795_, _14863_, _14856_);
  or _65839_ (_14864_, _14080_, \oc8051_golden_model_1.IRAM[0] [4]);
  and _65840_ (_14865_, _14864_, _14073_);
  nor _65841_ (_14866_, _09185_, _09180_);
  nor _65842_ (_14867_, _14866_, _09186_);
  or _65843_ (_14868_, _14867_, _07069_);
  and _65844_ (_14869_, _08292_, _08270_);
  nor _65845_ (_14870_, _08292_, _08270_);
  or _65846_ (_14871_, _14870_, _14869_);
  or _65847_ (_14872_, _14871_, _08286_);
  nand _65848_ (_14873_, _08581_, _08272_);
  nor _65849_ (_14874_, _08581_, _08272_);
  not _65850_ (_14875_, _14874_);
  and _65851_ (_14876_, _14875_, _14873_);
  and _65852_ (_14877_, _14876_, _08752_);
  nand _65853_ (_14878_, _12718_, _12716_);
  nand _65854_ (_14879_, _12717_, _10606_);
  and _65855_ (_14880_, _14879_, _06991_);
  and _65856_ (_14881_, _14880_, _14878_);
  nor _65857_ (_14882_, _12717_, _12716_);
  or _65858_ (_14883_, _14882_, _08378_);
  or _65859_ (_14884_, _14878_, _08380_);
  and _65860_ (_14885_, _08493_, _08272_);
  nor _65861_ (_14886_, _08493_, _08272_);
  or _65862_ (_14887_, _14886_, _14885_);
  or _65863_ (_14888_, _14887_, _08381_);
  and _65864_ (_14889_, _09180_, _06948_);
  or _65865_ (_14890_, _14871_, _08383_);
  nor _65866_ (_14891_, _06943_, _09880_);
  and _65867_ (_14892_, _11921_, _06943_);
  or _65868_ (_14893_, _14892_, _14891_);
  or _65869_ (_14894_, _14893_, _08384_);
  and _65870_ (_14895_, _14894_, _06949_);
  and _65871_ (_14896_, _14895_, _14890_);
  or _65872_ (_14897_, _14896_, _06955_);
  or _65873_ (_14898_, _14897_, _14889_);
  and _65874_ (_14899_, _14898_, _14888_);
  or _65875_ (_14900_, _14899_, _06953_);
  and _65876_ (_14901_, _14900_, _14884_);
  or _65877_ (_14902_, _14901_, _07272_);
  nor _65878_ (_14903_, _11921_, _05690_);
  nor _65879_ (_14904_, _14903_, _06963_);
  and _65880_ (_14905_, _14904_, _14902_);
  and _65881_ (_14906_, _09158_, _06963_);
  or _65882_ (_14907_, _14906_, _06975_);
  or _65883_ (_14908_, _14907_, _14905_);
  and _65884_ (_14909_, _14908_, _14883_);
  or _65885_ (_14910_, _14909_, _06038_);
  nand _65886_ (_14911_, _08272_, _06038_);
  and _65887_ (_14912_, _14911_, _06036_);
  and _65888_ (_14913_, _14912_, _14910_);
  not _65889_ (_14914_, _12719_);
  and _65890_ (_14915_, _14878_, _14914_);
  and _65891_ (_14916_, _14915_, _06035_);
  or _65892_ (_14917_, _14916_, _14913_);
  and _65893_ (_14918_, _14917_, _05686_);
  or _65894_ (_14919_, _11922_, _05686_);
  nand _65895_ (_14920_, _14919_, _06233_);
  or _65896_ (_14921_, _14920_, _14918_);
  nand _65897_ (_14922_, _08272_, _06573_);
  and _65898_ (_14923_, _14922_, _14921_);
  or _65899_ (_14924_, _14923_, _06992_);
  and _65900_ (_14925_, _09180_, _06053_);
  nand _65901_ (_14926_, _08225_, _06992_);
  or _65902_ (_14927_, _14926_, _14925_);
  and _65903_ (_14928_, _14927_, _07308_);
  and _65904_ (_14929_, _14928_, _14924_);
  or _65905_ (_14930_, _14929_, _14881_);
  and _65906_ (_14931_, _14930_, _05673_);
  or _65907_ (_14932_, _11922_, _05673_);
  nand _65908_ (_14933_, _14932_, _07009_);
  or _65909_ (_14934_, _14933_, _14931_);
  nand _65910_ (_14935_, _08270_, _08541_);
  and _65911_ (_14936_, _14935_, _14934_);
  or _65912_ (_14937_, _14936_, _07013_);
  or _65913_ (_14938_, _09180_, _07231_);
  and _65914_ (_14939_, _14938_, _08545_);
  and _65915_ (_14940_, _14939_, _14937_);
  nor _65916_ (_14941_, _08549_, _08270_);
  and _65917_ (_14942_, _08650_, \oc8051_golden_model_1.B [4]);
  and _65918_ (_14943_, _08654_, \oc8051_golden_model_1.ACC [4]);
  or _65919_ (_14944_, _14943_, _14942_);
  and _65920_ (_14945_, _08702_, \oc8051_golden_model_1.TL0 [4]);
  and _65921_ (_14946_, _08704_, \oc8051_golden_model_1.PSW [4]);
  or _65922_ (_14947_, _14946_, _14945_);
  or _65923_ (_14948_, _14947_, _14944_);
  and _65924_ (_14949_, _08680_, \oc8051_golden_model_1.TCON [4]);
  and _65925_ (_14950_, _08668_, \oc8051_golden_model_1.SCON [4]);
  or _65926_ (_14951_, _14950_, _14949_);
  and _65927_ (_14952_, _08660_, \oc8051_golden_model_1.P0 [4]);
  and _65928_ (_14953_, _08677_, \oc8051_golden_model_1.SBUF [4]);
  or _65929_ (_14954_, _14953_, _14952_);
  or _65930_ (_14955_, _14954_, _14951_);
  and _65931_ (_14956_, _08687_, \oc8051_golden_model_1.P2 [4]);
  and _65932_ (_14957_, _08690_, \oc8051_golden_model_1.IP [4]);
  or _65933_ (_14958_, _14957_, _14956_);
  and _65934_ (_14959_, _08693_, \oc8051_golden_model_1.IE [4]);
  and _65935_ (_14960_, _08695_, \oc8051_golden_model_1.P3 [4]);
  or _65936_ (_14961_, _14960_, _14959_);
  or _65937_ (_14962_, _14961_, _14958_);
  and _65938_ (_14963_, _08675_, \oc8051_golden_model_1.TMOD [4]);
  and _65939_ (_14964_, _08682_, \oc8051_golden_model_1.P1 [4]);
  or _65940_ (_14965_, _14964_, _14963_);
  or _65941_ (_14966_, _14965_, _14962_);
  or _65942_ (_14967_, _14966_, _14955_);
  or _65943_ (_14968_, _14967_, _14948_);
  and _65944_ (_14969_, _08728_, \oc8051_golden_model_1.DPL [4]);
  and _65945_ (_14970_, _08719_, \oc8051_golden_model_1.SP [4]);
  and _65946_ (_14971_, _08723_, \oc8051_golden_model_1.DPH [4]);
  or _65947_ (_14972_, _14971_, _14970_);
  or _65948_ (_14973_, _14972_, _14969_);
  and _65949_ (_14974_, _08716_, \oc8051_golden_model_1.TL1 [4]);
  and _65950_ (_14975_, _08725_, \oc8051_golden_model_1.TH1 [4]);
  or _65951_ (_14976_, _14975_, _14974_);
  and _65952_ (_14977_, _08732_, \oc8051_golden_model_1.PCON [4]);
  and _65953_ (_14978_, _08712_, \oc8051_golden_model_1.TH0 [4]);
  or _65954_ (_14979_, _14978_, _14977_);
  or _65955_ (_14980_, _14979_, _14976_);
  or _65956_ (_14981_, _14980_, _14973_);
  or _65957_ (_14982_, _14981_, _14968_);
  or _65958_ (_14983_, _14982_, _14941_);
  and _65959_ (_14984_, _14983_, _07010_);
  or _65960_ (_14985_, _14984_, _08743_);
  or _65961_ (_14986_, _14985_, _14940_);
  and _65962_ (_14987_, _08743_, _06758_);
  nor _65963_ (_14988_, _14987_, _06021_);
  and _65964_ (_14989_, _14988_, _14986_);
  and _65965_ (_14990_, _08665_, _06021_);
  or _65966_ (_14991_, _14990_, _05724_);
  or _65967_ (_14992_, _14991_, _14989_);
  and _65968_ (_14993_, _11922_, _05724_);
  nor _65969_ (_14994_, _14993_, _08752_);
  and _65970_ (_14995_, _14994_, _14992_);
  or _65971_ (_14996_, _14995_, _14877_);
  and _65972_ (_14997_, _14996_, _08765_);
  and _65973_ (_14998_, _10986_, _08757_);
  or _65974_ (_14999_, _14998_, _14997_);
  and _65975_ (_15000_, _14999_, _08764_);
  and _65976_ (_15001_, _14874_, _08301_);
  or _65977_ (_15002_, _15001_, _15000_);
  and _65978_ (_15003_, _15002_, _08300_);
  and _65979_ (_15004_, _10983_, _07031_);
  or _65980_ (_15005_, _15004_, _05736_);
  or _65981_ (_15006_, _15005_, _15003_);
  and _65982_ (_15007_, _11922_, _05736_);
  nor _65983_ (_15008_, _15007_, _08778_);
  and _65984_ (_15009_, _15008_, _15006_);
  and _65985_ (_15010_, _14873_, _08778_);
  or _65986_ (_15011_, _15010_, _08783_);
  or _65987_ (_15012_, _15011_, _15009_);
  nand _65988_ (_15013_, _10985_, _08783_);
  and _65989_ (_15014_, _15013_, _05734_);
  and _65990_ (_15015_, _15014_, _15012_);
  nand _65991_ (_15016_, _11921_, _05732_);
  nand _65992_ (_15017_, _15016_, _08286_);
  or _65993_ (_15018_, _15017_, _15015_);
  and _65994_ (_15019_, _15018_, _14872_);
  or _65995_ (_15020_, _15019_, _07210_);
  and _65996_ (_15021_, _10394_, _05495_);
  not _65997_ (_15022_, _15021_);
  or _65998_ (_15023_, _14871_, _07211_);
  and _65999_ (_15024_, _15023_, _15022_);
  and _66000_ (_15025_, _15024_, _15020_);
  nor _66001_ (_15026_, _09123_, _08937_);
  or _66002_ (_15027_, _15026_, _09124_);
  or _66003_ (_15028_, _15027_, _06712_);
  and _66004_ (_15029_, _15028_, _07051_);
  or _66005_ (_15030_, _15029_, _15025_);
  not _66006_ (_15031_, _06712_);
  or _66007_ (_15032_, _15027_, _15031_);
  and _66008_ (_15033_, _15032_, _08797_);
  and _66009_ (_15034_, _15033_, _15030_);
  and _66010_ (_15035_, _14887_, _07050_);
  or _66011_ (_15036_, _15035_, _06127_);
  or _66012_ (_15037_, _15036_, _15034_);
  nand _66013_ (_15038_, _12075_, _06127_);
  and _66014_ (_15039_, _15038_, _12766_);
  and _66015_ (_15040_, _15039_, _15037_);
  and _66016_ (_15041_, _11921_, _05752_);
  or _66017_ (_15042_, _15041_, _07058_);
  or _66018_ (_15043_, _15042_, _15040_);
  or _66019_ (_15044_, _14882_, _07295_);
  and _66020_ (_15045_, _15044_, _09154_);
  and _66021_ (_15046_, _15045_, _15043_);
  nor _66022_ (_15047_, _09164_, _09158_);
  nor _66023_ (_15048_, _15047_, _09165_);
  and _66024_ (_15049_, _15048_, _14235_);
  or _66025_ (_15050_, _15049_, _07068_);
  or _66026_ (_15051_, _15050_, _15046_);
  and _66027_ (_15052_, _15051_, _14868_);
  or _66028_ (_15053_, _15052_, _07067_);
  nor _66029_ (_15054_, _08273_, _08179_);
  nor _66030_ (_15055_, _15054_, _08274_);
  or _66031_ (_15056_, _15055_, _07232_);
  and _66032_ (_15057_, _15056_, _07304_);
  and _66033_ (_15058_, _15057_, _15053_);
  or _66034_ (_15059_, _15058_, _14254_);
  and _66035_ (_15060_, _15059_, _14865_);
  and _66036_ (_15061_, _12032_, _06127_);
  not _66037_ (_15062_, _11884_);
  nor _66038_ (_15063_, _15062_, _06127_);
  or _66039_ (_15064_, _15063_, _15061_);
  and _66040_ (_15065_, _15064_, _14460_);
  and _66041_ (_15066_, _15065_, _01336_);
  and _66042_ (_15067_, _15066_, _42882_);
  and _66043_ (_15068_, _15067_, _14459_);
  or _66044_ (_40797_, _15068_, _15060_);
  or _66045_ (_15069_, _14080_, \oc8051_golden_model_1.IRAM[0] [5]);
  and _66046_ (_15070_, _15069_, _14073_);
  nor _66047_ (_15071_, _08612_, _07979_);
  and _66048_ (_15072_, _15071_, _08301_);
  nand _66049_ (_15073_, _12640_, _12638_);
  nand _66050_ (_15074_, _12639_, _10606_);
  and _66051_ (_15075_, _15074_, _06991_);
  and _66052_ (_15076_, _15075_, _15073_);
  nor _66053_ (_15077_, _12639_, _12638_);
  or _66054_ (_15078_, _15077_, _08378_);
  or _66055_ (_15079_, _15073_, _08380_);
  or _66056_ (_15080_, _09179_, _06949_);
  nor _66057_ (_15081_, _14869_, _07977_);
  or _66058_ (_15082_, _15081_, _08293_);
  and _66059_ (_15083_, _15082_, _08384_);
  nand _66060_ (_15084_, _11917_, _06943_);
  or _66061_ (_15085_, _06943_, \oc8051_golden_model_1.ACC [5]);
  and _66062_ (_15086_, _15085_, _15084_);
  and _66063_ (_15087_, _15086_, _08383_);
  or _66064_ (_15088_, _15087_, _06948_);
  or _66065_ (_15089_, _15088_, _15083_);
  and _66066_ (_15090_, _15089_, _15080_);
  or _66067_ (_15091_, _15090_, _06955_);
  nor _66068_ (_15092_, _14885_, _07979_);
  or _66069_ (_15093_, _15092_, _08494_);
  or _66070_ (_15094_, _15093_, _08381_);
  and _66071_ (_15095_, _15094_, _15091_);
  or _66072_ (_15096_, _15095_, _06953_);
  and _66073_ (_15097_, _15096_, _15079_);
  or _66074_ (_15098_, _15097_, _07272_);
  nor _66075_ (_15099_, _11916_, _05690_);
  nor _66076_ (_15100_, _15099_, _06963_);
  and _66077_ (_15101_, _15100_, _15098_);
  and _66078_ (_15102_, _09157_, _06963_);
  or _66079_ (_15103_, _15102_, _06975_);
  or _66080_ (_15104_, _15103_, _15101_);
  and _66081_ (_15105_, _15104_, _15078_);
  or _66082_ (_15106_, _15105_, _06038_);
  nand _66083_ (_15107_, _07979_, _06038_);
  and _66084_ (_15108_, _15107_, _06036_);
  and _66085_ (_15109_, _15108_, _15106_);
  not _66086_ (_15110_, _12641_);
  and _66087_ (_15111_, _15073_, _15110_);
  and _66088_ (_15112_, _15111_, _06035_);
  or _66089_ (_15113_, _15112_, _15109_);
  and _66090_ (_15114_, _15113_, _05686_);
  or _66091_ (_15115_, _11917_, _05686_);
  nand _66092_ (_15116_, _15115_, _06233_);
  or _66093_ (_15117_, _15116_, _15114_);
  nand _66094_ (_15118_, _07979_, _06573_);
  and _66095_ (_15119_, _15118_, _15117_);
  or _66096_ (_15120_, _15119_, _06992_);
  and _66097_ (_15121_, _09179_, _06053_);
  nand _66098_ (_15122_, _07932_, _06992_);
  or _66099_ (_15123_, _15122_, _15121_);
  and _66100_ (_15124_, _15123_, _07308_);
  and _66101_ (_15125_, _15124_, _15120_);
  or _66102_ (_15126_, _15125_, _15076_);
  and _66103_ (_15127_, _15126_, _05673_);
  or _66104_ (_15128_, _11917_, _05673_);
  nand _66105_ (_15129_, _15128_, _07009_);
  or _66106_ (_15130_, _15129_, _15127_);
  nand _66107_ (_15131_, _07977_, _08541_);
  and _66108_ (_15132_, _15131_, _15130_);
  or _66109_ (_15133_, _15132_, _07013_);
  or _66110_ (_15134_, _09179_, _07231_);
  and _66111_ (_15135_, _15134_, _08545_);
  and _66112_ (_15136_, _15135_, _15133_);
  nor _66113_ (_15137_, _08549_, _07977_);
  and _66114_ (_15138_, _08675_, \oc8051_golden_model_1.TMOD [5]);
  and _66115_ (_15139_, _08668_, \oc8051_golden_model_1.SCON [5]);
  or _66116_ (_15140_, _15139_, _15138_);
  and _66117_ (_15141_, _08702_, \oc8051_golden_model_1.TL0 [5]);
  and _66118_ (_15142_, _08650_, \oc8051_golden_model_1.B [5]);
  or _66119_ (_15143_, _15142_, _15141_);
  or _66120_ (_15144_, _15143_, _15140_);
  and _66121_ (_15145_, _08660_, \oc8051_golden_model_1.P0 [5]);
  and _66122_ (_15146_, _08680_, \oc8051_golden_model_1.TCON [5]);
  or _66123_ (_15147_, _15146_, _15145_);
  and _66124_ (_15148_, _08682_, \oc8051_golden_model_1.P1 [5]);
  and _66125_ (_15149_, _08704_, \oc8051_golden_model_1.PSW [5]);
  or _66126_ (_15150_, _15149_, _15148_);
  or _66127_ (_15151_, _15150_, _15147_);
  and _66128_ (_15152_, _08693_, \oc8051_golden_model_1.IE [5]);
  and _66129_ (_15153_, _08690_, \oc8051_golden_model_1.IP [5]);
  or _66130_ (_15154_, _15153_, _15152_);
  and _66131_ (_15155_, _08687_, \oc8051_golden_model_1.P2 [5]);
  and _66132_ (_15156_, _08695_, \oc8051_golden_model_1.P3 [5]);
  or _66133_ (_15157_, _15156_, _15155_);
  or _66134_ (_15158_, _15157_, _15154_);
  and _66135_ (_15159_, _08677_, \oc8051_golden_model_1.SBUF [5]);
  and _66136_ (_15160_, _08654_, \oc8051_golden_model_1.ACC [5]);
  or _66137_ (_15161_, _15160_, _15159_);
  or _66138_ (_15162_, _15161_, _15158_);
  or _66139_ (_15163_, _15162_, _15151_);
  or _66140_ (_15164_, _15163_, _15144_);
  and _66141_ (_15165_, _08712_, \oc8051_golden_model_1.TH0 [5]);
  and _66142_ (_15166_, _08723_, \oc8051_golden_model_1.DPH [5]);
  and _66143_ (_15167_, _08725_, \oc8051_golden_model_1.TH1 [5]);
  or _66144_ (_15168_, _15167_, _15166_);
  or _66145_ (_15169_, _15168_, _15165_);
  and _66146_ (_15170_, _08732_, \oc8051_golden_model_1.PCON [5]);
  and _66147_ (_15171_, _08716_, \oc8051_golden_model_1.TL1 [5]);
  or _66148_ (_15172_, _15171_, _15170_);
  and _66149_ (_15173_, _08728_, \oc8051_golden_model_1.DPL [5]);
  and _66150_ (_15174_, _08719_, \oc8051_golden_model_1.SP [5]);
  or _66151_ (_15175_, _15174_, _15173_);
  or _66152_ (_15176_, _15175_, _15172_);
  or _66153_ (_15177_, _15176_, _15169_);
  or _66154_ (_15178_, _15177_, _15164_);
  or _66155_ (_15179_, _15178_, _15137_);
  and _66156_ (_15180_, _15179_, _07010_);
  or _66157_ (_15181_, _15180_, _08743_);
  or _66158_ (_15182_, _15181_, _15136_);
  and _66159_ (_15183_, _08743_, _06359_);
  nor _66160_ (_15184_, _15183_, _06021_);
  and _66161_ (_15185_, _15184_, _15182_);
  and _66162_ (_15186_, _08652_, _06021_);
  or _66163_ (_15187_, _15186_, _05724_);
  or _66164_ (_15188_, _15187_, _15185_);
  and _66165_ (_15189_, _11917_, _05724_);
  nor _66166_ (_15190_, _15189_, _08752_);
  and _66167_ (_15191_, _15190_, _15188_);
  not _66168_ (_15192_, _15071_);
  nand _66169_ (_15194_, _08612_, _07979_);
  and _66170_ (_15195_, _15194_, _15192_);
  and _66171_ (_15196_, _15195_, _08752_);
  or _66172_ (_15197_, _15196_, _08757_);
  or _66173_ (_15198_, _15197_, _15191_);
  or _66174_ (_15199_, _12306_, _08765_);
  and _66175_ (_15200_, _15199_, _08764_);
  and _66176_ (_15201_, _15200_, _15198_);
  or _66177_ (_15202_, _15201_, _15072_);
  and _66178_ (_15203_, _15202_, _08300_);
  and _66179_ (_15204_, _10981_, _07031_);
  or _66180_ (_15205_, _15204_, _05736_);
  or _66181_ (_15206_, _15205_, _15203_);
  and _66182_ (_15207_, _11917_, _05736_);
  nor _66183_ (_15208_, _15207_, _08778_);
  and _66184_ (_15209_, _15208_, _15206_);
  and _66185_ (_15210_, _15194_, _08778_);
  or _66186_ (_15211_, _15210_, _08783_);
  or _66187_ (_15212_, _15211_, _15209_);
  nand _66188_ (_15213_, _10982_, _08783_);
  and _66189_ (_15214_, _15213_, _05734_);
  and _66190_ (_15215_, _15214_, _15212_);
  nand _66191_ (_15216_, _11916_, _05732_);
  nand _66192_ (_15217_, _15216_, _08287_);
  or _66193_ (_15218_, _15217_, _15215_);
  or _66194_ (_15219_, _15082_, _08287_);
  and _66195_ (_15220_, _15219_, _15022_);
  and _66196_ (_15221_, _15220_, _15218_);
  nor _66197_ (_15222_, _09124_, _08888_);
  or _66198_ (_15223_, _15222_, _09125_);
  or _66199_ (_15224_, _15223_, _06712_);
  and _66200_ (_15225_, _15224_, _07051_);
  or _66201_ (_15226_, _15225_, _15221_);
  or _66202_ (_15227_, _15223_, _15031_);
  and _66203_ (_15228_, _15227_, _08797_);
  and _66204_ (_15229_, _15228_, _15226_);
  and _66205_ (_15230_, _15093_, _07050_);
  or _66206_ (_15231_, _15230_, _06127_);
  or _66207_ (_15232_, _15231_, _15229_);
  nand _66208_ (_15233_, _12070_, _06127_);
  and _66209_ (_15234_, _15233_, _12766_);
  and _66210_ (_15235_, _15234_, _15232_);
  and _66211_ (_15236_, _11916_, _05752_);
  or _66212_ (_15237_, _15236_, _07058_);
  or _66213_ (_15238_, _15237_, _15235_);
  or _66214_ (_15239_, _15077_, _07295_);
  and _66215_ (_15240_, _15239_, _09154_);
  and _66216_ (_15241_, _15240_, _15238_);
  or _66217_ (_15242_, _09165_, _09157_);
  nor _66218_ (_15243_, _09166_, _09154_);
  and _66219_ (_15244_, _15243_, _15242_);
  or _66220_ (_15245_, _15244_, _15241_);
  and _66221_ (_15246_, _15245_, _07069_);
  or _66222_ (_15247_, _09186_, _09179_);
  nor _66223_ (_15248_, _09187_, _07069_);
  and _66224_ (_15249_, _15248_, _15247_);
  or _66225_ (_15250_, _15249_, _07067_);
  or _66226_ (_15251_, _15250_, _15246_);
  nor _66227_ (_15252_, _08274_, _07980_);
  nor _66228_ (_15253_, _15252_, _08275_);
  or _66229_ (_15254_, _15253_, _07232_);
  and _66230_ (_15255_, _15254_, _07304_);
  and _66231_ (_15256_, _15255_, _15251_);
  or _66232_ (_15257_, _15256_, _14254_);
  and _66233_ (_15258_, _15257_, _15070_);
  not _66234_ (_15259_, _11880_);
  nor _66235_ (_15260_, _15259_, _06127_);
  and _66236_ (_15261_, _12027_, _06127_);
  or _66237_ (_15262_, _15261_, _15260_);
  and _66238_ (_15263_, _15262_, _14460_);
  and _66239_ (_15264_, _15263_, _01336_);
  and _66240_ (_15265_, _15264_, _42882_);
  and _66241_ (_15266_, _15265_, _14459_);
  or _66242_ (_40798_, _15266_, _15258_);
  or _66243_ (_15267_, _14080_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _66244_ (_15268_, _15267_, _14073_);
  nor _66245_ (_15269_, _09166_, _09156_);
  nor _66246_ (_15270_, _15269_, _09167_);
  and _66247_ (_15271_, _15270_, _14235_);
  nor _66248_ (_15272_, _09125_, _08843_);
  or _66249_ (_15273_, _15272_, _09126_);
  and _66250_ (_15274_, _15273_, _07051_);
  nor _66251_ (_15275_, _08293_, _07883_);
  or _66252_ (_15276_, _15275_, _08294_);
  or _66253_ (_15277_, _15276_, _08286_);
  nor _66254_ (_15278_, _12691_, _12690_);
  or _66255_ (_15279_, _15278_, _08378_);
  nand _66256_ (_15280_, _12692_, _12690_);
  or _66257_ (_15281_, _15280_, _08380_);
  or _66258_ (_15282_, _09178_, _06949_);
  and _66259_ (_15283_, _15276_, _08384_);
  nand _66260_ (_15284_, _11909_, _06943_);
  or _66261_ (_15285_, _06943_, \oc8051_golden_model_1.ACC [6]);
  and _66262_ (_15286_, _15285_, _15284_);
  and _66263_ (_15287_, _15286_, _08383_);
  or _66264_ (_15288_, _15287_, _06948_);
  or _66265_ (_15289_, _15288_, _15283_);
  and _66266_ (_15290_, _15289_, _15282_);
  or _66267_ (_15291_, _15290_, _06955_);
  nor _66268_ (_15292_, _08494_, _07885_);
  or _66269_ (_15293_, _15292_, _08495_);
  or _66270_ (_15294_, _15293_, _08381_);
  and _66271_ (_15295_, _15294_, _15291_);
  or _66272_ (_15296_, _15295_, _06953_);
  and _66273_ (_15297_, _15296_, _15281_);
  or _66274_ (_15298_, _15297_, _07272_);
  nor _66275_ (_15299_, _11908_, _05690_);
  nor _66276_ (_15300_, _15299_, _06963_);
  and _66277_ (_15301_, _15300_, _15298_);
  and _66278_ (_15302_, _09156_, _06963_);
  or _66279_ (_15303_, _15302_, _06975_);
  or _66280_ (_15304_, _15303_, _15301_);
  and _66281_ (_15305_, _15304_, _15279_);
  or _66282_ (_15306_, _15305_, _06038_);
  nand _66283_ (_15307_, _07885_, _06038_);
  and _66284_ (_15308_, _15307_, _06036_);
  and _66285_ (_15309_, _15308_, _15306_);
  not _66286_ (_15310_, _12693_);
  and _66287_ (_15311_, _15280_, _15310_);
  and _66288_ (_15312_, _15311_, _06035_);
  or _66289_ (_15313_, _15312_, _15309_);
  and _66290_ (_15314_, _15313_, _05686_);
  or _66291_ (_15315_, _11909_, _05686_);
  nand _66292_ (_15316_, _15315_, _06233_);
  or _66293_ (_15317_, _15316_, _15314_);
  nand _66294_ (_15318_, _07885_, _06573_);
  and _66295_ (_15319_, _15318_, _15317_);
  or _66296_ (_15320_, _15319_, _06992_);
  and _66297_ (_15321_, _09178_, _06053_);
  nand _66298_ (_15322_, _07838_, _06992_);
  or _66299_ (_15323_, _15322_, _15321_);
  and _66300_ (_15324_, _15323_, _07308_);
  and _66301_ (_15325_, _15324_, _15320_);
  nand _66302_ (_15326_, _12691_, _10606_);
  and _66303_ (_15327_, _15326_, _06991_);
  and _66304_ (_15328_, _15327_, _15280_);
  or _66305_ (_15329_, _15328_, _15325_);
  and _66306_ (_15330_, _15329_, _05673_);
  or _66307_ (_15331_, _11909_, _05673_);
  nand _66308_ (_15332_, _15331_, _07009_);
  or _66309_ (_15333_, _15332_, _15330_);
  nand _66310_ (_15334_, _07883_, _08541_);
  and _66311_ (_15335_, _15334_, _15333_);
  or _66312_ (_15336_, _15335_, _07013_);
  or _66313_ (_15337_, _09178_, _07231_);
  and _66314_ (_15338_, _15337_, _08545_);
  and _66315_ (_15339_, _15338_, _15336_);
  nor _66316_ (_15340_, _08549_, _07883_);
  and _66317_ (_15341_, _08654_, \oc8051_golden_model_1.ACC [6]);
  and _66318_ (_15342_, _08650_, \oc8051_golden_model_1.B [6]);
  or _66319_ (_15343_, _15342_, _15341_);
  and _66320_ (_15344_, _08702_, \oc8051_golden_model_1.TL0 [6]);
  and _66321_ (_15345_, _08677_, \oc8051_golden_model_1.SBUF [6]);
  or _66322_ (_15346_, _15345_, _15344_);
  or _66323_ (_15347_, _15346_, _15343_);
  and _66324_ (_15348_, _08660_, \oc8051_golden_model_1.P0 [6]);
  and _66325_ (_15349_, _08675_, \oc8051_golden_model_1.TMOD [6]);
  or _66326_ (_15350_, _15349_, _15348_);
  and _66327_ (_15351_, _08682_, \oc8051_golden_model_1.P1 [6]);
  and _66328_ (_15352_, _08668_, \oc8051_golden_model_1.SCON [6]);
  or _66329_ (_15353_, _15352_, _15351_);
  or _66330_ (_15354_, _15353_, _15350_);
  and _66331_ (_15355_, _08695_, \oc8051_golden_model_1.P3 [6]);
  and _66332_ (_15356_, _08690_, \oc8051_golden_model_1.IP [6]);
  or _66333_ (_15357_, _15356_, _15355_);
  and _66334_ (_15358_, _08687_, \oc8051_golden_model_1.P2 [6]);
  and _66335_ (_15359_, _08693_, \oc8051_golden_model_1.IE [6]);
  or _66336_ (_15360_, _15359_, _15358_);
  or _66337_ (_15361_, _15360_, _15357_);
  and _66338_ (_15362_, _08680_, \oc8051_golden_model_1.TCON [6]);
  and _66339_ (_15363_, _08704_, \oc8051_golden_model_1.PSW [6]);
  or _66340_ (_15364_, _15363_, _15362_);
  or _66341_ (_15365_, _15364_, _15361_);
  or _66342_ (_15366_, _15365_, _15354_);
  or _66343_ (_15367_, _15366_, _15347_);
  and _66344_ (_15368_, _08716_, \oc8051_golden_model_1.TL1 [6]);
  and _66345_ (_15369_, _08728_, \oc8051_golden_model_1.DPL [6]);
  and _66346_ (_15370_, _08723_, \oc8051_golden_model_1.DPH [6]);
  or _66347_ (_15371_, _15370_, _15369_);
  or _66348_ (_15372_, _15371_, _15368_);
  and _66349_ (_15373_, _08712_, \oc8051_golden_model_1.TH0 [6]);
  and _66350_ (_15374_, _08725_, \oc8051_golden_model_1.TH1 [6]);
  or _66351_ (_15375_, _15374_, _15373_);
  and _66352_ (_15376_, _08732_, \oc8051_golden_model_1.PCON [6]);
  and _66353_ (_15377_, _08719_, \oc8051_golden_model_1.SP [6]);
  or _66354_ (_15378_, _15377_, _15376_);
  or _66355_ (_15379_, _15378_, _15375_);
  or _66356_ (_15380_, _15379_, _15372_);
  or _66357_ (_15381_, _15380_, _15367_);
  or _66358_ (_15382_, _15381_, _15340_);
  and _66359_ (_15383_, _15382_, _07010_);
  or _66360_ (_15384_, _15383_, _08743_);
  or _66361_ (_15385_, _15384_, _15339_);
  and _66362_ (_15386_, _08743_, _06084_);
  nor _66363_ (_15387_, _15386_, _06021_);
  and _66364_ (_15388_, _15387_, _15385_);
  not _66365_ (_15389_, _08647_);
  and _66366_ (_15390_, _15389_, _06021_);
  or _66367_ (_15391_, _15390_, _05724_);
  or _66368_ (_15392_, _15391_, _15388_);
  and _66369_ (_15393_, _11909_, _05724_);
  nor _66370_ (_15394_, _15393_, _08752_);
  and _66371_ (_15395_, _15394_, _15392_);
  nand _66372_ (_15396_, _08647_, _07885_);
  nor _66373_ (_15397_, _08647_, _07885_);
  not _66374_ (_15398_, _15397_);
  and _66375_ (_15399_, _15398_, _15396_);
  and _66376_ (_15400_, _15399_, _08752_);
  or _66377_ (_15401_, _15400_, _15395_);
  and _66378_ (_15402_, _15401_, _08765_);
  and _66379_ (_15403_, _10980_, _08757_);
  or _66380_ (_15404_, _15403_, _15402_);
  and _66381_ (_15405_, _15404_, _08764_);
  and _66382_ (_15406_, _15397_, _08301_);
  or _66383_ (_15407_, _15406_, _15405_);
  and _66384_ (_15408_, _15407_, _08300_);
  and _66385_ (_15409_, _10977_, _07031_);
  or _66386_ (_15410_, _15409_, _05736_);
  or _66387_ (_15411_, _15410_, _15408_);
  and _66388_ (_15412_, _11909_, _05736_);
  nor _66389_ (_15413_, _15412_, _08778_);
  and _66390_ (_15414_, _15413_, _15411_);
  and _66391_ (_15415_, _15396_, _08778_);
  or _66392_ (_15416_, _15415_, _08783_);
  or _66393_ (_15417_, _15416_, _15414_);
  nand _66394_ (_15418_, _10979_, _08783_);
  and _66395_ (_15419_, _15418_, _05734_);
  and _66396_ (_15420_, _15419_, _15417_);
  nand _66397_ (_15421_, _11908_, _05732_);
  nand _66398_ (_15422_, _15421_, _08286_);
  or _66399_ (_15423_, _15422_, _15420_);
  and _66400_ (_15424_, _15423_, _15277_);
  or _66401_ (_15425_, _15424_, _07210_);
  or _66402_ (_15426_, _15276_, _07211_);
  and _66403_ (_15427_, _15426_, _07052_);
  and _66404_ (_15428_, _15427_, _15425_);
  or _66405_ (_15429_, _15428_, _15274_);
  and _66406_ (_15430_, _15429_, _08797_);
  and _66407_ (_15431_, _15293_, _07050_);
  or _66408_ (_15432_, _15431_, _06127_);
  or _66409_ (_15433_, _15432_, _15430_);
  nand _66410_ (_15434_, _12063_, _06127_);
  and _66411_ (_15435_, _15434_, _12766_);
  and _66412_ (_15436_, _15435_, _15433_);
  and _66413_ (_15437_, _11908_, _05752_);
  or _66414_ (_15438_, _15437_, _07058_);
  or _66415_ (_15439_, _15438_, _15436_);
  or _66416_ (_15440_, _15278_, _07295_);
  and _66417_ (_15441_, _15440_, _09154_);
  and _66418_ (_15442_, _15441_, _15439_);
  or _66419_ (_15443_, _15442_, _15271_);
  and _66420_ (_15444_, _15443_, _07069_);
  or _66421_ (_15445_, _09187_, _09178_);
  nor _66422_ (_15446_, _09188_, _07069_);
  and _66423_ (_15447_, _15446_, _15445_);
  or _66424_ (_15448_, _15447_, _07067_);
  or _66425_ (_15449_, _15448_, _15444_);
  nor _66426_ (_15450_, _08275_, _07886_);
  nor _66427_ (_15451_, _15450_, _08276_);
  or _66428_ (_15452_, _15451_, _07232_);
  and _66429_ (_15453_, _15452_, _07304_);
  and _66430_ (_15454_, _15453_, _15449_);
  or _66431_ (_15455_, _15454_, _14254_);
  and _66432_ (_15456_, _15455_, _15268_);
  not _66433_ (_15457_, _11875_);
  nor _66434_ (_15458_, _15457_, _06127_);
  and _66435_ (_15459_, _12020_, _06127_);
  or _66436_ (_15460_, _15459_, _15458_);
  and _66437_ (_15461_, _15460_, _14460_);
  and _66438_ (_15462_, _15461_, _01336_);
  and _66439_ (_15463_, _15462_, _42882_);
  and _66440_ (_15464_, _15463_, _14459_);
  or _66441_ (_40799_, _15464_, _15456_);
  nand _66442_ (_15465_, _14080_, _09196_);
  or _66443_ (_15466_, _14080_, \oc8051_golden_model_1.IRAM[0] [7]);
  and _66444_ (_15467_, _15466_, _14073_);
  and _66445_ (_15468_, _15467_, _15465_);
  and _66446_ (_15469_, _14072_, _09229_);
  or _66447_ (_40800_, _15469_, _15468_);
  nand _66448_ (_15470_, _14071_, _07356_);
  or _66449_ (_15471_, _15470_, _14068_);
  and _66450_ (_15472_, _14077_, _07229_);
  and _66451_ (_15473_, _15472_, _14076_);
  and _66452_ (_15474_, _15473_, _14247_);
  or _66453_ (_15475_, _15473_, _06880_);
  nand _66454_ (_15476_, _15475_, _15470_);
  or _66455_ (_15477_, _15476_, _15474_);
  and _66456_ (_40801_, _15477_, _15471_);
  not _66457_ (_15478_, _15473_);
  or _66458_ (_15479_, _15478_, _14436_);
  or _66459_ (_15480_, _15473_, \oc8051_golden_model_1.IRAM[1] [1]);
  and _66460_ (_15481_, _15480_, _15470_);
  and _66461_ (_15482_, _15481_, _15479_);
  and _66462_ (_15483_, _14447_, _14443_);
  and _66463_ (_15484_, _15483_, _14457_);
  and _66464_ (_15485_, _15484_, _14467_);
  or _66465_ (_40802_, _15485_, _15482_);
  or _66466_ (_15486_, _15478_, _14660_);
  or _66467_ (_15487_, _15473_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _66468_ (_15488_, _15487_, _15470_);
  and _66469_ (_15489_, _15488_, _15486_);
  and _66470_ (_15490_, _15484_, _14669_);
  or _66471_ (_40803_, _15490_, _15489_);
  or _66472_ (_15491_, _15478_, _14852_);
  or _66473_ (_15492_, _15473_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _66474_ (_15493_, _15492_, _15470_);
  and _66475_ (_15494_, _15493_, _15491_);
  and _66476_ (_15495_, _15484_, _14862_);
  or _66477_ (_40805_, _15495_, _15494_);
  or _66478_ (_15496_, _15478_, _15058_);
  or _66479_ (_15497_, _15473_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _66480_ (_15498_, _15497_, _15470_);
  and _66481_ (_15499_, _15498_, _15496_);
  and _66482_ (_15500_, _15484_, _15067_);
  or _66483_ (_40806_, _15500_, _15499_);
  or _66484_ (_15501_, _15478_, _15256_);
  or _66485_ (_15502_, _15473_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _66486_ (_15503_, _15502_, _15470_);
  and _66487_ (_15504_, _15503_, _15501_);
  and _66488_ (_15505_, _15484_, _15265_);
  or _66489_ (_40807_, _15505_, _15504_);
  or _66490_ (_15506_, _15478_, _15454_);
  or _66491_ (_15507_, _15473_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _66492_ (_15508_, _15507_, _15470_);
  and _66493_ (_15509_, _15508_, _15506_);
  and _66494_ (_15510_, _15484_, _15463_);
  or _66495_ (_40808_, _15510_, _15509_);
  and _66496_ (_15511_, _15473_, _09197_);
  or _66497_ (_15512_, _15473_, _07740_);
  nand _66498_ (_15513_, _15512_, _15470_);
  or _66499_ (_15514_, _15513_, _15511_);
  or _66500_ (_15515_, _15470_, _09229_);
  and _66501_ (_40809_, _15515_, _15514_);
  and _66502_ (_15516_, _14068_, _07628_);
  and _66503_ (_15517_, _14071_, _08399_);
  not _66504_ (_15518_, _15517_);
  or _66505_ (_15519_, _15518_, _15516_);
  and _66506_ (_15520_, _07306_, _07074_);
  and _66507_ (_15521_, _15520_, _14076_);
  and _66508_ (_15522_, _15521_, _14247_);
  nor _66509_ (_15523_, _15521_, _06888_);
  or _66510_ (_15524_, _15523_, _15517_);
  or _66511_ (_15525_, _15524_, _15522_);
  and _66512_ (_40813_, _15525_, _15519_);
  not _66513_ (_15526_, _15521_);
  or _66514_ (_15527_, _15526_, _14436_);
  or _66515_ (_15528_, _15521_, \oc8051_golden_model_1.IRAM[2] [1]);
  and _66516_ (_15529_, _15528_, _15518_);
  and _66517_ (_15530_, _15529_, _15527_);
  and _66518_ (_15531_, _14464_, _07628_);
  and _66519_ (_15532_, _15531_, _15517_);
  or _66520_ (_40814_, _15532_, _15530_);
  or _66521_ (_15533_, _15526_, _14660_);
  or _66522_ (_15534_, _15521_, \oc8051_golden_model_1.IRAM[2] [2]);
  and _66523_ (_15535_, _15534_, _15518_);
  and _66524_ (_15536_, _15535_, _15533_);
  and _66525_ (_15537_, _14666_, _07628_);
  and _66526_ (_15538_, _15537_, _15517_);
  or _66527_ (_40815_, _15538_, _15536_);
  or _66528_ (_15539_, _15526_, _14852_);
  or _66529_ (_15540_, _15521_, \oc8051_golden_model_1.IRAM[2] [3]);
  and _66530_ (_15541_, _15540_, _15518_);
  and _66531_ (_15542_, _15541_, _15539_);
  and _66532_ (_15543_, _14859_, _07628_);
  and _66533_ (_15544_, _15543_, _15517_);
  or _66534_ (_40816_, _15544_, _15542_);
  or _66535_ (_15545_, _15526_, _15058_);
  or _66536_ (_15546_, _15521_, \oc8051_golden_model_1.IRAM[2] [4]);
  and _66537_ (_15547_, _15546_, _15518_);
  and _66538_ (_15548_, _15547_, _15545_);
  and _66539_ (_15549_, _15064_, _07628_);
  and _66540_ (_15550_, _15549_, _15517_);
  or _66541_ (_40818_, _15550_, _15548_);
  or _66542_ (_15551_, _15526_, _15256_);
  or _66543_ (_15552_, _15521_, \oc8051_golden_model_1.IRAM[2] [5]);
  and _66544_ (_15553_, _15552_, _15518_);
  and _66545_ (_15554_, _15553_, _15551_);
  and _66546_ (_15555_, _15262_, _07628_);
  and _66547_ (_15556_, _15555_, _15517_);
  or _66548_ (_40819_, _15556_, _15554_);
  or _66549_ (_15557_, _15526_, _15454_);
  or _66550_ (_15558_, _15521_, \oc8051_golden_model_1.IRAM[2] [6]);
  and _66551_ (_15559_, _15558_, _15518_);
  and _66552_ (_15560_, _15559_, _15557_);
  and _66553_ (_15561_, _15460_, _07628_);
  and _66554_ (_15562_, _15561_, _15517_);
  or _66555_ (_40820_, _15562_, _15560_);
  or _66556_ (_15563_, _15526_, _09197_);
  or _66557_ (_15564_, _15521_, \oc8051_golden_model_1.IRAM[2] [7]);
  and _66558_ (_15565_, _15564_, _15518_);
  and _66559_ (_15566_, _15565_, _15563_);
  and _66560_ (_15567_, _15517_, _09230_);
  or _66561_ (_40821_, _15567_, _15566_);
  and _66562_ (_15568_, _14071_, _07080_);
  not _66563_ (_15569_, _15568_);
  or _66564_ (_15570_, _15569_, _15516_);
  and _66565_ (_15571_, _14076_, _07307_);
  and _66566_ (_15572_, _15571_, _14247_);
  nor _66567_ (_15573_, _15571_, _06885_);
  or _66568_ (_15574_, _15573_, _15568_);
  or _66569_ (_15575_, _15574_, _15572_);
  and _66570_ (_40823_, _15575_, _15570_);
  or _66571_ (_15576_, _15571_, \oc8051_golden_model_1.IRAM[3] [1]);
  and _66572_ (_15577_, _15576_, _15569_);
  not _66573_ (_15578_, _15571_);
  or _66574_ (_15579_, _15578_, _14436_);
  and _66575_ (_15580_, _15579_, _15577_);
  and _66576_ (_15581_, _15568_, _15531_);
  or _66577_ (_40824_, _15581_, _15580_);
  or _66578_ (_15582_, _15571_, \oc8051_golden_model_1.IRAM[3] [2]);
  and _66579_ (_15583_, _15582_, _15569_);
  or _66580_ (_15584_, _15578_, _14660_);
  and _66581_ (_15585_, _15584_, _15583_);
  and _66582_ (_15586_, _15568_, _15537_);
  or _66583_ (_40825_, _15586_, _15585_);
  or _66584_ (_15587_, _15571_, \oc8051_golden_model_1.IRAM[3] [3]);
  and _66585_ (_15588_, _15587_, _15569_);
  or _66586_ (_15589_, _15578_, _14852_);
  and _66587_ (_15590_, _15589_, _15588_);
  and _66588_ (_15591_, _15568_, _15543_);
  or _66589_ (_40827_, _15591_, _15590_);
  or _66590_ (_15592_, _15571_, \oc8051_golden_model_1.IRAM[3] [4]);
  and _66591_ (_15593_, _15592_, _15569_);
  or _66592_ (_15594_, _15578_, _15058_);
  and _66593_ (_15595_, _15594_, _15593_);
  and _66594_ (_15596_, _15568_, _15549_);
  or _66595_ (_40828_, _15596_, _15595_);
  or _66596_ (_15597_, _15571_, \oc8051_golden_model_1.IRAM[3] [5]);
  and _66597_ (_15598_, _15597_, _15569_);
  or _66598_ (_15599_, _15578_, _15256_);
  and _66599_ (_15600_, _15599_, _15598_);
  and _66600_ (_15601_, _15568_, _15555_);
  or _66601_ (_40829_, _15601_, _15600_);
  or _66602_ (_15602_, _15571_, \oc8051_golden_model_1.IRAM[3] [6]);
  and _66603_ (_15603_, _15602_, _15569_);
  or _66604_ (_15604_, _15578_, _15454_);
  and _66605_ (_15605_, _15604_, _15603_);
  and _66606_ (_15606_, _15568_, _15561_);
  or _66607_ (_40830_, _15606_, _15605_);
  or _66608_ (_15607_, _15571_, \oc8051_golden_model_1.IRAM[3] [7]);
  and _66609_ (_15608_, _15607_, _15569_);
  or _66610_ (_15609_, _15578_, _09197_);
  and _66611_ (_15610_, _15609_, _15608_);
  and _66612_ (_15611_, _15568_, _09230_);
  or _66613_ (_40831_, _15611_, _15610_);
  and _66614_ (_15612_, _07628_, _07622_);
  and _66615_ (_15613_, _15612_, _14453_);
  and _66616_ (_15614_, _15613_, _07081_);
  not _66617_ (_15615_, _15614_);
  and _66618_ (_15616_, _07615_, _07476_);
  and _66619_ (_15617_, _15616_, _14078_);
  or _66620_ (_15618_, _15617_, \oc8051_golden_model_1.IRAM[4] [0]);
  not _66621_ (_15619_, _15617_);
  or _66622_ (_15620_, _15619_, _14247_);
  and _66623_ (_15621_, _15620_, _15618_);
  and _66624_ (_15622_, _15621_, _15615_);
  and _66625_ (_15623_, _15614_, _15516_);
  or _66626_ (_40835_, _15623_, _15622_);
  or _66627_ (_15624_, _15619_, _14436_);
  or _66628_ (_15625_, _15617_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _66629_ (_15626_, _15625_, _15615_);
  and _66630_ (_15627_, _15626_, _15624_);
  and _66631_ (_15628_, _15614_, _15531_);
  or _66632_ (_40836_, _15628_, _15627_);
  or _66633_ (_15629_, _15619_, _14660_);
  or _66634_ (_15630_, _15617_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _66635_ (_15631_, _15630_, _15615_);
  and _66636_ (_15632_, _15631_, _15629_);
  and _66637_ (_15633_, _15614_, _15537_);
  or _66638_ (_40837_, _15633_, _15632_);
  or _66639_ (_15634_, _15619_, _14852_);
  or _66640_ (_15635_, _15617_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _66641_ (_15636_, _15635_, _15615_);
  and _66642_ (_15637_, _15636_, _15634_);
  and _66643_ (_15638_, _15614_, _15543_);
  or _66644_ (_40838_, _15638_, _15637_);
  or _66645_ (_15639_, _15619_, _15058_);
  or _66646_ (_15640_, _15617_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _66647_ (_15641_, _15640_, _15615_);
  and _66648_ (_15642_, _15641_, _15639_);
  and _66649_ (_15643_, _15614_, _15549_);
  or _66650_ (_40841_, _15643_, _15642_);
  or _66651_ (_15644_, _15619_, _15256_);
  or _66652_ (_15645_, _15617_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _66653_ (_15646_, _15645_, _15615_);
  and _66654_ (_15647_, _15646_, _15644_);
  and _66655_ (_15648_, _15614_, _15555_);
  or _66656_ (_40842_, _15648_, _15647_);
  or _66657_ (_15649_, _15619_, _15454_);
  or _66658_ (_15650_, _15617_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _66659_ (_15651_, _15650_, _15615_);
  and _66660_ (_15652_, _15651_, _15649_);
  and _66661_ (_15653_, _15614_, _15561_);
  or _66662_ (_40843_, _15653_, _15652_);
  or _66663_ (_15654_, _15619_, _09197_);
  or _66664_ (_15655_, _15617_, \oc8051_golden_model_1.IRAM[4] [7]);
  and _66665_ (_15656_, _15655_, _15615_);
  and _66666_ (_15657_, _15656_, _15654_);
  and _66667_ (_15658_, _15614_, _09230_);
  or _66668_ (_40844_, _15658_, _15657_);
  and _66669_ (_15659_, _15616_, _15472_);
  not _66670_ (_15660_, _15659_);
  or _66671_ (_15661_, _15660_, _14247_);
  and _66672_ (_15662_, _15613_, _07356_);
  not _66673_ (_15663_, _15662_);
  or _66674_ (_15664_, _15659_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _66675_ (_15665_, _15664_, _15663_);
  and _66676_ (_15666_, _15665_, _15661_);
  and _66677_ (_15667_, _15662_, _15516_);
  or _66678_ (_40848_, _15667_, _15666_);
  or _66679_ (_15668_, _15660_, _14436_);
  or _66680_ (_15669_, _15659_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _66681_ (_15670_, _15669_, _15663_);
  and _66682_ (_15671_, _15670_, _15668_);
  and _66683_ (_15672_, _15662_, _15531_);
  or _66684_ (_40849_, _15672_, _15671_);
  or _66685_ (_15673_, _15660_, _14660_);
  or _66686_ (_15674_, _15659_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _66687_ (_15675_, _15674_, _15663_);
  and _66688_ (_15676_, _15675_, _15673_);
  and _66689_ (_15677_, _15662_, _15537_);
  or _66690_ (_40850_, _15677_, _15676_);
  or _66691_ (_15678_, _15660_, _14852_);
  or _66692_ (_15679_, _15659_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _66693_ (_15680_, _15679_, _15663_);
  and _66694_ (_15681_, _15680_, _15678_);
  and _66695_ (_15682_, _15662_, _15543_);
  or _66696_ (_40851_, _15682_, _15681_);
  or _66697_ (_15683_, _15660_, _15058_);
  or _66698_ (_15684_, _15659_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _66699_ (_15685_, _15684_, _15663_);
  and _66700_ (_15686_, _15685_, _15683_);
  and _66701_ (_15687_, _15662_, _15549_);
  or _66702_ (_40853_, _15687_, _15686_);
  or _66703_ (_15688_, _15660_, _15256_);
  or _66704_ (_15689_, _15659_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _66705_ (_15690_, _15689_, _15663_);
  and _66706_ (_15691_, _15690_, _15688_);
  and _66707_ (_15692_, _15662_, _15555_);
  or _66708_ (_40854_, _15692_, _15691_);
  or _66709_ (_15693_, _15660_, _15454_);
  or _66710_ (_15694_, _15659_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _66711_ (_15695_, _15694_, _15663_);
  and _66712_ (_15696_, _15695_, _15693_);
  and _66713_ (_15697_, _15662_, _15561_);
  or _66714_ (_40855_, _15697_, _15696_);
  or _66715_ (_15698_, _15660_, _09197_);
  or _66716_ (_15699_, _15659_, \oc8051_golden_model_1.IRAM[5] [7]);
  and _66717_ (_15700_, _15699_, _15663_);
  and _66718_ (_15701_, _15700_, _15698_);
  and _66719_ (_15702_, _15662_, _09230_);
  or _66720_ (_40856_, _15702_, _15701_);
  and _66721_ (_15703_, _15613_, _08399_);
  not _66722_ (_15704_, _15703_);
  and _66723_ (_15705_, _15616_, _15520_);
  or _66724_ (_15706_, _15705_, \oc8051_golden_model_1.IRAM[6] [0]);
  not _66725_ (_15707_, _15705_);
  or _66726_ (_15708_, _15707_, _14247_);
  and _66727_ (_15709_, _15708_, _15706_);
  and _66728_ (_15710_, _15709_, _15704_);
  and _66729_ (_15711_, _15703_, _15516_);
  or _66730_ (_40860_, _15711_, _15710_);
  or _66731_ (_15712_, _15707_, _14436_);
  or _66732_ (_15713_, _15705_, \oc8051_golden_model_1.IRAM[6] [1]);
  and _66733_ (_15714_, _15713_, _15704_);
  and _66734_ (_15715_, _15714_, _15712_);
  and _66735_ (_15716_, _15703_, _15531_);
  or _66736_ (_40861_, _15716_, _15715_);
  or _66737_ (_15717_, _15707_, _14660_);
  or _66738_ (_15718_, _15705_, \oc8051_golden_model_1.IRAM[6] [2]);
  and _66739_ (_15719_, _15718_, _15704_);
  and _66740_ (_15720_, _15719_, _15717_);
  and _66741_ (_15721_, _15703_, _15537_);
  or _66742_ (_40862_, _15721_, _15720_);
  or _66743_ (_15722_, _15707_, _14852_);
  or _66744_ (_15723_, _15705_, \oc8051_golden_model_1.IRAM[6] [3]);
  and _66745_ (_15724_, _15723_, _15704_);
  and _66746_ (_15725_, _15724_, _15722_);
  and _66747_ (_15726_, _15703_, _15543_);
  or _66748_ (_40863_, _15726_, _15725_);
  or _66749_ (_15727_, _15707_, _15058_);
  or _66750_ (_15728_, _15705_, \oc8051_golden_model_1.IRAM[6] [4]);
  and _66751_ (_15729_, _15728_, _15704_);
  and _66752_ (_15730_, _15729_, _15727_);
  and _66753_ (_15731_, _15703_, _15549_);
  or _66754_ (_40864_, _15731_, _15730_);
  or _66755_ (_15732_, _15707_, _15256_);
  or _66756_ (_15733_, _15705_, \oc8051_golden_model_1.IRAM[6] [5]);
  and _66757_ (_15734_, _15733_, _15704_);
  and _66758_ (_15735_, _15734_, _15732_);
  and _66759_ (_15736_, _15703_, _15555_);
  or _66760_ (_40865_, _15736_, _15735_);
  or _66761_ (_15737_, _15707_, _15454_);
  or _66762_ (_15738_, _15705_, \oc8051_golden_model_1.IRAM[6] [6]);
  and _66763_ (_15739_, _15738_, _15704_);
  and _66764_ (_15740_, _15739_, _15737_);
  and _66765_ (_15741_, _15703_, _15561_);
  or _66766_ (_40866_, _15741_, _15740_);
  and _66767_ (_15742_, _15705_, _09197_);
  nor _66768_ (_15743_, _15705_, _07751_);
  or _66769_ (_15744_, _15743_, _15703_);
  or _66770_ (_15745_, _15744_, _15742_);
  or _66771_ (_15746_, _15704_, _09230_);
  and _66772_ (_40867_, _15746_, _15745_);
  and _66773_ (_15747_, _15613_, _07080_);
  not _66774_ (_15748_, _15747_);
  or _66775_ (_15749_, _15748_, _15516_);
  and _66776_ (_15750_, _15616_, _07307_);
  and _66777_ (_15751_, _15750_, _14247_);
  nor _66778_ (_15752_, _15750_, _06895_);
  or _66779_ (_15753_, _15752_, _15747_);
  or _66780_ (_15754_, _15753_, _15751_);
  and _66781_ (_40872_, _15754_, _15749_);
  or _66782_ (_15755_, _15750_, \oc8051_golden_model_1.IRAM[7] [1]);
  and _66783_ (_15756_, _15755_, _15748_);
  not _66784_ (_15757_, _15750_);
  or _66785_ (_15758_, _15757_, _14436_);
  and _66786_ (_15759_, _15758_, _15756_);
  and _66787_ (_15760_, _15747_, _15531_);
  or _66788_ (_40873_, _15760_, _15759_);
  or _66789_ (_15761_, _15750_, \oc8051_golden_model_1.IRAM[7] [2]);
  and _66790_ (_15762_, _15761_, _15748_);
  or _66791_ (_15763_, _15757_, _14660_);
  and _66792_ (_15764_, _15763_, _15762_);
  and _66793_ (_15765_, _15747_, _15537_);
  or _66794_ (_40874_, _15765_, _15764_);
  or _66795_ (_15766_, _15750_, \oc8051_golden_model_1.IRAM[7] [3]);
  and _66796_ (_15767_, _15766_, _15748_);
  or _66797_ (_15768_, _15757_, _14852_);
  and _66798_ (_15769_, _15768_, _15767_);
  and _66799_ (_15770_, _15747_, _15543_);
  or _66800_ (_40876_, _15770_, _15769_);
  or _66801_ (_15771_, _15750_, \oc8051_golden_model_1.IRAM[7] [4]);
  and _66802_ (_15772_, _15771_, _15748_);
  or _66803_ (_15773_, _15757_, _15058_);
  and _66804_ (_15774_, _15773_, _15772_);
  and _66805_ (_15775_, _15747_, _15549_);
  or _66806_ (_40877_, _15775_, _15774_);
  or _66807_ (_15776_, _15750_, \oc8051_golden_model_1.IRAM[7] [5]);
  and _66808_ (_15777_, _15776_, _15748_);
  or _66809_ (_15778_, _15757_, _15256_);
  and _66810_ (_15779_, _15778_, _15777_);
  and _66811_ (_15780_, _15747_, _15555_);
  or _66812_ (_40878_, _15780_, _15779_);
  or _66813_ (_15781_, _15750_, \oc8051_golden_model_1.IRAM[7] [6]);
  and _66814_ (_15782_, _15781_, _15748_);
  or _66815_ (_15783_, _15757_, _15454_);
  and _66816_ (_15784_, _15783_, _15782_);
  and _66817_ (_15785_, _15747_, _15561_);
  or _66818_ (_40879_, _15785_, _15784_);
  or _66819_ (_15786_, _15750_, \oc8051_golden_model_1.IRAM[7] [7]);
  and _66820_ (_15787_, _15786_, _15748_);
  or _66821_ (_15788_, _15757_, _09197_);
  and _66822_ (_15789_, _15788_, _15787_);
  and _66823_ (_15790_, _15747_, _09230_);
  or _66824_ (_40880_, _15790_, _15789_);
  and _66825_ (_15791_, _14075_, _07614_);
  and _66826_ (_15792_, _15791_, _14078_);
  or _66827_ (_15793_, _15792_, \oc8051_golden_model_1.IRAM[8] [0]);
  not _66828_ (_15794_, _15792_);
  or _66829_ (_15795_, _15794_, _14247_);
  and _66830_ (_15796_, _15795_, _15793_);
  and _66831_ (_15797_, _07629_, _14449_);
  and _66832_ (_15798_, _15797_, _07081_);
  or _66833_ (_15799_, _15798_, _15796_);
  not _66834_ (_15800_, _15798_);
  or _66835_ (_15801_, _15800_, _15516_);
  and _66836_ (_40884_, _15801_, _15799_);
  or _66837_ (_15802_, _15794_, _14436_);
  or _66838_ (_15803_, _15792_, \oc8051_golden_model_1.IRAM[8] [1]);
  and _66839_ (_15804_, _15803_, _15800_);
  and _66840_ (_15805_, _15804_, _15802_);
  and _66841_ (_15806_, _15798_, _15531_);
  or _66842_ (_40885_, _15806_, _15805_);
  or _66843_ (_15807_, _15794_, _14660_);
  or _66844_ (_15808_, _15792_, \oc8051_golden_model_1.IRAM[8] [2]);
  and _66845_ (_15809_, _15808_, _15800_);
  and _66846_ (_15810_, _15809_, _15807_);
  and _66847_ (_15811_, _15798_, _15537_);
  or _66848_ (_40886_, _15811_, _15810_);
  or _66849_ (_15812_, _15794_, _14852_);
  or _66850_ (_15813_, _15792_, \oc8051_golden_model_1.IRAM[8] [3]);
  and _66851_ (_15814_, _15813_, _15800_);
  and _66852_ (_15815_, _15814_, _15812_);
  and _66853_ (_15816_, _15798_, _15543_);
  or _66854_ (_40887_, _15816_, _15815_);
  or _66855_ (_15817_, _15794_, _15058_);
  or _66856_ (_15818_, _15792_, \oc8051_golden_model_1.IRAM[8] [4]);
  and _66857_ (_15819_, _15818_, _15800_);
  and _66858_ (_15820_, _15819_, _15817_);
  and _66859_ (_15821_, _15798_, _15549_);
  or _66860_ (_40889_, _15821_, _15820_);
  or _66861_ (_15822_, _15794_, _15256_);
  or _66862_ (_15823_, _15792_, \oc8051_golden_model_1.IRAM[8] [5]);
  and _66863_ (_15824_, _15823_, _15800_);
  and _66864_ (_15825_, _15824_, _15822_);
  and _66865_ (_15826_, _15798_, _15555_);
  or _66866_ (_40890_, _15826_, _15825_);
  or _66867_ (_15827_, _15794_, _15454_);
  or _66868_ (_15828_, _15792_, \oc8051_golden_model_1.IRAM[8] [6]);
  and _66869_ (_15829_, _15828_, _15800_);
  and _66870_ (_15830_, _15829_, _15827_);
  and _66871_ (_15831_, _15798_, _15561_);
  or _66872_ (_40891_, _15831_, _15830_);
  or _66873_ (_15832_, _15794_, _09197_);
  or _66874_ (_15833_, _15792_, \oc8051_golden_model_1.IRAM[8] [7]);
  and _66875_ (_15834_, _15833_, _15800_);
  and _66876_ (_15835_, _15834_, _15832_);
  and _66877_ (_15836_, _15798_, _09230_);
  or _66878_ (_40892_, _15836_, _15835_);
  and _66879_ (_15837_, _15791_, _15472_);
  or _66880_ (_15838_, _15837_, \oc8051_golden_model_1.IRAM[9] [0]);
  not _66881_ (_15839_, _15837_);
  or _66882_ (_15840_, _15839_, _14247_);
  and _66883_ (_15841_, _15840_, _15838_);
  and _66884_ (_15842_, _15797_, _07356_);
  or _66885_ (_15843_, _15842_, _15841_);
  not _66886_ (_15844_, _15842_);
  or _66887_ (_15845_, _15844_, _15516_);
  and _66888_ (_40896_, _15845_, _15843_);
  or _66889_ (_15846_, _15839_, _14436_);
  or _66890_ (_15847_, _15837_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _66891_ (_15848_, _15847_, _15844_);
  and _66892_ (_15849_, _15848_, _15846_);
  and _66893_ (_15850_, _15842_, _15531_);
  or _66894_ (_40897_, _15850_, _15849_);
  or _66895_ (_15851_, _15839_, _14660_);
  or _66896_ (_15852_, _15837_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _66897_ (_15853_, _15852_, _15844_);
  and _66898_ (_15854_, _15853_, _15851_);
  and _66899_ (_15855_, _15842_, _15537_);
  or _66900_ (_40898_, _15855_, _15854_);
  or _66901_ (_15856_, _15839_, _14852_);
  or _66902_ (_15857_, _15837_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _66903_ (_15858_, _15857_, _15844_);
  and _66904_ (_15859_, _15858_, _15856_);
  and _66905_ (_15860_, _15842_, _15543_);
  or _66906_ (_40899_, _15860_, _15859_);
  or _66907_ (_15861_, _15839_, _15058_);
  or _66908_ (_15862_, _15837_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _66909_ (_15863_, _15862_, _15844_);
  and _66910_ (_15864_, _15863_, _15861_);
  and _66911_ (_15865_, _15842_, _15549_);
  or _66912_ (_40901_, _15865_, _15864_);
  or _66913_ (_15866_, _15839_, _15256_);
  or _66914_ (_15867_, _15837_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _66915_ (_15868_, _15867_, _15844_);
  and _66916_ (_15869_, _15868_, _15866_);
  and _66917_ (_15870_, _15842_, _15555_);
  or _66918_ (_40902_, _15870_, _15869_);
  or _66919_ (_15871_, _15839_, _15454_);
  or _66920_ (_15872_, _15837_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _66921_ (_15873_, _15872_, _15844_);
  and _66922_ (_15874_, _15873_, _15871_);
  and _66923_ (_15875_, _15842_, _15561_);
  or _66924_ (_40903_, _15875_, _15874_);
  nor _66925_ (_15876_, _15839_, _09197_);
  nor _66926_ (_15877_, _15837_, \oc8051_golden_model_1.IRAM[9] [7]);
  or _66927_ (_15878_, _15877_, _15876_);
  nor _66928_ (_15879_, _15878_, _15842_);
  and _66929_ (_15880_, _15842_, _09230_);
  or _66930_ (_40904_, _15880_, _15879_);
  and _66931_ (_15881_, _15791_, _15520_);
  not _66932_ (_15882_, _15881_);
  or _66933_ (_15883_, _15882_, _14247_);
  and _66934_ (_15884_, _15797_, _08399_);
  not _66935_ (_15885_, _15884_);
  or _66936_ (_15886_, _15881_, \oc8051_golden_model_1.IRAM[10] [0]);
  and _66937_ (_15887_, _15886_, _15885_);
  and _66938_ (_15888_, _15887_, _15883_);
  and _66939_ (_15889_, _15884_, _15516_);
  or _66940_ (_40908_, _15889_, _15888_);
  or _66941_ (_15890_, _15882_, _14436_);
  or _66942_ (_15891_, _15881_, \oc8051_golden_model_1.IRAM[10] [1]);
  and _66943_ (_15892_, _15891_, _15885_);
  and _66944_ (_15893_, _15892_, _15890_);
  and _66945_ (_15894_, _15884_, _15531_);
  or _66946_ (_40909_, _15894_, _15893_);
  or _66947_ (_15895_, _15882_, _14660_);
  or _66948_ (_15896_, _15881_, \oc8051_golden_model_1.IRAM[10] [2]);
  and _66949_ (_15897_, _15896_, _15885_);
  and _66950_ (_15898_, _15897_, _15895_);
  and _66951_ (_15899_, _15884_, _15537_);
  or _66952_ (_40910_, _15899_, _15898_);
  or _66953_ (_15900_, _15882_, _14852_);
  or _66954_ (_15901_, _15881_, \oc8051_golden_model_1.IRAM[10] [3]);
  and _66955_ (_15902_, _15901_, _15885_);
  and _66956_ (_15903_, _15902_, _15900_);
  and _66957_ (_15904_, _15884_, _15543_);
  or _66958_ (_40912_, _15904_, _15903_);
  or _66959_ (_15905_, _15882_, _15058_);
  or _66960_ (_15906_, _15881_, \oc8051_golden_model_1.IRAM[10] [4]);
  and _66961_ (_15907_, _15906_, _15885_);
  and _66962_ (_15908_, _15907_, _15905_);
  and _66963_ (_15909_, _15884_, _15549_);
  or _66964_ (_40913_, _15909_, _15908_);
  or _66965_ (_15910_, _15882_, _15256_);
  or _66966_ (_15911_, _15881_, \oc8051_golden_model_1.IRAM[10] [5]);
  and _66967_ (_15912_, _15911_, _15885_);
  and _66968_ (_15913_, _15912_, _15910_);
  and _66969_ (_15914_, _15884_, _15555_);
  or _66970_ (_40914_, _15914_, _15913_);
  or _66971_ (_15915_, _15882_, _15454_);
  or _66972_ (_15916_, _15881_, \oc8051_golden_model_1.IRAM[10] [6]);
  and _66973_ (_15917_, _15916_, _15885_);
  and _66974_ (_15918_, _15917_, _15915_);
  and _66975_ (_15919_, _15884_, _15561_);
  or _66976_ (_40915_, _15919_, _15918_);
  or _66977_ (_15920_, _15882_, _09197_);
  or _66978_ (_15921_, _15881_, \oc8051_golden_model_1.IRAM[10] [7]);
  and _66979_ (_15922_, _15921_, _15885_);
  and _66980_ (_15923_, _15922_, _15920_);
  and _66981_ (_15924_, _15884_, _09230_);
  or _66982_ (_40916_, _15924_, _15923_);
  not _66983_ (_15925_, _07229_);
  and _66984_ (_15926_, _14077_, _15925_);
  and _66985_ (_15927_, _15791_, _15926_);
  nor _66986_ (_15928_, _15927_, \oc8051_golden_model_1.IRAM[11] [0]);
  not _66987_ (_15929_, _15927_);
  nor _66988_ (_15930_, _15929_, _14247_);
  or _66989_ (_15931_, _15930_, _15928_);
  and _66990_ (_15932_, _15797_, _07080_);
  not _66991_ (_15933_, _15932_);
  nand _66992_ (_15934_, _15933_, _15931_);
  or _66993_ (_15935_, _15933_, _15516_);
  and _66994_ (_40919_, _15935_, _15934_);
  or _66995_ (_15936_, _15927_, \oc8051_golden_model_1.IRAM[11] [1]);
  and _66996_ (_15937_, _15936_, _15933_);
  or _66997_ (_15938_, _15929_, _14436_);
  and _66998_ (_15939_, _15938_, _15937_);
  and _66999_ (_15940_, _15932_, _15531_);
  or _67000_ (_40920_, _15940_, _15939_);
  or _67001_ (_15941_, _15927_, \oc8051_golden_model_1.IRAM[11] [2]);
  and _67002_ (_15942_, _15941_, _15933_);
  or _67003_ (_15943_, _15929_, _14660_);
  and _67004_ (_15944_, _15943_, _15942_);
  and _67005_ (_15945_, _15932_, _15537_);
  or _67006_ (_40921_, _15945_, _15944_);
  or _67007_ (_15946_, _15927_, \oc8051_golden_model_1.IRAM[11] [3]);
  and _67008_ (_15947_, _15946_, _15933_);
  or _67009_ (_15948_, _15929_, _14852_);
  and _67010_ (_15949_, _15948_, _15947_);
  and _67011_ (_15950_, _15932_, _15543_);
  or _67012_ (_40924_, _15950_, _15949_);
  or _67013_ (_15951_, _15927_, \oc8051_golden_model_1.IRAM[11] [4]);
  and _67014_ (_15952_, _15951_, _15933_);
  or _67015_ (_15953_, _15929_, _15058_);
  and _67016_ (_15954_, _15953_, _15952_);
  and _67017_ (_15955_, _15932_, _15549_);
  or _67018_ (_40925_, _15955_, _15954_);
  or _67019_ (_15956_, _15927_, \oc8051_golden_model_1.IRAM[11] [5]);
  and _67020_ (_15957_, _15956_, _15933_);
  or _67021_ (_15958_, _15929_, _15256_);
  and _67022_ (_15959_, _15958_, _15957_);
  and _67023_ (_15960_, _15932_, _15555_);
  or _67024_ (_40926_, _15960_, _15959_);
  or _67025_ (_15961_, _15927_, \oc8051_golden_model_1.IRAM[11] [6]);
  and _67026_ (_15962_, _15961_, _15933_);
  or _67027_ (_15963_, _15929_, _15454_);
  and _67028_ (_15964_, _15963_, _15962_);
  and _67029_ (_15965_, _15932_, _15561_);
  or _67030_ (_40927_, _15965_, _15964_);
  or _67031_ (_15966_, _15927_, \oc8051_golden_model_1.IRAM[11] [7]);
  and _67032_ (_15967_, _15966_, _15933_);
  or _67033_ (_15968_, _15929_, _09197_);
  and _67034_ (_15969_, _15968_, _15967_);
  and _67035_ (_15970_, _15932_, _09230_);
  or _67036_ (_40928_, _15970_, _15969_);
  not _67037_ (_15971_, _07614_);
  and _67038_ (_15972_, _14075_, _15971_);
  and _67039_ (_15973_, _14078_, _15972_);
  not _67040_ (_15974_, _15973_);
  or _67041_ (_15975_, _15974_, _14247_);
  or _67042_ (_15976_, _15973_, \oc8051_golden_model_1.IRAM[12] [0]);
  and _67043_ (_15977_, _15976_, _15975_);
  and _67044_ (_15978_, _07630_, _07081_);
  or _67045_ (_15979_, _15978_, _15977_);
  not _67046_ (_15980_, _15978_);
  or _67047_ (_15981_, _15980_, _15516_);
  and _67048_ (_40932_, _15981_, _15979_);
  and _67049_ (_15982_, _14078_, _07617_);
  or _67050_ (_15983_, _15982_, \oc8051_golden_model_1.IRAM[12] [1]);
  and _67051_ (_15984_, _15983_, _15980_);
  not _67052_ (_15985_, _15982_);
  or _67053_ (_15986_, _15985_, _14436_);
  and _67054_ (_15987_, _15986_, _15984_);
  and _67055_ (_15988_, _15978_, _15531_);
  or _67056_ (_40933_, _15988_, _15987_);
  or _67057_ (_15989_, _15982_, \oc8051_golden_model_1.IRAM[12] [2]);
  and _67058_ (_15990_, _15989_, _15980_);
  or _67059_ (_15991_, _15985_, _14660_);
  and _67060_ (_15992_, _15991_, _15990_);
  and _67061_ (_15993_, _15978_, _15537_);
  or _67062_ (_40934_, _15993_, _15992_);
  or _67063_ (_15994_, _15982_, \oc8051_golden_model_1.IRAM[12] [3]);
  and _67064_ (_15995_, _15994_, _15980_);
  or _67065_ (_15996_, _15985_, _14852_);
  and _67066_ (_15997_, _15996_, _15995_);
  and _67067_ (_15998_, _15978_, _15543_);
  or _67068_ (_40935_, _15998_, _15997_);
  or _67069_ (_15999_, _15982_, \oc8051_golden_model_1.IRAM[12] [4]);
  and _67070_ (_16000_, _15999_, _15980_);
  or _67071_ (_16001_, _15985_, _15058_);
  and _67072_ (_16002_, _16001_, _16000_);
  and _67073_ (_16003_, _15978_, _15549_);
  or _67074_ (_40936_, _16003_, _16002_);
  or _67075_ (_16004_, _15982_, \oc8051_golden_model_1.IRAM[12] [5]);
  and _67076_ (_16005_, _16004_, _15980_);
  or _67077_ (_16006_, _15985_, _15256_);
  and _67078_ (_16007_, _16006_, _16005_);
  and _67079_ (_16008_, _15978_, _15555_);
  or _67080_ (_40937_, _16008_, _16007_);
  or _67081_ (_16009_, _15982_, \oc8051_golden_model_1.IRAM[12] [6]);
  and _67082_ (_16010_, _16009_, _15980_);
  or _67083_ (_16011_, _15985_, _15454_);
  and _67084_ (_16012_, _16011_, _16010_);
  and _67085_ (_16013_, _15978_, _15561_);
  or _67086_ (_40939_, _16013_, _16012_);
  or _67087_ (_16014_, _15982_, \oc8051_golden_model_1.IRAM[12] [7]);
  and _67088_ (_16015_, _16014_, _15980_);
  or _67089_ (_16016_, _15985_, _09197_);
  and _67090_ (_16017_, _16016_, _16015_);
  and _67091_ (_16018_, _15978_, _09230_);
  or _67092_ (_40940_, _16018_, _16017_);
  and _67093_ (_16019_, _15472_, _15972_);
  not _67094_ (_16020_, _16019_);
  or _67095_ (_16021_, _16020_, _14247_);
  and _67096_ (_16022_, _07630_, _07356_);
  not _67097_ (_16023_, _16022_);
  or _67098_ (_16024_, _16019_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _67099_ (_16025_, _16024_, _16023_);
  and _67100_ (_16026_, _16025_, _16021_);
  and _67101_ (_16027_, _16022_, _15516_);
  or _67102_ (_40943_, _16027_, _16026_);
  and _67103_ (_16028_, _15472_, _07617_);
  or _67104_ (_16029_, _16028_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _67105_ (_16030_, _16029_, _16023_);
  not _67106_ (_16031_, _16028_);
  or _67107_ (_16032_, _16031_, _14436_);
  and _67108_ (_16033_, _16032_, _16030_);
  and _67109_ (_16034_, _16022_, _15531_);
  or _67110_ (_40945_, _16034_, _16033_);
  or _67111_ (_16035_, _16028_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _67112_ (_16036_, _16035_, _16023_);
  or _67113_ (_16037_, _16031_, _14660_);
  and _67114_ (_16038_, _16037_, _16036_);
  and _67115_ (_16039_, _16022_, _15537_);
  or _67116_ (_40946_, _16039_, _16038_);
  or _67117_ (_16040_, _16028_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _67118_ (_16041_, _16040_, _16023_);
  or _67119_ (_16042_, _16031_, _14852_);
  and _67120_ (_16043_, _16042_, _16041_);
  and _67121_ (_16044_, _16022_, _15543_);
  or _67122_ (_40947_, _16044_, _16043_);
  or _67123_ (_16045_, _16028_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _67124_ (_16046_, _16045_, _16023_);
  or _67125_ (_16047_, _16031_, _15058_);
  and _67126_ (_16048_, _16047_, _16046_);
  and _67127_ (_16049_, _16022_, _15549_);
  or _67128_ (_40948_, _16049_, _16048_);
  or _67129_ (_16050_, _16028_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _67130_ (_16051_, _16050_, _16023_);
  or _67131_ (_16052_, _16031_, _15256_);
  and _67132_ (_16053_, _16052_, _16051_);
  and _67133_ (_16054_, _16022_, _15555_);
  or _67134_ (_40949_, _16054_, _16053_);
  or _67135_ (_16055_, _16028_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _67136_ (_16056_, _16055_, _16023_);
  or _67137_ (_16057_, _16031_, _15454_);
  and _67138_ (_16058_, _16057_, _16056_);
  and _67139_ (_16059_, _16022_, _15561_);
  or _67140_ (_40951_, _16059_, _16058_);
  nor _67141_ (_16060_, _16019_, \oc8051_golden_model_1.IRAM[13] [7]);
  nor _67142_ (_16061_, _16020_, _09197_);
  or _67143_ (_16062_, _16061_, _16060_);
  nand _67144_ (_16063_, _16062_, _16023_);
  or _67145_ (_16064_, _16023_, _09230_);
  and _67146_ (_40952_, _16064_, _16063_);
  and _67147_ (_16065_, _15520_, _15972_);
  not _67148_ (_16066_, _16065_);
  or _67149_ (_16067_, _16066_, _14247_);
  and _67150_ (_16068_, _08399_, _07630_);
  not _67151_ (_16069_, _16068_);
  or _67152_ (_16070_, _16065_, \oc8051_golden_model_1.IRAM[14] [0]);
  and _67153_ (_16071_, _16070_, _16069_);
  and _67154_ (_16072_, _16071_, _16067_);
  and _67155_ (_16073_, _16068_, _15516_);
  or _67156_ (_40956_, _16073_, _16072_);
  and _67157_ (_16074_, _15520_, _07617_);
  or _67158_ (_16075_, _16074_, \oc8051_golden_model_1.IRAM[14] [1]);
  and _67159_ (_16076_, _16075_, _16069_);
  not _67160_ (_16077_, _16074_);
  or _67161_ (_16078_, _16077_, _14436_);
  and _67162_ (_16079_, _16078_, _16076_);
  and _67163_ (_16080_, _16068_, _15531_);
  or _67164_ (_40957_, _16080_, _16079_);
  or _67165_ (_16081_, _16074_, \oc8051_golden_model_1.IRAM[14] [2]);
  and _67166_ (_16082_, _16081_, _16069_);
  or _67167_ (_16083_, _16077_, _14660_);
  and _67168_ (_16084_, _16083_, _16082_);
  and _67169_ (_16085_, _16068_, _15537_);
  or _67170_ (_40958_, _16085_, _16084_);
  or _67171_ (_16086_, _16074_, \oc8051_golden_model_1.IRAM[14] [3]);
  and _67172_ (_16087_, _16086_, _16069_);
  or _67173_ (_16088_, _16077_, _14852_);
  and _67174_ (_16089_, _16088_, _16087_);
  and _67175_ (_16090_, _16068_, _15543_);
  or _67176_ (_40959_, _16090_, _16089_);
  or _67177_ (_16091_, _16074_, \oc8051_golden_model_1.IRAM[14] [4]);
  and _67178_ (_16092_, _16091_, _16069_);
  or _67179_ (_16093_, _16077_, _15058_);
  and _67180_ (_16094_, _16093_, _16092_);
  and _67181_ (_16095_, _16068_, _15549_);
  or _67182_ (_40960_, _16095_, _16094_);
  or _67183_ (_16096_, _16074_, \oc8051_golden_model_1.IRAM[14] [5]);
  and _67184_ (_16097_, _16096_, _16069_);
  or _67185_ (_16098_, _16077_, _15256_);
  and _67186_ (_16099_, _16098_, _16097_);
  and _67187_ (_16100_, _16068_, _15555_);
  or _67188_ (_40962_, _16100_, _16099_);
  or _67189_ (_16101_, _16074_, \oc8051_golden_model_1.IRAM[14] [6]);
  and _67190_ (_16102_, _16101_, _16069_);
  or _67191_ (_16103_, _16077_, _15454_);
  and _67192_ (_16104_, _16103_, _16102_);
  and _67193_ (_16105_, _16068_, _15561_);
  or _67194_ (_40963_, _16105_, _16104_);
  or _67195_ (_16106_, _16074_, \oc8051_golden_model_1.IRAM[14] [7]);
  and _67196_ (_16107_, _16106_, _16069_);
  or _67197_ (_16108_, _16077_, _09197_);
  and _67198_ (_16109_, _16108_, _16107_);
  and _67199_ (_16110_, _16068_, _09230_);
  or _67200_ (_40964_, _16110_, _16109_);
  nand _67201_ (_16111_, _15972_, _15926_);
  or _67202_ (_16112_, _14247_, _16111_);
  or _67203_ (_16113_, _07618_, \oc8051_golden_model_1.IRAM[15] [0]);
  and _67204_ (_16114_, _16113_, _07632_);
  and _67205_ (_16115_, _16114_, _16112_);
  and _67206_ (_16116_, _15516_, _07631_);
  or _67207_ (_40967_, _16116_, _16115_);
  or _67208_ (_16117_, _07618_, \oc8051_golden_model_1.IRAM[15] [1]);
  and _67209_ (_16118_, _16117_, _07632_);
  or _67210_ (_16119_, _14436_, _07634_);
  and _67211_ (_16120_, _16119_, _16118_);
  and _67212_ (_16121_, _15531_, _07631_);
  or _67213_ (_40968_, _16121_, _16120_);
  or _67214_ (_16122_, _07618_, \oc8051_golden_model_1.IRAM[15] [2]);
  and _67215_ (_16123_, _16122_, _07632_);
  or _67216_ (_16124_, _14660_, _07634_);
  and _67217_ (_16125_, _16124_, _16123_);
  and _67218_ (_16126_, _15537_, _07631_);
  or _67219_ (_40969_, _16126_, _16125_);
  or _67220_ (_16127_, _07618_, \oc8051_golden_model_1.IRAM[15] [3]);
  and _67221_ (_16128_, _16127_, _07632_);
  or _67222_ (_16129_, _14852_, _07634_);
  and _67223_ (_16130_, _16129_, _16128_);
  and _67224_ (_16131_, _15543_, _07631_);
  or _67225_ (_40970_, _16131_, _16130_);
  or _67226_ (_16132_, _07618_, \oc8051_golden_model_1.IRAM[15] [4]);
  and _67227_ (_16133_, _16132_, _07632_);
  or _67228_ (_16134_, _15058_, _07634_);
  and _67229_ (_16135_, _16134_, _16133_);
  and _67230_ (_16136_, _15549_, _07631_);
  or _67231_ (_40971_, _16136_, _16135_);
  or _67232_ (_16137_, _15256_, _07634_);
  or _67233_ (_16138_, _07618_, \oc8051_golden_model_1.IRAM[15] [5]);
  and _67234_ (_16139_, _16138_, _07632_);
  and _67235_ (_16140_, _16139_, _16137_);
  and _67236_ (_16141_, _15555_, _07631_);
  or _67237_ (_40972_, _16141_, _16140_);
  or _67238_ (_16142_, _15454_, _07634_);
  or _67239_ (_16143_, _07618_, \oc8051_golden_model_1.IRAM[15] [6]);
  and _67240_ (_16144_, _16143_, _07632_);
  and _67241_ (_16145_, _16144_, _16142_);
  and _67242_ (_16146_, _15561_, _07631_);
  or _67243_ (_40973_, _16146_, _16145_);
  nor _67244_ (_16147_, _01336_, _09877_);
  nor _67245_ (_16148_, _07698_, _09877_);
  and _67246_ (_16149_, _07698_, _08672_);
  or _67247_ (_16150_, _16149_, _16148_);
  or _67248_ (_16151_, _16150_, _06020_);
  and _67249_ (_16152_, _14186_, _07698_);
  or _67250_ (_16153_, _16152_, _16148_);
  and _67251_ (_16154_, _16153_, _09833_);
  nor _67252_ (_16155_, _08127_, _09258_);
  or _67253_ (_16156_, _16155_, _16148_);
  and _67254_ (_16157_, _16156_, _06102_);
  nor _67255_ (_16158_, _06938_, _09877_);
  and _67256_ (_16159_, _07698_, \oc8051_golden_model_1.ACC [0]);
  or _67257_ (_16160_, _16159_, _16148_);
  and _67258_ (_16161_, _16160_, _06938_);
  or _67259_ (_16162_, _16161_, _16158_);
  and _67260_ (_16163_, _16162_, _06954_);
  or _67261_ (_16164_, _16163_, _06043_);
  or _67262_ (_16165_, _16164_, _16157_);
  and _67263_ (_16166_, _14102_, _08361_);
  nor _67264_ (_16167_, _08361_, _09877_);
  or _67265_ (_16168_, _16167_, _06044_);
  or _67266_ (_16169_, _16168_, _16166_);
  and _67267_ (_16170_, _16169_, _16165_);
  or _67268_ (_16171_, _16170_, _06239_);
  and _67269_ (_16172_, _07698_, _06931_);
  or _67270_ (_16173_, _16172_, _16148_);
  or _67271_ (_16174_, _16173_, _06848_);
  and _67272_ (_16175_, _16174_, _16171_);
  or _67273_ (_16176_, _16175_, _06219_);
  or _67274_ (_16177_, _16160_, _06220_);
  and _67275_ (_16178_, _16177_, _06040_);
  and _67276_ (_16179_, _16178_, _16176_);
  and _67277_ (_16180_, _16148_, _06039_);
  or _67278_ (_16181_, _16180_, _06032_);
  or _67279_ (_16182_, _16181_, _16179_);
  or _67280_ (_16183_, _16156_, _06033_);
  and _67281_ (_16184_, _16183_, _16182_);
  or _67282_ (_16185_, _16184_, _09269_);
  nor _67283_ (_16186_, _09765_, _09763_);
  nor _67284_ (_16187_, _16186_, _09766_);
  or _67285_ (_16188_, _16187_, _09800_);
  and _67286_ (_16189_, _16188_, _06027_);
  and _67287_ (_16190_, _16189_, _16185_);
  and _67288_ (_16191_, _14132_, _08361_);
  or _67289_ (_16192_, _16191_, _16167_);
  and _67290_ (_16193_, _16192_, _06026_);
  or _67291_ (_16194_, _16193_, _09818_);
  or _67292_ (_16195_, _16194_, _16190_);
  and _67293_ (_16196_, _09120_, _07698_);
  or _67294_ (_16197_, _16148_, _07012_);
  or _67295_ (_16198_, _16197_, _16196_);
  or _67296_ (_16199_, _16173_, _09827_);
  and _67297_ (_16200_, _16199_, _05669_);
  and _67298_ (_16201_, _16200_, _16198_);
  and _67299_ (_16202_, _16201_, _16195_);
  or _67300_ (_16203_, _16202_, _16154_);
  and _67301_ (_16204_, _16203_, _09839_);
  nand _67302_ (_16205_, _10184_, _05758_);
  or _67303_ (_16206_, _10178_, _10133_);
  or _67304_ (_16207_, _10184_, _16206_);
  and _67305_ (_16208_, _16207_, _09832_);
  and _67306_ (_16209_, _16208_, _16205_);
  or _67307_ (_16210_, _16209_, _06019_);
  or _67308_ (_16211_, _16210_, _16204_);
  and _67309_ (_16212_, _16211_, _16151_);
  or _67310_ (_16213_, _16212_, _06112_);
  and _67311_ (_16214_, _14086_, _07698_);
  or _67312_ (_16215_, _16148_, _08751_);
  or _67313_ (_16216_, _16215_, _16214_);
  and _67314_ (_16217_, _16216_, _08756_);
  and _67315_ (_16218_, _16217_, _16213_);
  nor _67316_ (_16219_, _12302_, _09258_);
  or _67317_ (_16220_, _16219_, _16148_);
  nand _67318_ (_16221_, _10995_, _07698_);
  and _67319_ (_16222_, _16221_, _06284_);
  and _67320_ (_16223_, _16222_, _16220_);
  or _67321_ (_16224_, _16223_, _16218_);
  and _67322_ (_16225_, _16224_, _07032_);
  nand _67323_ (_16226_, _16150_, _06108_);
  nor _67324_ (_16227_, _16226_, _16155_);
  or _67325_ (_16228_, _16227_, _06277_);
  or _67326_ (_16229_, _16228_, _16225_);
  nor _67327_ (_16230_, _16148_, _06278_);
  nand _67328_ (_16231_, _16230_, _16221_);
  and _67329_ (_16232_, _16231_, _16229_);
  or _67330_ (_16233_, _16232_, _06130_);
  and _67331_ (_16234_, _14083_, _07698_);
  or _67332_ (_16235_, _16148_, _08777_);
  or _67333_ (_16236_, _16235_, _16234_);
  and _67334_ (_16237_, _16236_, _08782_);
  and _67335_ (_16238_, _16237_, _16233_);
  and _67336_ (_16239_, _16220_, _06292_);
  or _67337_ (_16240_, _16239_, _06316_);
  or _67338_ (_16241_, _16240_, _16238_);
  or _67339_ (_16242_, _16156_, _06718_);
  and _67340_ (_16243_, _16242_, _16241_);
  or _67341_ (_16244_, _16243_, _05652_);
  or _67342_ (_16245_, _16148_, _05653_);
  and _67343_ (_16246_, _16245_, _16244_);
  or _67344_ (_16247_, _16246_, _06047_);
  or _67345_ (_16248_, _16156_, _06048_);
  and _67346_ (_16249_, _16248_, _01336_);
  and _67347_ (_16250_, _16249_, _16247_);
  or _67348_ (_16251_, _16250_, _16147_);
  and _67349_ (_43324_, _16251_, _42882_);
  nor _67350_ (_16252_, _01336_, _09842_);
  nor _67351_ (_16253_, _07698_, _09842_);
  nor _67352_ (_16254_, _10993_, _09258_);
  or _67353_ (_16255_, _16254_, _16253_);
  or _67354_ (_16256_, _16255_, _08782_);
  nor _67355_ (_16257_, _08361_, _09842_);
  and _67356_ (_16258_, _14273_, _08361_);
  or _67357_ (_16259_, _16258_, _16257_);
  and _67358_ (_16260_, _16259_, _06039_);
  nor _67359_ (_16261_, _09258_, _07132_);
  or _67360_ (_16262_, _16261_, _16253_);
  or _67361_ (_16263_, _16262_, _06848_);
  or _67362_ (_16264_, _07698_, \oc8051_golden_model_1.B [1]);
  and _67363_ (_16265_, _14284_, _07698_);
  not _67364_ (_16266_, _16265_);
  and _67365_ (_16267_, _16266_, _16264_);
  or _67366_ (_16268_, _16267_, _06954_);
  and _67367_ (_16269_, _07698_, \oc8051_golden_model_1.ACC [1]);
  or _67368_ (_16270_, _16269_, _16253_);
  and _67369_ (_16271_, _16270_, _06938_);
  nor _67370_ (_16272_, _06938_, _09842_);
  or _67371_ (_16273_, _16272_, _06102_);
  or _67372_ (_16274_, _16273_, _16271_);
  and _67373_ (_16275_, _16274_, _06044_);
  and _67374_ (_16276_, _16275_, _16268_);
  and _67375_ (_16277_, _14266_, _08361_);
  or _67376_ (_16278_, _16277_, _16257_);
  and _67377_ (_16279_, _16278_, _06043_);
  or _67378_ (_16280_, _16279_, _06239_);
  or _67379_ (_16281_, _16280_, _16276_);
  and _67380_ (_16282_, _16281_, _16263_);
  or _67381_ (_16283_, _16282_, _06219_);
  or _67382_ (_16284_, _16270_, _06220_);
  and _67383_ (_16285_, _16284_, _06040_);
  and _67384_ (_16286_, _16285_, _16283_);
  or _67385_ (_16287_, _16286_, _16260_);
  and _67386_ (_16288_, _16287_, _06033_);
  and _67387_ (_16289_, _16277_, _14302_);
  or _67388_ (_16290_, _16289_, _16257_);
  and _67389_ (_16291_, _16290_, _06032_);
  or _67390_ (_16292_, _16291_, _09269_);
  or _67391_ (_16293_, _16292_, _16288_);
  nor _67392_ (_16294_, _09768_, _09699_);
  nor _67393_ (_16295_, _16294_, _09769_);
  or _67394_ (_16296_, _16295_, _09800_);
  and _67395_ (_16297_, _16296_, _06027_);
  and _67396_ (_16298_, _16297_, _16293_);
  or _67397_ (_16299_, _16257_, _14267_);
  and _67398_ (_16300_, _16299_, _06026_);
  and _67399_ (_16301_, _16300_, _16278_);
  or _67400_ (_16302_, _16301_, _09818_);
  or _67401_ (_16303_, _16302_, _16298_);
  and _67402_ (_16304_, _09075_, _07698_);
  or _67403_ (_16305_, _16253_, _07012_);
  or _67404_ (_16306_, _16305_, _16304_);
  or _67405_ (_16307_, _16262_, _09827_);
  and _67406_ (_16308_, _16307_, _05669_);
  and _67407_ (_16309_, _16308_, _16306_);
  and _67408_ (_16310_, _16309_, _16303_);
  or _67409_ (_16311_, _14367_, _09258_);
  and _67410_ (_16312_, _16264_, _09833_);
  and _67411_ (_16313_, _16312_, _16311_);
  or _67412_ (_16314_, _16313_, _09832_);
  or _67413_ (_16315_, _16314_, _16310_);
  nor _67414_ (_16316_, _10179_, _10177_);
  or _67415_ (_16317_, _16316_, _10180_);
  nor _67416_ (_16318_, _16317_, _10184_);
  and _67417_ (_16319_, _10184_, _10130_);
  or _67418_ (_16320_, _16319_, _16318_);
  or _67419_ (_16321_, _16320_, _09839_);
  and _67420_ (_16322_, _16321_, _06020_);
  and _67421_ (_16323_, _16322_, _16315_);
  nand _67422_ (_16324_, _07698_, _06832_);
  and _67423_ (_16325_, _16264_, _06019_);
  and _67424_ (_16326_, _16325_, _16324_);
  or _67425_ (_16327_, _16326_, _16323_);
  and _67426_ (_16328_, _16327_, _08751_);
  or _67427_ (_16329_, _14263_, _09258_);
  and _67428_ (_16330_, _16264_, _06112_);
  and _67429_ (_16331_, _16330_, _16329_);
  or _67430_ (_16332_, _16331_, _06284_);
  or _67431_ (_16333_, _16332_, _16328_);
  and _67432_ (_16334_, _10994_, _07698_);
  or _67433_ (_16335_, _16334_, _16253_);
  or _67434_ (_16336_, _16335_, _08756_);
  and _67435_ (_16337_, _16336_, _07032_);
  and _67436_ (_16338_, _16337_, _16333_);
  or _67437_ (_16339_, _14261_, _09258_);
  and _67438_ (_16340_, _16264_, _06108_);
  and _67439_ (_16341_, _16340_, _16339_);
  or _67440_ (_16342_, _16341_, _06277_);
  or _67441_ (_16343_, _16342_, _16338_);
  and _67442_ (_16344_, _16269_, _08078_);
  or _67443_ (_16345_, _16253_, _06278_);
  or _67444_ (_16346_, _16345_, _16344_);
  and _67445_ (_16347_, _16346_, _08777_);
  and _67446_ (_16348_, _16347_, _16343_);
  or _67447_ (_16349_, _16324_, _08078_);
  and _67448_ (_16350_, _16264_, _06130_);
  and _67449_ (_16351_, _16350_, _16349_);
  or _67450_ (_16352_, _16351_, _06292_);
  or _67451_ (_16353_, _16352_, _16348_);
  and _67452_ (_16354_, _16353_, _16256_);
  or _67453_ (_16355_, _16354_, _06316_);
  or _67454_ (_16356_, _16267_, _06718_);
  and _67455_ (_16357_, _16356_, _05653_);
  and _67456_ (_16358_, _16357_, _16355_);
  and _67457_ (_16359_, _16259_, _05652_);
  or _67458_ (_16360_, _16359_, _06047_);
  or _67459_ (_16361_, _16360_, _16358_);
  or _67460_ (_16362_, _16253_, _06048_);
  or _67461_ (_16363_, _16362_, _16265_);
  and _67462_ (_16364_, _16363_, _01336_);
  and _67463_ (_16365_, _16364_, _16361_);
  or _67464_ (_16366_, _16365_, _16252_);
  and _67465_ (_43325_, _16366_, _42882_);
  nor _67466_ (_16367_, _01336_, _10002_);
  nor _67467_ (_16368_, _07698_, _10002_);
  and _67468_ (_16369_, _07698_, _08730_);
  or _67469_ (_16370_, _16369_, _16368_);
  or _67470_ (_16371_, _16370_, _06020_);
  and _67471_ (_16372_, _14580_, _07698_);
  or _67472_ (_16373_, _16372_, _16368_);
  and _67473_ (_16374_, _16373_, _09833_);
  nor _67474_ (_16375_, _08361_, _10002_);
  and _67475_ (_16376_, _14479_, _08361_);
  or _67476_ (_16377_, _16376_, _16375_);
  and _67477_ (_16378_, _16377_, _06039_);
  and _67478_ (_16379_, _14493_, _07698_);
  or _67479_ (_16380_, _16379_, _16368_);
  and _67480_ (_16381_, _16380_, _06102_);
  nor _67481_ (_16382_, _06938_, _10002_);
  and _67482_ (_16383_, _07698_, \oc8051_golden_model_1.ACC [2]);
  or _67483_ (_16384_, _16383_, _16368_);
  and _67484_ (_16385_, _16384_, _06938_);
  or _67485_ (_16386_, _16385_, _16382_);
  and _67486_ (_16387_, _16386_, _06954_);
  or _67487_ (_16388_, _16387_, _06043_);
  or _67488_ (_16389_, _16388_, _16381_);
  and _67489_ (_16390_, _14497_, _08361_);
  or _67490_ (_16391_, _16390_, _16375_);
  or _67491_ (_16392_, _16391_, _06044_);
  and _67492_ (_16393_, _16392_, _06848_);
  and _67493_ (_16394_, _16393_, _16389_);
  nor _67494_ (_16395_, _09258_, _07530_);
  or _67495_ (_16396_, _16395_, _16368_);
  and _67496_ (_16397_, _16396_, _06239_);
  or _67497_ (_16398_, _16397_, _06219_);
  or _67498_ (_16399_, _16398_, _16394_);
  or _67499_ (_16400_, _16384_, _06220_);
  and _67500_ (_16401_, _16400_, _06040_);
  and _67501_ (_16402_, _16401_, _16399_);
  or _67502_ (_16403_, _16402_, _16378_);
  and _67503_ (_16404_, _16403_, _06033_);
  or _67504_ (_16405_, _16375_, _14512_);
  and _67505_ (_16406_, _16391_, _06032_);
  and _67506_ (_16407_, _16406_, _16405_);
  or _67507_ (_16408_, _16407_, _09269_);
  or _67508_ (_16409_, _16408_, _16404_);
  or _67509_ (_16410_, _09770_, _09652_);
  and _67510_ (_16411_, _16410_, _09771_);
  or _67511_ (_16412_, _16411_, _09800_);
  and _67512_ (_16413_, _16412_, _06027_);
  and _67513_ (_16414_, _16413_, _16409_);
  or _67514_ (_16415_, _16375_, _14525_);
  and _67515_ (_16416_, _16415_, _06026_);
  and _67516_ (_16417_, _16416_, _16391_);
  or _67517_ (_16418_, _16417_, _09818_);
  or _67518_ (_16419_, _16418_, _16414_);
  and _67519_ (_16420_, _09182_, _07698_);
  or _67520_ (_16421_, _16368_, _07012_);
  or _67521_ (_16422_, _16421_, _16420_);
  or _67522_ (_16423_, _16396_, _09827_);
  and _67523_ (_16424_, _16423_, _05669_);
  and _67524_ (_16425_, _16424_, _16422_);
  and _67525_ (_16426_, _16425_, _16419_);
  or _67526_ (_16427_, _16426_, _16374_);
  and _67527_ (_16428_, _16427_, _09839_);
  nor _67528_ (_16429_, _10180_, _10131_);
  not _67529_ (_16430_, _16429_);
  and _67530_ (_16431_, _16430_, _10124_);
  nor _67531_ (_16432_, _16430_, _10124_);
  nor _67532_ (_16433_, _16432_, _16431_);
  or _67533_ (_16434_, _16433_, _10184_);
  nand _67534_ (_16435_, _10184_, _10121_);
  and _67535_ (_16436_, _16435_, _09832_);
  and _67536_ (_16437_, _16436_, _16434_);
  or _67537_ (_16438_, _16437_, _06019_);
  or _67538_ (_16439_, _16438_, _16428_);
  and _67539_ (_16440_, _16439_, _16371_);
  or _67540_ (_16441_, _16440_, _06112_);
  and _67541_ (_16442_, _14596_, _07698_);
  or _67542_ (_16443_, _16442_, _16368_);
  or _67543_ (_16444_, _16443_, _08751_);
  and _67544_ (_16445_, _16444_, _08756_);
  and _67545_ (_16446_, _16445_, _16441_);
  and _67546_ (_16447_, _10991_, _07698_);
  or _67547_ (_16448_, _16447_, _16368_);
  and _67548_ (_16449_, _16448_, _06284_);
  or _67549_ (_16450_, _16449_, _16446_);
  and _67550_ (_16451_, _16450_, _07032_);
  or _67551_ (_16452_, _16368_, _08177_);
  and _67552_ (_16453_, _16370_, _06108_);
  and _67553_ (_16454_, _16453_, _16452_);
  or _67554_ (_16455_, _16454_, _16451_);
  and _67555_ (_16456_, _16455_, _06278_);
  and _67556_ (_16457_, _16384_, _06277_);
  and _67557_ (_16458_, _16457_, _16452_);
  or _67558_ (_16459_, _16458_, _06130_);
  or _67559_ (_16460_, _16459_, _16456_);
  and _67560_ (_16461_, _14593_, _07698_);
  or _67561_ (_16462_, _16368_, _08777_);
  or _67562_ (_16463_, _16462_, _16461_);
  and _67563_ (_16464_, _16463_, _08782_);
  and _67564_ (_16465_, _16464_, _16460_);
  nor _67565_ (_16466_, _10990_, _09258_);
  or _67566_ (_16467_, _16466_, _16368_);
  and _67567_ (_16468_, _16467_, _06292_);
  or _67568_ (_16469_, _16468_, _06316_);
  or _67569_ (_16470_, _16469_, _16465_);
  or _67570_ (_16471_, _16380_, _06718_);
  and _67571_ (_16472_, _16471_, _05653_);
  and _67572_ (_16473_, _16472_, _16470_);
  and _67573_ (_16474_, _16377_, _05652_);
  or _67574_ (_16475_, _16474_, _06047_);
  or _67575_ (_16476_, _16475_, _16473_);
  and _67576_ (_16477_, _14657_, _07698_);
  or _67577_ (_16478_, _16368_, _06048_);
  or _67578_ (_16479_, _16478_, _16477_);
  and _67579_ (_16480_, _16479_, _01336_);
  and _67580_ (_16481_, _16480_, _16476_);
  or _67581_ (_16482_, _16481_, _16367_);
  and _67582_ (_43326_, _16482_, _42882_);
  nor _67583_ (_16483_, _01336_, _09927_);
  nor _67584_ (_16484_, _07698_, _09927_);
  and _67585_ (_16485_, _07698_, _08662_);
  or _67586_ (_16486_, _16485_, _16484_);
  or _67587_ (_16487_, _16486_, _06020_);
  and _67588_ (_16488_, _14778_, _07698_);
  or _67589_ (_16489_, _16488_, _16484_);
  and _67590_ (_16490_, _16489_, _09833_);
  nor _67591_ (_16491_, _08361_, _09927_);
  and _67592_ (_16492_, _14683_, _08361_);
  or _67593_ (_16493_, _16492_, _16491_);
  or _67594_ (_16494_, _16491_, _14708_);
  and _67595_ (_16495_, _16494_, _16493_);
  or _67596_ (_16496_, _16495_, _06033_);
  and _67597_ (_16497_, _14672_, _07698_);
  or _67598_ (_16498_, _16497_, _16484_);
  or _67599_ (_16499_, _16498_, _06954_);
  and _67600_ (_16500_, _07698_, \oc8051_golden_model_1.ACC [3]);
  or _67601_ (_16501_, _16500_, _16484_);
  and _67602_ (_16502_, _16501_, _06938_);
  nor _67603_ (_16503_, _06938_, _09927_);
  or _67604_ (_16504_, _16503_, _06102_);
  or _67605_ (_16505_, _16504_, _16502_);
  and _67606_ (_16506_, _16505_, _06044_);
  and _67607_ (_16507_, _16506_, _16499_);
  and _67608_ (_16508_, _16493_, _06043_);
  or _67609_ (_16509_, _16508_, _06239_);
  or _67610_ (_16510_, _16509_, _16507_);
  nor _67611_ (_16511_, _09258_, _07353_);
  or _67612_ (_16512_, _16511_, _16484_);
  or _67613_ (_16513_, _16512_, _06848_);
  and _67614_ (_16514_, _16513_, _16510_);
  or _67615_ (_16515_, _16514_, _06219_);
  or _67616_ (_16516_, _16501_, _06220_);
  and _67617_ (_16517_, _16516_, _06040_);
  and _67618_ (_16518_, _16517_, _16515_);
  and _67619_ (_16519_, _14681_, _08361_);
  or _67620_ (_16520_, _16519_, _16491_);
  and _67621_ (_16521_, _16520_, _06039_);
  or _67622_ (_16522_, _16521_, _06032_);
  or _67623_ (_16523_, _16522_, _16518_);
  and _67624_ (_16524_, _16523_, _16496_);
  or _67625_ (_16525_, _16524_, _09269_);
  nor _67626_ (_16526_, _09773_, _09594_);
  nor _67627_ (_16527_, _16526_, _09774_);
  or _67628_ (_16528_, _16527_, _09800_);
  and _67629_ (_16529_, _16528_, _06027_);
  and _67630_ (_16530_, _16529_, _16525_);
  and _67631_ (_16531_, _14724_, _08361_);
  or _67632_ (_16532_, _16531_, _16491_);
  and _67633_ (_16533_, _16532_, _06026_);
  or _67634_ (_16534_, _16533_, _09818_);
  or _67635_ (_16535_, _16534_, _16530_);
  and _67636_ (_16536_, _09181_, _07698_);
  or _67637_ (_16537_, _16484_, _07012_);
  or _67638_ (_16538_, _16537_, _16536_);
  or _67639_ (_16539_, _16512_, _09827_);
  and _67640_ (_16540_, _16539_, _05669_);
  and _67641_ (_16541_, _16540_, _16538_);
  and _67642_ (_16542_, _16541_, _16535_);
  or _67643_ (_16543_, _16542_, _16490_);
  and _67644_ (_16544_, _16543_, _09839_);
  nor _67645_ (_16545_, _16431_, _10123_);
  nor _67646_ (_16546_, _16545_, _10115_);
  and _67647_ (_16547_, _16545_, _10115_);
  or _67648_ (_16548_, _16547_, _16546_);
  or _67649_ (_16549_, _16548_, _10184_);
  not _67650_ (_16550_, _10112_);
  nand _67651_ (_16551_, _10184_, _16550_);
  and _67652_ (_16552_, _16551_, _09832_);
  and _67653_ (_16553_, _16552_, _16549_);
  or _67654_ (_16554_, _16553_, _06019_);
  or _67655_ (_16555_, _16554_, _16544_);
  and _67656_ (_16556_, _16555_, _16487_);
  or _67657_ (_16557_, _16556_, _06112_);
  and _67658_ (_16558_, _14793_, _07698_);
  or _67659_ (_16559_, _16484_, _08751_);
  or _67660_ (_16560_, _16559_, _16558_);
  and _67661_ (_16561_, _16560_, _08756_);
  and _67662_ (_16562_, _16561_, _16557_);
  and _67663_ (_16563_, _12299_, _07698_);
  or _67664_ (_16564_, _16563_, _16484_);
  and _67665_ (_16565_, _16564_, _06284_);
  or _67666_ (_16566_, _16565_, _16562_);
  and _67667_ (_16567_, _16566_, _07032_);
  or _67668_ (_16568_, _16484_, _08029_);
  and _67669_ (_16569_, _16486_, _06108_);
  and _67670_ (_16570_, _16569_, _16568_);
  or _67671_ (_16571_, _16570_, _16567_);
  and _67672_ (_16572_, _16571_, _06278_);
  and _67673_ (_16573_, _16501_, _06277_);
  and _67674_ (_16574_, _16573_, _16568_);
  or _67675_ (_16575_, _16574_, _06130_);
  or _67676_ (_16576_, _16575_, _16572_);
  and _67677_ (_16577_, _14792_, _07698_);
  or _67678_ (_16578_, _16484_, _08777_);
  or _67679_ (_16579_, _16578_, _16577_);
  and _67680_ (_16580_, _16579_, _08782_);
  and _67681_ (_16581_, _16580_, _16576_);
  nor _67682_ (_16582_, _10988_, _09258_);
  or _67683_ (_16583_, _16582_, _16484_);
  and _67684_ (_16584_, _16583_, _06292_);
  or _67685_ (_16585_, _16584_, _06316_);
  or _67686_ (_16586_, _16585_, _16581_);
  or _67687_ (_16587_, _16498_, _06718_);
  and _67688_ (_16588_, _16587_, _05653_);
  and _67689_ (_16589_, _16588_, _16586_);
  and _67690_ (_16590_, _16520_, _05652_);
  or _67691_ (_16591_, _16590_, _06047_);
  or _67692_ (_16592_, _16591_, _16589_);
  and _67693_ (_16593_, _14849_, _07698_);
  or _67694_ (_16594_, _16484_, _06048_);
  or _67695_ (_16595_, _16594_, _16593_);
  and _67696_ (_16596_, _16595_, _01336_);
  and _67697_ (_16597_, _16596_, _16592_);
  or _67698_ (_16598_, _16597_, _16483_);
  and _67699_ (_43327_, _16598_, _42882_);
  nor _67700_ (_16599_, _01336_, _09854_);
  nor _67701_ (_16600_, _07698_, _09854_);
  and _67702_ (_16601_, _08665_, _07698_);
  or _67703_ (_16602_, _16601_, _16600_);
  or _67704_ (_16603_, _16602_, _06020_);
  and _67705_ (_16604_, _14983_, _07698_);
  or _67706_ (_16605_, _16604_, _16600_);
  and _67707_ (_16606_, _16605_, _09833_);
  nor _67708_ (_16607_, _08361_, _09854_);
  and _67709_ (_16608_, _14882_, _08361_);
  or _67710_ (_16609_, _16608_, _16607_);
  and _67711_ (_16610_, _16609_, _06039_);
  and _67712_ (_16611_, _14887_, _07698_);
  or _67713_ (_16612_, _16611_, _16600_);
  or _67714_ (_16613_, _16612_, _06954_);
  and _67715_ (_16614_, _07698_, \oc8051_golden_model_1.ACC [4]);
  or _67716_ (_16615_, _16614_, _16600_);
  and _67717_ (_16616_, _16615_, _06938_);
  nor _67718_ (_16617_, _06938_, _09854_);
  or _67719_ (_16618_, _16617_, _06102_);
  or _67720_ (_16619_, _16618_, _16616_);
  and _67721_ (_16620_, _16619_, _06044_);
  and _67722_ (_16621_, _16620_, _16613_);
  and _67723_ (_16622_, _14878_, _08361_);
  or _67724_ (_16623_, _16622_, _16607_);
  and _67725_ (_16624_, _16623_, _06043_);
  or _67726_ (_16625_, _16624_, _06239_);
  or _67727_ (_16626_, _16625_, _16621_);
  nor _67728_ (_16627_, _08270_, _09258_);
  or _67729_ (_16628_, _16627_, _16600_);
  or _67730_ (_16629_, _16628_, _06848_);
  and _67731_ (_16630_, _16629_, _16626_);
  or _67732_ (_16631_, _16630_, _06219_);
  or _67733_ (_16632_, _16615_, _06220_);
  and _67734_ (_16633_, _16632_, _06040_);
  and _67735_ (_16634_, _16633_, _16631_);
  or _67736_ (_16635_, _16634_, _16610_);
  and _67737_ (_16636_, _16635_, _06033_);
  or _67738_ (_16637_, _16607_, _14914_);
  and _67739_ (_16638_, _16623_, _06032_);
  and _67740_ (_16639_, _16638_, _16637_);
  or _67741_ (_16640_, _16639_, _09269_);
  or _67742_ (_16641_, _16640_, _16636_);
  or _67743_ (_16642_, _09777_, _09775_);
  and _67744_ (_16643_, _16642_, _09778_);
  or _67745_ (_16644_, _16643_, _09800_);
  and _67746_ (_16645_, _16644_, _06027_);
  and _67747_ (_16646_, _16645_, _16641_);
  or _67748_ (_16647_, _16607_, _14879_);
  and _67749_ (_16648_, _16647_, _06026_);
  and _67750_ (_16649_, _16648_, _16623_);
  or _67751_ (_16650_, _16649_, _09818_);
  or _67752_ (_16651_, _16650_, _16646_);
  and _67753_ (_16652_, _09180_, _07698_);
  or _67754_ (_16653_, _16600_, _07012_);
  or _67755_ (_16654_, _16653_, _16652_);
  or _67756_ (_16655_, _16628_, _09827_);
  and _67757_ (_16656_, _16655_, _05669_);
  and _67758_ (_16657_, _16656_, _16654_);
  and _67759_ (_16658_, _16657_, _16651_);
  or _67760_ (_16659_, _16658_, _16606_);
  and _67761_ (_16660_, _16659_, _09839_);
  nand _67762_ (_16661_, _10184_, _10147_);
  nor _67763_ (_16662_, _16545_, _10114_);
  or _67764_ (_16663_, _16662_, _10113_);
  nand _67765_ (_16664_, _16663_, _10150_);
  or _67766_ (_16665_, _16663_, _10150_);
  and _67767_ (_16666_, _16665_, _16664_);
  or _67768_ (_16667_, _16666_, _10184_);
  and _67769_ (_16668_, _16667_, _09832_);
  and _67770_ (_16669_, _16668_, _16661_);
  or _67771_ (_16670_, _16669_, _06019_);
  or _67772_ (_16671_, _16670_, _16660_);
  and _67773_ (_16672_, _16671_, _16603_);
  or _67774_ (_16673_, _16672_, _06112_);
  and _67775_ (_16674_, _14876_, _07698_);
  or _67776_ (_16675_, _16600_, _08751_);
  or _67777_ (_16676_, _16675_, _16674_);
  and _67778_ (_16677_, _16676_, _08756_);
  and _67779_ (_16678_, _16677_, _16673_);
  and _67780_ (_16679_, _10986_, _07698_);
  or _67781_ (_16680_, _16679_, _16600_);
  and _67782_ (_16681_, _16680_, _06284_);
  or _67783_ (_16682_, _16681_, _16678_);
  and _67784_ (_16683_, _16682_, _07032_);
  or _67785_ (_16684_, _16600_, _08273_);
  and _67786_ (_16685_, _16602_, _06108_);
  and _67787_ (_16686_, _16685_, _16684_);
  or _67788_ (_16687_, _16686_, _16683_);
  and _67789_ (_16688_, _16687_, _06278_);
  and _67790_ (_16689_, _16615_, _06277_);
  and _67791_ (_16690_, _16689_, _16684_);
  or _67792_ (_16691_, _16690_, _06130_);
  or _67793_ (_16692_, _16691_, _16688_);
  and _67794_ (_16693_, _14873_, _07698_);
  or _67795_ (_16694_, _16600_, _08777_);
  or _67796_ (_16695_, _16694_, _16693_);
  and _67797_ (_16696_, _16695_, _08782_);
  and _67798_ (_16697_, _16696_, _16692_);
  nor _67799_ (_16698_, _10985_, _09258_);
  or _67800_ (_16699_, _16698_, _16600_);
  and _67801_ (_16700_, _16699_, _06292_);
  or _67802_ (_16701_, _16700_, _06316_);
  or _67803_ (_16702_, _16701_, _16697_);
  or _67804_ (_16703_, _16612_, _06718_);
  and _67805_ (_16704_, _16703_, _05653_);
  and _67806_ (_16705_, _16704_, _16702_);
  and _67807_ (_16706_, _16609_, _05652_);
  or _67808_ (_16707_, _16706_, _06047_);
  or _67809_ (_16708_, _16707_, _16705_);
  and _67810_ (_16709_, _15055_, _07698_);
  or _67811_ (_16710_, _16600_, _06048_);
  or _67812_ (_16711_, _16710_, _16709_);
  and _67813_ (_16712_, _16711_, _01336_);
  and _67814_ (_16713_, _16712_, _16708_);
  or _67815_ (_16714_, _16713_, _16599_);
  and _67816_ (_43328_, _16714_, _42882_);
  nor _67817_ (_16715_, _01336_, _09855_);
  nor _67818_ (_16716_, _07698_, _09855_);
  and _67819_ (_16717_, _15179_, _07698_);
  or _67820_ (_16718_, _16717_, _16716_);
  and _67821_ (_16719_, _16718_, _09833_);
  nor _67822_ (_16720_, _08361_, _09855_);
  and _67823_ (_16721_, _15077_, _08361_);
  or _67824_ (_16722_, _16721_, _16720_);
  and _67825_ (_16723_, _16722_, _06039_);
  and _67826_ (_16724_, _15093_, _07698_);
  or _67827_ (_16725_, _16724_, _16716_);
  or _67828_ (_16726_, _16725_, _06954_);
  and _67829_ (_16727_, _07698_, \oc8051_golden_model_1.ACC [5]);
  or _67830_ (_16728_, _16727_, _16716_);
  and _67831_ (_16729_, _16728_, _06938_);
  nor _67832_ (_16730_, _06938_, _09855_);
  or _67833_ (_16731_, _16730_, _06102_);
  or _67834_ (_16732_, _16731_, _16729_);
  and _67835_ (_16733_, _16732_, _06044_);
  and _67836_ (_16734_, _16733_, _16726_);
  and _67837_ (_16735_, _15073_, _08361_);
  or _67838_ (_16736_, _16735_, _16720_);
  and _67839_ (_16737_, _16736_, _06043_);
  or _67840_ (_16738_, _16737_, _06239_);
  or _67841_ (_16739_, _16738_, _16734_);
  nor _67842_ (_16740_, _07977_, _09258_);
  or _67843_ (_16741_, _16740_, _16716_);
  or _67844_ (_16742_, _16741_, _06848_);
  and _67845_ (_16743_, _16742_, _16739_);
  or _67846_ (_16744_, _16743_, _06219_);
  or _67847_ (_16745_, _16728_, _06220_);
  and _67848_ (_16746_, _16745_, _06040_);
  and _67849_ (_16747_, _16746_, _16744_);
  or _67850_ (_16748_, _16747_, _16723_);
  and _67851_ (_16749_, _16748_, _06033_);
  or _67852_ (_16750_, _16720_, _15110_);
  and _67853_ (_16751_, _16736_, _06032_);
  and _67854_ (_16752_, _16751_, _16750_);
  or _67855_ (_16753_, _16752_, _09269_);
  or _67856_ (_16754_, _16753_, _16749_);
  or _67857_ (_16755_, _09465_, _09466_);
  and _67858_ (_16756_, _16755_, _09779_);
  nor _67859_ (_16757_, _16756_, _09780_);
  or _67860_ (_16758_, _16757_, _09800_);
  and _67861_ (_16759_, _16758_, _06027_);
  and _67862_ (_16760_, _16759_, _16754_);
  or _67863_ (_16761_, _16720_, _15074_);
  and _67864_ (_16762_, _16761_, _06026_);
  and _67865_ (_16763_, _16762_, _16736_);
  or _67866_ (_16764_, _16763_, _09818_);
  or _67867_ (_16765_, _16764_, _16760_);
  and _67868_ (_16766_, _09179_, _07698_);
  or _67869_ (_16767_, _16716_, _07012_);
  or _67870_ (_16768_, _16767_, _16766_);
  or _67871_ (_16769_, _16741_, _09827_);
  and _67872_ (_16770_, _16769_, _05669_);
  and _67873_ (_16771_, _16770_, _16768_);
  and _67874_ (_16772_, _16771_, _16765_);
  or _67875_ (_16773_, _16772_, _16719_);
  and _67876_ (_16774_, _16773_, _09839_);
  and _67877_ (_16775_, _10184_, _09832_);
  and _67878_ (_16776_, _16775_, _10157_);
  not _67879_ (_16777_, _10149_);
  and _67880_ (_16778_, _16664_, _16777_);
  nor _67881_ (_16779_, _16778_, _10160_);
  and _67882_ (_16780_, _16778_, _10160_);
  or _67883_ (_16781_, _16780_, _16779_);
  nor _67884_ (_16782_, _10184_, _09839_);
  and _67885_ (_16783_, _16782_, _16781_);
  or _67886_ (_16784_, _16783_, _16776_);
  or _67887_ (_16785_, _16784_, _16774_);
  and _67888_ (_16786_, _16785_, _06020_);
  and _67889_ (_16787_, _08652_, _07698_);
  or _67890_ (_16788_, _16787_, _16716_);
  and _67891_ (_16789_, _16788_, _06019_);
  or _67892_ (_16790_, _16789_, _06112_);
  or _67893_ (_16791_, _16790_, _16786_);
  and _67894_ (_16792_, _15195_, _07698_);
  or _67895_ (_16793_, _16716_, _08751_);
  or _67896_ (_16794_, _16793_, _16792_);
  and _67897_ (_16795_, _16794_, _08756_);
  and _67898_ (_16796_, _16795_, _16791_);
  and _67899_ (_16797_, _12306_, _07698_);
  or _67900_ (_16798_, _16797_, _16716_);
  and _67901_ (_16799_, _16798_, _06284_);
  or _67902_ (_16800_, _16799_, _16796_);
  and _67903_ (_16801_, _16800_, _07032_);
  or _67904_ (_16802_, _16716_, _07980_);
  and _67905_ (_16803_, _16788_, _06108_);
  and _67906_ (_16804_, _16803_, _16802_);
  or _67907_ (_16805_, _16804_, _16801_);
  and _67908_ (_16806_, _16805_, _06278_);
  and _67909_ (_16807_, _16728_, _06277_);
  and _67910_ (_16808_, _16807_, _16802_);
  or _67911_ (_16809_, _16808_, _06130_);
  or _67912_ (_16810_, _16809_, _16806_);
  and _67913_ (_16811_, _15194_, _07698_);
  or _67914_ (_16812_, _16716_, _08777_);
  or _67915_ (_16813_, _16812_, _16811_);
  and _67916_ (_16814_, _16813_, _08782_);
  and _67917_ (_16815_, _16814_, _16810_);
  nor _67918_ (_16816_, _10982_, _09258_);
  or _67919_ (_16817_, _16816_, _16716_);
  and _67920_ (_16818_, _16817_, _06292_);
  or _67921_ (_16819_, _16818_, _06316_);
  or _67922_ (_16820_, _16819_, _16815_);
  or _67923_ (_16821_, _16725_, _06718_);
  and _67924_ (_16822_, _16821_, _05653_);
  and _67925_ (_16823_, _16822_, _16820_);
  and _67926_ (_16824_, _16722_, _05652_);
  or _67927_ (_16825_, _16824_, _06047_);
  or _67928_ (_16826_, _16825_, _16823_);
  and _67929_ (_16827_, _15253_, _07698_);
  or _67930_ (_16828_, _16716_, _06048_);
  or _67931_ (_16829_, _16828_, _16827_);
  and _67932_ (_16830_, _16829_, _01336_);
  and _67933_ (_16831_, _16830_, _16826_);
  or _67934_ (_16832_, _16831_, _16715_);
  and _67935_ (_43329_, _16832_, _42882_);
  nor _67936_ (_16833_, _01336_, _10089_);
  nor _67937_ (_16834_, _07698_, _10089_);
  and _67938_ (_16835_, _15389_, _07698_);
  or _67939_ (_16836_, _16835_, _16834_);
  or _67940_ (_16837_, _16836_, _06020_);
  and _67941_ (_16838_, _15382_, _07698_);
  or _67942_ (_16839_, _16838_, _16834_);
  and _67943_ (_16840_, _16839_, _09833_);
  nor _67944_ (_16841_, _08361_, _10089_);
  and _67945_ (_16842_, _15278_, _08361_);
  or _67946_ (_16843_, _16842_, _16841_);
  and _67947_ (_16844_, _16843_, _06039_);
  and _67948_ (_16845_, _15293_, _07698_);
  or _67949_ (_16846_, _16845_, _16834_);
  or _67950_ (_16847_, _16846_, _06954_);
  and _67951_ (_16848_, _07698_, \oc8051_golden_model_1.ACC [6]);
  or _67952_ (_16849_, _16848_, _16834_);
  and _67953_ (_16850_, _16849_, _06938_);
  nor _67954_ (_16851_, _06938_, _10089_);
  or _67955_ (_16852_, _16851_, _06102_);
  or _67956_ (_16853_, _16852_, _16850_);
  and _67957_ (_16854_, _16853_, _06044_);
  and _67958_ (_16855_, _16854_, _16847_);
  and _67959_ (_16856_, _15280_, _08361_);
  or _67960_ (_16857_, _16856_, _16841_);
  and _67961_ (_16858_, _16857_, _06043_);
  or _67962_ (_16859_, _16858_, _06239_);
  or _67963_ (_16860_, _16859_, _16855_);
  nor _67964_ (_16861_, _07883_, _09258_);
  or _67965_ (_16862_, _16861_, _16834_);
  or _67966_ (_16863_, _16862_, _06848_);
  and _67967_ (_16864_, _16863_, _16860_);
  or _67968_ (_16865_, _16864_, _06219_);
  or _67969_ (_16866_, _16849_, _06220_);
  and _67970_ (_16867_, _16866_, _06040_);
  and _67971_ (_16868_, _16867_, _16865_);
  or _67972_ (_16869_, _16868_, _16844_);
  and _67973_ (_16870_, _16869_, _06033_);
  or _67974_ (_16871_, _16841_, _15310_);
  and _67975_ (_16872_, _16857_, _06032_);
  and _67976_ (_16873_, _16872_, _16871_);
  or _67977_ (_16874_, _16873_, _09269_);
  or _67978_ (_16875_, _16874_, _16870_);
  not _67979_ (_16876_, _09799_);
  or _67980_ (_16877_, _09797_, _09781_);
  and _67981_ (_16878_, _16877_, _16876_);
  or _67982_ (_16879_, _16878_, _09800_);
  and _67983_ (_16880_, _16879_, _06027_);
  and _67984_ (_16881_, _16880_, _16875_);
  or _67985_ (_16882_, _16841_, _15326_);
  and _67986_ (_16883_, _16882_, _06026_);
  and _67987_ (_16884_, _16883_, _16857_);
  or _67988_ (_16885_, _16884_, _09818_);
  or _67989_ (_16886_, _16885_, _16881_);
  and _67990_ (_16887_, _09178_, _07698_);
  or _67991_ (_16888_, _16834_, _07012_);
  or _67992_ (_16889_, _16888_, _16887_);
  or _67993_ (_16890_, _16862_, _09827_);
  and _67994_ (_16891_, _16890_, _05669_);
  and _67995_ (_16892_, _16891_, _16889_);
  and _67996_ (_16893_, _16892_, _16886_);
  or _67997_ (_16894_, _16893_, _16840_);
  and _67998_ (_16895_, _16894_, _09839_);
  nor _67999_ (_16896_, _16778_, _10158_);
  or _68000_ (_16897_, _16896_, _10159_);
  nor _68001_ (_16898_, _16897_, _10164_);
  and _68002_ (_16899_, _16897_, _10164_);
  or _68003_ (_16900_, _16899_, _16898_);
  or _68004_ (_16901_, _16900_, _10184_);
  nor _68005_ (_16902_, _10102_, _09839_);
  or _68006_ (_16903_, _16902_, _16782_);
  and _68007_ (_16904_, _16903_, _16901_);
  or _68008_ (_16905_, _16904_, _06019_);
  or _68009_ (_16906_, _16905_, _16895_);
  and _68010_ (_16907_, _16906_, _16837_);
  or _68011_ (_16908_, _16907_, _06112_);
  and _68012_ (_16909_, _15399_, _07698_);
  or _68013_ (_16910_, _16909_, _16834_);
  or _68014_ (_16911_, _16910_, _08751_);
  and _68015_ (_16912_, _16911_, _08756_);
  and _68016_ (_16913_, _16912_, _16908_);
  and _68017_ (_16914_, _10980_, _07698_);
  or _68018_ (_16915_, _16914_, _16834_);
  and _68019_ (_16916_, _16915_, _06284_);
  or _68020_ (_16917_, _16916_, _16913_);
  and _68021_ (_16918_, _16917_, _07032_);
  or _68022_ (_16919_, _16834_, _07886_);
  and _68023_ (_16920_, _16836_, _06108_);
  and _68024_ (_16921_, _16920_, _16919_);
  or _68025_ (_16922_, _16921_, _16918_);
  and _68026_ (_16923_, _16922_, _06278_);
  and _68027_ (_16924_, _16849_, _06277_);
  and _68028_ (_16925_, _16924_, _16919_);
  or _68029_ (_16926_, _16925_, _06130_);
  or _68030_ (_16927_, _16926_, _16923_);
  and _68031_ (_16928_, _15396_, _07698_);
  or _68032_ (_16929_, _16834_, _08777_);
  or _68033_ (_16930_, _16929_, _16928_);
  and _68034_ (_16931_, _16930_, _08782_);
  and _68035_ (_16932_, _16931_, _16927_);
  nor _68036_ (_16933_, _10979_, _09258_);
  or _68037_ (_16934_, _16933_, _16834_);
  and _68038_ (_16935_, _16934_, _06292_);
  or _68039_ (_16936_, _16935_, _06316_);
  or _68040_ (_16937_, _16936_, _16932_);
  or _68041_ (_16938_, _16846_, _06718_);
  and _68042_ (_16939_, _16938_, _05653_);
  and _68043_ (_16940_, _16939_, _16937_);
  and _68044_ (_16941_, _16843_, _05652_);
  or _68045_ (_16942_, _16941_, _06047_);
  or _68046_ (_16943_, _16942_, _16940_);
  and _68047_ (_16944_, _15451_, _07698_);
  or _68048_ (_16945_, _16834_, _06048_);
  or _68049_ (_16946_, _16945_, _16944_);
  and _68050_ (_16947_, _16946_, _01336_);
  and _68051_ (_16948_, _16947_, _16943_);
  or _68052_ (_16949_, _16948_, _16833_);
  and _68053_ (_43330_, _16949_, _42882_);
  nor _68054_ (_16950_, _01336_, _05758_);
  nand _68055_ (_16951_, _11015_, _08393_);
  nand _68056_ (_16952_, _12303_, _06051_);
  and _68057_ (_16953_, _16952_, _11050_);
  nor _68058_ (_16954_, _06931_, \oc8051_golden_model_1.ACC [0]);
  nor _68059_ (_16955_, _10913_, _16954_);
  not _68060_ (_16956_, _10890_);
  and _68061_ (_16957_, _16956_, _16955_);
  nor _68062_ (_16958_, _10285_, _05758_);
  or _68063_ (_16959_, _16958_, _10477_);
  or _68064_ (_16960_, _10794_, _16959_);
  and _68065_ (_16961_, _16960_, _12525_);
  nand _68066_ (_16962_, _10781_, _12321_);
  and _68067_ (_16963_, _14086_, _07701_);
  nor _68068_ (_16964_, _07701_, _05758_);
  or _68069_ (_16965_, _16964_, _08751_);
  or _68070_ (_16966_, _16965_, _16963_);
  nor _68071_ (_16967_, _09120_, \oc8051_golden_model_1.ACC [0]);
  nor _68072_ (_16968_, _10955_, _16967_);
  or _68073_ (_16969_, _10686_, _16968_);
  not _68074_ (_16970_, _06650_);
  and _68075_ (_16971_, _06133_, _05726_);
  not _68076_ (_16972_, _16971_);
  and _68077_ (_16973_, _10677_, _16955_);
  nor _68078_ (_16974_, _12322_, _10606_);
  and _68079_ (_16975_, _12322_, _10606_);
  or _68080_ (_16976_, _16975_, _16974_);
  or _68081_ (_16977_, _16976_, _10307_);
  not _68082_ (_16978_, _10378_);
  or _68083_ (_16979_, _16978_, _06931_);
  or _68084_ (_16980_, _10400_, _06931_);
  nor _68085_ (_16981_, _06530_, _05758_);
  and _68086_ (_16982_, _06530_, _05758_);
  nor _68087_ (_16983_, _16982_, _16981_);
  nand _68088_ (_16984_, _16983_, _10400_);
  and _68089_ (_16985_, _16984_, _10390_);
  and _68090_ (_16986_, _16985_, _16980_);
  and _68091_ (_16987_, _16986_, _06949_);
  or _68092_ (_16988_, _16987_, _09120_);
  or _68093_ (_16989_, _16986_, _10389_);
  and _68094_ (_16990_, _16989_, _05698_);
  or _68095_ (_16991_, _16990_, _06948_);
  and _68096_ (_16992_, _16991_, _06954_);
  and _68097_ (_16993_, _16992_, _16988_);
  nor _68098_ (_16994_, _08127_, _10439_);
  or _68099_ (_16995_, _16994_, _16964_);
  and _68100_ (_16996_, _16995_, _06102_);
  or _68101_ (_16997_, _16996_, _06043_);
  or _68102_ (_16998_, _16997_, _16993_);
  and _68103_ (_16999_, _14102_, _08359_);
  nor _68104_ (_17000_, _08359_, _05758_);
  or _68105_ (_17001_, _17000_, _06044_);
  or _68106_ (_17002_, _17001_, _16999_);
  and _68107_ (_17003_, _17002_, _06848_);
  and _68108_ (_17004_, _17003_, _16998_);
  and _68109_ (_17005_, _07701_, _06931_);
  or _68110_ (_17006_, _17005_, _16964_);
  and _68111_ (_17007_, _17006_, _06239_);
  or _68112_ (_17008_, _17007_, _10378_);
  or _68113_ (_17009_, _17008_, _17004_);
  and _68114_ (_17010_, _17009_, _16979_);
  or _68115_ (_17011_, _17010_, _06970_);
  or _68116_ (_17012_, _09120_, _06971_);
  and _68117_ (_17013_, _17012_, _06220_);
  and _68118_ (_17014_, _17013_, _17011_);
  and _68119_ (_17015_, _08127_, _06219_);
  or _68120_ (_17016_, _17015_, _10376_);
  or _68121_ (_17017_, _17016_, _17014_);
  nand _68122_ (_17018_, _10376_, _09880_);
  and _68123_ (_17019_, _17018_, _17017_);
  or _68124_ (_17020_, _17019_, _06039_);
  or _68125_ (_17021_, _16964_, _06040_);
  and _68126_ (_17022_, _17021_, _06033_);
  and _68127_ (_17023_, _17022_, _17020_);
  and _68128_ (_17024_, _16995_, _06032_);
  or _68129_ (_17025_, _17024_, _09269_);
  or _68130_ (_17026_, _17025_, _17023_);
  nand _68131_ (_17027_, \oc8051_golden_model_1.B [0], \oc8051_golden_model_1.ACC [0]);
  nand _68132_ (_17028_, _17027_, _09269_);
  and _68133_ (_17029_, _17028_, _10469_);
  and _68134_ (_17030_, _17029_, _17026_);
  and _68135_ (_17031_, _16959_, _10468_);
  or _68136_ (_17032_, _17031_, _12361_);
  or _68137_ (_17033_, _17032_, _17030_);
  nor _68138_ (_17034_, _10542_, _05758_);
  or _68139_ (_17035_, _17034_, _10543_);
  or _68140_ (_17036_, _17035_, _13935_);
  and _68141_ (_17037_, _17036_, _06267_);
  and _68142_ (_17038_, _17037_, _17033_);
  nor _68143_ (_17039_, _10353_, _05758_);
  or _68144_ (_17040_, _17039_, _10354_);
  or _68145_ (_17041_, _17040_, _10306_);
  and _68146_ (_17042_, _17041_, _12367_);
  or _68147_ (_17043_, _17042_, _17038_);
  and _68148_ (_17044_, _17043_, _16977_);
  or _68149_ (_17045_, _17044_, _05676_);
  nand _68150_ (_17046_, _06016_, _05676_);
  and _68151_ (_17047_, _17046_, _06027_);
  and _68152_ (_17048_, _17047_, _17045_);
  and _68153_ (_17049_, _14132_, _08359_);
  or _68154_ (_17050_, _17049_, _17000_);
  and _68155_ (_17051_, _17050_, _06026_);
  or _68156_ (_17052_, _17051_, _09818_);
  or _68157_ (_17053_, _17052_, _17048_);
  and _68158_ (_17054_, _09120_, _07701_);
  or _68159_ (_17055_, _16964_, _07012_);
  or _68160_ (_17056_, _17055_, _17054_);
  or _68161_ (_17057_, _17006_, _09827_);
  and _68162_ (_17058_, _17057_, _05669_);
  and _68163_ (_17059_, _17058_, _17056_);
  and _68164_ (_17060_, _17059_, _17053_);
  and _68165_ (_17061_, _14186_, _07701_);
  or _68166_ (_17062_, _17061_, _16964_);
  and _68167_ (_17063_, _17062_, _09833_);
  or _68168_ (_17064_, _17063_, _09832_);
  or _68169_ (_17065_, _17064_, _17060_);
  nor _68170_ (_17066_, _16775_, _05663_);
  and _68171_ (_17067_, _17066_, _17065_);
  nor _68172_ (_17068_, _06016_, _05664_);
  or _68173_ (_17069_, _17068_, _06019_);
  or _68174_ (_17070_, _17069_, _17067_);
  and _68175_ (_17071_, _07701_, _08672_);
  or _68176_ (_17072_, _17071_, _16964_);
  or _68177_ (_17073_, _17072_, _06020_);
  and _68178_ (_17074_, _17073_, _10662_);
  and _68179_ (_17075_, _17074_, _17070_);
  nor _68180_ (_17076_, _10662_, _06016_);
  or _68181_ (_17077_, _17076_, _10669_);
  or _68182_ (_17078_, _17077_, _17075_);
  or _68183_ (_17079_, _10675_, _16955_);
  and _68184_ (_17080_, _17079_, _10678_);
  and _68185_ (_17081_, _17080_, _17078_);
  or _68186_ (_17082_, _17081_, _16973_);
  and _68187_ (_17083_, _17082_, _16972_);
  and _68188_ (_17084_, _16971_, _16955_);
  or _68189_ (_17085_, _17084_, _17083_);
  and _68190_ (_17086_, _17085_, _16970_);
  and _68191_ (_17087_, _16955_, _06650_);
  or _68192_ (_17088_, _17087_, _10685_);
  or _68193_ (_17089_, _17088_, _17086_);
  and _68194_ (_17090_, _17089_, _16969_);
  or _68195_ (_17091_, _17090_, _06282_);
  nand _68196_ (_17092_, _12303_, _06282_);
  and _68197_ (_17093_, _17092_, _10699_);
  and _68198_ (_17094_, _17093_, _17091_);
  and _68199_ (_17095_, _10698_, _12322_);
  or _68200_ (_17096_, _17095_, _06112_);
  or _68201_ (_17097_, _17096_, _17094_);
  and _68202_ (_17098_, _17097_, _16966_);
  or _68203_ (_17099_, _17098_, _06284_);
  or _68204_ (_17100_, _16964_, _08756_);
  nand _68205_ (_17101_, _05735_, _05567_);
  and _68206_ (_17102_, _17101_, _17100_);
  and _68207_ (_17103_, _17102_, _17099_);
  not _68208_ (_17104_, _17101_);
  and _68209_ (_17105_, _17104_, _10913_);
  or _68210_ (_17106_, _17105_, _10731_);
  or _68211_ (_17107_, _17106_, _17103_);
  or _68212_ (_17108_, _10736_, _10955_);
  and _68213_ (_17109_, _17108_, _10735_);
  and _68214_ (_17110_, _17109_, _17107_);
  or _68215_ (_17111_, _10741_, _10995_);
  and _68216_ (_17112_, _17111_, _10743_);
  or _68217_ (_17113_, _17112_, _17110_);
  or _68218_ (_17114_, _10747_, _11036_);
  and _68219_ (_17115_, _17114_, _07032_);
  and _68220_ (_17116_, _17115_, _17113_);
  nand _68221_ (_17117_, _17072_, _06108_);
  nor _68222_ (_17118_, _17117_, _16994_);
  or _68223_ (_17119_, _17118_, _10752_);
  or _68224_ (_17120_, _17119_, _17116_);
  nand _68225_ (_17121_, _16954_, _10752_);
  and _68226_ (_17122_, _17121_, _10760_);
  and _68227_ (_17123_, _17122_, _17120_);
  nor _68228_ (_17124_, _10760_, _16954_);
  or _68229_ (_17125_, _17124_, _10767_);
  or _68230_ (_17126_, _17125_, _17123_);
  nand _68231_ (_17127_, _10767_, _16954_);
  and _68232_ (_17128_, _17127_, _06668_);
  and _68233_ (_17129_, _17128_, _17126_);
  nor _68234_ (_17130_, _16954_, _06668_);
  or _68235_ (_17131_, _17130_, _10775_);
  or _68236_ (_17132_, _17131_, _17129_);
  nand _68237_ (_17133_, _10775_, _16967_);
  and _68238_ (_17134_, _17133_, _06291_);
  and _68239_ (_17135_, _17134_, _17132_);
  not _68240_ (_17136_, _10781_);
  nand _68241_ (_17137_, _17136_, _12302_);
  and _68242_ (_17138_, _17137_, _11987_);
  or _68243_ (_17139_, _17138_, _17135_);
  and _68244_ (_17140_, _17139_, _16962_);
  or _68245_ (_17141_, _17140_, _06130_);
  and _68246_ (_17142_, _14083_, _07701_);
  or _68247_ (_17143_, _16964_, _08777_);
  or _68248_ (_17144_, _17143_, _17142_);
  and _68249_ (_17145_, _17144_, _10304_);
  and _68250_ (_17146_, _17145_, _17141_);
  or _68251_ (_17147_, _17146_, _16961_);
  or _68252_ (_17148_, _10796_, _17035_);
  and _68253_ (_17149_, _17148_, _17147_);
  or _68254_ (_17150_, _17149_, _06288_);
  or _68255_ (_17151_, _17040_, _06289_);
  and _68256_ (_17152_, _17151_, _10856_);
  and _68257_ (_17153_, _17152_, _17150_);
  and _68258_ (_17154_, _10824_, _16976_);
  or _68259_ (_17155_, _17154_, _10854_);
  or _68260_ (_17156_, _17155_, _17153_);
  nand _68261_ (_17157_, _10854_, _10606_);
  and _68262_ (_17158_, _17157_, _10890_);
  and _68263_ (_17159_, _17158_, _17156_);
  or _68264_ (_17160_, _17159_, _16957_);
  and _68265_ (_17161_, _17160_, _10934_);
  and _68266_ (_17162_, _10932_, _16968_);
  or _68267_ (_17163_, _17162_, _06051_);
  or _68268_ (_17164_, _17163_, _17161_);
  and _68269_ (_17165_, _17164_, _16953_);
  and _68270_ (_17166_, _10974_, _12322_);
  or _68271_ (_17167_, _17166_, _11015_);
  or _68272_ (_17168_, _17167_, _17165_);
  and _68273_ (_17169_, _17168_, _16951_);
  or _68274_ (_17170_, _17169_, _06316_);
  or _68275_ (_17171_, _16995_, _06718_);
  and _68276_ (_17172_, _17171_, _11060_);
  and _68277_ (_17173_, _17172_, _17170_);
  nor _68278_ (_17174_, _11064_, _05758_);
  nor _68279_ (_17175_, _17174_, _12756_);
  or _68280_ (_17176_, _17175_, _17173_);
  nand _68281_ (_17177_, _11064_, _05784_);
  and _68282_ (_17178_, _17177_, _05653_);
  and _68283_ (_17179_, _17178_, _17176_);
  and _68284_ (_17180_, _16964_, _05652_);
  or _68285_ (_17181_, _17180_, _06047_);
  or _68286_ (_17182_, _17181_, _17179_);
  or _68287_ (_17183_, _16995_, _06048_);
  and _68288_ (_17184_, _17183_, _11083_);
  and _68289_ (_17185_, _17184_, _17182_);
  nor _68290_ (_17186_, _11089_, _05758_);
  nor _68291_ (_17187_, _17186_, _12779_);
  or _68292_ (_17188_, _17187_, _17185_);
  nand _68293_ (_17189_, _11089_, _05784_);
  and _68294_ (_17190_, _17189_, _01336_);
  and _68295_ (_17191_, _17190_, _17188_);
  or _68296_ (_17192_, _17191_, _16950_);
  and _68297_ (_43332_, _17192_, _42882_);
  nor _68298_ (_17193_, _01336_, _05784_);
  nor _68299_ (_17194_, _10835_, _10834_);
  nor _68300_ (_17195_, _17194_, _10836_);
  or _68301_ (_17196_, _17195_, _06289_);
  and _68302_ (_17197_, _17196_, _10856_);
  and _68303_ (_17198_, _07701_, _06832_);
  and _68304_ (_17199_, _17198_, _08077_);
  nor _68305_ (_17200_, _07701_, \oc8051_golden_model_1.ACC [1]);
  or _68306_ (_17201_, _17200_, _08777_);
  or _68307_ (_17202_, _17201_, _17199_);
  and _68308_ (_17203_, _06460_, _05739_);
  nor _68309_ (_17204_, _06834_, _17203_);
  not _68310_ (_17205_, _10752_);
  or _68311_ (_17206_, _10736_, _10951_);
  nor _68312_ (_17207_, _10677_, _10669_);
  not _68313_ (_17208_, _17207_);
  and _68314_ (_17209_, _17208_, _10912_);
  or _68315_ (_17210_, _10092_, _09839_);
  not _68316_ (_17211_, _10954_);
  nor _68317_ (_17212_, _10536_, _05758_);
  or _68318_ (_17213_, _17212_, _10541_);
  nand _68319_ (_17214_, _17213_, _17211_);
  or _68320_ (_17215_, _17213_, _17211_);
  and _68321_ (_17216_, _17215_, _12361_);
  and _68322_ (_17217_, _17216_, _17214_);
  nand _68323_ (_17218_, _10378_, _07132_);
  nor _68324_ (_17219_, _10389_, _06948_);
  or _68325_ (_17220_, _17219_, _09075_);
  nor _68326_ (_17221_, _10400_, _07132_);
  nor _68327_ (_17222_, _06530_, _05784_);
  and _68328_ (_17223_, _06530_, _05784_);
  or _68329_ (_17224_, _17223_, _17222_);
  and _68330_ (_17225_, _17224_, _10400_);
  or _68331_ (_17226_, _17225_, _10389_);
  or _68332_ (_17227_, _17226_, _17221_);
  and _68333_ (_17228_, _17227_, _05698_);
  or _68334_ (_17229_, _17228_, _06948_);
  and _68335_ (_17230_, _17229_, _06954_);
  and _68336_ (_17231_, _17230_, _17220_);
  and _68337_ (_17232_, _14284_, _07701_);
  nor _68338_ (_17233_, _17232_, _17200_);
  and _68339_ (_17234_, _17233_, _06102_);
  or _68340_ (_17235_, _17234_, _10412_);
  or _68341_ (_17236_, _17235_, _17231_);
  nor _68342_ (_17237_, _10416_, \oc8051_golden_model_1.PSW [6]);
  nor _68343_ (_17238_, _17237_, \oc8051_golden_model_1.ACC [1]);
  and _68344_ (_17239_, _17237_, \oc8051_golden_model_1.ACC [1]);
  nor _68345_ (_17240_, _17239_, _17238_);
  nand _68346_ (_17241_, _17240_, _10412_);
  and _68347_ (_17242_, _17241_, _06244_);
  and _68348_ (_17243_, _17242_, _17236_);
  nor _68349_ (_17244_, _08359_, _05784_);
  and _68350_ (_17245_, _14266_, _08359_);
  nor _68351_ (_17246_, _17245_, _17244_);
  nor _68352_ (_17247_, _17246_, _06044_);
  nor _68353_ (_17248_, _07701_, _05784_);
  nor _68354_ (_17249_, _10439_, _07132_);
  or _68355_ (_17250_, _17249_, _17248_);
  and _68356_ (_17251_, _17250_, _06239_);
  or _68357_ (_17252_, _17251_, _10378_);
  or _68358_ (_17253_, _17252_, _17247_);
  or _68359_ (_17254_, _17253_, _17243_);
  and _68360_ (_17255_, _17254_, _17218_);
  or _68361_ (_17256_, _17255_, _06970_);
  or _68362_ (_17257_, _09075_, _06971_);
  and _68363_ (_17258_, _17257_, _06220_);
  and _68364_ (_17259_, _17258_, _17256_);
  nor _68365_ (_17260_, _08077_, _06220_);
  or _68366_ (_17261_, _17260_, _10376_);
  or _68367_ (_17262_, _17261_, _17259_);
  nand _68368_ (_17263_, _10376_, _09906_);
  and _68369_ (_17264_, _17263_, _17262_);
  or _68370_ (_17265_, _17264_, _06039_);
  and _68371_ (_17266_, _14273_, _08359_);
  or _68372_ (_17267_, _17266_, _17244_);
  or _68373_ (_17268_, _17267_, _06040_);
  and _68374_ (_17269_, _17268_, _06033_);
  nand _68375_ (_17270_, _17269_, _17265_);
  nor _68376_ (_17271_, _17244_, _14302_);
  or _68377_ (_17272_, _17246_, _06033_);
  or _68378_ (_17273_, _17272_, _17271_);
  and _68379_ (_17274_, _17273_, _17270_);
  nor _68380_ (_17275_, _17274_, _09269_);
  nor _68381_ (_17276_, _09744_, _09743_);
  nor _68382_ (_17277_, _17276_, _09745_);
  nand _68383_ (_17278_, _17277_, _09269_);
  nand _68384_ (_17279_, _17278_, _10469_);
  or _68385_ (_17280_, _17279_, _17275_);
  nor _68386_ (_17281_, _10234_, _05758_);
  or _68387_ (_17282_, _17281_, _10284_);
  nor _68388_ (_17283_, _17282_, _10912_);
  and _68389_ (_17284_, _17282_, _10912_);
  or _68390_ (_17285_, _17284_, _17283_);
  or _68391_ (_17286_, _17285_, _10469_);
  and _68392_ (_17287_, _17286_, _13935_);
  and _68393_ (_17288_, _17287_, _17280_);
  or _68394_ (_17289_, _17288_, _17217_);
  and _68395_ (_17290_, _17289_, _06267_);
  nor _68396_ (_17291_, _10308_, _05758_);
  or _68397_ (_17292_, _17291_, _10352_);
  and _68398_ (_17293_, _17292_, _10994_);
  nor _68399_ (_17294_, _17292_, _10994_);
  or _68400_ (_17295_, _17294_, _17293_);
  and _68401_ (_17296_, _17295_, _06261_);
  or _68402_ (_17297_, _17296_, _17290_);
  and _68403_ (_17298_, _17297_, _10307_);
  nor _68404_ (_17299_, _06016_, \oc8051_golden_model_1.ACC [0]);
  nor _68405_ (_17300_, _17299_, _11035_);
  and _68406_ (_17301_, _17299_, _11035_);
  or _68407_ (_17302_, _17301_, _17300_);
  nor _68408_ (_17303_, _16974_, _17302_);
  and _68409_ (_17304_, _12323_, \oc8051_golden_model_1.PSW [7]);
  or _68410_ (_17305_, _17304_, _17303_);
  and _68411_ (_17306_, _17305_, _10306_);
  or _68412_ (_17307_, _17306_, _05676_);
  or _68413_ (_17308_, _17307_, _17298_);
  nand _68414_ (_17309_, _06799_, _05676_);
  and _68415_ (_17310_, _17309_, _06027_);
  and _68416_ (_17311_, _17310_, _17308_);
  or _68417_ (_17312_, _17244_, _14267_);
  nand _68418_ (_17313_, _17312_, _06026_);
  nor _68419_ (_17314_, _17313_, _17246_);
  or _68420_ (_17315_, _17314_, _09818_);
  or _68421_ (_17316_, _17315_, _17311_);
  and _68422_ (_17317_, _09075_, _07701_);
  or _68423_ (_17318_, _17248_, _07012_);
  or _68424_ (_17319_, _17318_, _17317_);
  or _68425_ (_17320_, _17250_, _09827_);
  and _68426_ (_17321_, _17320_, _05669_);
  and _68427_ (_17322_, _17321_, _17319_);
  and _68428_ (_17323_, _17322_, _17316_);
  or _68429_ (_17324_, _14367_, _10439_);
  nor _68430_ (_17325_, _17200_, _05669_);
  and _68431_ (_17326_, _17325_, _17324_);
  or _68432_ (_17327_, _17326_, _09832_);
  or _68433_ (_17328_, _17327_, _17323_);
  and _68434_ (_17329_, _17328_, _17210_);
  or _68435_ (_17330_, _17329_, _05663_);
  nand _68436_ (_17331_, _06799_, _05663_);
  and _68437_ (_17332_, _17331_, _06020_);
  and _68438_ (_17333_, _17332_, _17330_);
  or _68439_ (_17334_, _17198_, _06020_);
  nor _68440_ (_17335_, _17334_, _17200_);
  or _68441_ (_17336_, _17335_, _10661_);
  or _68442_ (_17337_, _17336_, _17333_);
  nand _68443_ (_17338_, _10661_, _06799_);
  and _68444_ (_17339_, _17338_, _17207_);
  and _68445_ (_17340_, _17339_, _17337_);
  or _68446_ (_17341_, _17340_, _17209_);
  and _68447_ (_17342_, _17341_, _16972_);
  and _68448_ (_17343_, _16971_, _10912_);
  or _68449_ (_17344_, _17343_, _17342_);
  and _68450_ (_17345_, _17344_, _16970_);
  and _68451_ (_17346_, _10912_, _06650_);
  or _68452_ (_17347_, _17346_, _17345_);
  and _68453_ (_17348_, _17347_, _10686_);
  and _68454_ (_17349_, _10685_, _10954_);
  or _68455_ (_17350_, _17349_, _06282_);
  or _68456_ (_17351_, _17350_, _17348_);
  or _68457_ (_17352_, _10994_, _06283_);
  and _68458_ (_17353_, _17352_, _10699_);
  and _68459_ (_17354_, _17353_, _17351_);
  and _68460_ (_17355_, _10698_, _11035_);
  or _68461_ (_17356_, _17355_, _17354_);
  and _68462_ (_17357_, _17356_, _08751_);
  or _68463_ (_17358_, _14263_, _10439_);
  nor _68464_ (_17359_, _17200_, _08751_);
  and _68465_ (_17360_, _17359_, _17358_);
  or _68466_ (_17361_, _17360_, _06284_);
  or _68467_ (_17362_, _17361_, _17357_);
  or _68468_ (_17363_, _17248_, _08756_);
  and _68469_ (_17364_, _17363_, _17101_);
  and _68470_ (_17365_, _17364_, _17362_);
  and _68471_ (_17366_, _17104_, _10910_);
  or _68472_ (_17367_, _17366_, _10731_);
  or _68473_ (_17368_, _17367_, _17365_);
  and _68474_ (_17369_, _17368_, _17206_);
  or _68475_ (_17370_, _17369_, _06279_);
  or _68476_ (_17371_, _10992_, _10735_);
  and _68477_ (_17372_, _17371_, _10747_);
  and _68478_ (_17373_, _17372_, _17370_);
  and _68479_ (_17375_, _10741_, _11033_);
  or _68480_ (_17376_, _17375_, _17373_);
  and _68481_ (_17377_, _17376_, _07032_);
  or _68482_ (_17378_, _14261_, _10439_);
  nor _68483_ (_17379_, _17200_, _07032_);
  and _68484_ (_17380_, _17379_, _17378_);
  or _68485_ (_17381_, _17380_, _17377_);
  and _68486_ (_17382_, _17381_, _17205_);
  nor _68487_ (_17383_, _10911_, _17205_);
  nor _68488_ (_17384_, _17383_, _17382_);
  nand _68489_ (_17386_, _17384_, _17204_);
  not _68490_ (_17387_, _11991_);
  not _68491_ (_17388_, _17204_);
  nand _68492_ (_17389_, _17388_, _10911_);
  and _68493_ (_17390_, _17389_, _17387_);
  and _68494_ (_17391_, _17390_, _17386_);
  nor _68495_ (_17392_, _17387_, _10911_);
  or _68496_ (_17393_, _17392_, _10775_);
  or _68497_ (_17394_, _17393_, _17391_);
  not _68498_ (_17395_, _10775_);
  or _68499_ (_17397_, _17395_, _10952_);
  and _68500_ (_17398_, _17397_, _06291_);
  and _68501_ (_17399_, _17398_, _17394_);
  nor _68502_ (_17400_, _10993_, _06291_);
  or _68503_ (_17401_, _17400_, _10781_);
  or _68504_ (_17402_, _17401_, _17399_);
  nand _68505_ (_17403_, _10781_, _11034_);
  and _68506_ (_17404_, _17403_, _08777_);
  nand _68507_ (_17405_, _17404_, _17402_);
  and _68508_ (_17406_, _17405_, _17202_);
  or _68509_ (_17408_, _17406_, _10303_);
  and _68510_ (_17409_, _10794_, _06545_);
  not _68511_ (_17410_, _17409_);
  and _68512_ (_17411_, _10287_, _10283_);
  or _68513_ (_17412_, _10304_, _10288_);
  or _68514_ (_17413_, _17412_, _17411_);
  and _68515_ (_17414_, _17413_, _17410_);
  and _68516_ (_17415_, _17414_, _17408_);
  and _68517_ (_17416_, _06513_, _05731_);
  and _68518_ (_17417_, _10805_, _10803_);
  or _68519_ (_17419_, _17417_, _10806_);
  and _68520_ (_17420_, _17419_, _17409_);
  or _68521_ (_17421_, _17420_, _17416_);
  nor _68522_ (_17422_, _17421_, _17415_);
  not _68523_ (_17423_, _17416_);
  or _68524_ (_17424_, _17419_, _17423_);
  nand _68525_ (_17425_, _17424_, _06289_);
  or _68526_ (_17426_, _17425_, _17422_);
  and _68527_ (_17427_, _17426_, _17197_);
  or _68528_ (_17428_, _10865_, _10864_);
  nor _68529_ (_17430_, _10866_, _10856_);
  and _68530_ (_17431_, _17430_, _17428_);
  or _68531_ (_17432_, _17431_, _10854_);
  or _68532_ (_17433_, _17432_, _17427_);
  nand _68533_ (_17434_, _10854_, _05758_);
  and _68534_ (_17435_, _17434_, _10890_);
  and _68535_ (_17436_, _17435_, _17433_);
  and _68536_ (_17437_, _10394_, _05746_);
  or _68537_ (_17438_, _10913_, _10912_);
  nor _68538_ (_17439_, _10914_, _10890_);
  and _68539_ (_17440_, _17439_, _17438_);
  or _68540_ (_17441_, _17440_, _17437_);
  or _68541_ (_17442_, _17441_, _17436_);
  not _68542_ (_17443_, _06692_);
  nor _68543_ (_17444_, _10955_, _10954_);
  nor _68544_ (_17445_, _17444_, _10956_);
  and _68545_ (_17446_, _17445_, _17443_);
  or _68546_ (_17447_, _17446_, _10934_);
  and _68547_ (_17448_, _17447_, _17442_);
  and _68548_ (_17449_, _17445_, _06692_);
  or _68549_ (_17450_, _17449_, _10976_);
  or _68550_ (_17451_, _17450_, _17448_);
  nor _68551_ (_17452_, _10995_, _10994_);
  nor _68552_ (_17453_, _17452_, _10996_);
  or _68553_ (_17454_, _17453_, _06052_);
  nor _68554_ (_17455_, _11036_, _11035_);
  nor _68555_ (_17456_, _17455_, _11037_);
  or _68556_ (_17457_, _17456_, _11050_);
  and _68557_ (_17458_, _17457_, _11016_);
  and _68558_ (_17459_, _17458_, _17454_);
  and _68559_ (_17460_, _17459_, _17451_);
  and _68560_ (_17461_, _11015_, \oc8051_golden_model_1.ACC [0]);
  or _68561_ (_17462_, _17461_, _06316_);
  or _68562_ (_17463_, _17462_, _17460_);
  or _68563_ (_17464_, _17233_, _06718_);
  and _68564_ (_17465_, _17464_, _11060_);
  and _68565_ (_17466_, _17465_, _17463_);
  nor _68566_ (_17467_, \oc8051_golden_model_1.ACC [1], \oc8051_golden_model_1.ACC [0]);
  nor _68567_ (_17468_, _11090_, _17467_);
  nor _68568_ (_17469_, _17468_, _11060_);
  or _68569_ (_17470_, _17469_, _11064_);
  or _68570_ (_17471_, _17470_, _17466_);
  nand _68571_ (_17472_, _11064_, _09956_);
  and _68572_ (_17473_, _17472_, _05653_);
  and _68573_ (_17474_, _17473_, _17471_);
  and _68574_ (_17475_, _17267_, _05652_);
  or _68575_ (_17476_, _17475_, _06047_);
  or _68576_ (_17477_, _17476_, _17474_);
  or _68577_ (_17478_, _17232_, _17248_);
  or _68578_ (_17479_, _17478_, _06048_);
  and _68579_ (_17480_, _17479_, _11083_);
  and _68580_ (_17481_, _17480_, _17477_);
  and _68581_ (_17482_, _17468_, _11082_);
  or _68582_ (_17483_, _17482_, _11089_);
  or _68583_ (_17484_, _17483_, _17481_);
  nand _68584_ (_17485_, _11089_, _09956_);
  and _68585_ (_17486_, _17485_, _01336_);
  and _68586_ (_17487_, _17486_, _17484_);
  or _68587_ (_17488_, _17487_, _17193_);
  and _68588_ (_43333_, _17488_, _42882_);
  nor _68589_ (_17489_, _01336_, _09956_);
  nand _68590_ (_17490_, _11015_, _05784_);
  nor _68591_ (_17491_, _10998_, _10991_);
  nor _68592_ (_17492_, _17491_, _10999_);
  or _68593_ (_17493_, _17492_, _06052_);
  and _68594_ (_17494_, _17493_, _11050_);
  and _68595_ (_17495_, _10837_, _10346_);
  nor _68596_ (_17496_, _17495_, _10838_);
  or _68597_ (_17497_, _17496_, _06289_);
  and _68598_ (_17498_, _17497_, _10856_);
  and _68599_ (_17499_, _14596_, _07701_);
  nor _68600_ (_17500_, _07701_, _09956_);
  or _68601_ (_17501_, _17500_, _08751_);
  or _68602_ (_17502_, _17501_, _17499_);
  and _68603_ (_17503_, _06227_, _05726_);
  and _68604_ (_17504_, _10909_, _17503_);
  nand _68605_ (_17505_, _10378_, _07530_);
  or _68606_ (_17506_, _17219_, _09182_);
  nor _68607_ (_17507_, _10400_, _07530_);
  nor _68608_ (_17508_, _06530_, _09956_);
  and _68609_ (_17509_, _06530_, _09956_);
  or _68610_ (_17510_, _17509_, _17508_);
  and _68611_ (_17511_, _17510_, _10400_);
  or _68612_ (_17512_, _17511_, _10389_);
  or _68613_ (_17513_, _17512_, _17507_);
  and _68614_ (_17514_, _17513_, _05698_);
  or _68615_ (_17515_, _17514_, _06948_);
  and _68616_ (_17516_, _17515_, _06954_);
  and _68617_ (_17517_, _17516_, _17506_);
  and _68618_ (_17518_, _14493_, _07701_);
  or _68619_ (_17519_, _17518_, _17500_);
  and _68620_ (_17520_, _17519_, _06102_);
  or _68621_ (_17521_, _17520_, _10412_);
  or _68622_ (_17522_, _17521_, _17517_);
  nor _68623_ (_17523_, _17238_, _09956_);
  and _68624_ (_17524_, _10415_, \oc8051_golden_model_1.PSW [6]);
  nor _68625_ (_17525_, _17524_, _17523_);
  nand _68626_ (_17526_, _17525_, _10412_);
  and _68627_ (_17527_, _17526_, _06244_);
  and _68628_ (_17528_, _17527_, _17522_);
  nor _68629_ (_17529_, _08359_, _09956_);
  and _68630_ (_17530_, _14497_, _08359_);
  or _68631_ (_17531_, _17530_, _17529_);
  and _68632_ (_17532_, _17531_, _06043_);
  nor _68633_ (_17533_, _10439_, _07530_);
  or _68634_ (_17534_, _17533_, _17500_);
  and _68635_ (_17535_, _17534_, _06239_);
  or _68636_ (_17536_, _17535_, _10378_);
  or _68637_ (_17537_, _17536_, _17532_);
  or _68638_ (_17538_, _17537_, _17528_);
  and _68639_ (_17539_, _17538_, _17505_);
  or _68640_ (_17540_, _17539_, _06970_);
  or _68641_ (_17541_, _09182_, _06971_);
  and _68642_ (_17542_, _17541_, _06220_);
  and _68643_ (_17543_, _17542_, _17540_);
  nor _68644_ (_17544_, _08176_, _06220_);
  or _68645_ (_17545_, _17544_, _10376_);
  or _68646_ (_17546_, _17545_, _17543_);
  nand _68647_ (_17547_, _10376_, _09861_);
  and _68648_ (_17548_, _17547_, _17546_);
  or _68649_ (_17549_, _17548_, _06039_);
  and _68650_ (_17550_, _14479_, _08359_);
  or _68651_ (_17551_, _17550_, _17529_);
  or _68652_ (_17552_, _17551_, _06040_);
  and _68653_ (_17553_, _17552_, _06033_);
  and _68654_ (_17554_, _17553_, _17549_);
  or _68655_ (_17555_, _17529_, _14512_);
  and _68656_ (_17556_, _17531_, _06032_);
  and _68657_ (_17557_, _17556_, _17555_);
  or _68658_ (_17558_, _17557_, _09269_);
  or _68659_ (_17559_, _17558_, _17554_);
  nor _68660_ (_17560_, _09747_, _09745_);
  or _68661_ (_17561_, _17560_, _09748_);
  nand _68662_ (_17562_, _17561_, _09269_);
  and _68663_ (_17563_, _17562_, _10469_);
  and _68664_ (_17564_, _17563_, _17559_);
  and _68665_ (_17565_, _07132_, \oc8051_golden_model_1.ACC [1]);
  and _68666_ (_17566_, _06931_, _05758_);
  nor _68667_ (_17567_, _17566_, _10912_);
  nor _68668_ (_17568_, _17567_, _17565_);
  nor _68669_ (_17569_, _10909_, _17568_);
  and _68670_ (_17570_, _10909_, _17568_);
  nor _68671_ (_17571_, _17570_, _17569_);
  nor _68672_ (_17572_, _16955_, _10912_);
  and _68673_ (_17573_, _17572_, \oc8051_golden_model_1.PSW [7]);
  or _68674_ (_17574_, _17573_, _17571_);
  nand _68675_ (_17575_, _17573_, _17571_);
  and _68676_ (_17576_, _17575_, _10468_);
  and _68677_ (_17577_, _17576_, _17574_);
  or _68678_ (_17578_, _17577_, _12361_);
  or _68679_ (_17579_, _17578_, _17564_);
  and _68680_ (_17580_, _12150_, \oc8051_golden_model_1.ACC [1]);
  not _68681_ (_17581_, _17580_);
  and _68682_ (_17582_, _09120_, _05758_);
  or _68683_ (_17583_, _17582_, _10954_);
  and _68684_ (_17584_, _17583_, _17581_);
  nor _68685_ (_17585_, _10949_, _17584_);
  and _68686_ (_17586_, _10949_, _17584_);
  nor _68687_ (_17587_, _17586_, _17585_);
  nor _68688_ (_17588_, _16968_, _10954_);
  not _68689_ (_17589_, _17588_);
  or _68690_ (_17590_, _17589_, _17587_);
  and _68691_ (_17591_, _17590_, \oc8051_golden_model_1.PSW [7]);
  nor _68692_ (_17592_, _17587_, \oc8051_golden_model_1.PSW [7]);
  nor _68693_ (_17593_, _17592_, _17591_);
  and _68694_ (_17594_, _17589_, _17587_);
  or _68695_ (_17595_, _17594_, _13935_);
  or _68696_ (_17596_, _17595_, _17593_);
  and _68697_ (_17597_, _17596_, _06267_);
  and _68698_ (_17598_, _17597_, _17579_);
  and _68699_ (_17599_, _08077_, \oc8051_golden_model_1.ACC [1]);
  and _68700_ (_17600_, _08127_, _05758_);
  nor _68701_ (_17601_, _17600_, _13785_);
  nor _68702_ (_17602_, _17601_, _17599_);
  nor _68703_ (_17603_, _10991_, _17602_);
  and _68704_ (_17604_, _10991_, _17602_);
  nor _68705_ (_17605_, _17604_, _17603_);
  and _68706_ (_17606_, _12304_, \oc8051_golden_model_1.PSW [7]);
  not _68707_ (_17607_, _17606_);
  and _68708_ (_17608_, _17607_, _17605_);
  or _68709_ (_17609_, _17607_, _17605_);
  nand _68710_ (_17610_, _17609_, _10307_);
  or _68711_ (_17611_, _17610_, _17608_);
  and _68712_ (_17612_, _17611_, _12367_);
  or _68713_ (_17613_, _17612_, _17598_);
  nor _68714_ (_17614_, _17300_, _13874_);
  nor _68715_ (_17615_, _12318_, _17614_);
  and _68716_ (_17616_, _12318_, _17614_);
  nor _68717_ (_17617_, _17616_, _17615_);
  not _68718_ (_17618_, _17304_);
  or _68719_ (_17619_, _17618_, _17617_);
  nand _68720_ (_17620_, _17618_, _17617_);
  and _68721_ (_17621_, _17620_, _10306_);
  nand _68722_ (_17622_, _17621_, _17619_);
  and _68723_ (_17623_, _17622_, _17613_);
  or _68724_ (_17624_, _17623_, _05676_);
  nand _68725_ (_17625_, _06403_, _05676_);
  and _68726_ (_17626_, _17625_, _06027_);
  and _68727_ (_17627_, _17626_, _17624_);
  or _68728_ (_17628_, _17529_, _14525_);
  and _68729_ (_17629_, _17628_, _06026_);
  and _68730_ (_17630_, _17629_, _17531_);
  or _68731_ (_17631_, _17630_, _09818_);
  or _68732_ (_17632_, _17631_, _17627_);
  and _68733_ (_17633_, _09182_, _07701_);
  or _68734_ (_17634_, _17500_, _07012_);
  or _68735_ (_17635_, _17634_, _17633_);
  or _68736_ (_17636_, _17534_, _09827_);
  and _68737_ (_17637_, _17636_, _05669_);
  and _68738_ (_17638_, _17637_, _17635_);
  and _68739_ (_17639_, _17638_, _17632_);
  and _68740_ (_17640_, _14580_, _07701_);
  or _68741_ (_17641_, _17640_, _17500_);
  and _68742_ (_17642_, _17641_, _09833_);
  or _68743_ (_17643_, _17642_, _09832_);
  or _68744_ (_17644_, _17643_, _17639_);
  or _68745_ (_17645_, _10028_, _09839_);
  and _68746_ (_17646_, _17645_, _05664_);
  and _68747_ (_17647_, _17646_, _17644_);
  nor _68748_ (_17648_, _06403_, _05664_);
  or _68749_ (_17649_, _17648_, _06019_);
  or _68750_ (_17650_, _17649_, _17647_);
  and _68751_ (_17651_, _07701_, _08730_);
  or _68752_ (_17652_, _17651_, _17500_);
  or _68753_ (_17653_, _17652_, _06020_);
  and _68754_ (_17654_, _17653_, _10662_);
  and _68755_ (_17655_, _17654_, _17650_);
  and _68756_ (_17656_, _06094_, _05726_);
  nor _68757_ (_17657_, _10662_, _06403_);
  or _68758_ (_17658_, _17657_, _17656_);
  or _68759_ (_17659_, _17658_, _17655_);
  not _68760_ (_17660_, _17656_);
  or _68761_ (_17661_, _10909_, _17660_);
  and _68762_ (_17662_, _07266_, _05726_);
  not _68763_ (_17663_, _17662_);
  and _68764_ (_17664_, _17663_, _17661_);
  and _68765_ (_17665_, _17664_, _17659_);
  and _68766_ (_17666_, _06229_, _05726_);
  and _68767_ (_17667_, _17662_, _10909_);
  or _68768_ (_17668_, _17667_, _17666_);
  or _68769_ (_17669_, _17668_, _17665_);
  not _68770_ (_17670_, _17503_);
  not _68771_ (_17671_, _17666_);
  or _68772_ (_17672_, _10909_, _17671_);
  and _68773_ (_17673_, _17672_, _17670_);
  and _68774_ (_17674_, _17673_, _17669_);
  or _68775_ (_17675_, _17674_, _17504_);
  and _68776_ (_17676_, _17675_, _10687_);
  and _68777_ (_17677_, _10681_, _10909_);
  or _68778_ (_17678_, _17677_, _10685_);
  or _68779_ (_17679_, _17678_, _17676_);
  or _68780_ (_17680_, _10686_, _10949_);
  and _68781_ (_17681_, _17680_, _17679_);
  or _68782_ (_17682_, _17681_, _06282_);
  or _68783_ (_17683_, _10991_, _06283_);
  and _68784_ (_17684_, _17683_, _10699_);
  and _68785_ (_17685_, _17684_, _17682_);
  nor _68786_ (_17686_, _10699_, _11032_);
  or _68787_ (_17687_, _17686_, _06112_);
  or _68788_ (_17688_, _17687_, _17685_);
  and _68789_ (_17689_, _17688_, _17502_);
  or _68790_ (_17690_, _17689_, _06284_);
  or _68791_ (_17691_, _17500_, _08756_);
  and _68792_ (_17692_, _17691_, _17101_);
  and _68793_ (_17693_, _17692_, _17690_);
  and _68794_ (_17694_, _17104_, _10907_);
  or _68795_ (_17695_, _17694_, _10731_);
  or _68796_ (_17696_, _17695_, _17693_);
  or _68797_ (_17697_, _10736_, _10947_);
  and _68798_ (_17698_, _17697_, _10735_);
  and _68799_ (_17699_, _17698_, _17696_);
  or _68800_ (_17700_, _10741_, _10989_);
  and _68801_ (_17701_, _17700_, _10743_);
  or _68802_ (_17702_, _17701_, _17699_);
  or _68803_ (_17703_, _10747_, _11030_);
  and _68804_ (_17704_, _17703_, _07032_);
  and _68805_ (_17705_, _17704_, _17702_);
  nand _68806_ (_17706_, _17652_, _06108_);
  nor _68807_ (_17707_, _17706_, _10990_);
  or _68808_ (_17708_, _17707_, _10752_);
  or _68809_ (_17709_, _17708_, _17705_);
  nand _68810_ (_17710_, _10908_, _10752_);
  and _68811_ (_17711_, _17710_, _10760_);
  and _68812_ (_17712_, _17711_, _17709_);
  nor _68813_ (_17713_, _10760_, _10908_);
  or _68814_ (_17714_, _17713_, _10767_);
  or _68815_ (_17715_, _17714_, _17712_);
  nand _68816_ (_17716_, _10767_, _10908_);
  and _68817_ (_17717_, _17716_, _06668_);
  and _68818_ (_17718_, _17717_, _17715_);
  nor _68819_ (_17719_, _10908_, _06668_);
  or _68820_ (_17720_, _17719_, _10775_);
  or _68821_ (_17721_, _17720_, _17718_);
  nand _68822_ (_17722_, _10775_, _10948_);
  and _68823_ (_17723_, _17722_, _06291_);
  and _68824_ (_17724_, _17723_, _17721_);
  nand _68825_ (_17725_, _17136_, _10990_);
  and _68826_ (_17726_, _17725_, _11987_);
  or _68827_ (_17727_, _17726_, _17724_);
  nand _68828_ (_17728_, _10781_, _11031_);
  and _68829_ (_17729_, _17728_, _17727_);
  or _68830_ (_17730_, _17729_, _06130_);
  and _68831_ (_17731_, _14593_, _07701_);
  or _68832_ (_17732_, _17500_, _08777_);
  or _68833_ (_17733_, _17732_, _17731_);
  and _68834_ (_17734_, _17733_, _10304_);
  and _68835_ (_17735_, _17734_, _17730_);
  nand _68836_ (_17736_, _10289_, _10277_);
  nor _68837_ (_17737_, _10304_, _10290_);
  and _68838_ (_17738_, _17737_, _17736_);
  or _68839_ (_17739_, _17738_, _17409_);
  or _68840_ (_17740_, _17739_, _17735_);
  and _68841_ (_17741_, _10807_, _10534_);
  nor _68842_ (_17742_, _17741_, _10808_);
  or _68843_ (_17743_, _17742_, _17410_);
  and _68844_ (_17744_, _17743_, _17423_);
  and _68845_ (_17745_, _17744_, _17740_);
  nand _68846_ (_17746_, _17742_, _17416_);
  nand _68847_ (_17747_, _17746_, _06289_);
  or _68848_ (_17748_, _17747_, _17745_);
  and _68849_ (_17749_, _17748_, _17498_);
  nand _68850_ (_17750_, _10867_, _10604_);
  nor _68851_ (_17751_, _10868_, _10856_);
  and _68852_ (_17752_, _17751_, _17750_);
  or _68853_ (_17753_, _17752_, _10854_);
  or _68854_ (_17754_, _17753_, _17749_);
  nand _68855_ (_17755_, _10854_, _05784_);
  and _68856_ (_17756_, _17755_, _10890_);
  and _68857_ (_17757_, _17756_, _17754_);
  nor _68858_ (_17758_, _10916_, _10909_);
  nor _68859_ (_17759_, _17758_, _10917_);
  and _68860_ (_17760_, _17759_, _16956_);
  or _68861_ (_17761_, _17760_, _17437_);
  or _68862_ (_17762_, _17761_, _17757_);
  and _68863_ (_17763_, _10957_, _10950_);
  nor _68864_ (_17764_, _17763_, _10958_);
  and _68865_ (_17765_, _17764_, _17443_);
  or _68866_ (_17766_, _17765_, _10934_);
  and _68867_ (_17767_, _17766_, _17762_);
  and _68868_ (_17768_, _17764_, _06692_);
  or _68869_ (_17769_, _17768_, _06051_);
  or _68870_ (_17770_, _17769_, _17767_);
  and _68871_ (_17771_, _17770_, _17494_);
  nand _68872_ (_17772_, _11038_, _11032_);
  nor _68873_ (_17773_, _11039_, _11050_);
  and _68874_ (_17774_, _17773_, _17772_);
  or _68875_ (_17775_, _17774_, _11015_);
  or _68876_ (_17776_, _17775_, _17771_);
  and _68877_ (_17777_, _17776_, _17490_);
  or _68878_ (_17778_, _17777_, _06316_);
  or _68879_ (_17779_, _17519_, _06718_);
  and _68880_ (_17780_, _17779_, _11060_);
  and _68881_ (_17781_, _17780_, _17778_);
  nor _68882_ (_17782_, _17467_, _09956_);
  or _68883_ (_17783_, _17782_, _11065_);
  nor _68884_ (_17784_, _17783_, _11064_);
  nor _68885_ (_17785_, _17784_, _12756_);
  or _68886_ (_17786_, _17785_, _17781_);
  nand _68887_ (_17787_, _11064_, _10010_);
  and _68888_ (_17788_, _17787_, _05653_);
  and _68889_ (_17789_, _17788_, _17786_);
  and _68890_ (_17790_, _17551_, _05652_);
  or _68891_ (_17791_, _17790_, _06047_);
  or _68892_ (_17792_, _17791_, _17789_);
  and _68893_ (_17793_, _14657_, _07701_);
  or _68894_ (_17794_, _17793_, _17500_);
  or _68895_ (_17795_, _17794_, _06048_);
  and _68896_ (_17796_, _17795_, _11083_);
  and _68897_ (_17797_, _17796_, _17792_);
  nor _68898_ (_17798_, _11090_, \oc8051_golden_model_1.ACC [2]);
  nor _68899_ (_17799_, _17798_, _11091_);
  and _68900_ (_17800_, _17799_, _11082_);
  or _68901_ (_17801_, _17800_, _11089_);
  or _68902_ (_17802_, _17801_, _17797_);
  nand _68903_ (_17803_, _11089_, _10010_);
  and _68904_ (_17804_, _17803_, _01336_);
  and _68905_ (_17805_, _17804_, _17802_);
  or _68906_ (_17806_, _17805_, _17489_);
  and _68907_ (_43334_, _17806_, _42882_);
  nor _68908_ (_17807_, _01336_, _10010_);
  and _68909_ (_17808_, _10291_, _10271_);
  nor _68910_ (_17809_, _17808_, _10292_);
  or _68911_ (_17810_, _17809_, _10304_);
  nor _68912_ (_17811_, _17387_, _10906_);
  or _68913_ (_17812_, _17811_, _10775_);
  nand _68914_ (_17813_, _10906_, _06477_);
  or _68915_ (_17814_, _10987_, _10735_);
  and _68916_ (_17815_, _17814_, _10747_);
  and _68917_ (_17816_, _14793_, _07701_);
  nor _68918_ (_17817_, _07701_, _10010_);
  or _68919_ (_17818_, _17817_, _08751_);
  or _68920_ (_17819_, _17818_, _17816_);
  nor _68921_ (_17820_, _10945_, _10946_);
  or _68922_ (_17821_, _17820_, _06648_);
  nor _68923_ (_17822_, _10662_, _05983_);
  nand _68924_ (_17823_, _10378_, _07353_);
  nor _68925_ (_17824_, _08359_, _10010_);
  and _68926_ (_17825_, _14683_, _08359_);
  or _68927_ (_17826_, _17825_, _17824_);
  or _68928_ (_17827_, _17826_, _06044_);
  and _68929_ (_17828_, _17827_, _06848_);
  and _68930_ (_17829_, _14672_, _07701_);
  or _68931_ (_17830_, _17829_, _17817_);
  and _68932_ (_17831_, _17830_, _06102_);
  or _68933_ (_17832_, _17219_, _09181_);
  nor _68934_ (_17833_, _10400_, _07353_);
  nor _68935_ (_17834_, _06530_, _10010_);
  and _68936_ (_17835_, _06530_, _10010_);
  or _68937_ (_17836_, _17835_, _17834_);
  and _68938_ (_17837_, _17836_, _10400_);
  or _68939_ (_17838_, _17837_, _10389_);
  or _68940_ (_17839_, _17838_, _17833_);
  and _68941_ (_17840_, _17839_, _05698_);
  or _68942_ (_17841_, _17840_, _06948_);
  and _68943_ (_17842_, _17841_, _06954_);
  and _68944_ (_17843_, _17842_, _17832_);
  or _68945_ (_17844_, _17843_, _17831_);
  and _68946_ (_17845_, _17844_, _10413_);
  not _68947_ (_17846_, \oc8051_golden_model_1.PSW [6]);
  nor _68948_ (_17847_, _10415_, _17846_);
  nor _68949_ (_17848_, _17847_, \oc8051_golden_model_1.ACC [3]);
  nor _68950_ (_17849_, _17848_, _10416_);
  and _68951_ (_17850_, _17849_, _10412_);
  or _68952_ (_17851_, _17850_, _06043_);
  or _68953_ (_17852_, _17851_, _17845_);
  and _68954_ (_17853_, _17852_, _17828_);
  nor _68955_ (_17854_, _10439_, _07353_);
  or _68956_ (_17855_, _17854_, _17817_);
  and _68957_ (_17856_, _17855_, _06239_);
  or _68958_ (_17857_, _17856_, _10378_);
  or _68959_ (_17858_, _17857_, _17853_);
  and _68960_ (_17859_, _17858_, _17823_);
  or _68961_ (_17860_, _17859_, _06970_);
  or _68962_ (_17861_, _09181_, _06971_);
  and _68963_ (_17862_, _17861_, _06220_);
  and _68964_ (_17863_, _17862_, _17860_);
  nor _68965_ (_17864_, _08028_, _06220_);
  or _68966_ (_17865_, _17864_, _10376_);
  or _68967_ (_17866_, _17865_, _17863_);
  nand _68968_ (_17867_, _10376_, _08393_);
  and _68969_ (_17868_, _17867_, _17866_);
  or _68970_ (_17869_, _17868_, _06039_);
  and _68971_ (_17870_, _14681_, _08359_);
  or _68972_ (_17871_, _17870_, _17824_);
  or _68973_ (_17872_, _17871_, _06040_);
  and _68974_ (_17873_, _17872_, _06033_);
  and _68975_ (_17874_, _17873_, _17869_);
  or _68976_ (_17875_, _17824_, _14708_);
  and _68977_ (_17876_, _17826_, _06032_);
  and _68978_ (_17877_, _17876_, _17875_);
  or _68979_ (_17878_, _17877_, _17874_);
  and _68980_ (_17879_, _17878_, _09800_);
  or _68981_ (_17880_, _09750_, _09748_);
  nor _68982_ (_17881_, _09751_, _09800_);
  and _68983_ (_17882_, _17881_, _17880_);
  or _68984_ (_17883_, _17882_, _10468_);
  or _68985_ (_17884_, _17883_, _17879_);
  and _68986_ (_17885_, _07530_, \oc8051_golden_model_1.ACC [2]);
  nor _68987_ (_17886_, _17569_, _17885_);
  nor _68988_ (_17887_, _10905_, _10906_);
  and _68989_ (_17888_, _17887_, _17886_);
  nor _68990_ (_17889_, _17887_, _17886_);
  or _68991_ (_17890_, _17889_, _17888_);
  nor _68992_ (_17891_, _17890_, _10606_);
  and _68993_ (_17892_, _17890_, _10606_);
  nor _68994_ (_17893_, _17892_, _17891_);
  and _68995_ (_17894_, _17571_, \oc8051_golden_model_1.PSW [7]);
  nor _68996_ (_17895_, _17572_, _10606_);
  nor _68997_ (_17896_, _17895_, _17894_);
  not _68998_ (_17897_, _17896_);
  and _68999_ (_17898_, _17897_, _17893_);
  nor _69000_ (_17899_, _17897_, _17893_);
  nor _69001_ (_17900_, _17899_, _17898_);
  or _69002_ (_17901_, _17900_, _10469_);
  and _69003_ (_17902_, _17901_, _17884_);
  or _69004_ (_17903_, _17902_, _12361_);
  and _69005_ (_17904_, _09030_, \oc8051_golden_model_1.ACC [2]);
  nor _69006_ (_17905_, _17585_, _17904_);
  and _69007_ (_17906_, _17820_, _17905_);
  nor _69008_ (_17907_, _17820_, _17905_);
  or _69009_ (_17908_, _17907_, _17906_);
  or _69010_ (_17909_, _17908_, _10606_);
  nand _69011_ (_17910_, _17908_, _10606_);
  and _69012_ (_17911_, _17910_, _17909_);
  and _69013_ (_17912_, _17911_, _17591_);
  nor _69014_ (_17913_, _17911_, _17591_);
  nor _69015_ (_17914_, _17913_, _17912_);
  or _69016_ (_17915_, _17914_, _13935_);
  and _69017_ (_17916_, _17915_, _06267_);
  and _69018_ (_17917_, _17916_, _17903_);
  and _69019_ (_17918_, _12305_, \oc8051_golden_model_1.PSW [7]);
  and _69020_ (_17919_, _08176_, \oc8051_golden_model_1.ACC [2]);
  nor _69021_ (_17920_, _17603_, _17919_);
  nor _69022_ (_17921_, _12299_, _17920_);
  and _69023_ (_17922_, _12299_, _17920_);
  nor _69024_ (_17923_, _17922_, _17921_);
  and _69025_ (_17924_, _17609_, _17923_);
  or _69026_ (_17925_, _17924_, _10306_);
  or _69027_ (_17926_, _17925_, _17918_);
  and _69028_ (_17927_, _17926_, _12367_);
  or _69029_ (_17928_, _17927_, _17917_);
  and _69030_ (_17929_, _06403_, \oc8051_golden_model_1.ACC [2]);
  nor _69031_ (_17930_, _17615_, _17929_);
  nor _69032_ (_17931_, _12319_, _17930_);
  and _69033_ (_17932_, _12319_, _17930_);
  nor _69034_ (_17933_, _17932_, _17931_);
  and _69035_ (_17934_, _17619_, _17933_);
  nor _69036_ (_17935_, _17619_, _17933_);
  or _69037_ (_17936_, _17935_, _10307_);
  or _69038_ (_17937_, _17936_, _17934_);
  and _69039_ (_17938_, _17937_, _17928_);
  or _69040_ (_17939_, _17938_, _05676_);
  nand _69041_ (_17940_, _05983_, _05676_);
  and _69042_ (_17941_, _17940_, _06027_);
  and _69043_ (_17942_, _17941_, _17939_);
  and _69044_ (_17943_, _14724_, _08359_);
  or _69045_ (_17944_, _17943_, _17824_);
  and _69046_ (_17945_, _17944_, _06026_);
  or _69047_ (_17946_, _17945_, _09818_);
  or _69048_ (_17947_, _17946_, _17942_);
  and _69049_ (_17948_, _09181_, _07701_);
  or _69050_ (_17949_, _17817_, _07012_);
  or _69051_ (_17950_, _17949_, _17948_);
  or _69052_ (_17951_, _17855_, _09827_);
  and _69053_ (_17952_, _17951_, _05669_);
  and _69054_ (_17953_, _17952_, _17950_);
  and _69055_ (_17954_, _17953_, _17947_);
  and _69056_ (_17955_, _14778_, _07701_);
  or _69057_ (_17956_, _17955_, _17817_);
  and _69058_ (_17957_, _17956_, _09833_);
  or _69059_ (_17958_, _17957_, _09832_);
  or _69060_ (_17959_, _17958_, _17954_);
  or _69061_ (_17960_, _09976_, _09839_);
  and _69062_ (_17961_, _17960_, _05664_);
  and _69063_ (_17962_, _17961_, _17959_);
  nor _69064_ (_17963_, _05983_, _05664_);
  or _69065_ (_17964_, _17963_, _06019_);
  or _69066_ (_17965_, _17964_, _17962_);
  and _69067_ (_17966_, _07701_, _08662_);
  or _69068_ (_17967_, _17966_, _17817_);
  or _69069_ (_17968_, _17967_, _06020_);
  and _69070_ (_17969_, _17968_, _10662_);
  and _69071_ (_17970_, _17969_, _17965_);
  or _69072_ (_17971_, _17970_, _17822_);
  and _69073_ (_17972_, _17971_, _17660_);
  and _69074_ (_17973_, _17887_, _17656_);
  or _69075_ (_17974_, _17973_, _17972_);
  and _69076_ (_17975_, _17974_, _17663_);
  and _69077_ (_17976_, _17662_, _17887_);
  or _69078_ (_17977_, _17976_, _17975_);
  and _69079_ (_17978_, _17977_, _17671_);
  and _69080_ (_17979_, _17887_, _17666_);
  or _69081_ (_17980_, _17979_, _17978_);
  and _69082_ (_17981_, _17980_, _17670_);
  and _69083_ (_17982_, _17887_, _17503_);
  or _69084_ (_17983_, _17982_, _17981_);
  and _69085_ (_17984_, _17983_, _16972_);
  and _69086_ (_17985_, _16971_, _17887_);
  or _69087_ (_17986_, _17985_, _06650_);
  or _69088_ (_17987_, _17986_, _17984_);
  and _69089_ (_17988_, _10394_, _05726_);
  nor _69090_ (_17989_, _17887_, _16970_);
  nor _69091_ (_17990_, _17989_, _17988_);
  and _69092_ (_17991_, _17990_, _17987_);
  or _69093_ (_17992_, _17820_, _06647_);
  and _69094_ (_17993_, _17992_, _10685_);
  or _69095_ (_17994_, _17993_, _17991_);
  and _69096_ (_17995_, _17994_, _17821_);
  or _69097_ (_17996_, _17995_, _06282_);
  or _69098_ (_17997_, _12299_, _06283_);
  and _69099_ (_17999_, _17997_, _10699_);
  and _69100_ (_18000_, _17999_, _17996_);
  and _69101_ (_18001_, _10698_, _12319_);
  or _69102_ (_18002_, _18001_, _06112_);
  or _69103_ (_18003_, _18002_, _18000_);
  nand _69104_ (_18004_, _18003_, _17819_);
  and _69105_ (_18005_, _18004_, _08756_);
  nor _69106_ (_18006_, _17817_, _08756_);
  or _69107_ (_18007_, _18006_, _11996_);
  or _69108_ (_18008_, _18007_, _18005_);
  nor _69109_ (_18009_, _11999_, _11998_);
  nand _69110_ (_18010_, _11996_, _10905_);
  and _69111_ (_18011_, _18010_, _18009_);
  and _69112_ (_18012_, _18011_, _18008_);
  nor _69113_ (_18013_, _18009_, _10905_);
  or _69114_ (_18014_, _18013_, _18012_);
  and _69115_ (_18015_, _18014_, _10736_);
  nor _69116_ (_18016_, _10736_, _10945_);
  or _69117_ (_18017_, _18016_, _18015_);
  nand _69118_ (_18018_, _18017_, _10735_);
  and _69119_ (_18019_, _18018_, _17815_);
  and _69120_ (_18020_, _10741_, _11028_);
  or _69121_ (_18021_, _18020_, _18019_);
  and _69122_ (_18022_, _18021_, _07032_);
  nand _69123_ (_18023_, _17967_, _06108_);
  nor _69124_ (_18024_, _18023_, _10988_);
  or _69125_ (_18025_, _18024_, _06477_);
  or _69126_ (_18026_, _18025_, _18022_);
  and _69127_ (_18027_, _18026_, _17813_);
  or _69128_ (_18028_, _18027_, _06834_);
  nand _69129_ (_18029_, _10906_, _06834_);
  and _69130_ (_18030_, _18029_, _17387_);
  and _69131_ (_18031_, _18030_, _18028_);
  or _69132_ (_18032_, _18031_, _17812_);
  nand _69133_ (_18033_, _10775_, _10946_);
  and _69134_ (_18034_, _18033_, _06291_);
  and _69135_ (_18035_, _18034_, _18032_);
  nor _69136_ (_18036_, _10988_, _06291_);
  or _69137_ (_18037_, _18036_, _10781_);
  or _69138_ (_18038_, _18037_, _18035_);
  nand _69139_ (_18039_, _10781_, _11029_);
  and _69140_ (_18040_, _18039_, _08777_);
  and _69141_ (_18041_, _18040_, _18038_);
  and _69142_ (_18042_, _14792_, _07701_);
  or _69143_ (_18043_, _18042_, _17817_);
  and _69144_ (_18044_, _18043_, _06130_);
  or _69145_ (_18045_, _18044_, _10303_);
  or _69146_ (_18046_, _18045_, _18041_);
  and _69147_ (_18047_, _18046_, _17810_);
  or _69148_ (_18048_, _18047_, _10794_);
  and _69149_ (_18049_, _10809_, _10528_);
  nor _69150_ (_18050_, _18049_, _10810_);
  or _69151_ (_18051_, _18050_, _10796_);
  and _69152_ (_18052_, _18051_, _06289_);
  and _69153_ (_18053_, _18052_, _18048_);
  and _69154_ (_18054_, _10839_, _10341_);
  nor _69155_ (_18055_, _18054_, _10840_);
  or _69156_ (_18056_, _18055_, _10824_);
  and _69157_ (_18057_, _18056_, _10826_);
  or _69158_ (_18058_, _18057_, _18053_);
  and _69159_ (_18059_, _10869_, _10598_);
  nor _69160_ (_18060_, _18059_, _10870_);
  or _69161_ (_18061_, _18060_, _10856_);
  and _69162_ (_18062_, _18061_, _10855_);
  and _69163_ (_18063_, _18062_, _18058_);
  nand _69164_ (_18064_, _10854_, \oc8051_golden_model_1.ACC [2]);
  nand _69165_ (_18065_, _18064_, _10889_);
  or _69166_ (_18066_, _18065_, _18063_);
  nor _69167_ (_18067_, _10918_, _17887_);
  and _69168_ (_18068_, _10918_, _17887_);
  or _69169_ (_18069_, _18068_, _18067_);
  or _69170_ (_18070_, _18069_, _10889_);
  and _69171_ (_18071_, _18070_, _10886_);
  and _69172_ (_18072_, _18071_, _18066_);
  and _69173_ (_18073_, _18069_, _10885_);
  or _69174_ (_18074_, _18073_, _10932_);
  or _69175_ (_18075_, _18074_, _18072_);
  and _69176_ (_18076_, _10959_, _17820_);
  nor _69177_ (_18077_, _10959_, _17820_);
  or _69178_ (_18078_, _18077_, _18076_);
  or _69179_ (_18079_, _18078_, _10934_);
  and _69180_ (_18080_, _18079_, _06052_);
  and _69181_ (_18081_, _18080_, _18075_);
  and _69182_ (_18082_, _11000_, _12299_);
  nor _69183_ (_18083_, _11000_, _12299_);
  or _69184_ (_18084_, _18083_, _18082_);
  and _69185_ (_18085_, _18084_, _06051_);
  or _69186_ (_18086_, _18085_, _10974_);
  or _69187_ (_18087_, _18086_, _18081_);
  and _69188_ (_18088_, _11040_, _12319_);
  nor _69189_ (_18089_, _11040_, _12319_);
  or _69190_ (_18090_, _18089_, _18088_);
  or _69191_ (_18091_, _18090_, _11050_);
  and _69192_ (_18092_, _18091_, _11016_);
  and _69193_ (_18093_, _18092_, _18087_);
  and _69194_ (_18094_, _11015_, \oc8051_golden_model_1.ACC [2]);
  or _69195_ (_18095_, _18094_, _06316_);
  or _69196_ (_18096_, _18095_, _18093_);
  or _69197_ (_18097_, _17830_, _06718_);
  and _69198_ (_18098_, _18097_, _11060_);
  and _69199_ (_18099_, _18098_, _18096_);
  nor _69200_ (_18100_, _11065_, _10010_);
  or _69201_ (_18101_, _18100_, _11066_);
  and _69202_ (_18102_, _18101_, _11059_);
  or _69203_ (_18103_, _18102_, _11064_);
  or _69204_ (_18104_, _18103_, _18099_);
  nand _69205_ (_18105_, _11064_, _09880_);
  and _69206_ (_18106_, _18105_, _05653_);
  and _69207_ (_18107_, _18106_, _18104_);
  and _69208_ (_18108_, _17871_, _05652_);
  or _69209_ (_18109_, _18108_, _06047_);
  or _69210_ (_18110_, _18109_, _18107_);
  and _69211_ (_18111_, _14849_, _07701_);
  or _69212_ (_18112_, _17817_, _06048_);
  or _69213_ (_18113_, _18112_, _18111_);
  and _69214_ (_18114_, _18113_, _11083_);
  and _69215_ (_18115_, _18114_, _18110_);
  nor _69216_ (_18116_, _11091_, \oc8051_golden_model_1.ACC [3]);
  nor _69217_ (_18117_, _18116_, _11092_);
  and _69218_ (_18118_, _18117_, _11082_);
  or _69219_ (_18119_, _18118_, _11089_);
  or _69220_ (_18120_, _18119_, _18115_);
  nand _69221_ (_18121_, _11089_, _09880_);
  and _69222_ (_18122_, _18121_, _01336_);
  and _69223_ (_18123_, _18122_, _18120_);
  or _69224_ (_18124_, _18123_, _17807_);
  and _69225_ (_43335_, _18124_, _42882_);
  nor _69226_ (_18125_, _01336_, _09880_);
  not _69227_ (_18126_, _17437_);
  or _69228_ (_18127_, _10961_, _10944_);
  and _69229_ (_18128_, _18127_, _10962_);
  or _69230_ (_18129_, _18128_, _18126_);
  and _69231_ (_18130_, _14876_, _07701_);
  nor _69232_ (_18131_, _07701_, _09880_);
  or _69233_ (_18132_, _18131_, _08751_);
  or _69234_ (_18133_, _18132_, _18130_);
  or _69235_ (_18134_, _10686_, _10944_);
  and _69236_ (_18135_, _06095_, _05661_);
  and _69237_ (_18136_, _18135_, _05726_);
  not _69238_ (_18137_, _17909_);
  or _69239_ (_18138_, _17912_, _18137_);
  and _69240_ (_18139_, _09181_, _10010_);
  or _69241_ (_18140_, _09181_, _10010_);
  and _69242_ (_18141_, _18140_, _17905_);
  or _69243_ (_18142_, _18141_, _18139_);
  nor _69244_ (_18143_, _10944_, _18142_);
  and _69245_ (_18144_, _10944_, _18142_);
  or _69246_ (_18145_, _18144_, _18143_);
  or _69247_ (_18146_, _18145_, _10606_);
  nand _69248_ (_18147_, _18145_, _10606_);
  and _69249_ (_18148_, _18147_, _18146_);
  and _69250_ (_18149_, _18148_, _18138_);
  nor _69251_ (_18150_, _18148_, _18138_);
  nor _69252_ (_18151_, _18150_, _18149_);
  or _69253_ (_18152_, _18151_, _13935_);
  nand _69254_ (_18153_, _10378_, _08270_);
  nor _69255_ (_18154_, _08359_, _09880_);
  and _69256_ (_18155_, _14878_, _08359_);
  or _69257_ (_18156_, _18155_, _18154_);
  or _69258_ (_18157_, _18156_, _06044_);
  and _69259_ (_18158_, _18157_, _06848_);
  and _69260_ (_18159_, _14887_, _07701_);
  or _69261_ (_18160_, _18159_, _18131_);
  and _69262_ (_18161_, _18160_, _06102_);
  or _69263_ (_18162_, _10390_, _09180_);
  nor _69264_ (_18163_, _10400_, _08270_);
  or _69265_ (_18164_, _06530_, \oc8051_golden_model_1.ACC [4]);
  nand _69266_ (_18165_, _06530_, \oc8051_golden_model_1.ACC [4]);
  and _69267_ (_18166_, _18165_, _18164_);
  and _69268_ (_18167_, _18166_, _10400_);
  or _69269_ (_18168_, _18167_, _10389_);
  or _69270_ (_18169_, _18168_, _18163_);
  and _69271_ (_18170_, _18169_, _10408_);
  and _69272_ (_18171_, _18170_, _18162_);
  or _69273_ (_18172_, _18171_, _18161_);
  and _69274_ (_18173_, _18172_, _10413_);
  nor _69275_ (_18174_, _10416_, \oc8051_golden_model_1.ACC [4]);
  nor _69276_ (_18175_, _18174_, _10417_);
  and _69277_ (_18176_, _18175_, _10412_);
  or _69278_ (_18177_, _18176_, _06043_);
  or _69279_ (_18178_, _18177_, _18173_);
  and _69280_ (_18179_, _18178_, _18158_);
  nor _69281_ (_18180_, _08270_, _10439_);
  or _69282_ (_18181_, _18180_, _18131_);
  and _69283_ (_18182_, _18181_, _06239_);
  or _69284_ (_18183_, _18182_, _10378_);
  or _69285_ (_18184_, _18183_, _18179_);
  and _69286_ (_18185_, _18184_, _18153_);
  or _69287_ (_18186_, _18185_, _06970_);
  or _69288_ (_18187_, _09180_, _06971_);
  and _69289_ (_18189_, _18187_, _06220_);
  and _69290_ (_18190_, _18189_, _18186_);
  nor _69291_ (_18191_, _08272_, _06220_);
  or _69292_ (_18192_, _18191_, _10376_);
  or _69293_ (_18193_, _18192_, _18190_);
  nand _69294_ (_18194_, _10376_, _05758_);
  and _69295_ (_18195_, _18194_, _18193_);
  or _69296_ (_18196_, _18195_, _06039_);
  and _69297_ (_18197_, _14882_, _08359_);
  or _69298_ (_18198_, _18197_, _18154_);
  or _69299_ (_18200_, _18198_, _06040_);
  and _69300_ (_18201_, _18200_, _06033_);
  and _69301_ (_18202_, _18201_, _18196_);
  or _69302_ (_18203_, _18154_, _14914_);
  and _69303_ (_18204_, _18156_, _06032_);
  and _69304_ (_18205_, _18204_, _18203_);
  or _69305_ (_18206_, _18205_, _09269_);
  or _69306_ (_18207_, _18206_, _18202_);
  nor _69307_ (_18208_, _09753_, _09751_);
  nor _69308_ (_18209_, _18208_, _09754_);
  or _69309_ (_18211_, _18209_, _09800_);
  and _69310_ (_18212_, _18211_, _10469_);
  and _69311_ (_18213_, _18212_, _18207_);
  or _69312_ (_18214_, _17898_, _17891_);
  nor _69313_ (_18215_, _07353_, \oc8051_golden_model_1.ACC [3]);
  nand _69314_ (_18216_, _07353_, \oc8051_golden_model_1.ACC [3]);
  and _69315_ (_18217_, _18216_, _17886_);
  or _69316_ (_18218_, _18217_, _18215_);
  nor _69317_ (_18219_, _10904_, _18218_);
  and _69318_ (_18220_, _10904_, _18218_);
  nor _69319_ (_18222_, _18220_, _18219_);
  and _69320_ (_18223_, _18222_, \oc8051_golden_model_1.PSW [7]);
  nor _69321_ (_18224_, _18222_, \oc8051_golden_model_1.PSW [7]);
  nor _69322_ (_18225_, _18224_, _18223_);
  or _69323_ (_18226_, _18225_, _18214_);
  and _69324_ (_18227_, _18225_, _18214_);
  nor _69325_ (_18228_, _18227_, _10469_);
  and _69326_ (_18229_, _18228_, _18226_);
  or _69327_ (_18230_, _18229_, _12361_);
  or _69328_ (_18231_, _18230_, _18213_);
  and _69329_ (_18233_, _18231_, _18152_);
  or _69330_ (_18234_, _18233_, _06261_);
  nor _69331_ (_18235_, _12305_, _10606_);
  or _69332_ (_18236_, _17920_, _13781_);
  and _69333_ (_18237_, _18236_, _13780_);
  nor _69334_ (_18238_, _10986_, _18237_);
  and _69335_ (_18239_, _10986_, _18237_);
  nor _69336_ (_18240_, _18239_, _18238_);
  and _69337_ (_18241_, _18240_, \oc8051_golden_model_1.PSW [7]);
  nor _69338_ (_18242_, _18240_, \oc8051_golden_model_1.PSW [7]);
  nor _69339_ (_18244_, _18242_, _18241_);
  and _69340_ (_18245_, _18244_, _18235_);
  nor _69341_ (_18246_, _18244_, _18235_);
  nor _69342_ (_18247_, _18246_, _18245_);
  or _69343_ (_18248_, _18247_, _06267_);
  and _69344_ (_18249_, _18248_, _10307_);
  and _69345_ (_18250_, _18249_, _18234_);
  nor _69346_ (_18251_, _12324_, _10606_);
  or _69347_ (_18252_, _17930_, _13880_);
  and _69348_ (_18253_, _18252_, _13879_);
  nor _69349_ (_18255_, _11027_, _18253_);
  and _69350_ (_18256_, _11027_, _18253_);
  nor _69351_ (_18257_, _18256_, _18255_);
  and _69352_ (_18258_, _18257_, \oc8051_golden_model_1.PSW [7]);
  nor _69353_ (_18259_, _18257_, \oc8051_golden_model_1.PSW [7]);
  nor _69354_ (_18260_, _18259_, _18258_);
  or _69355_ (_18261_, _18260_, _18251_);
  and _69356_ (_18262_, _18260_, _18251_);
  nor _69357_ (_18263_, _18262_, _10307_);
  and _69358_ (_18264_, _18263_, _18261_);
  or _69359_ (_18266_, _18264_, _05676_);
  or _69360_ (_18267_, _18266_, _18250_);
  nand _69361_ (_18268_, _06758_, _05676_);
  and _69362_ (_18269_, _18268_, _06027_);
  and _69363_ (_18270_, _18269_, _18267_);
  or _69364_ (_18271_, _18154_, _14879_);
  and _69365_ (_18272_, _18271_, _06026_);
  and _69366_ (_18273_, _18272_, _18156_);
  or _69367_ (_18274_, _18273_, _09818_);
  or _69368_ (_18275_, _18274_, _18270_);
  and _69369_ (_18277_, _09180_, _07701_);
  or _69370_ (_18278_, _18131_, _07012_);
  or _69371_ (_18279_, _18278_, _18277_);
  or _69372_ (_18280_, _18181_, _09827_);
  and _69373_ (_18281_, _18280_, _05669_);
  and _69374_ (_18282_, _18281_, _18279_);
  and _69375_ (_18283_, _18282_, _18275_);
  and _69376_ (_18284_, _14983_, _07701_);
  or _69377_ (_18285_, _18284_, _18131_);
  and _69378_ (_18286_, _18285_, _09833_);
  or _69379_ (_18288_, _18286_, _09832_);
  or _69380_ (_18289_, _18288_, _18283_);
  or _69381_ (_18290_, _09924_, _09839_);
  and _69382_ (_18291_, _18290_, _05664_);
  and _69383_ (_18292_, _18291_, _18289_);
  nor _69384_ (_18293_, _06758_, _05664_);
  or _69385_ (_18294_, _18293_, _06019_);
  or _69386_ (_18295_, _18294_, _18292_);
  and _69387_ (_18296_, _08665_, _07701_);
  or _69388_ (_18297_, _18296_, _18131_);
  or _69389_ (_18299_, _18297_, _06020_);
  and _69390_ (_18300_, _18299_, _10662_);
  and _69391_ (_18301_, _18300_, _18295_);
  nor _69392_ (_18302_, _10662_, _06758_);
  or _69393_ (_18303_, _18302_, _17656_);
  or _69394_ (_18304_, _18303_, _18301_);
  not _69395_ (_18305_, _06649_);
  or _69396_ (_18306_, _10904_, _17660_);
  and _69397_ (_18307_, _18306_, _18305_);
  and _69398_ (_18308_, _18307_, _18304_);
  and _69399_ (_18310_, _06098_, _05726_);
  and _69400_ (_18311_, _10904_, _06649_);
  or _69401_ (_18312_, _18311_, _18310_);
  or _69402_ (_18313_, _18312_, _18308_);
  and _69403_ (_18314_, _06136_, _05726_);
  not _69404_ (_18315_, _18314_);
  not _69405_ (_18316_, _18310_);
  or _69406_ (_18317_, _10904_, _18316_);
  and _69407_ (_18318_, _18317_, _18315_);
  and _69408_ (_18319_, _18318_, _18313_);
  and _69409_ (_18321_, _10904_, _18314_);
  or _69410_ (_18322_, _18321_, _17666_);
  or _69411_ (_18323_, _18322_, _18319_);
  or _69412_ (_18324_, _10904_, _17671_);
  nand _69413_ (_18325_, _18324_, _18323_);
  nor _69414_ (_18326_, _18325_, _18136_);
  and _69415_ (_18327_, _18136_, _10904_);
  or _69416_ (_18328_, _18327_, _10685_);
  or _69417_ (_18329_, _18328_, _18326_);
  and _69418_ (_18330_, _18329_, _18134_);
  or _69419_ (_18332_, _18330_, _06282_);
  or _69420_ (_18333_, _10986_, _06283_);
  and _69421_ (_18334_, _18333_, _10699_);
  and _69422_ (_18335_, _18334_, _18332_);
  nor _69423_ (_18336_, _10699_, _11026_);
  or _69424_ (_18337_, _18336_, _06112_);
  or _69425_ (_18338_, _18337_, _18335_);
  nand _69426_ (_18339_, _18338_, _18133_);
  and _69427_ (_18340_, _18339_, _08756_);
  nor _69428_ (_18341_, _18131_, _08756_);
  or _69429_ (_18343_, _18341_, _11996_);
  or _69430_ (_18344_, _18343_, _18340_);
  and _69431_ (_18345_, _18135_, _05735_);
  or _69432_ (_18346_, _18345_, _10901_);
  nand _69433_ (_18347_, _18346_, _17104_);
  and _69434_ (_18348_, _18347_, _18344_);
  and _69435_ (_18349_, _18345_, _10903_);
  or _69436_ (_18350_, _18349_, _10731_);
  nor _69437_ (_18351_, _18350_, _18348_);
  nor _69438_ (_18352_, _10736_, _10942_);
  or _69439_ (_18354_, _18352_, _06279_);
  or _69440_ (_18355_, _18354_, _18351_);
  or _69441_ (_18356_, _10983_, _10735_);
  and _69442_ (_18357_, _18356_, _10747_);
  and _69443_ (_18358_, _18357_, _18355_);
  and _69444_ (_18359_, _10741_, _11023_);
  or _69445_ (_18360_, _18359_, _18358_);
  and _69446_ (_18361_, _18360_, _07032_);
  nand _69447_ (_18362_, _18297_, _06108_);
  nor _69448_ (_18363_, _18362_, _10985_);
  or _69449_ (_18364_, _18363_, _10752_);
  or _69450_ (_18365_, _18364_, _18361_);
  or _69451_ (_18366_, _10902_, _17205_);
  and _69452_ (_18367_, _18366_, _10760_);
  and _69453_ (_18368_, _18367_, _18365_);
  and _69454_ (_18369_, _10759_, _10902_);
  or _69455_ (_18370_, _18369_, _10767_);
  or _69456_ (_18371_, _18370_, _18368_);
  or _69457_ (_18372_, _10766_, _10902_);
  and _69458_ (_18373_, _18372_, _06668_);
  and _69459_ (_18375_, _18373_, _18371_);
  and _69460_ (_18376_, _10902_, _06667_);
  or _69461_ (_18377_, _18376_, _10775_);
  or _69462_ (_18378_, _18377_, _18375_);
  or _69463_ (_18379_, _17395_, _10943_);
  and _69464_ (_18380_, _18379_, _06291_);
  and _69465_ (_18381_, _18380_, _18378_);
  nor _69466_ (_18382_, _10985_, _06291_);
  or _69467_ (_18383_, _18382_, _10781_);
  or _69468_ (_18384_, _18383_, _18381_);
  nand _69469_ (_18386_, _10781_, _11025_);
  and _69470_ (_18387_, _18386_, _18384_);
  or _69471_ (_18388_, _18387_, _06130_);
  and _69472_ (_18389_, _14873_, _07701_);
  or _69473_ (_18390_, _18131_, _08777_);
  or _69474_ (_18391_, _18390_, _18389_);
  and _69475_ (_18392_, _18391_, _10304_);
  and _69476_ (_18393_, _18392_, _18388_);
  or _69477_ (_18394_, _10293_, _10265_);
  and _69478_ (_18395_, _10303_, _10294_);
  and _69479_ (_18397_, _18395_, _18394_);
  or _69480_ (_18398_, _18397_, _17409_);
  or _69481_ (_18399_, _18398_, _18393_);
  or _69482_ (_18400_, _10811_, _10521_);
  and _69483_ (_18401_, _18400_, _10812_);
  or _69484_ (_18402_, _18401_, _17410_);
  and _69485_ (_18403_, _18402_, _17423_);
  and _69486_ (_18404_, _18403_, _18399_);
  and _69487_ (_18405_, _18401_, _17416_);
  or _69488_ (_18406_, _18405_, _06288_);
  or _69489_ (_18408_, _18406_, _18404_);
  or _69490_ (_18409_, _10841_, _10335_);
  and _69491_ (_18410_, _18409_, _10842_);
  or _69492_ (_18411_, _18410_, _06289_);
  and _69493_ (_18412_, _18411_, _10856_);
  and _69494_ (_18413_, _18412_, _18408_);
  or _69495_ (_18414_, _10871_, _10592_);
  and _69496_ (_18415_, _18414_, _10872_);
  and _69497_ (_18416_, _18415_, _10824_);
  or _69498_ (_18417_, _18416_, _10854_);
  or _69499_ (_18419_, _18417_, _18413_);
  nand _69500_ (_18420_, _10854_, _10010_);
  and _69501_ (_18421_, _18420_, _10890_);
  and _69502_ (_18422_, _18421_, _18419_);
  or _69503_ (_18423_, _10920_, _10904_);
  nor _69504_ (_18424_, _10921_, _10890_);
  and _69505_ (_18425_, _18424_, _18423_);
  or _69506_ (_18426_, _18425_, _17437_);
  or _69507_ (_18427_, _18426_, _18422_);
  and _69508_ (_18428_, _18427_, _18129_);
  or _69509_ (_18430_, _18428_, _06692_);
  or _69510_ (_18431_, _18128_, _17443_);
  and _69511_ (_18432_, _18431_, _10975_);
  and _69512_ (_18433_, _18432_, _18430_);
  or _69513_ (_18434_, _11002_, _10986_);
  and _69514_ (_18435_, _11003_, _06051_);
  and _69515_ (_18436_, _18435_, _18434_);
  or _69516_ (_18437_, _11042_, _11027_);
  and _69517_ (_18438_, _11043_, _10974_);
  and _69518_ (_18439_, _18438_, _18437_);
  or _69519_ (_18441_, _18439_, _11015_);
  or _69520_ (_18442_, _18441_, _18436_);
  or _69521_ (_18443_, _18442_, _18433_);
  nand _69522_ (_18444_, _11015_, _10010_);
  and _69523_ (_18445_, _18444_, _18443_);
  or _69524_ (_18446_, _18445_, _06316_);
  or _69525_ (_18447_, _18160_, _06718_);
  and _69526_ (_18448_, _18447_, _11060_);
  and _69527_ (_18449_, _18448_, _18446_);
  nor _69528_ (_18450_, _11066_, _09880_);
  or _69529_ (_18452_, _18450_, _11067_);
  and _69530_ (_18453_, _18452_, _11059_);
  or _69531_ (_18454_, _18453_, _11064_);
  or _69532_ (_18455_, _18454_, _18449_);
  nand _69533_ (_18456_, _11064_, _09906_);
  and _69534_ (_18457_, _18456_, _05653_);
  and _69535_ (_18458_, _18457_, _18455_);
  and _69536_ (_18459_, _18198_, _05652_);
  or _69537_ (_18460_, _18459_, _06047_);
  or _69538_ (_18461_, _18460_, _18458_);
  and _69539_ (_18463_, _15055_, _07701_);
  or _69540_ (_18464_, _18131_, _06048_);
  or _69541_ (_18465_, _18464_, _18463_);
  and _69542_ (_18466_, _18465_, _11083_);
  and _69543_ (_18467_, _18466_, _18461_);
  nor _69544_ (_18468_, _11092_, \oc8051_golden_model_1.ACC [4]);
  nor _69545_ (_18469_, _18468_, _11093_);
  and _69546_ (_18470_, _18469_, _11082_);
  or _69547_ (_18471_, _18470_, _11089_);
  or _69548_ (_18472_, _18471_, _18467_);
  nand _69549_ (_18474_, _11089_, _09906_);
  and _69550_ (_18475_, _18474_, _01336_);
  and _69551_ (_18476_, _18475_, _18472_);
  or _69552_ (_18477_, _18476_, _18125_);
  and _69553_ (_43336_, _18477_, _42882_);
  nor _69554_ (_18478_, _01336_, _09906_);
  and _69555_ (_18479_, _10295_, _10259_);
  nor _69556_ (_18480_, _18479_, _10296_);
  or _69557_ (_18481_, _18480_, _10304_);
  and _69558_ (_18482_, _15195_, _07701_);
  nor _69559_ (_18484_, _07701_, _09906_);
  or _69560_ (_18485_, _18484_, _08751_);
  or _69561_ (_18486_, _18485_, _18482_);
  and _69562_ (_18487_, _10677_, _10899_);
  and _69563_ (_18488_, _08937_, \oc8051_golden_model_1.ACC [4]);
  nor _69564_ (_18489_, _18143_, _18488_);
  or _69565_ (_18490_, _10941_, _18489_);
  nand _69566_ (_18491_, _10941_, _18489_);
  and _69567_ (_18492_, _18491_, _18490_);
  or _69568_ (_18493_, _18492_, _10606_);
  nand _69569_ (_18495_, _18492_, _10606_);
  and _69570_ (_18496_, _18495_, _18493_);
  not _69571_ (_18497_, _18146_);
  or _69572_ (_18498_, _18149_, _18497_);
  nand _69573_ (_18499_, _18498_, _18496_);
  or _69574_ (_18500_, _18498_, _18496_);
  and _69575_ (_18501_, _18500_, _18499_);
  or _69576_ (_18502_, _18501_, _13935_);
  nand _69577_ (_18503_, _10378_, _07977_);
  or _69578_ (_18504_, _10390_, _09179_);
  nor _69579_ (_18506_, _10400_, _07977_);
  or _69580_ (_18507_, _06530_, \oc8051_golden_model_1.ACC [5]);
  nand _69581_ (_18508_, _06530_, \oc8051_golden_model_1.ACC [5]);
  and _69582_ (_18509_, _18508_, _18507_);
  and _69583_ (_18510_, _18509_, _10400_);
  or _69584_ (_18511_, _18510_, _10389_);
  or _69585_ (_18512_, _18511_, _18506_);
  and _69586_ (_18513_, _18512_, _10408_);
  and _69587_ (_18514_, _18513_, _18504_);
  and _69588_ (_18515_, _15093_, _07701_);
  or _69589_ (_18517_, _18515_, _18484_);
  and _69590_ (_18518_, _18517_, _06102_);
  or _69591_ (_18519_, _18518_, _10412_);
  or _69592_ (_18520_, _18519_, _18514_);
  nor _69593_ (_18521_, _10431_, _10424_);
  nand _69594_ (_18522_, _10431_, _10424_);
  nand _69595_ (_18523_, _18522_, _10412_);
  or _69596_ (_18524_, _18523_, _18521_);
  and _69597_ (_18525_, _18524_, _06244_);
  and _69598_ (_18526_, _18525_, _18520_);
  nor _69599_ (_18528_, _08359_, _09906_);
  and _69600_ (_18529_, _15073_, _08359_);
  or _69601_ (_18530_, _18529_, _18528_);
  and _69602_ (_18531_, _18530_, _06043_);
  nor _69603_ (_18532_, _07977_, _10439_);
  or _69604_ (_18533_, _18532_, _18484_);
  and _69605_ (_18534_, _18533_, _06239_);
  or _69606_ (_18535_, _18534_, _10378_);
  or _69607_ (_18536_, _18535_, _18531_);
  or _69608_ (_18537_, _18536_, _18526_);
  and _69609_ (_18539_, _18537_, _18503_);
  or _69610_ (_18540_, _18539_, _06970_);
  or _69611_ (_18541_, _09179_, _06971_);
  and _69612_ (_18542_, _18541_, _06220_);
  and _69613_ (_18543_, _18542_, _18540_);
  nor _69614_ (_18544_, _07979_, _06220_);
  or _69615_ (_18545_, _18544_, _10376_);
  or _69616_ (_18546_, _18545_, _18543_);
  nand _69617_ (_18547_, _10376_, _05784_);
  and _69618_ (_18548_, _18547_, _18546_);
  or _69619_ (_18550_, _18548_, _06039_);
  and _69620_ (_18551_, _15077_, _08359_);
  or _69621_ (_18552_, _18551_, _18528_);
  or _69622_ (_18553_, _18552_, _06040_);
  and _69623_ (_18554_, _18553_, _06033_);
  and _69624_ (_18555_, _18554_, _18550_);
  or _69625_ (_18556_, _18528_, _15110_);
  and _69626_ (_18557_, _18530_, _06032_);
  and _69627_ (_18558_, _18557_, _18556_);
  or _69628_ (_18559_, _18558_, _18555_);
  and _69629_ (_18561_, _18559_, _09800_);
  or _69630_ (_18562_, _09756_, _09754_);
  nor _69631_ (_18563_, _09757_, _09800_);
  and _69632_ (_18564_, _18563_, _18562_);
  or _69633_ (_18565_, _18564_, _10468_);
  or _69634_ (_18566_, _18565_, _18561_);
  and _69635_ (_18567_, _08270_, \oc8051_golden_model_1.ACC [4]);
  nor _69636_ (_18568_, _18219_, _18567_);
  and _69637_ (_18569_, _10900_, _18568_);
  nor _69638_ (_18570_, _10900_, _18568_);
  nor _69639_ (_18572_, _18570_, _18569_);
  nor _69640_ (_18573_, _18572_, _10606_);
  and _69641_ (_18574_, _18572_, _10606_);
  nor _69642_ (_18575_, _18574_, _18573_);
  nor _69643_ (_18576_, _18227_, _18223_);
  not _69644_ (_18577_, _18576_);
  and _69645_ (_18578_, _18577_, _18575_);
  nor _69646_ (_18579_, _18577_, _18575_);
  nor _69647_ (_18580_, _18579_, _18578_);
  or _69648_ (_18581_, _18580_, _10469_);
  and _69649_ (_18583_, _18581_, _18566_);
  or _69650_ (_18584_, _18583_, _12361_);
  and _69651_ (_18585_, _18584_, _06267_);
  and _69652_ (_18586_, _18585_, _18502_);
  and _69653_ (_18587_, _08272_, \oc8051_golden_model_1.ACC [4]);
  nor _69654_ (_18588_, _18238_, _18587_);
  nor _69655_ (_18589_, _12306_, _18588_);
  and _69656_ (_18590_, _12306_, _18588_);
  nor _69657_ (_18591_, _18590_, _18589_);
  and _69658_ (_18592_, _18591_, \oc8051_golden_model_1.PSW [7]);
  nor _69659_ (_18594_, _18591_, \oc8051_golden_model_1.PSW [7]);
  nor _69660_ (_18595_, _18594_, _18592_);
  nor _69661_ (_18596_, _18245_, _18241_);
  not _69662_ (_18597_, _18596_);
  or _69663_ (_18598_, _18597_, _18595_);
  and _69664_ (_18599_, _18597_, _18595_);
  nor _69665_ (_18600_, _18599_, _06267_);
  and _69666_ (_18601_, _18600_, _18598_);
  or _69667_ (_18602_, _18601_, _18586_);
  and _69668_ (_18603_, _18602_, _10307_);
  and _69669_ (_18605_, _06758_, \oc8051_golden_model_1.ACC [4]);
  nor _69670_ (_18606_, _18255_, _18605_);
  nor _69671_ (_18607_, _12325_, _18606_);
  and _69672_ (_18608_, _12325_, _18606_);
  nor _69673_ (_18609_, _18608_, _18607_);
  and _69674_ (_18610_, _18609_, \oc8051_golden_model_1.PSW [7]);
  nor _69675_ (_18611_, _18609_, \oc8051_golden_model_1.PSW [7]);
  nor _69676_ (_18612_, _18611_, _18610_);
  nor _69677_ (_18613_, _18262_, _18258_);
  not _69678_ (_18614_, _18613_);
  or _69679_ (_18616_, _18614_, _18612_);
  and _69680_ (_18617_, _18614_, _18612_);
  nor _69681_ (_18618_, _18617_, _10307_);
  and _69682_ (_18619_, _18618_, _18616_);
  or _69683_ (_18620_, _18619_, _05676_);
  or _69684_ (_18621_, _18620_, _18603_);
  nand _69685_ (_18622_, _06359_, _05676_);
  and _69686_ (_18623_, _18622_, _06027_);
  and _69687_ (_18624_, _18623_, _18621_);
  or _69688_ (_18625_, _18528_, _15074_);
  and _69689_ (_18627_, _18625_, _06026_);
  and _69690_ (_18628_, _18627_, _18530_);
  or _69691_ (_18629_, _18628_, _09818_);
  or _69692_ (_18630_, _18629_, _18624_);
  and _69693_ (_18631_, _09179_, _07701_);
  or _69694_ (_18632_, _18484_, _07012_);
  or _69695_ (_18633_, _18632_, _18631_);
  or _69696_ (_18634_, _18533_, _09827_);
  and _69697_ (_18635_, _18634_, _05669_);
  and _69698_ (_18636_, _18635_, _18633_);
  and _69699_ (_18638_, _18636_, _18630_);
  and _69700_ (_18639_, _15179_, _07701_);
  or _69701_ (_18640_, _18639_, _18484_);
  and _69702_ (_18641_, _18640_, _09833_);
  or _69703_ (_18642_, _18641_, _09832_);
  or _69704_ (_18643_, _18642_, _18638_);
  or _69705_ (_18644_, _09894_, _09839_);
  and _69706_ (_18645_, _18644_, _05664_);
  and _69707_ (_18646_, _18645_, _18643_);
  nor _69708_ (_18647_, _06359_, _05664_);
  or _69709_ (_18649_, _18647_, _06019_);
  or _69710_ (_18650_, _18649_, _18646_);
  and _69711_ (_18651_, _08652_, _07701_);
  or _69712_ (_18652_, _18651_, _18484_);
  or _69713_ (_18653_, _18652_, _06020_);
  and _69714_ (_18654_, _18653_, _10662_);
  and _69715_ (_18655_, _18654_, _18650_);
  nor _69716_ (_18656_, _10662_, _06359_);
  or _69717_ (_18657_, _18656_, _17656_);
  or _69718_ (_18658_, _18657_, _18655_);
  or _69719_ (_18659_, _10899_, _17660_);
  and _69720_ (_18660_, _18659_, _18658_);
  and _69721_ (_18661_, _18660_, _18305_);
  and _69722_ (_18662_, _10899_, _06649_);
  or _69723_ (_18663_, _18662_, _18310_);
  or _69724_ (_18664_, _18663_, _18661_);
  or _69725_ (_18665_, _10899_, _18316_);
  and _69726_ (_18666_, _18665_, _10678_);
  and _69727_ (_18667_, _18666_, _18664_);
  or _69728_ (_18668_, _18667_, _18487_);
  and _69729_ (_18671_, _18668_, _16972_);
  and _69730_ (_18672_, _16971_, _10899_);
  or _69731_ (_18673_, _18672_, _18671_);
  and _69732_ (_18674_, _18673_, _16970_);
  and _69733_ (_18675_, _10899_, _06650_);
  or _69734_ (_18676_, _18675_, _18674_);
  and _69735_ (_18677_, _18676_, _10686_);
  nor _69736_ (_18678_, _10686_, _10941_);
  or _69737_ (_18679_, _18678_, _06282_);
  or _69738_ (_18680_, _18679_, _18677_);
  or _69739_ (_18682_, _12306_, _06283_);
  and _69740_ (_18683_, _18682_, _10699_);
  and _69741_ (_18684_, _18683_, _18680_);
  and _69742_ (_18685_, _10698_, _12325_);
  or _69743_ (_18686_, _18685_, _06112_);
  or _69744_ (_18687_, _18686_, _18684_);
  and _69745_ (_18688_, _18687_, _18486_);
  or _69746_ (_18689_, _18688_, _06284_);
  or _69747_ (_18690_, _18484_, _08756_);
  and _69748_ (_18691_, _18690_, _11997_);
  and _69749_ (_18692_, _18691_, _18689_);
  or _69750_ (_18693_, _18345_, _10897_);
  and _69751_ (_18694_, _18693_, _17104_);
  or _69752_ (_18695_, _18694_, _18692_);
  or _69753_ (_18696_, _18009_, _10897_);
  and _69754_ (_18697_, _18696_, _18695_);
  or _69755_ (_18698_, _18697_, _10731_);
  or _69756_ (_18699_, _10736_, _10939_);
  and _69757_ (_18700_, _18699_, _10735_);
  and _69758_ (_18701_, _18700_, _18698_);
  or _69759_ (_18704_, _10741_, _10981_);
  and _69760_ (_18705_, _18704_, _10743_);
  or _69761_ (_18706_, _18705_, _18701_);
  or _69762_ (_18707_, _10747_, _11021_);
  and _69763_ (_18708_, _18707_, _07032_);
  and _69764_ (_18709_, _18708_, _18706_);
  nand _69765_ (_18710_, _18652_, _06108_);
  nor _69766_ (_18711_, _18710_, _10982_);
  or _69767_ (_18712_, _18711_, _10752_);
  or _69768_ (_18713_, _18712_, _18709_);
  and _69769_ (_18715_, _10898_, _10752_);
  nor _69770_ (_18716_, _18715_, _17203_);
  and _69771_ (_18717_, _18716_, _18713_);
  not _69772_ (_18718_, _10898_);
  nand _69773_ (_18719_, _18718_, _17203_);
  nor _69774_ (_18720_, _10765_, _06834_);
  nand _69775_ (_18721_, _18720_, _18719_);
  or _69776_ (_18722_, _18721_, _18717_);
  or _69777_ (_18723_, _18720_, _18718_);
  and _69778_ (_18724_, _18723_, _06668_);
  and _69779_ (_18725_, _18724_, _18722_);
  nor _69780_ (_18726_, _10898_, _06668_);
  or _69781_ (_18727_, _18726_, _10775_);
  or _69782_ (_18728_, _18727_, _18725_);
  nand _69783_ (_18729_, _10775_, _09906_);
  or _69784_ (_18730_, _18729_, _09179_);
  and _69785_ (_18731_, _18730_, _06291_);
  and _69786_ (_18732_, _18731_, _18728_);
  nand _69787_ (_18733_, _17136_, _10982_);
  and _69788_ (_18734_, _18733_, _11987_);
  or _69789_ (_18737_, _18734_, _18732_);
  nand _69790_ (_18738_, _10781_, _11022_);
  and _69791_ (_18739_, _18738_, _08777_);
  and _69792_ (_18740_, _18739_, _18737_);
  and _69793_ (_18741_, _15194_, _07701_);
  or _69794_ (_18742_, _18741_, _18484_);
  and _69795_ (_18743_, _18742_, _06130_);
  or _69796_ (_18744_, _18743_, _10303_);
  or _69797_ (_18745_, _18744_, _18740_);
  and _69798_ (_18746_, _18745_, _18481_);
  or _69799_ (_18748_, _18746_, _10794_);
  and _69800_ (_18749_, _10813_, _10518_);
  nor _69801_ (_18750_, _18749_, _10814_);
  or _69802_ (_18751_, _18750_, _10796_);
  and _69803_ (_18752_, _18751_, _06289_);
  and _69804_ (_18753_, _18752_, _18748_);
  and _69805_ (_18754_, _10843_, _10329_);
  nor _69806_ (_18755_, _18754_, _10844_);
  or _69807_ (_18756_, _18755_, _10824_);
  and _69808_ (_18757_, _18756_, _10826_);
  or _69809_ (_18758_, _18757_, _18753_);
  and _69810_ (_18759_, _10873_, _10589_);
  nor _69811_ (_18760_, _18759_, _10874_);
  or _69812_ (_18761_, _18760_, _10856_);
  and _69813_ (_18762_, _18761_, _10855_);
  and _69814_ (_18763_, _18762_, _18758_);
  and _69815_ (_18764_, _10854_, \oc8051_golden_model_1.ACC [4]);
  or _69816_ (_18765_, _18764_, _10887_);
  or _69817_ (_18766_, _18765_, _18763_);
  nor _69818_ (_18767_, _10885_, _06691_);
  not _69819_ (_18770_, _18767_);
  nor _69820_ (_18771_, _06136_, _06229_);
  nor _69821_ (_18772_, _18771_, _06841_);
  or _69822_ (_18773_, _18772_, _18770_);
  not _69823_ (_18774_, _18773_);
  and _69824_ (_18775_, _10922_, _10900_);
  nor _69825_ (_18776_, _18775_, _10923_);
  and _69826_ (_18777_, _18776_, _18774_);
  or _69827_ (_18778_, _18777_, _10890_);
  and _69828_ (_18779_, _18778_, _18766_);
  and _69829_ (_18781_, _18776_, _18773_);
  or _69830_ (_18782_, _18781_, _10932_);
  or _69831_ (_18783_, _18782_, _18779_);
  and _69832_ (_18784_, _10963_, _10941_);
  nor _69833_ (_18785_, _18784_, _10964_);
  or _69834_ (_18786_, _18785_, _10934_);
  and _69835_ (_18787_, _18786_, _06052_);
  and _69836_ (_18788_, _18787_, _18783_);
  and _69837_ (_18789_, _11004_, _12306_);
  nor _69838_ (_18790_, _11004_, _12306_);
  or _69839_ (_18791_, _18790_, _18789_);
  and _69840_ (_18792_, _18791_, _06051_);
  or _69841_ (_18793_, _18792_, _10974_);
  or _69842_ (_18794_, _18793_, _18788_);
  and _69843_ (_18795_, _11044_, _12325_);
  nor _69844_ (_18796_, _11044_, _12325_);
  or _69845_ (_18797_, _18796_, _11050_);
  or _69846_ (_18798_, _18797_, _18795_);
  and _69847_ (_18799_, _18798_, _11016_);
  and _69848_ (_18800_, _18799_, _18794_);
  and _69849_ (_18803_, _11015_, \oc8051_golden_model_1.ACC [4]);
  or _69850_ (_18804_, _18803_, _06316_);
  or _69851_ (_18805_, _18804_, _18800_);
  or _69852_ (_18806_, _18517_, _06718_);
  and _69853_ (_18807_, _18806_, _11060_);
  and _69854_ (_18808_, _18807_, _18805_);
  nor _69855_ (_18809_, _11067_, _09906_);
  or _69856_ (_18810_, _18809_, _11068_);
  nor _69857_ (_18811_, _18810_, _11064_);
  nor _69858_ (_18812_, _18811_, _12756_);
  or _69859_ (_18814_, _18812_, _18808_);
  nand _69860_ (_18815_, _11064_, _09861_);
  and _69861_ (_18816_, _18815_, _05653_);
  and _69862_ (_18817_, _18816_, _18814_);
  and _69863_ (_18818_, _18552_, _05652_);
  or _69864_ (_18819_, _18818_, _06047_);
  or _69865_ (_18820_, _18819_, _18817_);
  and _69866_ (_18821_, _15253_, _07701_);
  or _69867_ (_18822_, _18484_, _06048_);
  or _69868_ (_18823_, _18822_, _18821_);
  and _69869_ (_18824_, _18823_, _11083_);
  and _69870_ (_18825_, _18824_, _18820_);
  nor _69871_ (_18826_, _11093_, \oc8051_golden_model_1.ACC [5]);
  nor _69872_ (_18827_, _18826_, _11094_);
  and _69873_ (_18828_, _18827_, _11082_);
  or _69874_ (_18829_, _18828_, _11089_);
  or _69875_ (_18830_, _18829_, _18825_);
  nand _69876_ (_18831_, _11089_, _09861_);
  and _69877_ (_18832_, _18831_, _01336_);
  and _69878_ (_18833_, _18832_, _18830_);
  or _69879_ (_18836_, _18833_, _18478_);
  and _69880_ (_43338_, _18836_, _42882_);
  nor _69881_ (_18837_, _01336_, _09861_);
  nand _69882_ (_18838_, _11015_, _09906_);
  or _69883_ (_18839_, _11006_, _10980_);
  and _69884_ (_18840_, _18839_, _11007_);
  or _69885_ (_18841_, _18840_, _06052_);
  and _69886_ (_18842_, _18841_, _11050_);
  nor _69887_ (_18843_, _10845_, _10368_);
  nor _69888_ (_18844_, _18843_, _10846_);
  or _69889_ (_18846_, _18844_, _06289_);
  and _69890_ (_18847_, _18846_, _10856_);
  or _69891_ (_18848_, _10893_, _10722_);
  and _69892_ (_18849_, _15399_, _07701_);
  nor _69893_ (_18850_, _07701_, _09861_);
  or _69894_ (_18851_, _18850_, _08751_);
  or _69895_ (_18852_, _18851_, _18849_);
  and _69896_ (_18853_, _10669_, _10896_);
  and _69897_ (_18854_, _15382_, _07701_);
  or _69898_ (_18855_, _18854_, _18850_);
  and _69899_ (_18856_, _18855_, _09833_);
  or _69900_ (_18857_, _09179_, _09906_);
  and _69901_ (_18858_, _09179_, _09906_);
  or _69902_ (_18859_, _18489_, _18858_);
  and _69903_ (_18860_, _18859_, _18857_);
  nor _69904_ (_18861_, _18860_, _10938_);
  and _69905_ (_18862_, _18860_, _10938_);
  nor _69906_ (_18863_, _18862_, _18861_);
  and _69907_ (_18864_, _18499_, _18493_);
  and _69908_ (_18865_, _18864_, \oc8051_golden_model_1.PSW [7]);
  or _69909_ (_18868_, _18865_, _18863_);
  nand _69910_ (_18869_, _18865_, _18863_);
  and _69911_ (_18870_, _18869_, _12361_);
  and _69912_ (_18871_, _18870_, _18868_);
  nand _69913_ (_18872_, _10378_, _07883_);
  or _69914_ (_18873_, _10390_, _09178_);
  nor _69915_ (_18874_, _10400_, _07883_);
  nor _69916_ (_18875_, _06530_, _09861_);
  and _69917_ (_18876_, _06530_, _09861_);
  or _69918_ (_18877_, _18876_, _18875_);
  and _69919_ (_18879_, _18877_, _10400_);
  or _69920_ (_18880_, _18879_, _10389_);
  or _69921_ (_18881_, _18880_, _18874_);
  and _69922_ (_18882_, _18881_, _10408_);
  and _69923_ (_18883_, _18882_, _18873_);
  and _69924_ (_18884_, _15293_, _07701_);
  or _69925_ (_18885_, _18884_, _18850_);
  and _69926_ (_18886_, _18885_, _06102_);
  or _69927_ (_18887_, _18886_, _10412_);
  or _69928_ (_18888_, _18887_, _18883_);
  not _69929_ (_18890_, _10426_);
  and _69930_ (_18891_, _18521_, _18890_);
  or _69931_ (_18892_, _18521_, _18890_);
  nand _69932_ (_18893_, _18892_, _10412_);
  or _69933_ (_18894_, _18893_, _18891_);
  and _69934_ (_18895_, _18894_, _06244_);
  and _69935_ (_18896_, _18895_, _18888_);
  nor _69936_ (_18897_, _08359_, _09861_);
  and _69937_ (_18898_, _15280_, _08359_);
  or _69938_ (_18899_, _18898_, _18897_);
  and _69939_ (_18901_, _18899_, _06043_);
  nor _69940_ (_18902_, _07883_, _10439_);
  or _69941_ (_18903_, _18902_, _18850_);
  and _69942_ (_18904_, _18903_, _06239_);
  or _69943_ (_18905_, _18904_, _10378_);
  or _69944_ (_18906_, _18905_, _18901_);
  or _69945_ (_18907_, _18906_, _18896_);
  and _69946_ (_18908_, _18907_, _18872_);
  or _69947_ (_18909_, _18908_, _06970_);
  or _69948_ (_18910_, _09178_, _06971_);
  and _69949_ (_18912_, _18910_, _06220_);
  and _69950_ (_18913_, _18912_, _18909_);
  nor _69951_ (_18914_, _07885_, _06220_);
  or _69952_ (_18915_, _18914_, _10376_);
  or _69953_ (_18916_, _18915_, _18913_);
  nand _69954_ (_18917_, _10376_, _09956_);
  and _69955_ (_18918_, _18917_, _18916_);
  or _69956_ (_18919_, _18918_, _06039_);
  and _69957_ (_18920_, _15278_, _08359_);
  or _69958_ (_18921_, _18920_, _18897_);
  or _69959_ (_18923_, _18921_, _06040_);
  and _69960_ (_18924_, _18923_, _06033_);
  and _69961_ (_18925_, _18924_, _18919_);
  or _69962_ (_18926_, _18897_, _15310_);
  and _69963_ (_18927_, _18899_, _06032_);
  and _69964_ (_18928_, _18927_, _18926_);
  or _69965_ (_18929_, _18928_, _09269_);
  or _69966_ (_18930_, _18929_, _18925_);
  nor _69967_ (_18931_, _09759_, _09757_);
  nor _69968_ (_18932_, _18931_, _09760_);
  or _69969_ (_18934_, _18932_, _09800_);
  and _69970_ (_18935_, _18934_, _10469_);
  and _69971_ (_18936_, _18935_, _18930_);
  nand _69972_ (_18937_, _07977_, \oc8051_golden_model_1.ACC [5]);
  nor _69973_ (_18938_, _07977_, \oc8051_golden_model_1.ACC [5]);
  or _69974_ (_18939_, _18568_, _18938_);
  and _69975_ (_18940_, _18939_, _18937_);
  nor _69976_ (_18941_, _18940_, _10896_);
  and _69977_ (_18942_, _18940_, _10896_);
  nor _69978_ (_18943_, _18942_, _18941_);
  nor _69979_ (_18945_, _18578_, _18573_);
  and _69980_ (_18946_, _18945_, \oc8051_golden_model_1.PSW [7]);
  nand _69981_ (_18947_, _18946_, _18943_);
  or _69982_ (_18948_, _18946_, _18943_);
  and _69983_ (_18949_, _18948_, _10468_);
  and _69984_ (_18950_, _18949_, _18947_);
  or _69985_ (_18951_, _18950_, _18936_);
  and _69986_ (_18952_, _18951_, _13935_);
  or _69987_ (_18953_, _18952_, _06261_);
  or _69988_ (_18954_, _18953_, _18871_);
  or _69989_ (_18956_, _18588_, _13769_);
  and _69990_ (_18957_, _18956_, _13768_);
  nor _69991_ (_18958_, _18957_, _10980_);
  and _69992_ (_18959_, _18957_, _10980_);
  nor _69993_ (_18960_, _18959_, _18958_);
  nor _69994_ (_18961_, _18599_, _18592_);
  and _69995_ (_18962_, _18961_, \oc8051_golden_model_1.PSW [7]);
  not _69996_ (_18963_, _18962_);
  nor _69997_ (_18964_, _18963_, _18960_);
  and _69998_ (_18965_, _18963_, _18960_);
  or _69999_ (_18967_, _18965_, _18964_);
  or _70000_ (_18968_, _18967_, _06267_);
  and _70001_ (_18969_, _18968_, _10307_);
  and _70002_ (_18970_, _18969_, _18954_);
  or _70003_ (_18971_, _18606_, _13887_);
  and _70004_ (_18972_, _18971_, _13886_);
  nor _70005_ (_18973_, _18972_, _11020_);
  and _70006_ (_18974_, _18972_, _11020_);
  nor _70007_ (_18975_, _18974_, _18973_);
  nor _70008_ (_18976_, _18617_, _18610_);
  and _70009_ (_18978_, _18976_, \oc8051_golden_model_1.PSW [7]);
  or _70010_ (_18979_, _18978_, _18975_);
  nand _70011_ (_18980_, _18978_, _18975_);
  and _70012_ (_18981_, _18980_, _10306_);
  and _70013_ (_18982_, _18981_, _18979_);
  or _70014_ (_18983_, _18982_, _05676_);
  or _70015_ (_18984_, _18983_, _18970_);
  nand _70016_ (_18985_, _06084_, _05676_);
  and _70017_ (_18986_, _18985_, _06027_);
  and _70018_ (_18987_, _18986_, _18984_);
  or _70019_ (_18989_, _18897_, _15326_);
  and _70020_ (_18990_, _18989_, _06026_);
  and _70021_ (_18991_, _18990_, _18899_);
  or _70022_ (_18992_, _18991_, _09818_);
  or _70023_ (_18993_, _18992_, _18987_);
  and _70024_ (_18994_, _09178_, _07701_);
  or _70025_ (_18995_, _18850_, _07012_);
  or _70026_ (_18996_, _18995_, _18994_);
  or _70027_ (_18997_, _18903_, _09827_);
  and _70028_ (_18998_, _18997_, _05669_);
  and _70029_ (_19000_, _18998_, _18996_);
  and _70030_ (_19001_, _19000_, _18993_);
  or _70031_ (_19002_, _19001_, _18856_);
  and _70032_ (_19003_, _19002_, _12389_);
  nor _70033_ (_19004_, _06084_, _05664_);
  not _70034_ (_19005_, _09866_);
  nor _70035_ (_19006_, _19005_, _09862_);
  and _70036_ (_19007_, _19006_, _05662_);
  and _70037_ (_19008_, _19007_, _09832_);
  or _70038_ (_19009_, _19008_, _19004_);
  or _70039_ (_19011_, _19009_, _19003_);
  and _70040_ (_19012_, _19011_, _06020_);
  and _70041_ (_19013_, _15389_, _07701_);
  or _70042_ (_19014_, _19013_, _18850_);
  and _70043_ (_19015_, _19014_, _06019_);
  or _70044_ (_19016_, _19015_, _10661_);
  or _70045_ (_19017_, _19016_, _19012_);
  nand _70046_ (_19018_, _10661_, _06084_);
  and _70047_ (_19019_, _19018_, _10675_);
  and _70048_ (_19020_, _19019_, _19017_);
  or _70049_ (_19022_, _19020_, _18853_);
  and _70050_ (_19023_, _19022_, _18315_);
  and _70051_ (_19024_, _10896_, _18314_);
  or _70052_ (_19025_, _19024_, _19023_);
  and _70053_ (_19026_, _19025_, _17671_);
  and _70054_ (_19027_, _10896_, _17666_);
  or _70055_ (_19028_, _19027_, _19026_);
  and _70056_ (_19029_, _19028_, _17670_);
  and _70057_ (_19030_, _10896_, _17503_);
  or _70058_ (_19031_, _19030_, _19029_);
  and _70059_ (_19033_, _19031_, _16972_);
  and _70060_ (_19034_, _16971_, _10896_);
  or _70061_ (_19035_, _19034_, _19033_);
  and _70062_ (_19036_, _19035_, _16970_);
  and _70063_ (_19037_, _10896_, _06650_);
  or _70064_ (_19038_, _19037_, _19036_);
  and _70065_ (_19039_, _19038_, _10686_);
  and _70066_ (_19040_, _10685_, _10938_);
  or _70067_ (_19041_, _19040_, _06282_);
  or _70068_ (_19042_, _19041_, _19039_);
  or _70069_ (_19044_, _10980_, _06283_);
  and _70070_ (_19045_, _19044_, _10699_);
  and _70071_ (_19046_, _19045_, _19042_);
  and _70072_ (_19047_, _10698_, _11020_);
  or _70073_ (_19048_, _19047_, _06112_);
  or _70074_ (_19049_, _19048_, _19046_);
  and _70075_ (_19050_, _19049_, _18852_);
  or _70076_ (_19051_, _19050_, _06284_);
  or _70077_ (_19052_, _18850_, _08756_);
  and _70078_ (_19053_, _06093_, _05735_);
  not _70079_ (_19055_, _19053_);
  and _70080_ (_19056_, _19055_, _10725_);
  and _70081_ (_19057_, _19056_, _19052_);
  and _70082_ (_19058_, _19057_, _19051_);
  or _70083_ (_19059_, _10893_, _10721_);
  and _70084_ (_19060_, _19059_, _17104_);
  or _70085_ (_19061_, _19060_, _19058_);
  and _70086_ (_19062_, _19061_, _18848_);
  or _70087_ (_19063_, _19062_, _10731_);
  or _70088_ (_19064_, _10736_, _10935_);
  and _70089_ (_19066_, _19064_, _10735_);
  and _70090_ (_19067_, _19066_, _19063_);
  and _70091_ (_19068_, _10977_, _06279_);
  or _70092_ (_19069_, _19068_, _10741_);
  or _70093_ (_19070_, _19069_, _19067_);
  or _70094_ (_19071_, _10747_, _11017_);
  and _70095_ (_19072_, _19071_, _07032_);
  and _70096_ (_19073_, _19072_, _19070_);
  nand _70097_ (_19074_, _19014_, _06108_);
  nor _70098_ (_19075_, _19074_, _10979_);
  or _70099_ (_19077_, _19075_, _10752_);
  or _70100_ (_19078_, _19077_, _19073_);
  or _70101_ (_19079_, _10895_, _17205_);
  and _70102_ (_19080_, _19079_, _10760_);
  and _70103_ (_19081_, _19080_, _19078_);
  and _70104_ (_19082_, _10759_, _10895_);
  or _70105_ (_19083_, _19082_, _10767_);
  or _70106_ (_19084_, _19083_, _19081_);
  or _70107_ (_19085_, _10766_, _10895_);
  and _70108_ (_19086_, _19085_, _06668_);
  and _70109_ (_19088_, _19086_, _19084_);
  and _70110_ (_19089_, _10895_, _06667_);
  or _70111_ (_19090_, _19089_, _10775_);
  or _70112_ (_19091_, _19090_, _19088_);
  or _70113_ (_19092_, _17395_, _10936_);
  and _70114_ (_19093_, _19092_, _06291_);
  and _70115_ (_19094_, _19093_, _19091_);
  nor _70116_ (_19095_, _10979_, _06291_);
  or _70117_ (_19096_, _19095_, _10781_);
  or _70118_ (_19097_, _19096_, _19094_);
  nand _70119_ (_19099_, _10781_, _11019_);
  and _70120_ (_19100_, _19099_, _19097_);
  or _70121_ (_19101_, _19100_, _06130_);
  and _70122_ (_19102_, _15396_, _07701_);
  or _70123_ (_19103_, _18850_, _08777_);
  or _70124_ (_19104_, _19103_, _19102_);
  and _70125_ (_19105_, _19104_, _10304_);
  and _70126_ (_19106_, _19105_, _19101_);
  or _70127_ (_19107_, _10297_, _10253_);
  nor _70128_ (_19108_, _10304_, _10298_);
  and _70129_ (_19110_, _19108_, _19107_);
  or _70130_ (_19111_, _19110_, _17409_);
  or _70131_ (_19112_, _19111_, _19106_);
  or _70132_ (_19113_, _10815_, _10554_);
  and _70133_ (_19114_, _19113_, _10816_);
  or _70134_ (_19115_, _19114_, _17410_);
  and _70135_ (_19116_, _19115_, _17423_);
  and _70136_ (_19117_, _19116_, _19112_);
  nand _70137_ (_19118_, _19114_, _17416_);
  nand _70138_ (_19119_, _19118_, _06289_);
  or _70139_ (_19121_, _19119_, _19117_);
  and _70140_ (_19122_, _19121_, _18847_);
  or _70141_ (_19123_, _10875_, _10626_);
  and _70142_ (_19124_, _10876_, _10824_);
  and _70143_ (_19125_, _19124_, _19123_);
  or _70144_ (_19126_, _19125_, _10854_);
  or _70145_ (_19127_, _19126_, _19122_);
  nand _70146_ (_19128_, _10854_, _09906_);
  and _70147_ (_19129_, _19128_, _10890_);
  and _70148_ (_19130_, _19129_, _19127_);
  or _70149_ (_19132_, _10924_, _10896_);
  and _70150_ (_19133_, _19132_, _10925_);
  and _70151_ (_19134_, _19133_, _16956_);
  or _70152_ (_19135_, _19134_, _17437_);
  or _70153_ (_19136_, _19135_, _19130_);
  nor _70154_ (_19137_, _10965_, _10938_);
  nor _70155_ (_19138_, _19137_, _10966_);
  and _70156_ (_19139_, _19138_, _17443_);
  or _70157_ (_19140_, _19139_, _10934_);
  and _70158_ (_19141_, _19140_, _19136_);
  and _70159_ (_19143_, _19138_, _06692_);
  or _70160_ (_19144_, _19143_, _06051_);
  or _70161_ (_19145_, _19144_, _19141_);
  and _70162_ (_19146_, _19145_, _18842_);
  or _70163_ (_19147_, _11046_, _11020_);
  and _70164_ (_19148_, _11047_, _10974_);
  and _70165_ (_19149_, _19148_, _19147_);
  or _70166_ (_19150_, _19149_, _11015_);
  or _70167_ (_19151_, _19150_, _19146_);
  and _70168_ (_19152_, _19151_, _18838_);
  or _70169_ (_19154_, _19152_, _06316_);
  or _70170_ (_19155_, _18885_, _06718_);
  and _70171_ (_19156_, _19155_, _11060_);
  and _70172_ (_19157_, _19156_, _19154_);
  nor _70173_ (_19158_, _11068_, _09861_);
  or _70174_ (_19159_, _19158_, _11069_);
  and _70175_ (_19160_, _19159_, _11059_);
  or _70176_ (_19161_, _19160_, _11064_);
  or _70177_ (_19162_, _19161_, _19157_);
  nand _70178_ (_19163_, _11064_, _08393_);
  and _70179_ (_19165_, _19163_, _05653_);
  and _70180_ (_19166_, _19165_, _19162_);
  and _70181_ (_19167_, _18921_, _05652_);
  or _70182_ (_19168_, _19167_, _06047_);
  or _70183_ (_19169_, _19168_, _19166_);
  and _70184_ (_19170_, _15451_, _07701_);
  or _70185_ (_19171_, _18850_, _06048_);
  or _70186_ (_19172_, _19171_, _19170_);
  and _70187_ (_19173_, _19172_, _11083_);
  and _70188_ (_19174_, _19173_, _19169_);
  nor _70189_ (_19176_, _11094_, \oc8051_golden_model_1.ACC [6]);
  nor _70190_ (_19177_, _19176_, _11095_);
  and _70191_ (_19178_, _19177_, _11082_);
  or _70192_ (_19179_, _19178_, _11089_);
  or _70193_ (_19180_, _19179_, _19174_);
  nand _70194_ (_19181_, _11089_, _08393_);
  and _70195_ (_19182_, _19181_, _01336_);
  and _70196_ (_19183_, _19182_, _19180_);
  or _70197_ (_19184_, _19183_, _18837_);
  and _70198_ (_43339_, _19184_, _42882_);
  not _70199_ (_19186_, \oc8051_golden_model_1.PCON [0]);
  nor _70200_ (_19187_, _01336_, _19186_);
  nand _70201_ (_19188_, _10995_, _07641_);
  nor _70202_ (_19189_, _07641_, _19186_);
  nor _70203_ (_19190_, _19189_, _06278_);
  nand _70204_ (_19191_, _19190_, _19188_);
  and _70205_ (_19192_, _09120_, _07641_);
  or _70206_ (_19193_, _19189_, _07012_);
  or _70207_ (_19194_, _19193_, _19192_);
  and _70208_ (_19195_, _07641_, _06931_);
  nor _70209_ (_19197_, _19195_, _19189_);
  nand _70210_ (_19198_, _19197_, _09815_);
  nor _70211_ (_19199_, _08127_, _11109_);
  or _70212_ (_19200_, _19199_, _19189_);
  or _70213_ (_19201_, _19200_, _06954_);
  and _70214_ (_19202_, _07641_, \oc8051_golden_model_1.ACC [0]);
  nor _70215_ (_19203_, _19202_, _19189_);
  nor _70216_ (_19204_, _19203_, _06939_);
  nor _70217_ (_19205_, _06938_, _19186_);
  or _70218_ (_19206_, _19205_, _06102_);
  or _70219_ (_19208_, _19206_, _19204_);
  and _70220_ (_19209_, _19208_, _06848_);
  and _70221_ (_19210_, _19209_, _19201_);
  nor _70222_ (_19211_, _19197_, _06848_);
  or _70223_ (_19212_, _19211_, _19210_);
  nand _70224_ (_19213_, _19212_, _06220_);
  or _70225_ (_19214_, _19203_, _06220_);
  and _70226_ (_19215_, _19214_, _09817_);
  nand _70227_ (_19216_, _19215_, _19213_);
  and _70228_ (_19217_, _19216_, _19198_);
  and _70229_ (_19219_, _19217_, _19194_);
  or _70230_ (_19220_, _19219_, _09833_);
  and _70231_ (_19221_, _14186_, _07641_);
  or _70232_ (_19222_, _19221_, _19189_);
  or _70233_ (_19223_, _19222_, _05669_);
  and _70234_ (_19224_, _19223_, _06020_);
  and _70235_ (_19225_, _19224_, _19220_);
  and _70236_ (_19226_, _07641_, _08672_);
  or _70237_ (_19227_, _19226_, _19189_);
  and _70238_ (_19228_, _19227_, _06019_);
  or _70239_ (_19230_, _19228_, _06112_);
  or _70240_ (_19231_, _19230_, _19225_);
  and _70241_ (_19232_, _14086_, _07641_);
  or _70242_ (_19233_, _19189_, _08751_);
  or _70243_ (_19234_, _19233_, _19232_);
  and _70244_ (_19235_, _19234_, _08756_);
  and _70245_ (_19236_, _19235_, _19231_);
  nor _70246_ (_19237_, _12302_, _11109_);
  or _70247_ (_19238_, _19237_, _19189_);
  and _70248_ (_19239_, _19188_, _06284_);
  and _70249_ (_19241_, _19239_, _19238_);
  or _70250_ (_19242_, _19241_, _19236_);
  and _70251_ (_19243_, _19242_, _07032_);
  nand _70252_ (_19244_, _19227_, _06108_);
  nor _70253_ (_19245_, _19244_, _19199_);
  or _70254_ (_19246_, _19245_, _06277_);
  or _70255_ (_19247_, _19246_, _19243_);
  and _70256_ (_19248_, _19247_, _19191_);
  or _70257_ (_19249_, _19248_, _06130_);
  and _70258_ (_19250_, _14083_, _07641_);
  or _70259_ (_19252_, _19189_, _08777_);
  or _70260_ (_19253_, _19252_, _19250_);
  and _70261_ (_19254_, _19253_, _08782_);
  and _70262_ (_19255_, _19254_, _19249_);
  not _70263_ (_19256_, _06408_);
  and _70264_ (_19257_, _19238_, _06292_);
  or _70265_ (_19258_, _19257_, _19256_);
  or _70266_ (_19259_, _19258_, _19255_);
  or _70267_ (_19260_, _19200_, _06408_);
  and _70268_ (_19261_, _19260_, _01336_);
  and _70269_ (_19263_, _19261_, _19259_);
  or _70270_ (_19264_, _19263_, _19187_);
  and _70271_ (_43340_, _19264_, _42882_);
  not _70272_ (_19265_, \oc8051_golden_model_1.PCON [1]);
  nor _70273_ (_19266_, _01336_, _19265_);
  and _70274_ (_19267_, _09075_, _07641_);
  nor _70275_ (_19268_, _07641_, _19265_);
  or _70276_ (_19269_, _19268_, _07012_);
  or _70277_ (_19270_, _19269_, _19267_);
  or _70278_ (_19271_, _07641_, \oc8051_golden_model_1.PCON [1]);
  and _70279_ (_19273_, _14284_, _07641_);
  not _70280_ (_19274_, _19273_);
  and _70281_ (_19275_, _19274_, _19271_);
  or _70282_ (_19276_, _19275_, _06954_);
  and _70283_ (_19277_, _07641_, \oc8051_golden_model_1.ACC [1]);
  or _70284_ (_19278_, _19277_, _19268_);
  and _70285_ (_19279_, _19278_, _06938_);
  nor _70286_ (_19280_, _06938_, _19265_);
  or _70287_ (_19281_, _19280_, _06102_);
  or _70288_ (_19282_, _19281_, _19279_);
  and _70289_ (_19284_, _19282_, _06848_);
  and _70290_ (_19285_, _19284_, _19276_);
  nor _70291_ (_19286_, _11109_, _07132_);
  or _70292_ (_19287_, _19286_, _19268_);
  and _70293_ (_19288_, _19287_, _06239_);
  or _70294_ (_19289_, _19288_, _19285_);
  and _70295_ (_19290_, _19289_, _06220_);
  and _70296_ (_19291_, _19278_, _06219_);
  or _70297_ (_19292_, _19291_, _09818_);
  or _70298_ (_19293_, _19292_, _19290_);
  or _70299_ (_19295_, _19287_, _09827_);
  and _70300_ (_19296_, _19295_, _05669_);
  and _70301_ (_19297_, _19296_, _19293_);
  and _70302_ (_19298_, _19297_, _19270_);
  or _70303_ (_19299_, _14367_, _11109_);
  and _70304_ (_19300_, _19271_, _09833_);
  and _70305_ (_19301_, _19300_, _19299_);
  or _70306_ (_19302_, _19301_, _19298_);
  and _70307_ (_19303_, _19302_, _06020_);
  nand _70308_ (_19304_, _07641_, _06832_);
  and _70309_ (_19306_, _19271_, _06019_);
  and _70310_ (_19307_, _19306_, _19304_);
  or _70311_ (_19308_, _19307_, _19303_);
  and _70312_ (_19309_, _19308_, _08751_);
  or _70313_ (_19310_, _14263_, _11109_);
  and _70314_ (_19311_, _19271_, _06112_);
  and _70315_ (_19312_, _19311_, _19310_);
  or _70316_ (_19313_, _19312_, _06284_);
  or _70317_ (_19314_, _19313_, _19309_);
  and _70318_ (_19315_, _10994_, _07641_);
  or _70319_ (_19317_, _19315_, _19268_);
  or _70320_ (_19318_, _19317_, _08756_);
  and _70321_ (_19319_, _19318_, _07032_);
  and _70322_ (_19320_, _19319_, _19314_);
  or _70323_ (_19321_, _14261_, _11109_);
  and _70324_ (_19322_, _19271_, _06108_);
  and _70325_ (_19323_, _19322_, _19321_);
  or _70326_ (_19324_, _19323_, _06277_);
  or _70327_ (_19325_, _19324_, _19320_);
  and _70328_ (_19326_, _19277_, _08078_);
  or _70329_ (_19328_, _19268_, _06278_);
  or _70330_ (_19329_, _19328_, _19326_);
  and _70331_ (_19330_, _19329_, _08777_);
  and _70332_ (_19331_, _19330_, _19325_);
  or _70333_ (_19332_, _19304_, _08078_);
  and _70334_ (_19333_, _19271_, _06130_);
  and _70335_ (_19334_, _19333_, _19332_);
  or _70336_ (_19335_, _19334_, _06292_);
  or _70337_ (_19336_, _19335_, _19331_);
  nor _70338_ (_19337_, _10993_, _11109_);
  or _70339_ (_19339_, _19337_, _19268_);
  or _70340_ (_19340_, _19339_, _08782_);
  and _70341_ (_19341_, _19340_, _06718_);
  and _70342_ (_19342_, _19341_, _19336_);
  and _70343_ (_19343_, _19275_, _06316_);
  or _70344_ (_19344_, _19343_, _06047_);
  or _70345_ (_19345_, _19344_, _19342_);
  or _70346_ (_19346_, _19268_, _06048_);
  or _70347_ (_19347_, _19346_, _19273_);
  and _70348_ (_19348_, _19347_, _01336_);
  and _70349_ (_19350_, _19348_, _19345_);
  or _70350_ (_19351_, _19350_, _19266_);
  and _70351_ (_43342_, _19351_, _42882_);
  not _70352_ (_19352_, \oc8051_golden_model_1.PCON [2]);
  nor _70353_ (_19353_, _01336_, _19352_);
  and _70354_ (_19354_, _09182_, _07641_);
  nor _70355_ (_19355_, _07641_, _19352_);
  or _70356_ (_19356_, _19355_, _07012_);
  or _70357_ (_19357_, _19356_, _19354_);
  nor _70358_ (_19358_, _11109_, _07530_);
  nor _70359_ (_19360_, _19358_, _19355_);
  nand _70360_ (_19361_, _19360_, _09815_);
  and _70361_ (_19362_, _14493_, _07641_);
  or _70362_ (_19363_, _19362_, _19355_);
  or _70363_ (_19364_, _19363_, _06954_);
  and _70364_ (_19365_, _07641_, \oc8051_golden_model_1.ACC [2]);
  nor _70365_ (_19366_, _19365_, _19355_);
  nor _70366_ (_19367_, _19366_, _06939_);
  nor _70367_ (_19368_, _06938_, _19352_);
  or _70368_ (_19369_, _19368_, _06102_);
  or _70369_ (_19371_, _19369_, _19367_);
  and _70370_ (_19372_, _19371_, _06848_);
  and _70371_ (_19373_, _19372_, _19364_);
  nor _70372_ (_19374_, _19360_, _06848_);
  or _70373_ (_19375_, _19374_, _19373_);
  nand _70374_ (_19376_, _19375_, _06220_);
  or _70375_ (_19377_, _19366_, _06220_);
  and _70376_ (_19378_, _19377_, _09817_);
  nand _70377_ (_19379_, _19378_, _19376_);
  and _70378_ (_19380_, _19379_, _19361_);
  and _70379_ (_19382_, _19380_, _19357_);
  or _70380_ (_19383_, _19382_, _09833_);
  and _70381_ (_19384_, _14580_, _07641_);
  or _70382_ (_19385_, _19384_, _19355_);
  or _70383_ (_19386_, _19385_, _05669_);
  and _70384_ (_19387_, _19386_, _06020_);
  and _70385_ (_19388_, _19387_, _19383_);
  and _70386_ (_19389_, _07641_, _08730_);
  or _70387_ (_19390_, _19389_, _19355_);
  and _70388_ (_19391_, _19390_, _06019_);
  or _70389_ (_19393_, _19391_, _06112_);
  or _70390_ (_19394_, _19393_, _19388_);
  and _70391_ (_19395_, _14596_, _07641_);
  or _70392_ (_19396_, _19355_, _08751_);
  or _70393_ (_19397_, _19396_, _19395_);
  and _70394_ (_19398_, _19397_, _08756_);
  and _70395_ (_19399_, _19398_, _19394_);
  and _70396_ (_19400_, _10991_, _07641_);
  or _70397_ (_19401_, _19400_, _19355_);
  and _70398_ (_19402_, _19401_, _06284_);
  or _70399_ (_19404_, _19402_, _19399_);
  and _70400_ (_19405_, _19404_, _07032_);
  or _70401_ (_19406_, _19355_, _08177_);
  and _70402_ (_19407_, _19390_, _06108_);
  and _70403_ (_19408_, _19407_, _19406_);
  or _70404_ (_19409_, _19408_, _19405_);
  and _70405_ (_19410_, _19409_, _06278_);
  nor _70406_ (_19411_, _19366_, _06278_);
  and _70407_ (_19412_, _19411_, _19406_);
  or _70408_ (_19413_, _19412_, _06130_);
  or _70409_ (_19415_, _19413_, _19410_);
  and _70410_ (_19416_, _14593_, _07641_);
  or _70411_ (_19417_, _19355_, _08777_);
  or _70412_ (_19418_, _19417_, _19416_);
  and _70413_ (_19419_, _19418_, _08782_);
  and _70414_ (_19420_, _19419_, _19415_);
  nor _70415_ (_19421_, _10990_, _11109_);
  or _70416_ (_19422_, _19421_, _19355_);
  and _70417_ (_19423_, _19422_, _06292_);
  or _70418_ (_19424_, _19423_, _19420_);
  and _70419_ (_19426_, _19424_, _06718_);
  and _70420_ (_19427_, _19363_, _06316_);
  or _70421_ (_19428_, _19427_, _06047_);
  or _70422_ (_19429_, _19428_, _19426_);
  and _70423_ (_19430_, _14657_, _07641_);
  or _70424_ (_19431_, _19355_, _06048_);
  or _70425_ (_19432_, _19431_, _19430_);
  and _70426_ (_19433_, _19432_, _01336_);
  and _70427_ (_19434_, _19433_, _19429_);
  or _70428_ (_19435_, _19434_, _19353_);
  and _70429_ (_43343_, _19435_, _42882_);
  not _70430_ (_19437_, \oc8051_golden_model_1.PCON [3]);
  nor _70431_ (_19438_, _01336_, _19437_);
  nor _70432_ (_19439_, _07641_, _19437_);
  or _70433_ (_19440_, _19439_, _08029_);
  and _70434_ (_19441_, _07641_, _08662_);
  or _70435_ (_19442_, _19441_, _19439_);
  and _70436_ (_19443_, _19442_, _06108_);
  and _70437_ (_19444_, _19443_, _19440_);
  and _70438_ (_19445_, _09181_, _07641_);
  or _70439_ (_19447_, _19439_, _07012_);
  or _70440_ (_19448_, _19447_, _19445_);
  nor _70441_ (_19449_, _11109_, _07353_);
  nor _70442_ (_19450_, _19449_, _19439_);
  nand _70443_ (_19451_, _19450_, _09815_);
  and _70444_ (_19452_, _14672_, _07641_);
  or _70445_ (_19453_, _19452_, _19439_);
  or _70446_ (_19454_, _19453_, _06954_);
  and _70447_ (_19455_, _07641_, \oc8051_golden_model_1.ACC [3]);
  nor _70448_ (_19456_, _19455_, _19439_);
  nor _70449_ (_19458_, _19456_, _06939_);
  nor _70450_ (_19459_, _06938_, _19437_);
  or _70451_ (_19460_, _19459_, _06102_);
  or _70452_ (_19461_, _19460_, _19458_);
  and _70453_ (_19462_, _19461_, _06848_);
  and _70454_ (_19463_, _19462_, _19454_);
  nor _70455_ (_19464_, _19450_, _06848_);
  or _70456_ (_19465_, _19464_, _19463_);
  nand _70457_ (_19466_, _19465_, _06220_);
  or _70458_ (_19467_, _19456_, _06220_);
  and _70459_ (_19469_, _19467_, _09817_);
  nand _70460_ (_19470_, _19469_, _19466_);
  and _70461_ (_19471_, _19470_, _19451_);
  and _70462_ (_19472_, _19471_, _19448_);
  or _70463_ (_19473_, _19472_, _09833_);
  and _70464_ (_19474_, _14778_, _07641_);
  or _70465_ (_19475_, _19474_, _19439_);
  or _70466_ (_19476_, _19475_, _05669_);
  and _70467_ (_19477_, _19476_, _06020_);
  and _70468_ (_19478_, _19477_, _19473_);
  and _70469_ (_19480_, _19442_, _06019_);
  or _70470_ (_19481_, _19480_, _06112_);
  or _70471_ (_19482_, _19481_, _19478_);
  and _70472_ (_19483_, _14793_, _07641_);
  or _70473_ (_19484_, _19483_, _19439_);
  or _70474_ (_19485_, _19484_, _08751_);
  and _70475_ (_19486_, _19485_, _08756_);
  and _70476_ (_19487_, _19486_, _19482_);
  and _70477_ (_19488_, _12299_, _07641_);
  or _70478_ (_19489_, _19488_, _19439_);
  and _70479_ (_19491_, _19489_, _06284_);
  or _70480_ (_19492_, _19491_, _19487_);
  and _70481_ (_19493_, _19492_, _07032_);
  or _70482_ (_19494_, _19493_, _19444_);
  and _70483_ (_19495_, _19494_, _06278_);
  nor _70484_ (_19496_, _19456_, _06278_);
  and _70485_ (_19497_, _19496_, _19440_);
  or _70486_ (_19498_, _19497_, _06130_);
  or _70487_ (_19499_, _19498_, _19495_);
  and _70488_ (_19500_, _14792_, _07641_);
  or _70489_ (_19502_, _19439_, _08777_);
  or _70490_ (_19503_, _19502_, _19500_);
  and _70491_ (_19504_, _19503_, _08782_);
  and _70492_ (_19505_, _19504_, _19499_);
  nor _70493_ (_19506_, _10988_, _11109_);
  or _70494_ (_19507_, _19506_, _19439_);
  and _70495_ (_19508_, _19507_, _06292_);
  or _70496_ (_19509_, _19508_, _19505_);
  and _70497_ (_19510_, _19509_, _06718_);
  and _70498_ (_19511_, _19453_, _06316_);
  or _70499_ (_19513_, _19511_, _06047_);
  or _70500_ (_19514_, _19513_, _19510_);
  and _70501_ (_19515_, _14849_, _07641_);
  or _70502_ (_19516_, _19439_, _06048_);
  or _70503_ (_19517_, _19516_, _19515_);
  and _70504_ (_19518_, _19517_, _01336_);
  and _70505_ (_19519_, _19518_, _19514_);
  or _70506_ (_19520_, _19519_, _19438_);
  and _70507_ (_43344_, _19520_, _42882_);
  not _70508_ (_19521_, \oc8051_golden_model_1.PCON [4]);
  nor _70509_ (_19523_, _01336_, _19521_);
  nor _70510_ (_19524_, _07641_, _19521_);
  or _70511_ (_19525_, _19524_, _08273_);
  and _70512_ (_19526_, _08665_, _07641_);
  or _70513_ (_19527_, _19526_, _19524_);
  and _70514_ (_19528_, _19527_, _06108_);
  and _70515_ (_19529_, _19528_, _19525_);
  or _70516_ (_19530_, _19527_, _06020_);
  and _70517_ (_19531_, _14887_, _07641_);
  or _70518_ (_19532_, _19531_, _19524_);
  or _70519_ (_19534_, _19532_, _06954_);
  and _70520_ (_19535_, _07641_, \oc8051_golden_model_1.ACC [4]);
  or _70521_ (_19536_, _19535_, _19524_);
  and _70522_ (_19537_, _19536_, _06938_);
  nor _70523_ (_19538_, _06938_, _19521_);
  or _70524_ (_19539_, _19538_, _06102_);
  or _70525_ (_19540_, _19539_, _19537_);
  and _70526_ (_19541_, _19540_, _06848_);
  and _70527_ (_19542_, _19541_, _19534_);
  nor _70528_ (_19543_, _08270_, _11109_);
  or _70529_ (_19545_, _19543_, _19524_);
  and _70530_ (_19546_, _19545_, _06239_);
  or _70531_ (_19547_, _19546_, _19542_);
  and _70532_ (_19548_, _19547_, _06220_);
  and _70533_ (_19549_, _19536_, _06219_);
  or _70534_ (_19550_, _19549_, _09818_);
  or _70535_ (_19551_, _19550_, _19548_);
  and _70536_ (_19552_, _09180_, _07641_);
  or _70537_ (_19553_, _19524_, _07012_);
  or _70538_ (_19554_, _19553_, _19552_);
  or _70539_ (_19556_, _19545_, _09827_);
  and _70540_ (_19557_, _19556_, _05669_);
  and _70541_ (_19558_, _19557_, _19554_);
  and _70542_ (_19559_, _19558_, _19551_);
  and _70543_ (_19560_, _14983_, _07641_);
  or _70544_ (_19561_, _19560_, _19524_);
  and _70545_ (_19562_, _19561_, _09833_);
  or _70546_ (_19563_, _19562_, _06019_);
  or _70547_ (_19564_, _19563_, _19559_);
  and _70548_ (_19565_, _19564_, _19530_);
  or _70549_ (_19567_, _19565_, _06112_);
  and _70550_ (_19568_, _14876_, _07641_);
  or _70551_ (_19569_, _19524_, _08751_);
  or _70552_ (_19570_, _19569_, _19568_);
  and _70553_ (_19571_, _19570_, _08756_);
  and _70554_ (_19572_, _19571_, _19567_);
  and _70555_ (_19573_, _10986_, _07641_);
  or _70556_ (_19574_, _19573_, _19524_);
  and _70557_ (_19575_, _19574_, _06284_);
  or _70558_ (_19576_, _19575_, _19572_);
  and _70559_ (_19578_, _19576_, _07032_);
  or _70560_ (_19579_, _19578_, _19529_);
  and _70561_ (_19580_, _19579_, _06278_);
  and _70562_ (_19581_, _19536_, _06277_);
  and _70563_ (_19582_, _19581_, _19525_);
  or _70564_ (_19583_, _19582_, _06130_);
  or _70565_ (_19584_, _19583_, _19580_);
  and _70566_ (_19585_, _14873_, _07641_);
  or _70567_ (_19586_, _19524_, _08777_);
  or _70568_ (_19587_, _19586_, _19585_);
  and _70569_ (_19589_, _19587_, _08782_);
  and _70570_ (_19590_, _19589_, _19584_);
  nor _70571_ (_19591_, _10985_, _11109_);
  or _70572_ (_19592_, _19591_, _19524_);
  and _70573_ (_19593_, _19592_, _06292_);
  or _70574_ (_19594_, _19593_, _19590_);
  and _70575_ (_19595_, _19594_, _06718_);
  and _70576_ (_19596_, _19532_, _06316_);
  or _70577_ (_19597_, _19596_, _06047_);
  or _70578_ (_19598_, _19597_, _19595_);
  and _70579_ (_19600_, _15055_, _07641_);
  or _70580_ (_19601_, _19524_, _06048_);
  or _70581_ (_19602_, _19601_, _19600_);
  and _70582_ (_19603_, _19602_, _01336_);
  and _70583_ (_19604_, _19603_, _19598_);
  or _70584_ (_19605_, _19604_, _19523_);
  and _70585_ (_43345_, _19605_, _42882_);
  not _70586_ (_19606_, \oc8051_golden_model_1.PCON [5]);
  nor _70587_ (_19607_, _01336_, _19606_);
  nor _70588_ (_19608_, _07641_, _19606_);
  and _70589_ (_19610_, _08652_, _07641_);
  or _70590_ (_19611_, _19610_, _19608_);
  or _70591_ (_19612_, _19611_, _06020_);
  and _70592_ (_19613_, _15093_, _07641_);
  or _70593_ (_19614_, _19613_, _19608_);
  or _70594_ (_19615_, _19614_, _06954_);
  and _70595_ (_19616_, _07641_, \oc8051_golden_model_1.ACC [5]);
  or _70596_ (_19617_, _19616_, _19608_);
  and _70597_ (_19618_, _19617_, _06938_);
  nor _70598_ (_19619_, _06938_, _19606_);
  or _70599_ (_19621_, _19619_, _06102_);
  or _70600_ (_19622_, _19621_, _19618_);
  and _70601_ (_19623_, _19622_, _06848_);
  and _70602_ (_19624_, _19623_, _19615_);
  nor _70603_ (_19625_, _07977_, _11109_);
  or _70604_ (_19626_, _19625_, _19608_);
  and _70605_ (_19627_, _19626_, _06239_);
  or _70606_ (_19628_, _19627_, _19624_);
  and _70607_ (_19629_, _19628_, _06220_);
  and _70608_ (_19630_, _19617_, _06219_);
  or _70609_ (_19632_, _19630_, _09818_);
  or _70610_ (_19633_, _19632_, _19629_);
  and _70611_ (_19634_, _09179_, _07641_);
  or _70612_ (_19635_, _19608_, _07012_);
  or _70613_ (_19636_, _19635_, _19634_);
  or _70614_ (_19637_, _19626_, _09827_);
  and _70615_ (_19638_, _19637_, _05669_);
  and _70616_ (_19639_, _19638_, _19636_);
  and _70617_ (_19640_, _19639_, _19633_);
  and _70618_ (_19641_, _15179_, _07641_);
  or _70619_ (_19643_, _19641_, _19608_);
  and _70620_ (_19644_, _19643_, _09833_);
  or _70621_ (_19645_, _19644_, _06019_);
  or _70622_ (_19646_, _19645_, _19640_);
  and _70623_ (_19647_, _19646_, _19612_);
  or _70624_ (_19648_, _19647_, _06112_);
  and _70625_ (_19649_, _15195_, _07641_);
  or _70626_ (_19650_, _19649_, _19608_);
  or _70627_ (_19651_, _19650_, _08751_);
  and _70628_ (_19652_, _19651_, _08756_);
  and _70629_ (_19654_, _19652_, _19648_);
  and _70630_ (_19655_, _12306_, _07641_);
  or _70631_ (_19656_, _19655_, _19608_);
  and _70632_ (_19657_, _19656_, _06284_);
  or _70633_ (_19658_, _19657_, _19654_);
  and _70634_ (_19659_, _19658_, _07032_);
  or _70635_ (_19660_, _19608_, _07980_);
  and _70636_ (_19661_, _19611_, _06108_);
  and _70637_ (_19662_, _19661_, _19660_);
  or _70638_ (_19663_, _19662_, _19659_);
  and _70639_ (_19665_, _19663_, _06278_);
  and _70640_ (_19666_, _19617_, _06277_);
  and _70641_ (_19667_, _19666_, _19660_);
  or _70642_ (_19668_, _19667_, _06130_);
  or _70643_ (_19669_, _19668_, _19665_);
  and _70644_ (_19670_, _15194_, _07641_);
  or _70645_ (_19671_, _19608_, _08777_);
  or _70646_ (_19672_, _19671_, _19670_);
  and _70647_ (_19673_, _19672_, _08782_);
  and _70648_ (_19674_, _19673_, _19669_);
  nor _70649_ (_19676_, _10982_, _11109_);
  or _70650_ (_19677_, _19676_, _19608_);
  and _70651_ (_19678_, _19677_, _06292_);
  or _70652_ (_19679_, _19678_, _19674_);
  and _70653_ (_19680_, _19679_, _06718_);
  and _70654_ (_19681_, _19614_, _06316_);
  or _70655_ (_19682_, _19681_, _06047_);
  or _70656_ (_19683_, _19682_, _19680_);
  and _70657_ (_19684_, _15253_, _07641_);
  or _70658_ (_19685_, _19608_, _06048_);
  or _70659_ (_19687_, _19685_, _19684_);
  and _70660_ (_19688_, _19687_, _01336_);
  and _70661_ (_19689_, _19688_, _19683_);
  or _70662_ (_19690_, _19689_, _19607_);
  and _70663_ (_43346_, _19690_, _42882_);
  not _70664_ (_19691_, \oc8051_golden_model_1.PCON [6]);
  nor _70665_ (_19692_, _01336_, _19691_);
  nor _70666_ (_19693_, _07641_, _19691_);
  and _70667_ (_19694_, _15389_, _07641_);
  or _70668_ (_19695_, _19694_, _19693_);
  or _70669_ (_19697_, _19695_, _06020_);
  and _70670_ (_19698_, _15293_, _07641_);
  or _70671_ (_19699_, _19698_, _19693_);
  or _70672_ (_19700_, _19699_, _06954_);
  and _70673_ (_19701_, _07641_, \oc8051_golden_model_1.ACC [6]);
  or _70674_ (_19702_, _19701_, _19693_);
  and _70675_ (_19703_, _19702_, _06938_);
  nor _70676_ (_19704_, _06938_, _19691_);
  or _70677_ (_19705_, _19704_, _06102_);
  or _70678_ (_19706_, _19705_, _19703_);
  and _70679_ (_19708_, _19706_, _06848_);
  and _70680_ (_19709_, _19708_, _19700_);
  nor _70681_ (_19710_, _07883_, _11109_);
  or _70682_ (_19711_, _19710_, _19693_);
  and _70683_ (_19712_, _19711_, _06239_);
  or _70684_ (_19713_, _19712_, _19709_);
  and _70685_ (_19714_, _19713_, _06220_);
  and _70686_ (_19715_, _19702_, _06219_);
  or _70687_ (_19716_, _19715_, _09818_);
  or _70688_ (_19717_, _19716_, _19714_);
  and _70689_ (_19719_, _09178_, _07641_);
  or _70690_ (_19720_, _19693_, _07012_);
  or _70691_ (_19721_, _19720_, _19719_);
  or _70692_ (_19722_, _19711_, _09827_);
  and _70693_ (_19723_, _19722_, _05669_);
  and _70694_ (_19724_, _19723_, _19721_);
  and _70695_ (_19725_, _19724_, _19717_);
  and _70696_ (_19726_, _15382_, _07641_);
  or _70697_ (_19727_, _19726_, _19693_);
  and _70698_ (_19728_, _19727_, _09833_);
  or _70699_ (_19730_, _19728_, _06019_);
  or _70700_ (_19731_, _19730_, _19725_);
  and _70701_ (_19732_, _19731_, _19697_);
  or _70702_ (_19733_, _19732_, _06112_);
  and _70703_ (_19734_, _15399_, _07641_);
  or _70704_ (_19735_, _19734_, _19693_);
  or _70705_ (_19736_, _19735_, _08751_);
  and _70706_ (_19737_, _19736_, _08756_);
  and _70707_ (_19738_, _19737_, _19733_);
  and _70708_ (_19739_, _10980_, _07641_);
  or _70709_ (_19741_, _19739_, _19693_);
  and _70710_ (_19742_, _19741_, _06284_);
  or _70711_ (_19743_, _19742_, _19738_);
  and _70712_ (_19744_, _19743_, _07032_);
  or _70713_ (_19745_, _19693_, _07886_);
  and _70714_ (_19746_, _19695_, _06108_);
  and _70715_ (_19747_, _19746_, _19745_);
  or _70716_ (_19748_, _19747_, _19744_);
  and _70717_ (_19749_, _19748_, _06278_);
  and _70718_ (_19750_, _19702_, _06277_);
  and _70719_ (_19752_, _19750_, _19745_);
  or _70720_ (_19753_, _19752_, _06130_);
  or _70721_ (_19754_, _19753_, _19749_);
  and _70722_ (_19755_, _15396_, _07641_);
  or _70723_ (_19756_, _19693_, _08777_);
  or _70724_ (_19757_, _19756_, _19755_);
  and _70725_ (_19758_, _19757_, _08782_);
  and _70726_ (_19759_, _19758_, _19754_);
  nor _70727_ (_19760_, _10979_, _11109_);
  or _70728_ (_19761_, _19760_, _19693_);
  and _70729_ (_19763_, _19761_, _06292_);
  or _70730_ (_19764_, _19763_, _19759_);
  and _70731_ (_19765_, _19764_, _06718_);
  and _70732_ (_19766_, _19699_, _06316_);
  or _70733_ (_19767_, _19766_, _06047_);
  or _70734_ (_19768_, _19767_, _19765_);
  and _70735_ (_19769_, _15451_, _07641_);
  or _70736_ (_19770_, _19693_, _06048_);
  or _70737_ (_19771_, _19770_, _19769_);
  and _70738_ (_19772_, _19771_, _01336_);
  and _70739_ (_19774_, _19772_, _19768_);
  or _70740_ (_19775_, _19774_, _19692_);
  and _70741_ (_43347_, _19775_, _42882_);
  not _70742_ (_19776_, \oc8051_golden_model_1.TMOD [0]);
  nor _70743_ (_19777_, _01336_, _19776_);
  nand _70744_ (_19778_, _10995_, _07653_);
  nor _70745_ (_19779_, _07653_, _19776_);
  nor _70746_ (_19780_, _19779_, _06278_);
  nand _70747_ (_19781_, _19780_, _19778_);
  and _70748_ (_19782_, _09120_, _07653_);
  or _70749_ (_19784_, _19779_, _07012_);
  or _70750_ (_19785_, _19784_, _19782_);
  and _70751_ (_19786_, _07653_, _06931_);
  nor _70752_ (_19787_, _19786_, _19779_);
  nand _70753_ (_19788_, _19787_, _09815_);
  nor _70754_ (_19789_, _08127_, _11185_);
  or _70755_ (_19790_, _19789_, _19779_);
  or _70756_ (_19791_, _19790_, _06954_);
  and _70757_ (_19792_, _07653_, \oc8051_golden_model_1.ACC [0]);
  nor _70758_ (_19793_, _19792_, _19779_);
  nor _70759_ (_19795_, _19793_, _06939_);
  nor _70760_ (_19796_, _06938_, _19776_);
  or _70761_ (_19797_, _19796_, _06102_);
  or _70762_ (_19798_, _19797_, _19795_);
  and _70763_ (_19799_, _19798_, _06848_);
  and _70764_ (_19800_, _19799_, _19791_);
  nor _70765_ (_19801_, _19787_, _06848_);
  or _70766_ (_19802_, _19801_, _19800_);
  nand _70767_ (_19803_, _19802_, _06220_);
  or _70768_ (_19804_, _19793_, _06220_);
  and _70769_ (_19806_, _19804_, _09817_);
  nand _70770_ (_19807_, _19806_, _19803_);
  and _70771_ (_19808_, _19807_, _19788_);
  and _70772_ (_19809_, _19808_, _19785_);
  or _70773_ (_19810_, _19809_, _09833_);
  and _70774_ (_19811_, _14186_, _07653_);
  or _70775_ (_19812_, _19811_, _19779_);
  or _70776_ (_19813_, _19812_, _05669_);
  and _70777_ (_19814_, _19813_, _06020_);
  and _70778_ (_19815_, _19814_, _19810_);
  and _70779_ (_19817_, _07653_, _08672_);
  or _70780_ (_19818_, _19817_, _19779_);
  and _70781_ (_19819_, _19818_, _06019_);
  or _70782_ (_19820_, _19819_, _06112_);
  or _70783_ (_19821_, _19820_, _19815_);
  and _70784_ (_19822_, _14086_, _07653_);
  or _70785_ (_19823_, _19779_, _08751_);
  or _70786_ (_19824_, _19823_, _19822_);
  and _70787_ (_19825_, _19824_, _08756_);
  and _70788_ (_19826_, _19825_, _19821_);
  nor _70789_ (_19828_, _12302_, _11185_);
  or _70790_ (_19829_, _19828_, _19779_);
  and _70791_ (_19830_, _19778_, _06284_);
  and _70792_ (_19831_, _19830_, _19829_);
  or _70793_ (_19832_, _19831_, _19826_);
  and _70794_ (_19833_, _19832_, _07032_);
  nand _70795_ (_19834_, _19818_, _06108_);
  nor _70796_ (_19835_, _19834_, _19789_);
  or _70797_ (_19836_, _19835_, _06277_);
  or _70798_ (_19837_, _19836_, _19833_);
  and _70799_ (_19839_, _19837_, _19781_);
  or _70800_ (_19840_, _19839_, _06130_);
  and _70801_ (_19841_, _14083_, _07653_);
  or _70802_ (_19842_, _19779_, _08777_);
  or _70803_ (_19843_, _19842_, _19841_);
  and _70804_ (_19844_, _19843_, _08782_);
  and _70805_ (_19845_, _19844_, _19840_);
  and _70806_ (_19846_, _19829_, _06292_);
  or _70807_ (_19847_, _19846_, _19256_);
  or _70808_ (_19848_, _19847_, _19845_);
  or _70809_ (_19850_, _19790_, _06408_);
  and _70810_ (_19851_, _19850_, _01336_);
  and _70811_ (_19852_, _19851_, _19848_);
  or _70812_ (_19853_, _19852_, _19777_);
  and _70813_ (_43349_, _19853_, _42882_);
  and _70814_ (_19854_, _01340_, \oc8051_golden_model_1.TMOD [1]);
  or _70815_ (_19855_, _14367_, _11185_);
  or _70816_ (_19856_, _07653_, \oc8051_golden_model_1.TMOD [1]);
  and _70817_ (_19857_, _19856_, _09833_);
  and _70818_ (_19858_, _19857_, _19855_);
  and _70819_ (_19861_, _09075_, _07653_);
  and _70820_ (_19862_, _11185_, \oc8051_golden_model_1.TMOD [1]);
  or _70821_ (_19863_, _19862_, _07012_);
  or _70822_ (_19864_, _19863_, _19861_);
  and _70823_ (_19865_, _14284_, _07653_);
  not _70824_ (_19866_, _19865_);
  and _70825_ (_19867_, _19866_, _19856_);
  or _70826_ (_19868_, _19867_, _06954_);
  and _70827_ (_19869_, _07653_, \oc8051_golden_model_1.ACC [1]);
  or _70828_ (_19870_, _19869_, _19862_);
  and _70829_ (_19873_, _19870_, _06938_);
  and _70830_ (_19874_, _06939_, \oc8051_golden_model_1.TMOD [1]);
  or _70831_ (_19875_, _19874_, _06102_);
  or _70832_ (_19876_, _19875_, _19873_);
  and _70833_ (_19877_, _19876_, _06848_);
  and _70834_ (_19878_, _19877_, _19868_);
  nor _70835_ (_19879_, _11185_, _07132_);
  or _70836_ (_19880_, _19879_, _19862_);
  and _70837_ (_19881_, _19880_, _06239_);
  or _70838_ (_19882_, _19881_, _19878_);
  and _70839_ (_19885_, _19882_, _06220_);
  and _70840_ (_19886_, _19870_, _06219_);
  or _70841_ (_19887_, _19886_, _09818_);
  or _70842_ (_19888_, _19887_, _19885_);
  or _70843_ (_19889_, _19880_, _09827_);
  and _70844_ (_19890_, _19889_, _05669_);
  and _70845_ (_19891_, _19890_, _19888_);
  and _70846_ (_19892_, _19891_, _19864_);
  or _70847_ (_19893_, _19892_, _19858_);
  and _70848_ (_19894_, _19893_, _06020_);
  nand _70849_ (_19897_, _07653_, _06832_);
  and _70850_ (_19898_, _19856_, _06019_);
  and _70851_ (_19899_, _19898_, _19897_);
  or _70852_ (_19900_, _19899_, _19894_);
  and _70853_ (_19901_, _19900_, _08751_);
  or _70854_ (_19902_, _14263_, _11185_);
  and _70855_ (_19903_, _19856_, _06112_);
  and _70856_ (_19904_, _19903_, _19902_);
  or _70857_ (_19905_, _19904_, _06284_);
  or _70858_ (_19906_, _19905_, _19901_);
  and _70859_ (_19909_, _10994_, _07653_);
  or _70860_ (_19910_, _19909_, _19862_);
  or _70861_ (_19911_, _19910_, _08756_);
  and _70862_ (_19912_, _19911_, _07032_);
  and _70863_ (_19913_, _19912_, _19906_);
  or _70864_ (_19914_, _14261_, _11185_);
  and _70865_ (_19915_, _19856_, _06108_);
  and _70866_ (_19916_, _19915_, _19914_);
  or _70867_ (_19917_, _19916_, _06277_);
  or _70868_ (_19918_, _19917_, _19913_);
  and _70869_ (_19921_, _19869_, _08078_);
  or _70870_ (_19922_, _19862_, _06278_);
  or _70871_ (_19923_, _19922_, _19921_);
  and _70872_ (_19924_, _19923_, _08777_);
  and _70873_ (_19925_, _19924_, _19918_);
  or _70874_ (_19926_, _19897_, _08078_);
  and _70875_ (_19927_, _19856_, _06130_);
  and _70876_ (_19928_, _19927_, _19926_);
  or _70877_ (_19929_, _19928_, _06292_);
  or _70878_ (_19930_, _19929_, _19925_);
  nor _70879_ (_19933_, _10993_, _11185_);
  or _70880_ (_19934_, _19933_, _19862_);
  or _70881_ (_19935_, _19934_, _08782_);
  and _70882_ (_19936_, _19935_, _06718_);
  and _70883_ (_19937_, _19936_, _19930_);
  and _70884_ (_19938_, _19867_, _06316_);
  or _70885_ (_19939_, _19938_, _06047_);
  or _70886_ (_19940_, _19939_, _19937_);
  or _70887_ (_19941_, _19862_, _06048_);
  or _70888_ (_19942_, _19941_, _19865_);
  and _70889_ (_19944_, _19942_, _01336_);
  and _70890_ (_19945_, _19944_, _19940_);
  or _70891_ (_19946_, _19945_, _19854_);
  and _70892_ (_43350_, _19946_, _42882_);
  not _70893_ (_19947_, \oc8051_golden_model_1.TMOD [2]);
  nor _70894_ (_19948_, _01336_, _19947_);
  nor _70895_ (_19949_, _07653_, _19947_);
  or _70896_ (_19950_, _19949_, _08177_);
  and _70897_ (_19951_, _07653_, _08730_);
  or _70898_ (_19952_, _19951_, _19949_);
  and _70899_ (_19954_, _19952_, _06108_);
  and _70900_ (_19955_, _19954_, _19950_);
  and _70901_ (_19956_, _09182_, _07653_);
  or _70902_ (_19957_, _19949_, _07012_);
  or _70903_ (_19958_, _19957_, _19956_);
  nor _70904_ (_19959_, _11185_, _07530_);
  nor _70905_ (_19960_, _19959_, _19949_);
  nand _70906_ (_19961_, _19960_, _09815_);
  and _70907_ (_19962_, _14493_, _07653_);
  or _70908_ (_19963_, _19962_, _19949_);
  or _70909_ (_19965_, _19963_, _06954_);
  and _70910_ (_19966_, _07653_, \oc8051_golden_model_1.ACC [2]);
  nor _70911_ (_19967_, _19966_, _19949_);
  nor _70912_ (_19968_, _19967_, _06939_);
  nor _70913_ (_19969_, _06938_, _19947_);
  or _70914_ (_19970_, _19969_, _06102_);
  or _70915_ (_19971_, _19970_, _19968_);
  and _70916_ (_19972_, _19971_, _06848_);
  and _70917_ (_19973_, _19972_, _19965_);
  nor _70918_ (_19974_, _19960_, _06848_);
  or _70919_ (_19976_, _19974_, _19973_);
  nand _70920_ (_19977_, _19976_, _06220_);
  or _70921_ (_19978_, _19967_, _06220_);
  and _70922_ (_19979_, _19978_, _09817_);
  nand _70923_ (_19980_, _19979_, _19977_);
  and _70924_ (_19981_, _19980_, _19961_);
  and _70925_ (_19982_, _19981_, _19958_);
  or _70926_ (_19983_, _19982_, _09833_);
  and _70927_ (_19984_, _14580_, _07653_);
  or _70928_ (_19985_, _19984_, _19949_);
  or _70929_ (_19987_, _19985_, _05669_);
  and _70930_ (_19988_, _19987_, _06020_);
  and _70931_ (_19989_, _19988_, _19983_);
  and _70932_ (_19990_, _19952_, _06019_);
  or _70933_ (_19991_, _19990_, _06112_);
  or _70934_ (_19992_, _19991_, _19989_);
  and _70935_ (_19993_, _14596_, _07653_);
  or _70936_ (_19994_, _19993_, _19949_);
  or _70937_ (_19995_, _19994_, _08751_);
  and _70938_ (_19996_, _19995_, _08756_);
  and _70939_ (_19998_, _19996_, _19992_);
  and _70940_ (_19999_, _10991_, _07653_);
  or _70941_ (_20000_, _19999_, _19949_);
  and _70942_ (_20001_, _20000_, _06284_);
  or _70943_ (_20002_, _20001_, _19998_);
  and _70944_ (_20003_, _20002_, _07032_);
  or _70945_ (_20004_, _20003_, _19955_);
  and _70946_ (_20005_, _20004_, _06278_);
  nor _70947_ (_20006_, _19967_, _06278_);
  and _70948_ (_20007_, _20006_, _19950_);
  or _70949_ (_20009_, _20007_, _06130_);
  or _70950_ (_20010_, _20009_, _20005_);
  and _70951_ (_20011_, _14593_, _07653_);
  or _70952_ (_20012_, _19949_, _08777_);
  or _70953_ (_20013_, _20012_, _20011_);
  and _70954_ (_20014_, _20013_, _08782_);
  and _70955_ (_20015_, _20014_, _20010_);
  nor _70956_ (_20016_, _10990_, _11185_);
  or _70957_ (_20017_, _20016_, _19949_);
  and _70958_ (_20018_, _20017_, _06292_);
  or _70959_ (_20020_, _20018_, _20015_);
  and _70960_ (_20021_, _20020_, _06718_);
  and _70961_ (_20022_, _19963_, _06316_);
  or _70962_ (_20023_, _20022_, _06047_);
  or _70963_ (_20024_, _20023_, _20021_);
  and _70964_ (_20025_, _14657_, _07653_);
  or _70965_ (_20026_, _19949_, _06048_);
  or _70966_ (_20027_, _20026_, _20025_);
  and _70967_ (_20028_, _20027_, _01336_);
  and _70968_ (_20029_, _20028_, _20024_);
  or _70969_ (_20031_, _20029_, _19948_);
  and _70970_ (_43351_, _20031_, _42882_);
  and _70971_ (_20032_, _01340_, \oc8051_golden_model_1.TMOD [3]);
  and _70972_ (_20033_, _11185_, \oc8051_golden_model_1.TMOD [3]);
  or _70973_ (_20034_, _20033_, _08029_);
  and _70974_ (_20035_, _07653_, _08662_);
  or _70975_ (_20036_, _20035_, _20033_);
  and _70976_ (_20037_, _20036_, _06108_);
  and _70977_ (_20038_, _20037_, _20034_);
  or _70978_ (_20039_, _20036_, _06020_);
  and _70979_ (_20041_, _09181_, _07653_);
  or _70980_ (_20042_, _20033_, _07012_);
  or _70981_ (_20043_, _20042_, _20041_);
  and _70982_ (_20044_, _14672_, _07653_);
  or _70983_ (_20045_, _20044_, _20033_);
  or _70984_ (_20046_, _20045_, _06954_);
  and _70985_ (_20047_, _07653_, \oc8051_golden_model_1.ACC [3]);
  or _70986_ (_20048_, _20047_, _20033_);
  and _70987_ (_20049_, _20048_, _06938_);
  and _70988_ (_20050_, _06939_, \oc8051_golden_model_1.TMOD [3]);
  or _70989_ (_20052_, _20050_, _06102_);
  or _70990_ (_20053_, _20052_, _20049_);
  and _70991_ (_20054_, _20053_, _06848_);
  and _70992_ (_20055_, _20054_, _20046_);
  nor _70993_ (_20056_, _11185_, _07353_);
  or _70994_ (_20057_, _20056_, _20033_);
  and _70995_ (_20058_, _20057_, _06239_);
  or _70996_ (_20059_, _20058_, _20055_);
  and _70997_ (_20060_, _20059_, _06220_);
  and _70998_ (_20061_, _20048_, _06219_);
  or _70999_ (_20063_, _20061_, _09818_);
  or _71000_ (_20064_, _20063_, _20060_);
  or _71001_ (_20065_, _20057_, _09827_);
  and _71002_ (_20066_, _20065_, _05669_);
  and _71003_ (_20067_, _20066_, _20064_);
  and _71004_ (_20068_, _20067_, _20043_);
  and _71005_ (_20069_, _14778_, _07653_);
  or _71006_ (_20070_, _20069_, _20033_);
  and _71007_ (_20071_, _20070_, _09833_);
  or _71008_ (_20072_, _20071_, _06019_);
  or _71009_ (_20074_, _20072_, _20068_);
  and _71010_ (_20075_, _20074_, _20039_);
  or _71011_ (_20076_, _20075_, _06112_);
  and _71012_ (_20077_, _14793_, _07653_);
  or _71013_ (_20078_, _20033_, _08751_);
  or _71014_ (_20079_, _20078_, _20077_);
  and _71015_ (_20080_, _20079_, _08756_);
  and _71016_ (_20081_, _20080_, _20076_);
  and _71017_ (_20082_, _12299_, _07653_);
  or _71018_ (_20083_, _20082_, _20033_);
  and _71019_ (_20085_, _20083_, _06284_);
  or _71020_ (_20086_, _20085_, _20081_);
  and _71021_ (_20087_, _20086_, _07032_);
  or _71022_ (_20088_, _20087_, _20038_);
  and _71023_ (_20089_, _20088_, _06278_);
  and _71024_ (_20090_, _20048_, _06277_);
  and _71025_ (_20091_, _20090_, _20034_);
  or _71026_ (_20092_, _20091_, _06130_);
  or _71027_ (_20093_, _20092_, _20089_);
  and _71028_ (_20094_, _14792_, _07653_);
  or _71029_ (_20096_, _20033_, _08777_);
  or _71030_ (_20097_, _20096_, _20094_);
  and _71031_ (_20098_, _20097_, _08782_);
  and _71032_ (_20099_, _20098_, _20093_);
  nor _71033_ (_20100_, _10988_, _11185_);
  or _71034_ (_20101_, _20100_, _20033_);
  and _71035_ (_20102_, _20101_, _06292_);
  or _71036_ (_20103_, _20102_, _20099_);
  and _71037_ (_20104_, _20103_, _06718_);
  and _71038_ (_20105_, _20045_, _06316_);
  or _71039_ (_20107_, _20105_, _06047_);
  or _71040_ (_20108_, _20107_, _20104_);
  and _71041_ (_20109_, _14849_, _07653_);
  or _71042_ (_20110_, _20033_, _06048_);
  or _71043_ (_20111_, _20110_, _20109_);
  and _71044_ (_20112_, _20111_, _01336_);
  and _71045_ (_20113_, _20112_, _20108_);
  or _71046_ (_20114_, _20113_, _20032_);
  and _71047_ (_43352_, _20114_, _42882_);
  and _71048_ (_20115_, _01340_, \oc8051_golden_model_1.TMOD [4]);
  and _71049_ (_20117_, _11185_, \oc8051_golden_model_1.TMOD [4]);
  and _71050_ (_20118_, _08665_, _07653_);
  or _71051_ (_20119_, _20118_, _20117_);
  or _71052_ (_20120_, _20119_, _06020_);
  and _71053_ (_20121_, _14887_, _07653_);
  or _71054_ (_20122_, _20121_, _20117_);
  or _71055_ (_20123_, _20122_, _06954_);
  and _71056_ (_20124_, _07653_, \oc8051_golden_model_1.ACC [4]);
  or _71057_ (_20125_, _20124_, _20117_);
  and _71058_ (_20126_, _20125_, _06938_);
  and _71059_ (_20128_, _06939_, \oc8051_golden_model_1.TMOD [4]);
  or _71060_ (_20129_, _20128_, _06102_);
  or _71061_ (_20130_, _20129_, _20126_);
  and _71062_ (_20131_, _20130_, _06848_);
  and _71063_ (_20132_, _20131_, _20123_);
  nor _71064_ (_20133_, _08270_, _11185_);
  or _71065_ (_20134_, _20133_, _20117_);
  and _71066_ (_20135_, _20134_, _06239_);
  or _71067_ (_20136_, _20135_, _20132_);
  and _71068_ (_20137_, _20136_, _06220_);
  and _71069_ (_20139_, _20125_, _06219_);
  or _71070_ (_20140_, _20139_, _09818_);
  or _71071_ (_20141_, _20140_, _20137_);
  and _71072_ (_20142_, _09180_, _07653_);
  or _71073_ (_20143_, _20117_, _07012_);
  or _71074_ (_20144_, _20143_, _20142_);
  or _71075_ (_20145_, _20134_, _09827_);
  and _71076_ (_20146_, _20145_, _05669_);
  and _71077_ (_20147_, _20146_, _20144_);
  and _71078_ (_20148_, _20147_, _20141_);
  and _71079_ (_20150_, _14983_, _07653_);
  or _71080_ (_20151_, _20150_, _20117_);
  and _71081_ (_20152_, _20151_, _09833_);
  or _71082_ (_20153_, _20152_, _06019_);
  or _71083_ (_20154_, _20153_, _20148_);
  and _71084_ (_20155_, _20154_, _20120_);
  or _71085_ (_20156_, _20155_, _06112_);
  and _71086_ (_20157_, _14876_, _07653_);
  or _71087_ (_20158_, _20117_, _08751_);
  or _71088_ (_20159_, _20158_, _20157_);
  and _71089_ (_20161_, _20159_, _08756_);
  and _71090_ (_20162_, _20161_, _20156_);
  and _71091_ (_20163_, _10986_, _07653_);
  or _71092_ (_20164_, _20163_, _20117_);
  and _71093_ (_20165_, _20164_, _06284_);
  or _71094_ (_20166_, _20165_, _20162_);
  and _71095_ (_20167_, _20166_, _07032_);
  or _71096_ (_20168_, _20117_, _08273_);
  and _71097_ (_20169_, _20119_, _06108_);
  and _71098_ (_20170_, _20169_, _20168_);
  or _71099_ (_20172_, _20170_, _20167_);
  and _71100_ (_20173_, _20172_, _06278_);
  and _71101_ (_20174_, _20125_, _06277_);
  and _71102_ (_20175_, _20174_, _20168_);
  or _71103_ (_20176_, _20175_, _06130_);
  or _71104_ (_20177_, _20176_, _20173_);
  and _71105_ (_20178_, _14873_, _07653_);
  or _71106_ (_20179_, _20117_, _08777_);
  or _71107_ (_20180_, _20179_, _20178_);
  and _71108_ (_20181_, _20180_, _08782_);
  and _71109_ (_20183_, _20181_, _20177_);
  nor _71110_ (_20184_, _10985_, _11185_);
  or _71111_ (_20185_, _20184_, _20117_);
  and _71112_ (_20186_, _20185_, _06292_);
  or _71113_ (_20187_, _20186_, _20183_);
  and _71114_ (_20188_, _20187_, _06718_);
  and _71115_ (_20189_, _20122_, _06316_);
  or _71116_ (_20190_, _20189_, _06047_);
  or _71117_ (_20191_, _20190_, _20188_);
  and _71118_ (_20192_, _15055_, _07653_);
  or _71119_ (_20194_, _20117_, _06048_);
  or _71120_ (_20195_, _20194_, _20192_);
  and _71121_ (_20196_, _20195_, _01336_);
  and _71122_ (_20197_, _20196_, _20191_);
  or _71123_ (_20198_, _20197_, _20115_);
  and _71124_ (_43353_, _20198_, _42882_);
  and _71125_ (_20199_, _01340_, \oc8051_golden_model_1.TMOD [5]);
  and _71126_ (_20200_, _11185_, \oc8051_golden_model_1.TMOD [5]);
  or _71127_ (_20201_, _20200_, _07980_);
  and _71128_ (_20202_, _08652_, _07653_);
  or _71129_ (_20204_, _20202_, _20200_);
  and _71130_ (_20205_, _20204_, _06108_);
  and _71131_ (_20206_, _20205_, _20201_);
  or _71132_ (_20207_, _20204_, _06020_);
  and _71133_ (_20208_, _15093_, _07653_);
  or _71134_ (_20209_, _20208_, _20200_);
  or _71135_ (_20210_, _20209_, _06954_);
  and _71136_ (_20211_, _07653_, \oc8051_golden_model_1.ACC [5]);
  or _71137_ (_20212_, _20211_, _20200_);
  and _71138_ (_20213_, _20212_, _06938_);
  and _71139_ (_20215_, _06939_, \oc8051_golden_model_1.TMOD [5]);
  or _71140_ (_20216_, _20215_, _06102_);
  or _71141_ (_20217_, _20216_, _20213_);
  and _71142_ (_20218_, _20217_, _06848_);
  and _71143_ (_20219_, _20218_, _20210_);
  nor _71144_ (_20220_, _07977_, _11185_);
  or _71145_ (_20221_, _20220_, _20200_);
  and _71146_ (_20222_, _20221_, _06239_);
  or _71147_ (_20223_, _20222_, _20219_);
  and _71148_ (_20224_, _20223_, _06220_);
  and _71149_ (_20226_, _20212_, _06219_);
  or _71150_ (_20227_, _20226_, _09818_);
  or _71151_ (_20228_, _20227_, _20224_);
  and _71152_ (_20229_, _09179_, _07653_);
  or _71153_ (_20230_, _20200_, _07012_);
  or _71154_ (_20231_, _20230_, _20229_);
  or _71155_ (_20232_, _20221_, _09827_);
  and _71156_ (_20233_, _20232_, _05669_);
  and _71157_ (_20234_, _20233_, _20231_);
  and _71158_ (_20235_, _20234_, _20228_);
  and _71159_ (_20237_, _15179_, _07653_);
  or _71160_ (_20238_, _20237_, _20200_);
  and _71161_ (_20239_, _20238_, _09833_);
  or _71162_ (_20240_, _20239_, _06019_);
  or _71163_ (_20241_, _20240_, _20235_);
  and _71164_ (_20242_, _20241_, _20207_);
  or _71165_ (_20243_, _20242_, _06112_);
  and _71166_ (_20244_, _15195_, _07653_);
  or _71167_ (_20245_, _20244_, _20200_);
  or _71168_ (_20246_, _20245_, _08751_);
  and _71169_ (_20248_, _20246_, _08756_);
  and _71170_ (_20249_, _20248_, _20243_);
  and _71171_ (_20250_, _12306_, _07653_);
  or _71172_ (_20251_, _20250_, _20200_);
  and _71173_ (_20252_, _20251_, _06284_);
  or _71174_ (_20253_, _20252_, _20249_);
  and _71175_ (_20254_, _20253_, _07032_);
  or _71176_ (_20255_, _20254_, _20206_);
  and _71177_ (_20256_, _20255_, _06278_);
  and _71178_ (_20257_, _20212_, _06277_);
  and _71179_ (_20259_, _20257_, _20201_);
  or _71180_ (_20260_, _20259_, _06130_);
  or _71181_ (_20261_, _20260_, _20256_);
  and _71182_ (_20262_, _15194_, _07653_);
  or _71183_ (_20263_, _20200_, _08777_);
  or _71184_ (_20264_, _20263_, _20262_);
  and _71185_ (_20265_, _20264_, _08782_);
  and _71186_ (_20266_, _20265_, _20261_);
  nor _71187_ (_20267_, _10982_, _11185_);
  or _71188_ (_20268_, _20267_, _20200_);
  and _71189_ (_20270_, _20268_, _06292_);
  or _71190_ (_20271_, _20270_, _20266_);
  and _71191_ (_20272_, _20271_, _06718_);
  and _71192_ (_20273_, _20209_, _06316_);
  or _71193_ (_20274_, _20273_, _06047_);
  or _71194_ (_20275_, _20274_, _20272_);
  and _71195_ (_20276_, _15253_, _07653_);
  or _71196_ (_20277_, _20200_, _06048_);
  or _71197_ (_20278_, _20277_, _20276_);
  and _71198_ (_20279_, _20278_, _01336_);
  and _71199_ (_20281_, _20279_, _20275_);
  or _71200_ (_20282_, _20281_, _20199_);
  and _71201_ (_43354_, _20282_, _42882_);
  and _71202_ (_20283_, _01340_, \oc8051_golden_model_1.TMOD [6]);
  and _71203_ (_20284_, _11185_, \oc8051_golden_model_1.TMOD [6]);
  or _71204_ (_20285_, _20284_, _07886_);
  and _71205_ (_20286_, _15389_, _07653_);
  or _71206_ (_20287_, _20286_, _20284_);
  and _71207_ (_20288_, _20287_, _06108_);
  and _71208_ (_20289_, _20288_, _20285_);
  or _71209_ (_20291_, _20287_, _06020_);
  and _71210_ (_20292_, _15293_, _07653_);
  or _71211_ (_20293_, _20292_, _20284_);
  or _71212_ (_20294_, _20293_, _06954_);
  and _71213_ (_20295_, _07653_, \oc8051_golden_model_1.ACC [6]);
  or _71214_ (_20296_, _20295_, _20284_);
  and _71215_ (_20297_, _20296_, _06938_);
  and _71216_ (_20298_, _06939_, \oc8051_golden_model_1.TMOD [6]);
  or _71217_ (_20299_, _20298_, _06102_);
  or _71218_ (_20300_, _20299_, _20297_);
  and _71219_ (_20302_, _20300_, _06848_);
  and _71220_ (_20303_, _20302_, _20294_);
  nor _71221_ (_20304_, _07883_, _11185_);
  or _71222_ (_20305_, _20304_, _20284_);
  and _71223_ (_20306_, _20305_, _06239_);
  or _71224_ (_20307_, _20306_, _20303_);
  and _71225_ (_20308_, _20307_, _06220_);
  and _71226_ (_20309_, _20296_, _06219_);
  or _71227_ (_20310_, _20309_, _09818_);
  or _71228_ (_20311_, _20310_, _20308_);
  and _71229_ (_20313_, _09178_, _07653_);
  or _71230_ (_20314_, _20284_, _07012_);
  or _71231_ (_20315_, _20314_, _20313_);
  or _71232_ (_20316_, _20305_, _09827_);
  and _71233_ (_20317_, _20316_, _05669_);
  and _71234_ (_20318_, _20317_, _20315_);
  and _71235_ (_20319_, _20318_, _20311_);
  and _71236_ (_20320_, _15382_, _07653_);
  or _71237_ (_20321_, _20320_, _20284_);
  and _71238_ (_20322_, _20321_, _09833_);
  or _71239_ (_20324_, _20322_, _06019_);
  or _71240_ (_20325_, _20324_, _20319_);
  and _71241_ (_20326_, _20325_, _20291_);
  or _71242_ (_20327_, _20326_, _06112_);
  and _71243_ (_20328_, _15399_, _07653_);
  or _71244_ (_20329_, _20328_, _20284_);
  or _71245_ (_20330_, _20329_, _08751_);
  and _71246_ (_20331_, _20330_, _08756_);
  and _71247_ (_20332_, _20331_, _20327_);
  and _71248_ (_20333_, _10980_, _07653_);
  or _71249_ (_20335_, _20333_, _20284_);
  and _71250_ (_20336_, _20335_, _06284_);
  or _71251_ (_20337_, _20336_, _20332_);
  and _71252_ (_20338_, _20337_, _07032_);
  or _71253_ (_20339_, _20338_, _20289_);
  and _71254_ (_20340_, _20339_, _06278_);
  and _71255_ (_20341_, _20296_, _06277_);
  and _71256_ (_20342_, _20341_, _20285_);
  or _71257_ (_20343_, _20342_, _06130_);
  or _71258_ (_20344_, _20343_, _20340_);
  and _71259_ (_20346_, _15396_, _07653_);
  or _71260_ (_20347_, _20284_, _08777_);
  or _71261_ (_20348_, _20347_, _20346_);
  and _71262_ (_20349_, _20348_, _08782_);
  and _71263_ (_20350_, _20349_, _20344_);
  nor _71264_ (_20351_, _10979_, _11185_);
  or _71265_ (_20352_, _20351_, _20284_);
  and _71266_ (_20353_, _20352_, _06292_);
  or _71267_ (_20354_, _20353_, _20350_);
  and _71268_ (_20355_, _20354_, _06718_);
  and _71269_ (_20357_, _20293_, _06316_);
  or _71270_ (_20358_, _20357_, _06047_);
  or _71271_ (_20359_, _20358_, _20355_);
  and _71272_ (_20360_, _15451_, _07653_);
  or _71273_ (_20361_, _20284_, _06048_);
  or _71274_ (_20362_, _20361_, _20360_);
  and _71275_ (_20363_, _20362_, _01336_);
  and _71276_ (_20364_, _20363_, _20359_);
  or _71277_ (_20365_, _20364_, _20283_);
  and _71278_ (_43355_, _20365_, _42882_);
  not _71279_ (_20367_, \oc8051_golden_model_1.DPL [0]);
  nor _71280_ (_20368_, _01336_, _20367_);
  nand _71281_ (_20369_, _10995_, _07733_);
  nor _71282_ (_20370_, _07733_, _20367_);
  nor _71283_ (_20371_, _20370_, _06278_);
  nand _71284_ (_20372_, _20371_, _20369_);
  and _71285_ (_20373_, _09120_, _07733_);
  or _71286_ (_20374_, _20370_, _07012_);
  or _71287_ (_20375_, _20374_, _20373_);
  and _71288_ (_20376_, _07733_, _06931_);
  nor _71289_ (_20378_, _20376_, _20370_);
  nand _71290_ (_20379_, _20378_, _09815_);
  and _71291_ (_20380_, _07733_, \oc8051_golden_model_1.ACC [0]);
  nor _71292_ (_20381_, _20380_, _20370_);
  and _71293_ (_20382_, _20381_, _06219_);
  nor _71294_ (_20383_, _08127_, _11264_);
  or _71295_ (_20384_, _20383_, _20370_);
  or _71296_ (_20385_, _20384_, _06954_);
  nor _71297_ (_20386_, _20381_, _06939_);
  nor _71298_ (_20387_, _06938_, _20367_);
  or _71299_ (_20389_, _20387_, _06102_);
  or _71300_ (_20390_, _20389_, _20386_);
  and _71301_ (_20391_, _20390_, _06848_);
  nand _71302_ (_20392_, _20391_, _20385_);
  or _71303_ (_20393_, _20378_, _06848_);
  and _71304_ (_20394_, _20393_, _06220_);
  and _71305_ (_20395_, _20394_, _20392_);
  or _71306_ (_20396_, _20395_, _20382_);
  and _71307_ (_20397_, _20396_, _11291_);
  and _71308_ (_20398_, _11290_, \oc8051_golden_model_1.DPL [0]);
  or _71309_ (_20400_, _20398_, _06110_);
  or _71310_ (_20401_, _20400_, _20397_);
  or _71311_ (_20402_, _06633_, _06111_);
  and _71312_ (_20403_, _20402_, _09817_);
  nand _71313_ (_20404_, _20403_, _20401_);
  and _71314_ (_20405_, _20404_, _20379_);
  and _71315_ (_20406_, _20405_, _20375_);
  or _71316_ (_20407_, _20406_, _09833_);
  and _71317_ (_20408_, _14186_, _07733_);
  or _71318_ (_20409_, _20370_, _05669_);
  or _71319_ (_20411_, _20409_, _20408_);
  and _71320_ (_20412_, _20411_, _06020_);
  and _71321_ (_20413_, _20412_, _20407_);
  and _71322_ (_20414_, _07733_, _08672_);
  or _71323_ (_20415_, _20414_, _20370_);
  and _71324_ (_20416_, _20415_, _06019_);
  or _71325_ (_20417_, _20416_, _06112_);
  or _71326_ (_20418_, _20417_, _20413_);
  and _71327_ (_20419_, _14086_, _07733_);
  or _71328_ (_20420_, _20370_, _08751_);
  or _71329_ (_20422_, _20420_, _20419_);
  and _71330_ (_20423_, _20422_, _08756_);
  and _71331_ (_20424_, _20423_, _20418_);
  nor _71332_ (_20425_, _12302_, _11264_);
  or _71333_ (_20426_, _20425_, _20370_);
  and _71334_ (_20427_, _20369_, _06284_);
  and _71335_ (_20428_, _20427_, _20426_);
  or _71336_ (_20429_, _20428_, _20424_);
  and _71337_ (_20430_, _20429_, _07032_);
  nand _71338_ (_20431_, _20415_, _06108_);
  nor _71339_ (_20433_, _20431_, _20383_);
  or _71340_ (_20434_, _20433_, _06277_);
  or _71341_ (_20435_, _20434_, _20430_);
  and _71342_ (_20436_, _20435_, _20372_);
  or _71343_ (_20437_, _20436_, _06130_);
  and _71344_ (_20438_, _14083_, _07733_);
  or _71345_ (_20439_, _20370_, _08777_);
  or _71346_ (_20440_, _20439_, _20438_);
  and _71347_ (_20441_, _20440_, _08782_);
  and _71348_ (_20442_, _20441_, _20437_);
  and _71349_ (_20444_, _20426_, _06292_);
  or _71350_ (_20445_, _20444_, _19256_);
  or _71351_ (_20446_, _20445_, _20442_);
  or _71352_ (_20447_, _20384_, _06408_);
  and _71353_ (_20448_, _20447_, _01336_);
  and _71354_ (_20449_, _20448_, _20446_);
  or _71355_ (_20450_, _20449_, _20368_);
  and _71356_ (_43357_, _20450_, _42882_);
  not _71357_ (_20451_, \oc8051_golden_model_1.DPL [1]);
  nor _71358_ (_20452_, _01336_, _20451_);
  and _71359_ (_20454_, _09075_, _07733_);
  nor _71360_ (_20455_, _07733_, _20451_);
  or _71361_ (_20456_, _20455_, _07012_);
  or _71362_ (_20457_, _20456_, _20454_);
  or _71363_ (_20458_, _07733_, \oc8051_golden_model_1.DPL [1]);
  and _71364_ (_20459_, _14284_, _07733_);
  not _71365_ (_20460_, _20459_);
  and _71366_ (_20461_, _20460_, _20458_);
  or _71367_ (_20462_, _20461_, _06954_);
  and _71368_ (_20463_, _07733_, \oc8051_golden_model_1.ACC [1]);
  or _71369_ (_20465_, _20463_, _20455_);
  and _71370_ (_20466_, _20465_, _06938_);
  nor _71371_ (_20467_, _06938_, _20451_);
  or _71372_ (_20468_, _20467_, _06102_);
  or _71373_ (_20469_, _20468_, _20466_);
  and _71374_ (_20470_, _20469_, _06848_);
  and _71375_ (_20471_, _20470_, _20462_);
  nor _71376_ (_20472_, _11264_, _07132_);
  or _71377_ (_20473_, _20472_, _20455_);
  and _71378_ (_20474_, _20473_, _06239_);
  or _71379_ (_20476_, _20474_, _06219_);
  or _71380_ (_20477_, _20476_, _20471_);
  or _71381_ (_20478_, _20465_, _06220_);
  and _71382_ (_20479_, _20478_, _11291_);
  and _71383_ (_20480_, _20479_, _20477_);
  nor _71384_ (_20481_, \oc8051_golden_model_1.DPL [1], \oc8051_golden_model_1.DPL [0]);
  nor _71385_ (_20482_, _20481_, _11295_);
  and _71386_ (_20483_, _20482_, _11290_);
  or _71387_ (_20484_, _20483_, _20480_);
  and _71388_ (_20485_, _20484_, _06111_);
  nor _71389_ (_20487_, _06832_, _06111_);
  or _71390_ (_20488_, _20487_, _09818_);
  or _71391_ (_20489_, _20488_, _20485_);
  or _71392_ (_20490_, _20473_, _09827_);
  and _71393_ (_20491_, _20490_, _05669_);
  and _71394_ (_20492_, _20491_, _20489_);
  and _71395_ (_20493_, _20492_, _20457_);
  or _71396_ (_20494_, _14367_, _11264_);
  and _71397_ (_20495_, _20458_, _09833_);
  and _71398_ (_20496_, _20495_, _20494_);
  or _71399_ (_20498_, _20496_, _20493_);
  and _71400_ (_20499_, _20498_, _06020_);
  nand _71401_ (_20500_, _07733_, _06832_);
  and _71402_ (_20501_, _20458_, _06019_);
  and _71403_ (_20502_, _20501_, _20500_);
  or _71404_ (_20503_, _20502_, _20499_);
  and _71405_ (_20504_, _20503_, _08751_);
  or _71406_ (_20505_, _14263_, _11264_);
  and _71407_ (_20506_, _20458_, _06112_);
  and _71408_ (_20507_, _20506_, _20505_);
  or _71409_ (_20509_, _20507_, _06284_);
  or _71410_ (_20510_, _20509_, _20504_);
  nor _71411_ (_20511_, _10993_, _11264_);
  or _71412_ (_20512_, _20511_, _20455_);
  nand _71413_ (_20513_, _10992_, _07733_);
  and _71414_ (_20514_, _20513_, _20512_);
  or _71415_ (_20515_, _20514_, _08756_);
  and _71416_ (_20516_, _20515_, _07032_);
  and _71417_ (_20517_, _20516_, _20510_);
  or _71418_ (_20518_, _14261_, _11264_);
  and _71419_ (_20520_, _20458_, _06108_);
  and _71420_ (_20521_, _20520_, _20518_);
  or _71421_ (_20522_, _20521_, _06277_);
  or _71422_ (_20523_, _20522_, _20517_);
  nor _71423_ (_20524_, _20455_, _06278_);
  nand _71424_ (_20525_, _20524_, _20513_);
  and _71425_ (_20526_, _20525_, _08777_);
  and _71426_ (_20527_, _20526_, _20523_);
  or _71427_ (_20528_, _20500_, _08078_);
  and _71428_ (_20529_, _20458_, _06130_);
  and _71429_ (_20531_, _20529_, _20528_);
  or _71430_ (_20532_, _20531_, _06292_);
  or _71431_ (_20533_, _20532_, _20527_);
  or _71432_ (_20534_, _20512_, _08782_);
  and _71433_ (_20535_, _20534_, _06718_);
  and _71434_ (_20536_, _20535_, _20533_);
  and _71435_ (_20537_, _20461_, _06316_);
  or _71436_ (_20538_, _20537_, _06047_);
  or _71437_ (_20539_, _20538_, _20536_);
  or _71438_ (_20540_, _20455_, _06048_);
  or _71439_ (_20542_, _20540_, _20459_);
  and _71440_ (_20543_, _20542_, _01336_);
  and _71441_ (_20544_, _20543_, _20539_);
  or _71442_ (_20545_, _20544_, _20452_);
  and _71443_ (_43358_, _20545_, _42882_);
  not _71444_ (_20546_, \oc8051_golden_model_1.DPL [2]);
  nor _71445_ (_20547_, _01336_, _20546_);
  nor _71446_ (_20548_, _07733_, _20546_);
  or _71447_ (_20549_, _20548_, _08177_);
  and _71448_ (_20550_, _07733_, _08730_);
  or _71449_ (_20552_, _20550_, _20548_);
  and _71450_ (_20553_, _20552_, _06108_);
  and _71451_ (_20554_, _20553_, _20549_);
  or _71452_ (_20555_, _20552_, _06020_);
  and _71453_ (_20556_, _14493_, _07733_);
  or _71454_ (_20557_, _20556_, _20548_);
  or _71455_ (_20558_, _20557_, _06954_);
  and _71456_ (_20559_, _07733_, \oc8051_golden_model_1.ACC [2]);
  or _71457_ (_20560_, _20559_, _20548_);
  and _71458_ (_20561_, _20560_, _06938_);
  nor _71459_ (_20563_, _06938_, _20546_);
  or _71460_ (_20564_, _20563_, _06102_);
  or _71461_ (_20565_, _20564_, _20561_);
  and _71462_ (_20566_, _20565_, _06848_);
  and _71463_ (_20567_, _20566_, _20558_);
  nor _71464_ (_20568_, _11264_, _07530_);
  or _71465_ (_20569_, _20568_, _20548_);
  and _71466_ (_20570_, _20569_, _06239_);
  or _71467_ (_20571_, _20570_, _06219_);
  or _71468_ (_20572_, _20571_, _20567_);
  or _71469_ (_20574_, _20560_, _06220_);
  and _71470_ (_20575_, _20574_, _11291_);
  and _71471_ (_20576_, _20575_, _20572_);
  nor _71472_ (_20577_, _11295_, \oc8051_golden_model_1.DPL [2]);
  nor _71473_ (_20578_, _20577_, _11296_);
  and _71474_ (_20579_, _20578_, _11290_);
  or _71475_ (_20580_, _20579_, _20576_);
  and _71476_ (_20581_, _20580_, _06111_);
  nor _71477_ (_20582_, _06445_, _06111_);
  or _71478_ (_20583_, _20582_, _09818_);
  or _71479_ (_20585_, _20583_, _20581_);
  and _71480_ (_20586_, _09182_, _07733_);
  or _71481_ (_20587_, _20548_, _07012_);
  or _71482_ (_20588_, _20587_, _20586_);
  or _71483_ (_20589_, _20569_, _09827_);
  and _71484_ (_20590_, _20589_, _05669_);
  and _71485_ (_20591_, _20590_, _20588_);
  and _71486_ (_20592_, _20591_, _20585_);
  and _71487_ (_20593_, _14580_, _07733_);
  or _71488_ (_20594_, _20593_, _20548_);
  and _71489_ (_20596_, _20594_, _09833_);
  or _71490_ (_20597_, _20596_, _06019_);
  or _71491_ (_20598_, _20597_, _20592_);
  and _71492_ (_20599_, _20598_, _20555_);
  or _71493_ (_20600_, _20599_, _06112_);
  and _71494_ (_20601_, _14596_, _07733_);
  or _71495_ (_20602_, _20601_, _20548_);
  or _71496_ (_20603_, _20602_, _08751_);
  and _71497_ (_20604_, _20603_, _08756_);
  and _71498_ (_20605_, _20604_, _20600_);
  and _71499_ (_20607_, _10991_, _07733_);
  or _71500_ (_20608_, _20607_, _20548_);
  and _71501_ (_20609_, _20608_, _06284_);
  or _71502_ (_20610_, _20609_, _20605_);
  and _71503_ (_20611_, _20610_, _07032_);
  or _71504_ (_20612_, _20611_, _20554_);
  and _71505_ (_20613_, _20612_, _06278_);
  and _71506_ (_20614_, _20560_, _06277_);
  and _71507_ (_20615_, _20614_, _20549_);
  or _71508_ (_20616_, _20615_, _06130_);
  or _71509_ (_20618_, _20616_, _20613_);
  and _71510_ (_20619_, _14593_, _07733_);
  or _71511_ (_20620_, _20548_, _08777_);
  or _71512_ (_20621_, _20620_, _20619_);
  and _71513_ (_20622_, _20621_, _08782_);
  and _71514_ (_20623_, _20622_, _20618_);
  nor _71515_ (_20624_, _10990_, _11264_);
  or _71516_ (_20625_, _20624_, _20548_);
  and _71517_ (_20626_, _20625_, _06292_);
  or _71518_ (_20627_, _20626_, _20623_);
  and _71519_ (_20629_, _20627_, _06718_);
  and _71520_ (_20630_, _20557_, _06316_);
  or _71521_ (_20631_, _20630_, _06047_);
  or _71522_ (_20632_, _20631_, _20629_);
  and _71523_ (_20633_, _14657_, _07733_);
  or _71524_ (_20634_, _20548_, _06048_);
  or _71525_ (_20635_, _20634_, _20633_);
  and _71526_ (_20636_, _20635_, _01336_);
  and _71527_ (_20637_, _20636_, _20632_);
  or _71528_ (_20638_, _20637_, _20547_);
  and _71529_ (_43359_, _20638_, _42882_);
  not _71530_ (_20640_, \oc8051_golden_model_1.DPL [3]);
  nor _71531_ (_20641_, _01336_, _20640_);
  nor _71532_ (_20642_, _07733_, _20640_);
  or _71533_ (_20643_, _20642_, _08029_);
  and _71534_ (_20644_, _07733_, _08662_);
  or _71535_ (_20645_, _20644_, _20642_);
  and _71536_ (_20646_, _20645_, _06108_);
  and _71537_ (_20647_, _20646_, _20643_);
  or _71538_ (_20648_, _20645_, _06020_);
  and _71539_ (_20650_, _14672_, _07733_);
  or _71540_ (_20651_, _20650_, _20642_);
  or _71541_ (_20652_, _20651_, _06954_);
  and _71542_ (_20653_, _07733_, \oc8051_golden_model_1.ACC [3]);
  or _71543_ (_20654_, _20653_, _20642_);
  and _71544_ (_20655_, _20654_, _06938_);
  nor _71545_ (_20656_, _06938_, _20640_);
  or _71546_ (_20657_, _20656_, _06102_);
  or _71547_ (_20658_, _20657_, _20655_);
  and _71548_ (_20659_, _20658_, _06848_);
  and _71549_ (_20661_, _20659_, _20652_);
  nor _71550_ (_20662_, _11264_, _07353_);
  or _71551_ (_20663_, _20662_, _20642_);
  and _71552_ (_20664_, _20663_, _06239_);
  or _71553_ (_20665_, _20664_, _06219_);
  or _71554_ (_20666_, _20665_, _20661_);
  or _71555_ (_20667_, _20654_, _06220_);
  and _71556_ (_20668_, _20667_, _11291_);
  and _71557_ (_20669_, _20668_, _20666_);
  nor _71558_ (_20670_, _11296_, \oc8051_golden_model_1.DPL [3]);
  nor _71559_ (_20672_, _20670_, _11297_);
  and _71560_ (_20673_, _20672_, _11290_);
  or _71561_ (_20674_, _20673_, _20669_);
  and _71562_ (_20675_, _20674_, _06111_);
  nor _71563_ (_20676_, _06215_, _06111_);
  or _71564_ (_20677_, _20676_, _09818_);
  or _71565_ (_20678_, _20677_, _20675_);
  and _71566_ (_20679_, _09181_, _07733_);
  or _71567_ (_20680_, _20642_, _07012_);
  or _71568_ (_20681_, _20680_, _20679_);
  or _71569_ (_20683_, _20663_, _09827_);
  and _71570_ (_20684_, _20683_, _05669_);
  and _71571_ (_20685_, _20684_, _20681_);
  and _71572_ (_20686_, _20685_, _20678_);
  and _71573_ (_20687_, _14778_, _07733_);
  or _71574_ (_20688_, _20687_, _20642_);
  and _71575_ (_20689_, _20688_, _09833_);
  or _71576_ (_20690_, _20689_, _06019_);
  or _71577_ (_20691_, _20690_, _20686_);
  and _71578_ (_20692_, _20691_, _20648_);
  or _71579_ (_20694_, _20692_, _06112_);
  and _71580_ (_20695_, _14793_, _07733_);
  or _71581_ (_20696_, _20642_, _08751_);
  or _71582_ (_20697_, _20696_, _20695_);
  and _71583_ (_20698_, _20697_, _08756_);
  and _71584_ (_20699_, _20698_, _20694_);
  and _71585_ (_20700_, _12299_, _07733_);
  or _71586_ (_20701_, _20700_, _20642_);
  and _71587_ (_20702_, _20701_, _06284_);
  or _71588_ (_20703_, _20702_, _20699_);
  and _71589_ (_20705_, _20703_, _07032_);
  or _71590_ (_20706_, _20705_, _20647_);
  and _71591_ (_20707_, _20706_, _06278_);
  and _71592_ (_20708_, _20654_, _06277_);
  and _71593_ (_20709_, _20708_, _20643_);
  or _71594_ (_20710_, _20709_, _06130_);
  or _71595_ (_20711_, _20710_, _20707_);
  and _71596_ (_20712_, _14792_, _07733_);
  or _71597_ (_20713_, _20642_, _08777_);
  or _71598_ (_20714_, _20713_, _20712_);
  and _71599_ (_20716_, _20714_, _08782_);
  and _71600_ (_20717_, _20716_, _20711_);
  nor _71601_ (_20718_, _10988_, _11264_);
  or _71602_ (_20719_, _20718_, _20642_);
  and _71603_ (_20720_, _20719_, _06292_);
  or _71604_ (_20721_, _20720_, _20717_);
  and _71605_ (_20722_, _20721_, _06718_);
  and _71606_ (_20723_, _20651_, _06316_);
  or _71607_ (_20724_, _20723_, _06047_);
  or _71608_ (_20725_, _20724_, _20722_);
  and _71609_ (_20727_, _14849_, _07733_);
  or _71610_ (_20728_, _20642_, _06048_);
  or _71611_ (_20729_, _20728_, _20727_);
  and _71612_ (_20730_, _20729_, _01336_);
  and _71613_ (_20731_, _20730_, _20725_);
  or _71614_ (_20732_, _20731_, _20641_);
  and _71615_ (_43361_, _20732_, _42882_);
  not _71616_ (_20733_, \oc8051_golden_model_1.DPL [4]);
  nor _71617_ (_20734_, _01336_, _20733_);
  nor _71618_ (_20735_, _07733_, _20733_);
  or _71619_ (_20737_, _20735_, _08273_);
  and _71620_ (_20738_, _08665_, _07733_);
  or _71621_ (_20739_, _20738_, _20735_);
  and _71622_ (_20740_, _20739_, _06108_);
  and _71623_ (_20741_, _20740_, _20737_);
  or _71624_ (_20742_, _20739_, _06020_);
  and _71625_ (_20743_, _14887_, _07733_);
  or _71626_ (_20744_, _20743_, _20735_);
  or _71627_ (_20745_, _20744_, _06954_);
  and _71628_ (_20746_, _07733_, \oc8051_golden_model_1.ACC [4]);
  or _71629_ (_20748_, _20746_, _20735_);
  and _71630_ (_20749_, _20748_, _06938_);
  nor _71631_ (_20750_, _06938_, _20733_);
  or _71632_ (_20751_, _20750_, _06102_);
  or _71633_ (_20752_, _20751_, _20749_);
  and _71634_ (_20753_, _20752_, _06848_);
  and _71635_ (_20754_, _20753_, _20745_);
  nor _71636_ (_20755_, _08270_, _11264_);
  or _71637_ (_20756_, _20755_, _20735_);
  and _71638_ (_20757_, _20756_, _06239_);
  or _71639_ (_20758_, _20757_, _06219_);
  or _71640_ (_20759_, _20758_, _20754_);
  or _71641_ (_20760_, _20748_, _06220_);
  and _71642_ (_20761_, _20760_, _11291_);
  and _71643_ (_20762_, _20761_, _20759_);
  nor _71644_ (_20763_, _11297_, \oc8051_golden_model_1.DPL [4]);
  nor _71645_ (_20764_, _20763_, _11298_);
  and _71646_ (_20765_, _20764_, _11290_);
  or _71647_ (_20766_, _20765_, _20762_);
  and _71648_ (_20767_, _20766_, _06111_);
  nor _71649_ (_20769_, _08581_, _06111_);
  or _71650_ (_20770_, _20769_, _09818_);
  or _71651_ (_20771_, _20770_, _20767_);
  and _71652_ (_20772_, _09180_, _07733_);
  or _71653_ (_20773_, _20735_, _07012_);
  or _71654_ (_20774_, _20773_, _20772_);
  or _71655_ (_20775_, _20756_, _09827_);
  and _71656_ (_20776_, _20775_, _05669_);
  and _71657_ (_20777_, _20776_, _20774_);
  and _71658_ (_20778_, _20777_, _20771_);
  and _71659_ (_20781_, _14983_, _07733_);
  or _71660_ (_20782_, _20781_, _20735_);
  and _71661_ (_20783_, _20782_, _09833_);
  or _71662_ (_20784_, _20783_, _06019_);
  or _71663_ (_20785_, _20784_, _20778_);
  and _71664_ (_20786_, _20785_, _20742_);
  or _71665_ (_20787_, _20786_, _06112_);
  and _71666_ (_20788_, _14876_, _07733_);
  or _71667_ (_20789_, _20788_, _20735_);
  or _71668_ (_20790_, _20789_, _08751_);
  and _71669_ (_20792_, _20790_, _08756_);
  and _71670_ (_20793_, _20792_, _20787_);
  and _71671_ (_20794_, _10986_, _07733_);
  or _71672_ (_20795_, _20794_, _20735_);
  and _71673_ (_20796_, _20795_, _06284_);
  or _71674_ (_20797_, _20796_, _20793_);
  and _71675_ (_20798_, _20797_, _07032_);
  or _71676_ (_20799_, _20798_, _20741_);
  and _71677_ (_20800_, _20799_, _06278_);
  and _71678_ (_20801_, _20748_, _06277_);
  and _71679_ (_20802_, _20801_, _20737_);
  or _71680_ (_20803_, _20802_, _06130_);
  or _71681_ (_20804_, _20803_, _20800_);
  and _71682_ (_20805_, _14873_, _07733_);
  or _71683_ (_20806_, _20735_, _08777_);
  or _71684_ (_20807_, _20806_, _20805_);
  and _71685_ (_20808_, _20807_, _08782_);
  and _71686_ (_20809_, _20808_, _20804_);
  nor _71687_ (_20810_, _10985_, _11264_);
  or _71688_ (_20811_, _20810_, _20735_);
  and _71689_ (_20813_, _20811_, _06292_);
  or _71690_ (_20814_, _20813_, _20809_);
  and _71691_ (_20815_, _20814_, _06718_);
  and _71692_ (_20816_, _20744_, _06316_);
  or _71693_ (_20817_, _20816_, _06047_);
  or _71694_ (_20818_, _20817_, _20815_);
  and _71695_ (_20819_, _15055_, _07733_);
  or _71696_ (_20820_, _20735_, _06048_);
  or _71697_ (_20821_, _20820_, _20819_);
  and _71698_ (_20822_, _20821_, _01336_);
  and _71699_ (_20825_, _20822_, _20818_);
  or _71700_ (_20826_, _20825_, _20734_);
  and _71701_ (_43362_, _20826_, _42882_);
  not _71702_ (_20827_, \oc8051_golden_model_1.DPL [5]);
  nor _71703_ (_20828_, _01336_, _20827_);
  nor _71704_ (_20829_, _07733_, _20827_);
  and _71705_ (_20830_, _08652_, _07733_);
  or _71706_ (_20831_, _20830_, _20829_);
  or _71707_ (_20832_, _20831_, _06020_);
  and _71708_ (_20833_, _15093_, _07733_);
  or _71709_ (_20834_, _20833_, _20829_);
  or _71710_ (_20835_, _20834_, _06954_);
  and _71711_ (_20836_, _07733_, \oc8051_golden_model_1.ACC [5]);
  or _71712_ (_20837_, _20836_, _20829_);
  and _71713_ (_20838_, _20837_, _06938_);
  nor _71714_ (_20839_, _06938_, _20827_);
  or _71715_ (_20840_, _20839_, _06102_);
  or _71716_ (_20841_, _20840_, _20838_);
  and _71717_ (_20842_, _20841_, _06848_);
  and _71718_ (_20843_, _20842_, _20835_);
  nor _71719_ (_20845_, _07977_, _11264_);
  or _71720_ (_20846_, _20845_, _20829_);
  and _71721_ (_20847_, _20846_, _06239_);
  or _71722_ (_20848_, _20847_, _06219_);
  or _71723_ (_20849_, _20848_, _20843_);
  or _71724_ (_20850_, _20837_, _06220_);
  and _71725_ (_20851_, _20850_, _11291_);
  and _71726_ (_20852_, _20851_, _20849_);
  nor _71727_ (_20853_, _11298_, \oc8051_golden_model_1.DPL [5]);
  nor _71728_ (_20854_, _20853_, _11299_);
  and _71729_ (_20857_, _20854_, _11290_);
  or _71730_ (_20858_, _20857_, _20852_);
  and _71731_ (_20859_, _20858_, _06111_);
  nor _71732_ (_20860_, _08612_, _06111_);
  or _71733_ (_20861_, _20860_, _09818_);
  or _71734_ (_20862_, _20861_, _20859_);
  and _71735_ (_20863_, _09179_, _07733_);
  or _71736_ (_20864_, _20829_, _07012_);
  or _71737_ (_20865_, _20864_, _20863_);
  or _71738_ (_20866_, _20846_, _09827_);
  and _71739_ (_20868_, _20866_, _05669_);
  and _71740_ (_20869_, _20868_, _20865_);
  and _71741_ (_20870_, _20869_, _20862_);
  and _71742_ (_20871_, _15179_, _07733_);
  or _71743_ (_20872_, _20871_, _20829_);
  and _71744_ (_20873_, _20872_, _09833_);
  or _71745_ (_20874_, _20873_, _06019_);
  or _71746_ (_20875_, _20874_, _20870_);
  and _71747_ (_20876_, _20875_, _20832_);
  or _71748_ (_20877_, _20876_, _06112_);
  and _71749_ (_20879_, _15195_, _07733_);
  or _71750_ (_20880_, _20879_, _20829_);
  or _71751_ (_20881_, _20880_, _08751_);
  and _71752_ (_20882_, _20881_, _08756_);
  and _71753_ (_20883_, _20882_, _20877_);
  and _71754_ (_20884_, _12306_, _07733_);
  or _71755_ (_20885_, _20884_, _20829_);
  and _71756_ (_20886_, _20885_, _06284_);
  or _71757_ (_20887_, _20886_, _20883_);
  and _71758_ (_20888_, _20887_, _07032_);
  or _71759_ (_20890_, _20829_, _07980_);
  and _71760_ (_20891_, _20831_, _06108_);
  and _71761_ (_20892_, _20891_, _20890_);
  or _71762_ (_20893_, _20892_, _20888_);
  and _71763_ (_20894_, _20893_, _06278_);
  and _71764_ (_20895_, _20837_, _06277_);
  and _71765_ (_20896_, _20895_, _20890_);
  or _71766_ (_20897_, _20896_, _06130_);
  or _71767_ (_20898_, _20897_, _20894_);
  and _71768_ (_20899_, _15194_, _07733_);
  or _71769_ (_20900_, _20829_, _08777_);
  or _71770_ (_20901_, _20900_, _20899_);
  and _71771_ (_20902_, _20901_, _08782_);
  and _71772_ (_20903_, _20902_, _20898_);
  nor _71773_ (_20904_, _10982_, _11264_);
  or _71774_ (_20905_, _20904_, _20829_);
  and _71775_ (_20906_, _20905_, _06292_);
  or _71776_ (_20907_, _20906_, _20903_);
  and _71777_ (_20908_, _20907_, _06718_);
  and _71778_ (_20909_, _20834_, _06316_);
  or _71779_ (_20912_, _20909_, _06047_);
  or _71780_ (_20913_, _20912_, _20908_);
  and _71781_ (_20914_, _15253_, _07733_);
  or _71782_ (_20915_, _20829_, _06048_);
  or _71783_ (_20916_, _20915_, _20914_);
  and _71784_ (_20917_, _20916_, _01336_);
  and _71785_ (_20918_, _20917_, _20913_);
  or _71786_ (_20919_, _20918_, _20828_);
  and _71787_ (_43363_, _20919_, _42882_);
  not _71788_ (_20920_, \oc8051_golden_model_1.DPL [6]);
  nor _71789_ (_20922_, _01336_, _20920_);
  nor _71790_ (_20923_, _07733_, _20920_);
  and _71791_ (_20924_, _15389_, _07733_);
  or _71792_ (_20925_, _20924_, _20923_);
  or _71793_ (_20926_, _20925_, _06020_);
  and _71794_ (_20927_, _15293_, _07733_);
  or _71795_ (_20928_, _20927_, _20923_);
  or _71796_ (_20929_, _20928_, _06954_);
  and _71797_ (_20930_, _07733_, \oc8051_golden_model_1.ACC [6]);
  or _71798_ (_20931_, _20930_, _20923_);
  and _71799_ (_20933_, _20931_, _06938_);
  nor _71800_ (_20934_, _06938_, _20920_);
  or _71801_ (_20935_, _20934_, _06102_);
  or _71802_ (_20936_, _20935_, _20933_);
  and _71803_ (_20937_, _20936_, _06848_);
  and _71804_ (_20938_, _20937_, _20929_);
  nor _71805_ (_20939_, _07883_, _11264_);
  or _71806_ (_20940_, _20939_, _20923_);
  and _71807_ (_20941_, _20940_, _06239_);
  or _71808_ (_20942_, _20941_, _06219_);
  or _71809_ (_20944_, _20942_, _20938_);
  or _71810_ (_20945_, _20931_, _06220_);
  and _71811_ (_20946_, _20945_, _11291_);
  and _71812_ (_20947_, _20946_, _20944_);
  nor _71813_ (_20948_, _11299_, \oc8051_golden_model_1.DPL [6]);
  nor _71814_ (_20949_, _20948_, _11300_);
  and _71815_ (_20950_, _20949_, _11290_);
  or _71816_ (_20951_, _20950_, _20947_);
  and _71817_ (_20952_, _20951_, _06111_);
  nor _71818_ (_20953_, _08647_, _06111_);
  or _71819_ (_20955_, _20953_, _09818_);
  or _71820_ (_20956_, _20955_, _20952_);
  and _71821_ (_20957_, _09178_, _07733_);
  or _71822_ (_20958_, _20923_, _07012_);
  or _71823_ (_20959_, _20958_, _20957_);
  or _71824_ (_20960_, _20940_, _09827_);
  and _71825_ (_20961_, _20960_, _05669_);
  and _71826_ (_20962_, _20961_, _20959_);
  and _71827_ (_20963_, _20962_, _20956_);
  and _71828_ (_20964_, _15382_, _07733_);
  or _71829_ (_20966_, _20964_, _20923_);
  and _71830_ (_20967_, _20966_, _09833_);
  or _71831_ (_20968_, _20967_, _06019_);
  or _71832_ (_20969_, _20968_, _20963_);
  and _71833_ (_20970_, _20969_, _20926_);
  or _71834_ (_20971_, _20970_, _06112_);
  and _71835_ (_20972_, _15399_, _07733_);
  or _71836_ (_20973_, _20923_, _08751_);
  or _71837_ (_20974_, _20973_, _20972_);
  and _71838_ (_20975_, _20974_, _08756_);
  and _71839_ (_20977_, _20975_, _20971_);
  and _71840_ (_20978_, _10980_, _07733_);
  or _71841_ (_20979_, _20978_, _20923_);
  and _71842_ (_20980_, _20979_, _06284_);
  or _71843_ (_20981_, _20980_, _20977_);
  and _71844_ (_20982_, _20981_, _07032_);
  or _71845_ (_20983_, _20923_, _07886_);
  and _71846_ (_20984_, _20925_, _06108_);
  and _71847_ (_20985_, _20984_, _20983_);
  or _71848_ (_20986_, _20985_, _20982_);
  and _71849_ (_20988_, _20986_, _06278_);
  and _71850_ (_20989_, _20931_, _06277_);
  and _71851_ (_20990_, _20989_, _20983_);
  or _71852_ (_20991_, _20990_, _06130_);
  or _71853_ (_20992_, _20991_, _20988_);
  and _71854_ (_20993_, _15396_, _07733_);
  or _71855_ (_20994_, _20923_, _08777_);
  or _71856_ (_20995_, _20994_, _20993_);
  and _71857_ (_20996_, _20995_, _08782_);
  and _71858_ (_20997_, _20996_, _20992_);
  nor _71859_ (_20999_, _10979_, _11264_);
  or _71860_ (_21000_, _20999_, _20923_);
  and _71861_ (_21001_, _21000_, _06292_);
  or _71862_ (_21002_, _21001_, _20997_);
  and _71863_ (_21003_, _21002_, _06718_);
  and _71864_ (_21004_, _20928_, _06316_);
  or _71865_ (_21005_, _21004_, _06047_);
  or _71866_ (_21006_, _21005_, _21003_);
  and _71867_ (_21007_, _15451_, _07733_);
  or _71868_ (_21008_, _20923_, _06048_);
  or _71869_ (_21010_, _21008_, _21007_);
  and _71870_ (_21011_, _21010_, _01336_);
  and _71871_ (_21012_, _21011_, _21006_);
  or _71872_ (_21013_, _21012_, _20922_);
  and _71873_ (_43364_, _21013_, _42882_);
  not _71874_ (_21014_, \oc8051_golden_model_1.DPH [0]);
  nor _71875_ (_21015_, _01336_, _21014_);
  nor _71876_ (_21016_, _07802_, _21014_);
  and _71877_ (_21017_, _07802_, \oc8051_golden_model_1.ACC [0]);
  and _71878_ (_21018_, _21017_, _08127_);
  or _71879_ (_21020_, _21018_, _21016_);
  or _71880_ (_21021_, _21020_, _06278_);
  or _71881_ (_21022_, _21016_, _07012_);
  and _71882_ (_21023_, _09120_, _07802_);
  or _71883_ (_21024_, _21023_, _21022_);
  and _71884_ (_21025_, _07724_, _06931_);
  nor _71885_ (_21026_, _21025_, _21016_);
  nand _71886_ (_21027_, _21026_, _09815_);
  nor _71887_ (_21028_, _08127_, _11359_);
  or _71888_ (_21029_, _21028_, _21016_);
  or _71889_ (_21030_, _21029_, _06954_);
  nor _71890_ (_21031_, _21017_, _21016_);
  nor _71891_ (_21032_, _21031_, _06939_);
  nor _71892_ (_21033_, _06938_, _21014_);
  or _71893_ (_21034_, _21033_, _06102_);
  or _71894_ (_21035_, _21034_, _21032_);
  and _71895_ (_21036_, _21035_, _06848_);
  nand _71896_ (_21037_, _21036_, _21030_);
  or _71897_ (_21038_, _21026_, _06848_);
  and _71898_ (_21039_, _21038_, _06220_);
  and _71899_ (_21042_, _21039_, _21037_);
  and _71900_ (_21043_, _21031_, _06219_);
  or _71901_ (_21044_, _21043_, _11290_);
  or _71902_ (_21045_, _21044_, _21042_);
  nor _71903_ (_21046_, _11302_, \oc8051_golden_model_1.DPH [0]);
  or _71904_ (_21047_, _11388_, _11291_);
  or _71905_ (_21048_, _21047_, _21046_);
  and _71906_ (_21049_, _21048_, _21045_);
  or _71907_ (_21050_, _21049_, _06110_);
  or _71908_ (_21051_, _06111_, _06016_);
  and _71909_ (_21053_, _21051_, _09817_);
  nand _71910_ (_21054_, _21053_, _21050_);
  and _71911_ (_21055_, _21054_, _21027_);
  and _71912_ (_21056_, _21055_, _21024_);
  or _71913_ (_21057_, _21056_, _09833_);
  and _71914_ (_21058_, _14186_, _07724_);
  or _71915_ (_21059_, _21016_, _05669_);
  or _71916_ (_21060_, _21059_, _21058_);
  and _71917_ (_21061_, _21060_, _06020_);
  and _71918_ (_21062_, _21061_, _21057_);
  and _71919_ (_21064_, _07802_, _08672_);
  or _71920_ (_21065_, _21064_, _21016_);
  and _71921_ (_21066_, _21065_, _06019_);
  or _71922_ (_21067_, _21066_, _06112_);
  or _71923_ (_21068_, _21067_, _21062_);
  and _71924_ (_21069_, _14086_, _07724_);
  or _71925_ (_21070_, _21016_, _08751_);
  or _71926_ (_21071_, _21070_, _21069_);
  and _71927_ (_21072_, _21071_, _08756_);
  and _71928_ (_21073_, _21072_, _21068_);
  nor _71929_ (_21075_, _12302_, _11359_);
  or _71930_ (_21076_, _21075_, _21016_);
  nor _71931_ (_21077_, _21018_, _08756_);
  and _71932_ (_21078_, _21077_, _21076_);
  or _71933_ (_21079_, _21078_, _21073_);
  and _71934_ (_21080_, _21079_, _07032_);
  nand _71935_ (_21081_, _21065_, _06108_);
  nor _71936_ (_21082_, _21081_, _21028_);
  or _71937_ (_21083_, _21082_, _06277_);
  or _71938_ (_21084_, _21083_, _21080_);
  and _71939_ (_21086_, _21084_, _21021_);
  or _71940_ (_21087_, _21086_, _06130_);
  and _71941_ (_21088_, _14083_, _07724_);
  or _71942_ (_21089_, _21016_, _08777_);
  or _71943_ (_21090_, _21089_, _21088_);
  and _71944_ (_21091_, _21090_, _08782_);
  and _71945_ (_21092_, _21091_, _21087_);
  and _71946_ (_21093_, _21076_, _06292_);
  or _71947_ (_21094_, _21093_, _19256_);
  or _71948_ (_21095_, _21094_, _21092_);
  or _71949_ (_21097_, _21029_, _06408_);
  and _71950_ (_21098_, _21097_, _01336_);
  and _71951_ (_21099_, _21098_, _21095_);
  or _71952_ (_21100_, _21099_, _21015_);
  and _71953_ (_43366_, _21100_, _42882_);
  not _71954_ (_21101_, \oc8051_golden_model_1.DPH [1]);
  nor _71955_ (_21102_, _01336_, _21101_);
  or _71956_ (_21103_, _07802_, \oc8051_golden_model_1.DPH [1]);
  and _71957_ (_21104_, _21103_, _09833_);
  or _71958_ (_21105_, _14367_, _11359_);
  and _71959_ (_21107_, _21105_, _21104_);
  nor _71960_ (_21108_, _07802_, _21101_);
  nor _71961_ (_21109_, _11359_, _07132_);
  or _71962_ (_21110_, _21109_, _21108_);
  or _71963_ (_21111_, _21110_, _06848_);
  and _71964_ (_21112_, _14284_, _07724_);
  not _71965_ (_21113_, _21112_);
  and _71966_ (_21114_, _21113_, _21103_);
  and _71967_ (_21115_, _21114_, _06102_);
  nor _71968_ (_21116_, _06938_, _21101_);
  and _71969_ (_21118_, _07802_, \oc8051_golden_model_1.ACC [1]);
  or _71970_ (_21119_, _21118_, _21108_);
  and _71971_ (_21120_, _21119_, _06938_);
  or _71972_ (_21121_, _21120_, _21116_);
  and _71973_ (_21122_, _21121_, _06954_);
  or _71974_ (_21123_, _21122_, _06239_);
  or _71975_ (_21124_, _21123_, _21115_);
  and _71976_ (_21125_, _21124_, _21111_);
  or _71977_ (_21126_, _21125_, _06219_);
  or _71978_ (_21127_, _21119_, _06220_);
  and _71979_ (_21129_, _21127_, _11291_);
  and _71980_ (_21130_, _21129_, _21126_);
  or _71981_ (_21131_, _11388_, \oc8051_golden_model_1.DPH [1]);
  nand _71982_ (_21132_, _21131_, _11290_);
  nor _71983_ (_21133_, _21132_, _11389_);
  or _71984_ (_21134_, _21133_, _21130_);
  and _71985_ (_21135_, _21134_, _06111_);
  nor _71986_ (_21136_, _06799_, _06111_);
  or _71987_ (_21137_, _21136_, _09818_);
  or _71988_ (_21138_, _21137_, _21135_);
  or _71989_ (_21140_, _21108_, _07012_);
  and _71990_ (_21141_, _09075_, _07802_);
  or _71991_ (_21142_, _21141_, _21140_);
  or _71992_ (_21143_, _21110_, _09827_);
  and _71993_ (_21144_, _21143_, _05669_);
  and _71994_ (_21145_, _21144_, _21142_);
  and _71995_ (_21146_, _21145_, _21138_);
  or _71996_ (_21147_, _21146_, _21107_);
  and _71997_ (_21148_, _21147_, _06020_);
  and _71998_ (_21149_, _21103_, _06019_);
  nand _71999_ (_21151_, _07724_, _06832_);
  and _72000_ (_21152_, _21151_, _21149_);
  or _72001_ (_21153_, _21152_, _21148_);
  and _72002_ (_21154_, _21153_, _08751_);
  or _72003_ (_21155_, _14263_, _11359_);
  and _72004_ (_21156_, _21103_, _06112_);
  and _72005_ (_21157_, _21156_, _21155_);
  or _72006_ (_21158_, _21157_, _06284_);
  or _72007_ (_21159_, _21158_, _21154_);
  nor _72008_ (_21160_, _10993_, _11359_);
  or _72009_ (_21162_, _21160_, _21108_);
  nand _72010_ (_21163_, _10992_, _07724_);
  and _72011_ (_21164_, _21163_, _21162_);
  or _72012_ (_21165_, _21164_, _08756_);
  and _72013_ (_21166_, _21165_, _07032_);
  and _72014_ (_21167_, _21166_, _21159_);
  or _72015_ (_21168_, _14261_, _11359_);
  and _72016_ (_21169_, _21103_, _06108_);
  and _72017_ (_21170_, _21169_, _21168_);
  or _72018_ (_21171_, _21170_, _06277_);
  or _72019_ (_21173_, _21171_, _21167_);
  nor _72020_ (_21174_, _21108_, _06278_);
  nand _72021_ (_21175_, _21174_, _21163_);
  and _72022_ (_21176_, _21175_, _08777_);
  and _72023_ (_21177_, _21176_, _21173_);
  or _72024_ (_21178_, _21151_, _08078_);
  and _72025_ (_21179_, _21103_, _06130_);
  and _72026_ (_21180_, _21179_, _21178_);
  or _72027_ (_21181_, _21180_, _06292_);
  or _72028_ (_21182_, _21181_, _21177_);
  or _72029_ (_21184_, _21162_, _08782_);
  and _72030_ (_21185_, _21184_, _06718_);
  and _72031_ (_21186_, _21185_, _21182_);
  and _72032_ (_21187_, _21114_, _06316_);
  or _72033_ (_21188_, _21187_, _06047_);
  or _72034_ (_21189_, _21188_, _21186_);
  or _72035_ (_21190_, _21108_, _06048_);
  or _72036_ (_21191_, _21190_, _21112_);
  and _72037_ (_21192_, _21191_, _01336_);
  and _72038_ (_21193_, _21192_, _21189_);
  or _72039_ (_21195_, _21193_, _21102_);
  and _72040_ (_43367_, _21195_, _42882_);
  and _72041_ (_21196_, _01340_, \oc8051_golden_model_1.DPH [2]);
  and _72042_ (_21197_, _11359_, \oc8051_golden_model_1.DPH [2]);
  and _72043_ (_21198_, _07802_, _08730_);
  or _72044_ (_21199_, _21198_, _21197_);
  or _72045_ (_21200_, _21199_, _06020_);
  and _72046_ (_21201_, _14493_, _07724_);
  or _72047_ (_21202_, _21201_, _21197_);
  or _72048_ (_21203_, _21202_, _06954_);
  and _72049_ (_21204_, _07802_, \oc8051_golden_model_1.ACC [2]);
  or _72050_ (_21205_, _21204_, _21197_);
  and _72051_ (_21206_, _21205_, _06938_);
  and _72052_ (_21207_, _06939_, \oc8051_golden_model_1.DPH [2]);
  or _72053_ (_21208_, _21207_, _06102_);
  or _72054_ (_21209_, _21208_, _21206_);
  and _72055_ (_21210_, _21209_, _06848_);
  and _72056_ (_21211_, _21210_, _21203_);
  nor _72057_ (_21212_, _11359_, _07530_);
  or _72058_ (_21213_, _21212_, _21197_);
  and _72059_ (_21216_, _21213_, _06239_);
  or _72060_ (_21217_, _21216_, _06219_);
  or _72061_ (_21218_, _21217_, _21211_);
  or _72062_ (_21219_, _21205_, _06220_);
  and _72063_ (_21220_, _21219_, _11291_);
  and _72064_ (_21221_, _21220_, _21218_);
  or _72065_ (_21222_, _11389_, \oc8051_golden_model_1.DPH [2]);
  nor _72066_ (_21223_, _11390_, _11291_);
  and _72067_ (_21224_, _21223_, _21222_);
  or _72068_ (_21225_, _21224_, _21221_);
  and _72069_ (_21227_, _21225_, _06111_);
  nor _72070_ (_21228_, _06403_, _06111_);
  or _72071_ (_21229_, _21228_, _09818_);
  or _72072_ (_21230_, _21229_, _21227_);
  or _72073_ (_21231_, _21197_, _07012_);
  and _72074_ (_21232_, _09182_, _07802_);
  or _72075_ (_21233_, _21232_, _21231_);
  or _72076_ (_21234_, _21213_, _09827_);
  and _72077_ (_21235_, _21234_, _05669_);
  and _72078_ (_21236_, _21235_, _21233_);
  and _72079_ (_21238_, _21236_, _21230_);
  and _72080_ (_21239_, _14580_, _07724_);
  or _72081_ (_21240_, _21239_, _21197_);
  and _72082_ (_21241_, _21240_, _09833_);
  or _72083_ (_21242_, _21241_, _06019_);
  or _72084_ (_21243_, _21242_, _21238_);
  and _72085_ (_21244_, _21243_, _21200_);
  or _72086_ (_21245_, _21244_, _06112_);
  and _72087_ (_21246_, _14596_, _07724_);
  or _72088_ (_21247_, _21197_, _08751_);
  or _72089_ (_21249_, _21247_, _21246_);
  and _72090_ (_21250_, _21249_, _08756_);
  and _72091_ (_21251_, _21250_, _21245_);
  and _72092_ (_21252_, _10991_, _07802_);
  or _72093_ (_21253_, _21252_, _21197_);
  and _72094_ (_21254_, _21253_, _06284_);
  or _72095_ (_21255_, _21254_, _21251_);
  and _72096_ (_21256_, _21255_, _07032_);
  or _72097_ (_21257_, _21197_, _08177_);
  and _72098_ (_21258_, _21199_, _06108_);
  and _72099_ (_21260_, _21258_, _21257_);
  or _72100_ (_21261_, _21260_, _21256_);
  and _72101_ (_21262_, _21261_, _06278_);
  and _72102_ (_21263_, _21205_, _06277_);
  and _72103_ (_21264_, _21263_, _21257_);
  or _72104_ (_21265_, _21264_, _06130_);
  or _72105_ (_21266_, _21265_, _21262_);
  and _72106_ (_21267_, _14593_, _07724_);
  or _72107_ (_21268_, _21197_, _08777_);
  or _72108_ (_21269_, _21268_, _21267_);
  and _72109_ (_21271_, _21269_, _08782_);
  and _72110_ (_21272_, _21271_, _21266_);
  nor _72111_ (_21273_, _10990_, _11359_);
  or _72112_ (_21274_, _21273_, _21197_);
  and _72113_ (_21275_, _21274_, _06292_);
  or _72114_ (_21276_, _21275_, _21272_);
  and _72115_ (_21277_, _21276_, _06718_);
  and _72116_ (_21278_, _21202_, _06316_);
  or _72117_ (_21279_, _21278_, _06047_);
  or _72118_ (_21280_, _21279_, _21277_);
  and _72119_ (_21282_, _14657_, _07724_);
  or _72120_ (_21283_, _21197_, _06048_);
  or _72121_ (_21284_, _21283_, _21282_);
  and _72122_ (_21285_, _21284_, _01336_);
  and _72123_ (_21286_, _21285_, _21280_);
  or _72124_ (_21287_, _21286_, _21196_);
  and _72125_ (_43368_, _21287_, _42882_);
  and _72126_ (_21288_, _01340_, \oc8051_golden_model_1.DPH [3]);
  and _72127_ (_21289_, _11359_, \oc8051_golden_model_1.DPH [3]);
  or _72128_ (_21290_, _21289_, _08029_);
  and _72129_ (_21292_, _07802_, _08662_);
  or _72130_ (_21293_, _21292_, _21289_);
  and _72131_ (_21294_, _21293_, _06108_);
  and _72132_ (_21295_, _21294_, _21290_);
  or _72133_ (_21296_, _21293_, _06020_);
  and _72134_ (_21297_, _14672_, _07724_);
  or _72135_ (_21298_, _21297_, _21289_);
  or _72136_ (_21299_, _21298_, _06954_);
  and _72137_ (_21300_, _07802_, \oc8051_golden_model_1.ACC [3]);
  or _72138_ (_21301_, _21300_, _21289_);
  and _72139_ (_21303_, _21301_, _06938_);
  and _72140_ (_21304_, _06939_, \oc8051_golden_model_1.DPH [3]);
  or _72141_ (_21305_, _21304_, _06102_);
  or _72142_ (_21306_, _21305_, _21303_);
  and _72143_ (_21307_, _21306_, _06848_);
  and _72144_ (_21308_, _21307_, _21299_);
  nor _72145_ (_21309_, _11359_, _07353_);
  or _72146_ (_21310_, _21309_, _21289_);
  and _72147_ (_21311_, _21310_, _06239_);
  or _72148_ (_21312_, _21311_, _06219_);
  or _72149_ (_21314_, _21312_, _21308_);
  or _72150_ (_21315_, _21301_, _06220_);
  and _72151_ (_21316_, _21315_, _11291_);
  and _72152_ (_21317_, _21316_, _21314_);
  or _72153_ (_21318_, _11390_, \oc8051_golden_model_1.DPH [3]);
  nor _72154_ (_21319_, _11391_, _11291_);
  and _72155_ (_21320_, _21319_, _21318_);
  or _72156_ (_21321_, _21320_, _21317_);
  and _72157_ (_21322_, _21321_, _06111_);
  nor _72158_ (_21323_, _06111_, _05983_);
  or _72159_ (_21325_, _21323_, _09818_);
  or _72160_ (_21326_, _21325_, _21322_);
  or _72161_ (_21327_, _21289_, _07012_);
  and _72162_ (_21328_, _09181_, _07802_);
  or _72163_ (_21329_, _21328_, _21327_);
  or _72164_ (_21330_, _21310_, _09827_);
  and _72165_ (_21331_, _21330_, _05669_);
  and _72166_ (_21332_, _21331_, _21329_);
  and _72167_ (_21333_, _21332_, _21326_);
  and _72168_ (_21334_, _14778_, _07724_);
  or _72169_ (_21336_, _21334_, _21289_);
  and _72170_ (_21337_, _21336_, _09833_);
  or _72171_ (_21338_, _21337_, _06019_);
  or _72172_ (_21339_, _21338_, _21333_);
  and _72173_ (_21340_, _21339_, _21296_);
  or _72174_ (_21341_, _21340_, _06112_);
  and _72175_ (_21342_, _14793_, _07802_);
  or _72176_ (_21343_, _21342_, _21289_);
  or _72177_ (_21344_, _21343_, _08751_);
  and _72178_ (_21345_, _21344_, _08756_);
  and _72179_ (_21347_, _21345_, _21341_);
  and _72180_ (_21348_, _12299_, _07802_);
  or _72181_ (_21349_, _21348_, _21289_);
  and _72182_ (_21350_, _21349_, _06284_);
  or _72183_ (_21351_, _21350_, _21347_);
  and _72184_ (_21352_, _21351_, _07032_);
  or _72185_ (_21353_, _21352_, _21295_);
  and _72186_ (_21354_, _21353_, _06278_);
  and _72187_ (_21355_, _21301_, _06277_);
  and _72188_ (_21356_, _21355_, _21290_);
  or _72189_ (_21358_, _21356_, _06130_);
  or _72190_ (_21359_, _21358_, _21354_);
  and _72191_ (_21360_, _14792_, _07724_);
  or _72192_ (_21361_, _21289_, _08777_);
  or _72193_ (_21362_, _21361_, _21360_);
  and _72194_ (_21363_, _21362_, _08782_);
  and _72195_ (_21364_, _21363_, _21359_);
  nor _72196_ (_21365_, _10988_, _11359_);
  or _72197_ (_21366_, _21365_, _21289_);
  and _72198_ (_21367_, _21366_, _06292_);
  or _72199_ (_21369_, _21367_, _21364_);
  and _72200_ (_21370_, _21369_, _06718_);
  and _72201_ (_21371_, _21298_, _06316_);
  or _72202_ (_21372_, _21371_, _06047_);
  or _72203_ (_21373_, _21372_, _21370_);
  and _72204_ (_21374_, _14849_, _07724_);
  or _72205_ (_21375_, _21289_, _06048_);
  or _72206_ (_21376_, _21375_, _21374_);
  and _72207_ (_21377_, _21376_, _01336_);
  and _72208_ (_21378_, _21377_, _21373_);
  or _72209_ (_21380_, _21378_, _21288_);
  and _72210_ (_43369_, _21380_, _42882_);
  not _72211_ (_21381_, \oc8051_golden_model_1.DPH [4]);
  nor _72212_ (_21382_, _01336_, _21381_);
  nor _72213_ (_21383_, _07802_, _21381_);
  or _72214_ (_21384_, _21383_, _08273_);
  and _72215_ (_21385_, _08665_, _07802_);
  or _72216_ (_21386_, _21385_, _21383_);
  and _72217_ (_21387_, _21386_, _06108_);
  and _72218_ (_21388_, _21387_, _21384_);
  or _72219_ (_21390_, _21386_, _06020_);
  and _72220_ (_21391_, _14887_, _07724_);
  or _72221_ (_21392_, _21391_, _21383_);
  or _72222_ (_21393_, _21392_, _06954_);
  and _72223_ (_21394_, _07802_, \oc8051_golden_model_1.ACC [4]);
  or _72224_ (_21395_, _21394_, _21383_);
  and _72225_ (_21396_, _21395_, _06938_);
  nor _72226_ (_21397_, _06938_, _21381_);
  or _72227_ (_21398_, _21397_, _06102_);
  or _72228_ (_21399_, _21398_, _21396_);
  and _72229_ (_21400_, _21399_, _06848_);
  and _72230_ (_21401_, _21400_, _21393_);
  nor _72231_ (_21402_, _08270_, _11359_);
  or _72232_ (_21403_, _21402_, _21383_);
  and _72233_ (_21404_, _21403_, _06239_);
  or _72234_ (_21405_, _21404_, _06219_);
  or _72235_ (_21406_, _21405_, _21401_);
  or _72236_ (_21407_, _21395_, _06220_);
  and _72237_ (_21408_, _21407_, _11291_);
  and _72238_ (_21409_, _21408_, _21406_);
  or _72239_ (_21412_, _11391_, \oc8051_golden_model_1.DPH [4]);
  nor _72240_ (_21413_, _11392_, _11291_);
  and _72241_ (_21414_, _21413_, _21412_);
  or _72242_ (_21415_, _21414_, _21409_);
  and _72243_ (_21416_, _21415_, _06111_);
  nor _72244_ (_21417_, _06758_, _06111_);
  or _72245_ (_21418_, _21417_, _09818_);
  or _72246_ (_21419_, _21418_, _21416_);
  or _72247_ (_21420_, _21383_, _07012_);
  and _72248_ (_21421_, _09180_, _07802_);
  or _72249_ (_21423_, _21421_, _21420_);
  or _72250_ (_21424_, _21403_, _09827_);
  and _72251_ (_21425_, _21424_, _05669_);
  and _72252_ (_21426_, _21425_, _21423_);
  and _72253_ (_21427_, _21426_, _21419_);
  and _72254_ (_21428_, _14983_, _07724_);
  or _72255_ (_21429_, _21428_, _21383_);
  and _72256_ (_21430_, _21429_, _09833_);
  or _72257_ (_21431_, _21430_, _06019_);
  or _72258_ (_21432_, _21431_, _21427_);
  and _72259_ (_21434_, _21432_, _21390_);
  or _72260_ (_21435_, _21434_, _06112_);
  and _72261_ (_21436_, _14876_, _07802_);
  or _72262_ (_21437_, _21436_, _21383_);
  or _72263_ (_21438_, _21437_, _08751_);
  and _72264_ (_21439_, _21438_, _08756_);
  and _72265_ (_21440_, _21439_, _21435_);
  and _72266_ (_21441_, _10986_, _07802_);
  or _72267_ (_21442_, _21441_, _21383_);
  and _72268_ (_21443_, _21442_, _06284_);
  or _72269_ (_21445_, _21443_, _21440_);
  and _72270_ (_21446_, _21445_, _07032_);
  or _72271_ (_21447_, _21446_, _21388_);
  and _72272_ (_21448_, _21447_, _06278_);
  and _72273_ (_21449_, _21395_, _06277_);
  and _72274_ (_21450_, _21449_, _21384_);
  or _72275_ (_21451_, _21450_, _06130_);
  or _72276_ (_21452_, _21451_, _21448_);
  and _72277_ (_21453_, _14873_, _07724_);
  or _72278_ (_21454_, _21383_, _08777_);
  or _72279_ (_21456_, _21454_, _21453_);
  and _72280_ (_21457_, _21456_, _08782_);
  and _72281_ (_21458_, _21457_, _21452_);
  nor _72282_ (_21459_, _10985_, _11359_);
  or _72283_ (_21460_, _21459_, _21383_);
  and _72284_ (_21461_, _21460_, _06292_);
  or _72285_ (_21462_, _21461_, _21458_);
  and _72286_ (_21463_, _21462_, _06718_);
  and _72287_ (_21464_, _21392_, _06316_);
  or _72288_ (_21465_, _21464_, _06047_);
  or _72289_ (_21467_, _21465_, _21463_);
  and _72290_ (_21468_, _15055_, _07724_);
  or _72291_ (_21469_, _21383_, _06048_);
  or _72292_ (_21470_, _21469_, _21468_);
  and _72293_ (_21471_, _21470_, _01336_);
  and _72294_ (_21472_, _21471_, _21467_);
  or _72295_ (_21473_, _21472_, _21382_);
  and _72296_ (_43370_, _21473_, _42882_);
  and _72297_ (_21474_, _01340_, \oc8051_golden_model_1.DPH [5]);
  and _72298_ (_21475_, _11359_, \oc8051_golden_model_1.DPH [5]);
  and _72299_ (_21477_, _08652_, _07802_);
  or _72300_ (_21478_, _21477_, _21475_);
  or _72301_ (_21479_, _21478_, _06020_);
  and _72302_ (_21480_, _15093_, _07724_);
  or _72303_ (_21481_, _21480_, _21475_);
  or _72304_ (_21482_, _21481_, _06954_);
  and _72305_ (_21483_, _07802_, \oc8051_golden_model_1.ACC [5]);
  or _72306_ (_21484_, _21483_, _21475_);
  and _72307_ (_21485_, _21484_, _06938_);
  and _72308_ (_21486_, _06939_, \oc8051_golden_model_1.DPH [5]);
  or _72309_ (_21488_, _21486_, _06102_);
  or _72310_ (_21489_, _21488_, _21485_);
  and _72311_ (_21490_, _21489_, _06848_);
  and _72312_ (_21491_, _21490_, _21482_);
  nor _72313_ (_21492_, _07977_, _11359_);
  or _72314_ (_21493_, _21492_, _21475_);
  and _72315_ (_21494_, _21493_, _06239_);
  or _72316_ (_21495_, _21494_, _06219_);
  or _72317_ (_21496_, _21495_, _21491_);
  or _72318_ (_21497_, _21484_, _06220_);
  and _72319_ (_21499_, _21497_, _11291_);
  and _72320_ (_21500_, _21499_, _21496_);
  or _72321_ (_21501_, _11392_, \oc8051_golden_model_1.DPH [5]);
  nor _72322_ (_21502_, _11393_, _11291_);
  and _72323_ (_21503_, _21502_, _21501_);
  or _72324_ (_21504_, _21503_, _21500_);
  and _72325_ (_21505_, _21504_, _06111_);
  nor _72326_ (_21506_, _06359_, _06111_);
  or _72327_ (_21507_, _21506_, _09818_);
  or _72328_ (_21508_, _21507_, _21505_);
  or _72329_ (_21510_, _21475_, _07012_);
  and _72330_ (_21511_, _09179_, _07802_);
  or _72331_ (_21512_, _21511_, _21510_);
  or _72332_ (_21513_, _21493_, _09827_);
  and _72333_ (_21514_, _21513_, _05669_);
  and _72334_ (_21515_, _21514_, _21512_);
  and _72335_ (_21516_, _21515_, _21508_);
  and _72336_ (_21517_, _15179_, _07724_);
  or _72337_ (_21518_, _21517_, _21475_);
  and _72338_ (_21519_, _21518_, _09833_);
  or _72339_ (_21521_, _21519_, _06019_);
  or _72340_ (_21522_, _21521_, _21516_);
  and _72341_ (_21523_, _21522_, _21479_);
  or _72342_ (_21524_, _21523_, _06112_);
  and _72343_ (_21525_, _15195_, _07802_);
  or _72344_ (_21526_, _21525_, _21475_);
  or _72345_ (_21527_, _21526_, _08751_);
  and _72346_ (_21528_, _21527_, _08756_);
  and _72347_ (_21529_, _21528_, _21524_);
  and _72348_ (_21530_, _12306_, _07802_);
  or _72349_ (_21532_, _21530_, _21475_);
  and _72350_ (_21533_, _21532_, _06284_);
  or _72351_ (_21534_, _21533_, _21529_);
  and _72352_ (_21535_, _21534_, _07032_);
  or _72353_ (_21536_, _21475_, _07980_);
  and _72354_ (_21537_, _21478_, _06108_);
  and _72355_ (_21538_, _21537_, _21536_);
  or _72356_ (_21539_, _21538_, _21535_);
  and _72357_ (_21540_, _21539_, _06278_);
  and _72358_ (_21541_, _21484_, _06277_);
  and _72359_ (_21543_, _21541_, _21536_);
  or _72360_ (_21544_, _21543_, _06130_);
  or _72361_ (_21545_, _21544_, _21540_);
  and _72362_ (_21546_, _15194_, _07724_);
  or _72363_ (_21547_, _21475_, _08777_);
  or _72364_ (_21548_, _21547_, _21546_);
  and _72365_ (_21549_, _21548_, _08782_);
  and _72366_ (_21550_, _21549_, _21545_);
  nor _72367_ (_21551_, _10982_, _11359_);
  or _72368_ (_21552_, _21551_, _21475_);
  and _72369_ (_21554_, _21552_, _06292_);
  or _72370_ (_21555_, _21554_, _21550_);
  and _72371_ (_21556_, _21555_, _06718_);
  and _72372_ (_21557_, _21481_, _06316_);
  or _72373_ (_21558_, _21557_, _06047_);
  or _72374_ (_21559_, _21558_, _21556_);
  and _72375_ (_21560_, _15253_, _07724_);
  or _72376_ (_21561_, _21475_, _06048_);
  or _72377_ (_21562_, _21561_, _21560_);
  and _72378_ (_21563_, _21562_, _01336_);
  and _72379_ (_21565_, _21563_, _21559_);
  or _72380_ (_21566_, _21565_, _21474_);
  and _72381_ (_43371_, _21566_, _42882_);
  and _72382_ (_21567_, _01340_, \oc8051_golden_model_1.DPH [6]);
  and _72383_ (_21568_, _11359_, \oc8051_golden_model_1.DPH [6]);
  and _72384_ (_21569_, _15389_, _07802_);
  or _72385_ (_21570_, _21569_, _21568_);
  or _72386_ (_21571_, _21570_, _06020_);
  and _72387_ (_21572_, _15293_, _07724_);
  or _72388_ (_21573_, _21572_, _21568_);
  or _72389_ (_21575_, _21573_, _06954_);
  and _72390_ (_21576_, _07802_, \oc8051_golden_model_1.ACC [6]);
  or _72391_ (_21577_, _21576_, _21568_);
  and _72392_ (_21578_, _21577_, _06938_);
  and _72393_ (_21579_, _06939_, \oc8051_golden_model_1.DPH [6]);
  or _72394_ (_21580_, _21579_, _06102_);
  or _72395_ (_21581_, _21580_, _21578_);
  and _72396_ (_21582_, _21581_, _06848_);
  and _72397_ (_21583_, _21582_, _21575_);
  nor _72398_ (_21584_, _07883_, _11359_);
  or _72399_ (_21586_, _21584_, _21568_);
  and _72400_ (_21587_, _21586_, _06239_);
  or _72401_ (_21588_, _21587_, _06219_);
  or _72402_ (_21589_, _21588_, _21583_);
  or _72403_ (_21590_, _21577_, _06220_);
  and _72404_ (_21591_, _21590_, _11291_);
  and _72405_ (_21592_, _21591_, _21589_);
  or _72406_ (_21593_, _11393_, \oc8051_golden_model_1.DPH [6]);
  nor _72407_ (_21594_, _11394_, _11291_);
  and _72408_ (_21595_, _21594_, _21593_);
  or _72409_ (_21597_, _21595_, _21592_);
  and _72410_ (_21598_, _21597_, _06111_);
  nor _72411_ (_21599_, _06111_, _06084_);
  or _72412_ (_21600_, _21599_, _09818_);
  or _72413_ (_21601_, _21600_, _21598_);
  or _72414_ (_21602_, _21568_, _07012_);
  and _72415_ (_21603_, _09178_, _07802_);
  or _72416_ (_21604_, _21603_, _21602_);
  or _72417_ (_21605_, _21586_, _09827_);
  and _72418_ (_21606_, _21605_, _05669_);
  and _72419_ (_21608_, _21606_, _21604_);
  and _72420_ (_21609_, _21608_, _21601_);
  and _72421_ (_21610_, _15382_, _07724_);
  or _72422_ (_21611_, _21610_, _21568_);
  and _72423_ (_21612_, _21611_, _09833_);
  or _72424_ (_21613_, _21612_, _06019_);
  or _72425_ (_21614_, _21613_, _21609_);
  and _72426_ (_21615_, _21614_, _21571_);
  or _72427_ (_21616_, _21615_, _06112_);
  and _72428_ (_21617_, _15399_, _07724_);
  or _72429_ (_21619_, _21568_, _08751_);
  or _72430_ (_21620_, _21619_, _21617_);
  and _72431_ (_21621_, _21620_, _08756_);
  and _72432_ (_21622_, _21621_, _21616_);
  and _72433_ (_21623_, _10980_, _07802_);
  or _72434_ (_21624_, _21623_, _21568_);
  and _72435_ (_21625_, _21624_, _06284_);
  or _72436_ (_21626_, _21625_, _21622_);
  and _72437_ (_21627_, _21626_, _07032_);
  or _72438_ (_21628_, _21568_, _07886_);
  and _72439_ (_21630_, _21570_, _06108_);
  and _72440_ (_21631_, _21630_, _21628_);
  or _72441_ (_21632_, _21631_, _21627_);
  and _72442_ (_21633_, _21632_, _06278_);
  and _72443_ (_21634_, _21577_, _06277_);
  and _72444_ (_21635_, _21634_, _21628_);
  or _72445_ (_21636_, _21635_, _06130_);
  or _72446_ (_21637_, _21636_, _21633_);
  and _72447_ (_21638_, _15396_, _07724_);
  or _72448_ (_21639_, _21568_, _08777_);
  or _72449_ (_21641_, _21639_, _21638_);
  and _72450_ (_21642_, _21641_, _08782_);
  and _72451_ (_21643_, _21642_, _21637_);
  nor _72452_ (_21644_, _10979_, _11359_);
  or _72453_ (_21645_, _21644_, _21568_);
  and _72454_ (_21646_, _21645_, _06292_);
  or _72455_ (_21647_, _21646_, _21643_);
  and _72456_ (_21648_, _21647_, _06718_);
  and _72457_ (_21649_, _21573_, _06316_);
  or _72458_ (_21650_, _21649_, _06047_);
  or _72459_ (_21652_, _21650_, _21648_);
  and _72460_ (_21653_, _15451_, _07724_);
  or _72461_ (_21654_, _21568_, _06048_);
  or _72462_ (_21655_, _21654_, _21653_);
  and _72463_ (_21656_, _21655_, _01336_);
  and _72464_ (_21657_, _21656_, _21652_);
  or _72465_ (_21658_, _21657_, _21567_);
  and _72466_ (_43372_, _21658_, _42882_);
  not _72467_ (_21659_, \oc8051_golden_model_1.TL1 [0]);
  nor _72468_ (_21660_, _01336_, _21659_);
  nand _72469_ (_21662_, _10995_, _07667_);
  nor _72470_ (_21663_, _07667_, _21659_);
  nor _72471_ (_21664_, _21663_, _06278_);
  nand _72472_ (_21665_, _21664_, _21662_);
  and _72473_ (_21666_, _09120_, _07667_);
  or _72474_ (_21667_, _21663_, _07012_);
  or _72475_ (_21668_, _21667_, _21666_);
  and _72476_ (_21669_, _07667_, _06931_);
  nor _72477_ (_21670_, _21669_, _21663_);
  nand _72478_ (_21671_, _21670_, _09815_);
  nor _72479_ (_21673_, _08127_, _11451_);
  or _72480_ (_21674_, _21673_, _21663_);
  or _72481_ (_21675_, _21674_, _06954_);
  and _72482_ (_21676_, _07667_, \oc8051_golden_model_1.ACC [0]);
  nor _72483_ (_21677_, _21676_, _21663_);
  nor _72484_ (_21678_, _21677_, _06939_);
  nor _72485_ (_21679_, _06938_, _21659_);
  or _72486_ (_21680_, _21679_, _06102_);
  or _72487_ (_21681_, _21680_, _21678_);
  and _72488_ (_21682_, _21681_, _06848_);
  and _72489_ (_21684_, _21682_, _21675_);
  nor _72490_ (_21685_, _21670_, _06848_);
  or _72491_ (_21686_, _21685_, _21684_);
  nand _72492_ (_21687_, _21686_, _06220_);
  or _72493_ (_21688_, _21677_, _06220_);
  and _72494_ (_21689_, _21688_, _09817_);
  nand _72495_ (_21690_, _21689_, _21687_);
  and _72496_ (_21691_, _21690_, _21671_);
  and _72497_ (_21692_, _21691_, _21668_);
  or _72498_ (_21693_, _21692_, _09833_);
  and _72499_ (_21695_, _14186_, _07667_);
  or _72500_ (_21696_, _21663_, _05669_);
  or _72501_ (_21697_, _21696_, _21695_);
  and _72502_ (_21698_, _21697_, _06020_);
  and _72503_ (_21699_, _21698_, _21693_);
  and _72504_ (_21700_, _07667_, _08672_);
  or _72505_ (_21701_, _21700_, _21663_);
  and _72506_ (_21702_, _21701_, _06019_);
  or _72507_ (_21703_, _21702_, _06112_);
  or _72508_ (_21704_, _21703_, _21699_);
  and _72509_ (_21706_, _14086_, _07667_);
  or _72510_ (_21707_, _21663_, _08751_);
  or _72511_ (_21708_, _21707_, _21706_);
  and _72512_ (_21709_, _21708_, _08756_);
  and _72513_ (_21710_, _21709_, _21704_);
  nor _72514_ (_21711_, _12302_, _11451_);
  or _72515_ (_21712_, _21711_, _21663_);
  and _72516_ (_21713_, _21662_, _06284_);
  and _72517_ (_21714_, _21713_, _21712_);
  or _72518_ (_21715_, _21714_, _21710_);
  and _72519_ (_21717_, _21715_, _07032_);
  nand _72520_ (_21718_, _21701_, _06108_);
  nor _72521_ (_21719_, _21718_, _21673_);
  or _72522_ (_21720_, _21719_, _06277_);
  or _72523_ (_21721_, _21720_, _21717_);
  and _72524_ (_21722_, _21721_, _21665_);
  or _72525_ (_21723_, _21722_, _06130_);
  and _72526_ (_21724_, _14083_, _07667_);
  or _72527_ (_21725_, _21663_, _08777_);
  or _72528_ (_21726_, _21725_, _21724_);
  and _72529_ (_21728_, _21726_, _08782_);
  and _72530_ (_21729_, _21728_, _21723_);
  and _72531_ (_21730_, _21712_, _06292_);
  or _72532_ (_21731_, _21730_, _19256_);
  or _72533_ (_21732_, _21731_, _21729_);
  or _72534_ (_21733_, _21674_, _06408_);
  and _72535_ (_21734_, _21733_, _01336_);
  and _72536_ (_21735_, _21734_, _21732_);
  or _72537_ (_21736_, _21735_, _21660_);
  and _72538_ (_43374_, _21736_, _42882_);
  not _72539_ (_21738_, \oc8051_golden_model_1.TL1 [1]);
  nor _72540_ (_21739_, _01336_, _21738_);
  or _72541_ (_21740_, _14367_, _11451_);
  or _72542_ (_21741_, _07667_, \oc8051_golden_model_1.TL1 [1]);
  and _72543_ (_21742_, _21741_, _09833_);
  and _72544_ (_21743_, _21742_, _21740_);
  and _72545_ (_21744_, _09075_, _07667_);
  nor _72546_ (_21745_, _07667_, _21738_);
  or _72547_ (_21746_, _21745_, _07012_);
  or _72548_ (_21747_, _21746_, _21744_);
  and _72549_ (_21748_, _14284_, _07667_);
  not _72550_ (_21749_, _21748_);
  and _72551_ (_21750_, _21749_, _21741_);
  or _72552_ (_21751_, _21750_, _06954_);
  and _72553_ (_21752_, _07667_, \oc8051_golden_model_1.ACC [1]);
  or _72554_ (_21753_, _21752_, _21745_);
  and _72555_ (_21754_, _21753_, _06938_);
  nor _72556_ (_21755_, _06938_, _21738_);
  or _72557_ (_21756_, _21755_, _06102_);
  or _72558_ (_21757_, _21756_, _21754_);
  and _72559_ (_21760_, _21757_, _06848_);
  and _72560_ (_21761_, _21760_, _21751_);
  nor _72561_ (_21762_, _11451_, _07132_);
  or _72562_ (_21763_, _21762_, _21745_);
  and _72563_ (_21764_, _21763_, _06239_);
  or _72564_ (_21765_, _21764_, _21761_);
  and _72565_ (_21766_, _21765_, _06220_);
  and _72566_ (_21767_, _21753_, _06219_);
  or _72567_ (_21768_, _21767_, _09818_);
  or _72568_ (_21769_, _21768_, _21766_);
  or _72569_ (_21771_, _21763_, _09827_);
  and _72570_ (_21772_, _21771_, _05669_);
  and _72571_ (_21773_, _21772_, _21769_);
  and _72572_ (_21774_, _21773_, _21747_);
  or _72573_ (_21775_, _21774_, _21743_);
  and _72574_ (_21776_, _21775_, _06020_);
  nand _72575_ (_21777_, _07667_, _06832_);
  and _72576_ (_21778_, _21741_, _06019_);
  and _72577_ (_21779_, _21778_, _21777_);
  or _72578_ (_21780_, _21779_, _21776_);
  and _72579_ (_21782_, _21780_, _08751_);
  or _72580_ (_21783_, _14263_, _11451_);
  and _72581_ (_21784_, _21741_, _06112_);
  and _72582_ (_21785_, _21784_, _21783_);
  or _72583_ (_21786_, _21785_, _06284_);
  or _72584_ (_21787_, _21786_, _21782_);
  nor _72585_ (_21788_, _10993_, _11451_);
  or _72586_ (_21789_, _21788_, _21745_);
  nand _72587_ (_21790_, _10992_, _07667_);
  and _72588_ (_21791_, _21790_, _21789_);
  or _72589_ (_21793_, _21791_, _08756_);
  and _72590_ (_21794_, _21793_, _07032_);
  and _72591_ (_21795_, _21794_, _21787_);
  or _72592_ (_21796_, _14261_, _11451_);
  and _72593_ (_21797_, _21741_, _06108_);
  and _72594_ (_21798_, _21797_, _21796_);
  or _72595_ (_21799_, _21798_, _06277_);
  or _72596_ (_21800_, _21799_, _21795_);
  nor _72597_ (_21801_, _21745_, _06278_);
  nand _72598_ (_21802_, _21801_, _21790_);
  and _72599_ (_21804_, _21802_, _08777_);
  and _72600_ (_21805_, _21804_, _21800_);
  or _72601_ (_21806_, _21777_, _08078_);
  and _72602_ (_21807_, _21741_, _06130_);
  and _72603_ (_21808_, _21807_, _21806_);
  or _72604_ (_21809_, _21808_, _06292_);
  or _72605_ (_21810_, _21809_, _21805_);
  or _72606_ (_21811_, _21789_, _08782_);
  and _72607_ (_21812_, _21811_, _06718_);
  and _72608_ (_21813_, _21812_, _21810_);
  and _72609_ (_21815_, _21750_, _06316_);
  or _72610_ (_21816_, _21815_, _06047_);
  or _72611_ (_21817_, _21816_, _21813_);
  or _72612_ (_21818_, _21745_, _06048_);
  or _72613_ (_21819_, _21818_, _21748_);
  and _72614_ (_21820_, _21819_, _01336_);
  and _72615_ (_21821_, _21820_, _21817_);
  or _72616_ (_21822_, _21821_, _21739_);
  and _72617_ (_43375_, _21822_, _42882_);
  not _72618_ (_21823_, \oc8051_golden_model_1.TL1 [2]);
  nor _72619_ (_21825_, _01336_, _21823_);
  and _72620_ (_21826_, _09182_, _07667_);
  nor _72621_ (_21827_, _07667_, _21823_);
  or _72622_ (_21828_, _21827_, _07012_);
  or _72623_ (_21829_, _21828_, _21826_);
  nor _72624_ (_21830_, _11451_, _07530_);
  nor _72625_ (_21831_, _21830_, _21827_);
  nand _72626_ (_21832_, _21831_, _09815_);
  and _72627_ (_21833_, _14493_, _07667_);
  or _72628_ (_21834_, _21833_, _21827_);
  and _72629_ (_21836_, _21834_, _06102_);
  nor _72630_ (_21837_, _06938_, _21823_);
  and _72631_ (_21838_, _07667_, \oc8051_golden_model_1.ACC [2]);
  nor _72632_ (_21839_, _21838_, _21827_);
  nor _72633_ (_21840_, _21839_, _06939_);
  or _72634_ (_21841_, _21840_, _21837_);
  and _72635_ (_21842_, _21841_, _06954_);
  or _72636_ (_21843_, _21842_, _06239_);
  or _72637_ (_21844_, _21843_, _21836_);
  nand _72638_ (_21845_, _21831_, _06239_);
  and _72639_ (_21847_, _21845_, _06220_);
  nand _72640_ (_21848_, _21847_, _21844_);
  or _72641_ (_21849_, _21839_, _06220_);
  and _72642_ (_21850_, _21849_, _09817_);
  nand _72643_ (_21851_, _21850_, _21848_);
  and _72644_ (_21852_, _21851_, _21832_);
  and _72645_ (_21853_, _21852_, _21829_);
  or _72646_ (_21854_, _21853_, _09833_);
  and _72647_ (_21855_, _14580_, _07667_);
  or _72648_ (_21856_, _21855_, _21827_);
  or _72649_ (_21857_, _21856_, _05669_);
  and _72650_ (_21858_, _21857_, _06020_);
  and _72651_ (_21859_, _21858_, _21854_);
  and _72652_ (_21860_, _07667_, _08730_);
  or _72653_ (_21861_, _21860_, _21827_);
  and _72654_ (_21862_, _21861_, _06019_);
  or _72655_ (_21863_, _21862_, _06112_);
  or _72656_ (_21864_, _21863_, _21859_);
  and _72657_ (_21865_, _14596_, _07667_);
  or _72658_ (_21866_, _21827_, _08751_);
  or _72659_ (_21869_, _21866_, _21865_);
  and _72660_ (_21870_, _21869_, _08756_);
  and _72661_ (_21871_, _21870_, _21864_);
  and _72662_ (_21872_, _10991_, _07667_);
  or _72663_ (_21873_, _21872_, _21827_);
  and _72664_ (_21874_, _21873_, _06284_);
  or _72665_ (_21875_, _21874_, _21871_);
  and _72666_ (_21876_, _21875_, _07032_);
  or _72667_ (_21877_, _21827_, _08177_);
  and _72668_ (_21878_, _21861_, _06108_);
  and _72669_ (_21880_, _21878_, _21877_);
  or _72670_ (_21881_, _21880_, _21876_);
  and _72671_ (_21882_, _21881_, _06278_);
  nor _72672_ (_21883_, _21839_, _06278_);
  and _72673_ (_21884_, _21883_, _21877_);
  or _72674_ (_21885_, _21884_, _06130_);
  or _72675_ (_21886_, _21885_, _21882_);
  and _72676_ (_21887_, _14593_, _07667_);
  or _72677_ (_21888_, _21827_, _08777_);
  or _72678_ (_21889_, _21888_, _21887_);
  and _72679_ (_21891_, _21889_, _08782_);
  and _72680_ (_21892_, _21891_, _21886_);
  nor _72681_ (_21893_, _10990_, _11451_);
  or _72682_ (_21894_, _21893_, _21827_);
  and _72683_ (_21895_, _21894_, _06292_);
  or _72684_ (_21896_, _21895_, _21892_);
  and _72685_ (_21897_, _21896_, _06718_);
  and _72686_ (_21898_, _21834_, _06316_);
  or _72687_ (_21899_, _21898_, _06047_);
  or _72688_ (_21900_, _21899_, _21897_);
  and _72689_ (_21902_, _14657_, _07667_);
  or _72690_ (_21903_, _21827_, _06048_);
  or _72691_ (_21904_, _21903_, _21902_);
  and _72692_ (_21905_, _21904_, _01336_);
  and _72693_ (_21906_, _21905_, _21900_);
  or _72694_ (_21907_, _21906_, _21825_);
  and _72695_ (_43376_, _21907_, _42882_);
  not _72696_ (_21908_, \oc8051_golden_model_1.TL1 [3]);
  nor _72697_ (_21909_, _01336_, _21908_);
  and _72698_ (_21910_, _09181_, _07667_);
  nor _72699_ (_21912_, _07667_, _21908_);
  or _72700_ (_21913_, _21912_, _07012_);
  or _72701_ (_21914_, _21913_, _21910_);
  nor _72702_ (_21915_, _11451_, _07353_);
  nor _72703_ (_21916_, _21915_, _21912_);
  nand _72704_ (_21917_, _21916_, _09815_);
  and _72705_ (_21918_, _14672_, _07667_);
  or _72706_ (_21919_, _21918_, _21912_);
  or _72707_ (_21920_, _21919_, _06954_);
  and _72708_ (_21921_, _07667_, \oc8051_golden_model_1.ACC [3]);
  nor _72709_ (_21923_, _21921_, _21912_);
  nor _72710_ (_21924_, _21923_, _06939_);
  nor _72711_ (_21925_, _06938_, _21908_);
  or _72712_ (_21926_, _21925_, _06102_);
  or _72713_ (_21927_, _21926_, _21924_);
  and _72714_ (_21928_, _21927_, _06848_);
  and _72715_ (_21929_, _21928_, _21920_);
  nor _72716_ (_21930_, _21916_, _06848_);
  or _72717_ (_21931_, _21930_, _21929_);
  nand _72718_ (_21932_, _21931_, _06220_);
  or _72719_ (_21934_, _21923_, _06220_);
  and _72720_ (_21935_, _21934_, _09817_);
  nand _72721_ (_21936_, _21935_, _21932_);
  and _72722_ (_21937_, _21936_, _21917_);
  and _72723_ (_21938_, _21937_, _21914_);
  or _72724_ (_21939_, _21938_, _09833_);
  and _72725_ (_21940_, _14778_, _07667_);
  or _72726_ (_21941_, _21912_, _05669_);
  or _72727_ (_21942_, _21941_, _21940_);
  and _72728_ (_21943_, _21942_, _06020_);
  and _72729_ (_21945_, _21943_, _21939_);
  and _72730_ (_21946_, _07667_, _08662_);
  or _72731_ (_21947_, _21946_, _21912_);
  and _72732_ (_21948_, _21947_, _06019_);
  or _72733_ (_21949_, _21948_, _06112_);
  or _72734_ (_21950_, _21949_, _21945_);
  and _72735_ (_21951_, _14793_, _07667_);
  or _72736_ (_21952_, _21912_, _08751_);
  or _72737_ (_21953_, _21952_, _21951_);
  and _72738_ (_21954_, _21953_, _08756_);
  and _72739_ (_21956_, _21954_, _21950_);
  and _72740_ (_21957_, _12299_, _07667_);
  or _72741_ (_21958_, _21957_, _21912_);
  and _72742_ (_21959_, _21958_, _06284_);
  or _72743_ (_21960_, _21959_, _21956_);
  and _72744_ (_21961_, _21960_, _07032_);
  or _72745_ (_21962_, _21912_, _08029_);
  and _72746_ (_21963_, _21947_, _06108_);
  and _72747_ (_21964_, _21963_, _21962_);
  or _72748_ (_21965_, _21964_, _21961_);
  and _72749_ (_21967_, _21965_, _06278_);
  nor _72750_ (_21968_, _21923_, _06278_);
  and _72751_ (_21969_, _21968_, _21962_);
  or _72752_ (_21970_, _21969_, _06130_);
  or _72753_ (_21971_, _21970_, _21967_);
  and _72754_ (_21972_, _14792_, _07667_);
  or _72755_ (_21973_, _21912_, _08777_);
  or _72756_ (_21974_, _21973_, _21972_);
  and _72757_ (_21975_, _21974_, _08782_);
  and _72758_ (_21976_, _21975_, _21971_);
  nor _72759_ (_21978_, _10988_, _11451_);
  or _72760_ (_21979_, _21978_, _21912_);
  and _72761_ (_21980_, _21979_, _06292_);
  or _72762_ (_21981_, _21980_, _21976_);
  and _72763_ (_21982_, _21981_, _06718_);
  and _72764_ (_21983_, _21919_, _06316_);
  or _72765_ (_21984_, _21983_, _06047_);
  or _72766_ (_21985_, _21984_, _21982_);
  and _72767_ (_21986_, _14849_, _07667_);
  or _72768_ (_21987_, _21912_, _06048_);
  or _72769_ (_21989_, _21987_, _21986_);
  and _72770_ (_21990_, _21989_, _01336_);
  and _72771_ (_21991_, _21990_, _21985_);
  or _72772_ (_21992_, _21991_, _21909_);
  and _72773_ (_43377_, _21992_, _42882_);
  and _72774_ (_21993_, _01340_, \oc8051_golden_model_1.TL1 [4]);
  and _72775_ (_21994_, _11451_, \oc8051_golden_model_1.TL1 [4]);
  and _72776_ (_21995_, _08665_, _07667_);
  or _72777_ (_21996_, _21995_, _21994_);
  or _72778_ (_21997_, _21996_, _06020_);
  and _72779_ (_21999_, _14887_, _07667_);
  or _72780_ (_22000_, _21999_, _21994_);
  or _72781_ (_22001_, _22000_, _06954_);
  and _72782_ (_22002_, _07667_, \oc8051_golden_model_1.ACC [4]);
  or _72783_ (_22003_, _22002_, _21994_);
  and _72784_ (_22004_, _22003_, _06938_);
  and _72785_ (_22005_, _06939_, \oc8051_golden_model_1.TL1 [4]);
  or _72786_ (_22006_, _22005_, _06102_);
  or _72787_ (_22007_, _22006_, _22004_);
  and _72788_ (_22008_, _22007_, _06848_);
  and _72789_ (_22010_, _22008_, _22001_);
  nor _72790_ (_22011_, _08270_, _11451_);
  or _72791_ (_22012_, _22011_, _21994_);
  and _72792_ (_22013_, _22012_, _06239_);
  or _72793_ (_22014_, _22013_, _22010_);
  and _72794_ (_22015_, _22014_, _06220_);
  and _72795_ (_22016_, _22003_, _06219_);
  or _72796_ (_22017_, _22016_, _09818_);
  or _72797_ (_22018_, _22017_, _22015_);
  and _72798_ (_22019_, _09180_, _07667_);
  or _72799_ (_22021_, _21994_, _07012_);
  or _72800_ (_22022_, _22021_, _22019_);
  or _72801_ (_22023_, _22012_, _09827_);
  and _72802_ (_22024_, _22023_, _05669_);
  and _72803_ (_22025_, _22024_, _22022_);
  and _72804_ (_22026_, _22025_, _22018_);
  and _72805_ (_22027_, _14983_, _07667_);
  or _72806_ (_22028_, _22027_, _21994_);
  and _72807_ (_22029_, _22028_, _09833_);
  or _72808_ (_22030_, _22029_, _06019_);
  or _72809_ (_22032_, _22030_, _22026_);
  and _72810_ (_22033_, _22032_, _21997_);
  or _72811_ (_22034_, _22033_, _06112_);
  and _72812_ (_22035_, _14876_, _07667_);
  or _72813_ (_22036_, _21994_, _08751_);
  or _72814_ (_22037_, _22036_, _22035_);
  and _72815_ (_22038_, _22037_, _08756_);
  and _72816_ (_22039_, _22038_, _22034_);
  and _72817_ (_22040_, _10986_, _07667_);
  or _72818_ (_22041_, _22040_, _21994_);
  and _72819_ (_22043_, _22041_, _06284_);
  or _72820_ (_22044_, _22043_, _22039_);
  and _72821_ (_22045_, _22044_, _07032_);
  or _72822_ (_22046_, _21994_, _08273_);
  and _72823_ (_22047_, _21996_, _06108_);
  and _72824_ (_22048_, _22047_, _22046_);
  or _72825_ (_22049_, _22048_, _22045_);
  and _72826_ (_22050_, _22049_, _06278_);
  and _72827_ (_22051_, _22003_, _06277_);
  and _72828_ (_22052_, _22051_, _22046_);
  or _72829_ (_22054_, _22052_, _06130_);
  or _72830_ (_22055_, _22054_, _22050_);
  and _72831_ (_22056_, _14873_, _07667_);
  or _72832_ (_22057_, _21994_, _08777_);
  or _72833_ (_22058_, _22057_, _22056_);
  and _72834_ (_22059_, _22058_, _08782_);
  and _72835_ (_22060_, _22059_, _22055_);
  nor _72836_ (_22061_, _10985_, _11451_);
  or _72837_ (_22062_, _22061_, _21994_);
  and _72838_ (_22063_, _22062_, _06292_);
  or _72839_ (_22065_, _22063_, _22060_);
  and _72840_ (_22066_, _22065_, _06718_);
  and _72841_ (_22067_, _22000_, _06316_);
  or _72842_ (_22068_, _22067_, _06047_);
  or _72843_ (_22069_, _22068_, _22066_);
  and _72844_ (_22070_, _15055_, _07667_);
  or _72845_ (_22071_, _21994_, _06048_);
  or _72846_ (_22072_, _22071_, _22070_);
  and _72847_ (_22073_, _22072_, _01336_);
  and _72848_ (_22074_, _22073_, _22069_);
  or _72849_ (_22076_, _22074_, _21993_);
  and _72850_ (_43378_, _22076_, _42882_);
  and _72851_ (_22077_, _01340_, \oc8051_golden_model_1.TL1 [5]);
  and _72852_ (_22078_, _11451_, \oc8051_golden_model_1.TL1 [5]);
  and _72853_ (_22079_, _08652_, _07667_);
  or _72854_ (_22080_, _22079_, _22078_);
  or _72855_ (_22081_, _22080_, _06020_);
  and _72856_ (_22082_, _15093_, _07667_);
  or _72857_ (_22083_, _22082_, _22078_);
  or _72858_ (_22084_, _22083_, _06954_);
  and _72859_ (_22086_, _07667_, \oc8051_golden_model_1.ACC [5]);
  or _72860_ (_22087_, _22086_, _22078_);
  and _72861_ (_22088_, _22087_, _06938_);
  and _72862_ (_22089_, _06939_, \oc8051_golden_model_1.TL1 [5]);
  or _72863_ (_22090_, _22089_, _06102_);
  or _72864_ (_22091_, _22090_, _22088_);
  and _72865_ (_22092_, _22091_, _06848_);
  and _72866_ (_22093_, _22092_, _22084_);
  nor _72867_ (_22094_, _07977_, _11451_);
  or _72868_ (_22095_, _22094_, _22078_);
  and _72869_ (_22097_, _22095_, _06239_);
  or _72870_ (_22098_, _22097_, _22093_);
  and _72871_ (_22099_, _22098_, _06220_);
  and _72872_ (_22100_, _22087_, _06219_);
  or _72873_ (_22101_, _22100_, _09818_);
  or _72874_ (_22102_, _22101_, _22099_);
  and _72875_ (_22103_, _09179_, _07667_);
  or _72876_ (_22104_, _22078_, _07012_);
  or _72877_ (_22105_, _22104_, _22103_);
  or _72878_ (_22106_, _22095_, _09827_);
  and _72879_ (_22108_, _22106_, _05669_);
  and _72880_ (_22109_, _22108_, _22105_);
  and _72881_ (_22110_, _22109_, _22102_);
  and _72882_ (_22111_, _15179_, _07667_);
  or _72883_ (_22112_, _22111_, _22078_);
  and _72884_ (_22113_, _22112_, _09833_);
  or _72885_ (_22114_, _22113_, _06019_);
  or _72886_ (_22115_, _22114_, _22110_);
  and _72887_ (_22116_, _22115_, _22081_);
  or _72888_ (_22117_, _22116_, _06112_);
  and _72889_ (_22119_, _15195_, _07667_);
  or _72890_ (_22120_, _22119_, _22078_);
  or _72891_ (_22121_, _22120_, _08751_);
  and _72892_ (_22122_, _22121_, _08756_);
  and _72893_ (_22123_, _22122_, _22117_);
  and _72894_ (_22124_, _12306_, _07667_);
  or _72895_ (_22125_, _22124_, _22078_);
  and _72896_ (_22126_, _22125_, _06284_);
  or _72897_ (_22127_, _22126_, _22123_);
  and _72898_ (_22128_, _22127_, _07032_);
  or _72899_ (_22130_, _22078_, _07980_);
  and _72900_ (_22131_, _22080_, _06108_);
  and _72901_ (_22132_, _22131_, _22130_);
  or _72902_ (_22133_, _22132_, _22128_);
  and _72903_ (_22134_, _22133_, _06278_);
  and _72904_ (_22135_, _22087_, _06277_);
  and _72905_ (_22136_, _22135_, _22130_);
  or _72906_ (_22137_, _22136_, _06130_);
  or _72907_ (_22138_, _22137_, _22134_);
  and _72908_ (_22139_, _15194_, _07667_);
  or _72909_ (_22141_, _22078_, _08777_);
  or _72910_ (_22142_, _22141_, _22139_);
  and _72911_ (_22143_, _22142_, _08782_);
  and _72912_ (_22144_, _22143_, _22138_);
  nor _72913_ (_22145_, _10982_, _11451_);
  or _72914_ (_22146_, _22145_, _22078_);
  and _72915_ (_22147_, _22146_, _06292_);
  or _72916_ (_22148_, _22147_, _22144_);
  and _72917_ (_22149_, _22148_, _06718_);
  and _72918_ (_22150_, _22083_, _06316_);
  or _72919_ (_22152_, _22150_, _06047_);
  or _72920_ (_22153_, _22152_, _22149_);
  and _72921_ (_22154_, _15253_, _07667_);
  or _72922_ (_22155_, _22078_, _06048_);
  or _72923_ (_22156_, _22155_, _22154_);
  and _72924_ (_22157_, _22156_, _01336_);
  and _72925_ (_22158_, _22157_, _22153_);
  or _72926_ (_22159_, _22158_, _22077_);
  and _72927_ (_43380_, _22159_, _42882_);
  and _72928_ (_22160_, _01340_, \oc8051_golden_model_1.TL1 [6]);
  and _72929_ (_22162_, _11451_, \oc8051_golden_model_1.TL1 [6]);
  and _72930_ (_22163_, _15389_, _07667_);
  or _72931_ (_22164_, _22163_, _22162_);
  or _72932_ (_22165_, _22164_, _06020_);
  and _72933_ (_22166_, _15293_, _07667_);
  or _72934_ (_22167_, _22166_, _22162_);
  or _72935_ (_22168_, _22167_, _06954_);
  and _72936_ (_22169_, _07667_, \oc8051_golden_model_1.ACC [6]);
  or _72937_ (_22170_, _22169_, _22162_);
  and _72938_ (_22171_, _22170_, _06938_);
  and _72939_ (_22173_, _06939_, \oc8051_golden_model_1.TL1 [6]);
  or _72940_ (_22174_, _22173_, _06102_);
  or _72941_ (_22175_, _22174_, _22171_);
  and _72942_ (_22176_, _22175_, _06848_);
  and _72943_ (_22177_, _22176_, _22168_);
  nor _72944_ (_22178_, _07883_, _11451_);
  or _72945_ (_22179_, _22178_, _22162_);
  and _72946_ (_22180_, _22179_, _06239_);
  or _72947_ (_22181_, _22180_, _22177_);
  and _72948_ (_22182_, _22181_, _06220_);
  and _72949_ (_22184_, _22170_, _06219_);
  or _72950_ (_22185_, _22184_, _09818_);
  or _72951_ (_22186_, _22185_, _22182_);
  and _72952_ (_22187_, _09178_, _07667_);
  or _72953_ (_22188_, _22162_, _07012_);
  or _72954_ (_22189_, _22188_, _22187_);
  or _72955_ (_22190_, _22179_, _09827_);
  and _72956_ (_22191_, _22190_, _05669_);
  and _72957_ (_22192_, _22191_, _22189_);
  and _72958_ (_22193_, _22192_, _22186_);
  and _72959_ (_22195_, _15382_, _07667_);
  or _72960_ (_22196_, _22195_, _22162_);
  and _72961_ (_22197_, _22196_, _09833_);
  or _72962_ (_22198_, _22197_, _06019_);
  or _72963_ (_22199_, _22198_, _22193_);
  and _72964_ (_22200_, _22199_, _22165_);
  or _72965_ (_22201_, _22200_, _06112_);
  and _72966_ (_22202_, _15399_, _07667_);
  or _72967_ (_22203_, _22162_, _08751_);
  or _72968_ (_22204_, _22203_, _22202_);
  and _72969_ (_22206_, _22204_, _08756_);
  and _72970_ (_22207_, _22206_, _22201_);
  and _72971_ (_22208_, _10980_, _07667_);
  or _72972_ (_22209_, _22208_, _22162_);
  and _72973_ (_22210_, _22209_, _06284_);
  or _72974_ (_22211_, _22210_, _22207_);
  and _72975_ (_22212_, _22211_, _07032_);
  or _72976_ (_22213_, _22162_, _07886_);
  and _72977_ (_22214_, _22164_, _06108_);
  and _72978_ (_22215_, _22214_, _22213_);
  or _72979_ (_22218_, _22215_, _22212_);
  and _72980_ (_22219_, _22218_, _06278_);
  and _72981_ (_22220_, _22170_, _06277_);
  and _72982_ (_22221_, _22220_, _22213_);
  or _72983_ (_22222_, _22221_, _06130_);
  or _72984_ (_22223_, _22222_, _22219_);
  and _72985_ (_22224_, _15396_, _07667_);
  or _72986_ (_22225_, _22162_, _08777_);
  or _72987_ (_22226_, _22225_, _22224_);
  and _72988_ (_22227_, _22226_, _08782_);
  and _72989_ (_22229_, _22227_, _22223_);
  nor _72990_ (_22230_, _10979_, _11451_);
  or _72991_ (_22231_, _22230_, _22162_);
  and _72992_ (_22232_, _22231_, _06292_);
  or _72993_ (_22233_, _22232_, _22229_);
  and _72994_ (_22234_, _22233_, _06718_);
  and _72995_ (_22235_, _22167_, _06316_);
  or _72996_ (_22236_, _22235_, _06047_);
  or _72997_ (_22237_, _22236_, _22234_);
  and _72998_ (_22238_, _15451_, _07667_);
  or _72999_ (_22240_, _22162_, _06048_);
  or _73000_ (_22241_, _22240_, _22238_);
  and _73001_ (_22242_, _22241_, _01336_);
  and _73002_ (_22243_, _22242_, _22237_);
  or _73003_ (_22244_, _22243_, _22160_);
  and _73004_ (_43381_, _22244_, _42882_);
  not _73005_ (_22245_, \oc8051_golden_model_1.TL0 [0]);
  nor _73006_ (_22246_, _01336_, _22245_);
  nand _73007_ (_22247_, _10995_, _07659_);
  nor _73008_ (_22248_, _07659_, _22245_);
  nor _73009_ (_22250_, _22248_, _06278_);
  nand _73010_ (_22251_, _22250_, _22247_);
  and _73011_ (_22252_, _09120_, _07659_);
  or _73012_ (_22253_, _22248_, _07012_);
  or _73013_ (_22254_, _22253_, _22252_);
  and _73014_ (_22255_, _07659_, _06931_);
  nor _73015_ (_22256_, _22255_, _22248_);
  nand _73016_ (_22257_, _22256_, _09815_);
  nor _73017_ (_22258_, _08127_, _11528_);
  or _73018_ (_22259_, _22258_, _22248_);
  and _73019_ (_22261_, _22259_, _06102_);
  nor _73020_ (_22262_, _06938_, _22245_);
  and _73021_ (_22263_, _07659_, \oc8051_golden_model_1.ACC [0]);
  nor _73022_ (_22264_, _22263_, _22248_);
  nor _73023_ (_22265_, _22264_, _06939_);
  or _73024_ (_22266_, _22265_, _22262_);
  and _73025_ (_22267_, _22266_, _06954_);
  or _73026_ (_22268_, _22267_, _06239_);
  or _73027_ (_22269_, _22268_, _22261_);
  nand _73028_ (_22270_, _22256_, _06239_);
  and _73029_ (_22272_, _22270_, _06220_);
  nand _73030_ (_22273_, _22272_, _22269_);
  or _73031_ (_22274_, _22264_, _06220_);
  and _73032_ (_22275_, _22274_, _09817_);
  nand _73033_ (_22276_, _22275_, _22273_);
  and _73034_ (_22277_, _22276_, _22257_);
  and _73035_ (_22278_, _22277_, _22254_);
  or _73036_ (_22279_, _22278_, _09833_);
  and _73037_ (_22280_, _14186_, _07659_);
  or _73038_ (_22281_, _22248_, _05669_);
  or _73039_ (_22283_, _22281_, _22280_);
  and _73040_ (_22284_, _22283_, _06020_);
  and _73041_ (_22285_, _22284_, _22279_);
  and _73042_ (_22286_, _07659_, _08672_);
  or _73043_ (_22287_, _22286_, _22248_);
  and _73044_ (_22288_, _22287_, _06019_);
  or _73045_ (_22289_, _22288_, _06112_);
  or _73046_ (_22290_, _22289_, _22285_);
  and _73047_ (_22291_, _14086_, _07659_);
  or _73048_ (_22292_, _22291_, _22248_);
  or _73049_ (_22294_, _22292_, _08751_);
  and _73050_ (_22295_, _22294_, _08756_);
  and _73051_ (_22296_, _22295_, _22290_);
  nor _73052_ (_22297_, _12302_, _11528_);
  or _73053_ (_22298_, _22297_, _22248_);
  and _73054_ (_22299_, _22247_, _06284_);
  and _73055_ (_22300_, _22299_, _22298_);
  or _73056_ (_22301_, _22300_, _22296_);
  and _73057_ (_22302_, _22301_, _07032_);
  nand _73058_ (_22303_, _22287_, _06108_);
  nor _73059_ (_22304_, _22303_, _22258_);
  or _73060_ (_22305_, _22304_, _06277_);
  or _73061_ (_22306_, _22305_, _22302_);
  and _73062_ (_22307_, _22306_, _22251_);
  or _73063_ (_22308_, _22307_, _06130_);
  and _73064_ (_22309_, _14083_, _07659_);
  or _73065_ (_22310_, _22248_, _08777_);
  or _73066_ (_22311_, _22310_, _22309_);
  and _73067_ (_22312_, _22311_, _08782_);
  and _73068_ (_22313_, _22312_, _22308_);
  and _73069_ (_22316_, _22298_, _06292_);
  or _73070_ (_22317_, _22316_, _19256_);
  or _73071_ (_22318_, _22317_, _22313_);
  or _73072_ (_22319_, _22259_, _06408_);
  and _73073_ (_22320_, _22319_, _01336_);
  and _73074_ (_22321_, _22320_, _22318_);
  or _73075_ (_22322_, _22321_, _22246_);
  and _73076_ (_43382_, _22322_, _42882_);
  not _73077_ (_22323_, \oc8051_golden_model_1.TL0 [1]);
  nor _73078_ (_22324_, _01336_, _22323_);
  or _73079_ (_22326_, _14367_, _11528_);
  or _73080_ (_22327_, _07659_, \oc8051_golden_model_1.TL0 [1]);
  and _73081_ (_22328_, _22327_, _09833_);
  and _73082_ (_22329_, _22328_, _22326_);
  and _73083_ (_22330_, _09075_, _07659_);
  nor _73084_ (_22331_, _07659_, _22323_);
  or _73085_ (_22332_, _22331_, _07012_);
  or _73086_ (_22333_, _22332_, _22330_);
  and _73087_ (_22334_, _14284_, _07659_);
  not _73088_ (_22335_, _22334_);
  and _73089_ (_22337_, _22335_, _22327_);
  and _73090_ (_22338_, _22337_, _06102_);
  nor _73091_ (_22339_, _06938_, _22323_);
  and _73092_ (_22340_, _07659_, \oc8051_golden_model_1.ACC [1]);
  or _73093_ (_22341_, _22340_, _22331_);
  and _73094_ (_22342_, _22341_, _06938_);
  or _73095_ (_22343_, _22342_, _22339_);
  and _73096_ (_22344_, _22343_, _06954_);
  or _73097_ (_22345_, _22344_, _06239_);
  or _73098_ (_22346_, _22345_, _22338_);
  nor _73099_ (_22348_, _11528_, _07132_);
  or _73100_ (_22349_, _22348_, _22331_);
  or _73101_ (_22350_, _22349_, _06848_);
  and _73102_ (_22351_, _22350_, _06220_);
  and _73103_ (_22352_, _22351_, _22346_);
  and _73104_ (_22353_, _22341_, _06219_);
  or _73105_ (_22354_, _22353_, _09818_);
  or _73106_ (_22355_, _22354_, _22352_);
  or _73107_ (_22356_, _22349_, _09827_);
  and _73108_ (_22357_, _22356_, _05669_);
  and _73109_ (_22359_, _22357_, _22355_);
  and _73110_ (_22360_, _22359_, _22333_);
  or _73111_ (_22361_, _22360_, _22329_);
  and _73112_ (_22362_, _22361_, _06020_);
  nand _73113_ (_22363_, _07659_, _06832_);
  and _73114_ (_22364_, _22327_, _06019_);
  and _73115_ (_22365_, _22364_, _22363_);
  or _73116_ (_22366_, _22365_, _22362_);
  and _73117_ (_22367_, _22366_, _08751_);
  or _73118_ (_22368_, _14263_, _11528_);
  and _73119_ (_22370_, _22327_, _06112_);
  and _73120_ (_22371_, _22370_, _22368_);
  or _73121_ (_22372_, _22371_, _06284_);
  or _73122_ (_22373_, _22372_, _22367_);
  nor _73123_ (_22374_, _10993_, _11528_);
  or _73124_ (_22375_, _22374_, _22331_);
  nand _73125_ (_22376_, _10992_, _07659_);
  and _73126_ (_22377_, _22376_, _22375_);
  or _73127_ (_22378_, _22377_, _08756_);
  and _73128_ (_22379_, _22378_, _07032_);
  and _73129_ (_22381_, _22379_, _22373_);
  or _73130_ (_22382_, _14261_, _11528_);
  and _73131_ (_22383_, _22327_, _06108_);
  and _73132_ (_22384_, _22383_, _22382_);
  or _73133_ (_22385_, _22384_, _06277_);
  or _73134_ (_22386_, _22385_, _22381_);
  nor _73135_ (_22387_, _22331_, _06278_);
  nand _73136_ (_22388_, _22387_, _22376_);
  and _73137_ (_22389_, _22388_, _08777_);
  and _73138_ (_22390_, _22389_, _22386_);
  or _73139_ (_22392_, _22363_, _08078_);
  and _73140_ (_22393_, _22327_, _06130_);
  and _73141_ (_22394_, _22393_, _22392_);
  or _73142_ (_22395_, _22394_, _06292_);
  or _73143_ (_22396_, _22395_, _22390_);
  or _73144_ (_22397_, _22375_, _08782_);
  and _73145_ (_22398_, _22397_, _06718_);
  and _73146_ (_22399_, _22398_, _22396_);
  and _73147_ (_22400_, _22337_, _06316_);
  or _73148_ (_22401_, _22400_, _06047_);
  or _73149_ (_22403_, _22401_, _22399_);
  or _73150_ (_22404_, _22331_, _06048_);
  or _73151_ (_22405_, _22404_, _22334_);
  and _73152_ (_22406_, _22405_, _01336_);
  and _73153_ (_22407_, _22406_, _22403_);
  or _73154_ (_22408_, _22407_, _22324_);
  and _73155_ (_43384_, _22408_, _42882_);
  not _73156_ (_22409_, \oc8051_golden_model_1.TL0 [2]);
  nor _73157_ (_22410_, _01336_, _22409_);
  and _73158_ (_22411_, _09182_, _07659_);
  nor _73159_ (_22413_, _07659_, _22409_);
  or _73160_ (_22414_, _22413_, _07012_);
  or _73161_ (_22415_, _22414_, _22411_);
  nor _73162_ (_22416_, _11528_, _07530_);
  nor _73163_ (_22417_, _22416_, _22413_);
  nand _73164_ (_22418_, _22417_, _09815_);
  and _73165_ (_22419_, _14493_, _07659_);
  or _73166_ (_22420_, _22419_, _22413_);
  and _73167_ (_22421_, _22420_, _06102_);
  nor _73168_ (_22422_, _06938_, _22409_);
  and _73169_ (_22424_, _07659_, \oc8051_golden_model_1.ACC [2]);
  nor _73170_ (_22425_, _22424_, _22413_);
  nor _73171_ (_22426_, _22425_, _06939_);
  or _73172_ (_22427_, _22426_, _22422_);
  and _73173_ (_22428_, _22427_, _06954_);
  or _73174_ (_22429_, _22428_, _06239_);
  or _73175_ (_22430_, _22429_, _22421_);
  nand _73176_ (_22431_, _22417_, _06239_);
  and _73177_ (_22432_, _22431_, _06220_);
  nand _73178_ (_22433_, _22432_, _22430_);
  or _73179_ (_22435_, _22425_, _06220_);
  and _73180_ (_22436_, _22435_, _09817_);
  nand _73181_ (_22437_, _22436_, _22433_);
  and _73182_ (_22438_, _22437_, _22418_);
  and _73183_ (_22439_, _22438_, _22415_);
  or _73184_ (_22440_, _22439_, _09833_);
  and _73185_ (_22441_, _14580_, _07659_);
  or _73186_ (_22442_, _22441_, _22413_);
  or _73187_ (_22443_, _22442_, _05669_);
  and _73188_ (_22444_, _22443_, _06020_);
  and _73189_ (_22446_, _22444_, _22440_);
  and _73190_ (_22447_, _07659_, _08730_);
  or _73191_ (_22448_, _22447_, _22413_);
  and _73192_ (_22449_, _22448_, _06019_);
  or _73193_ (_22450_, _22449_, _06112_);
  or _73194_ (_22451_, _22450_, _22446_);
  and _73195_ (_22452_, _14596_, _07659_);
  or _73196_ (_22453_, _22413_, _08751_);
  or _73197_ (_22454_, _22453_, _22452_);
  and _73198_ (_22455_, _22454_, _08756_);
  and _73199_ (_22457_, _22455_, _22451_);
  and _73200_ (_22458_, _10991_, _07659_);
  or _73201_ (_22459_, _22458_, _22413_);
  and _73202_ (_22460_, _22459_, _06284_);
  or _73203_ (_22461_, _22460_, _22457_);
  and _73204_ (_22462_, _22461_, _07032_);
  or _73205_ (_22463_, _22413_, _08177_);
  and _73206_ (_22464_, _22448_, _06108_);
  and _73207_ (_22465_, _22464_, _22463_);
  or _73208_ (_22466_, _22465_, _22462_);
  and _73209_ (_22468_, _22466_, _06278_);
  nor _73210_ (_22469_, _22425_, _06278_);
  and _73211_ (_22470_, _22469_, _22463_);
  or _73212_ (_22471_, _22470_, _06130_);
  or _73213_ (_22472_, _22471_, _22468_);
  and _73214_ (_22473_, _14593_, _07659_);
  or _73215_ (_22474_, _22413_, _08777_);
  or _73216_ (_22475_, _22474_, _22473_);
  and _73217_ (_22476_, _22475_, _08782_);
  and _73218_ (_22477_, _22476_, _22472_);
  nor _73219_ (_22479_, _10990_, _11528_);
  or _73220_ (_22480_, _22479_, _22413_);
  and _73221_ (_22481_, _22480_, _06292_);
  or _73222_ (_22482_, _22481_, _22477_);
  and _73223_ (_22483_, _22482_, _06718_);
  and _73224_ (_22484_, _22420_, _06316_);
  or _73225_ (_22485_, _22484_, _06047_);
  or _73226_ (_22486_, _22485_, _22483_);
  and _73227_ (_22487_, _14657_, _07659_);
  or _73228_ (_22488_, _22413_, _06048_);
  or _73229_ (_22490_, _22488_, _22487_);
  and _73230_ (_22491_, _22490_, _01336_);
  and _73231_ (_22492_, _22491_, _22486_);
  or _73232_ (_22493_, _22492_, _22410_);
  and _73233_ (_43385_, _22493_, _42882_);
  not _73234_ (_22494_, \oc8051_golden_model_1.TL0 [3]);
  nor _73235_ (_22495_, _01336_, _22494_);
  and _73236_ (_22496_, _09181_, _07659_);
  nor _73237_ (_22497_, _07659_, _22494_);
  or _73238_ (_22498_, _22497_, _07012_);
  or _73239_ (_22500_, _22498_, _22496_);
  nor _73240_ (_22501_, _11528_, _07353_);
  nor _73241_ (_22502_, _22501_, _22497_);
  nand _73242_ (_22503_, _22502_, _09815_);
  and _73243_ (_22504_, _14672_, _07659_);
  or _73244_ (_22505_, _22504_, _22497_);
  or _73245_ (_22506_, _22505_, _06954_);
  and _73246_ (_22507_, _07659_, \oc8051_golden_model_1.ACC [3]);
  nor _73247_ (_22508_, _22507_, _22497_);
  nor _73248_ (_22509_, _22508_, _06939_);
  nor _73249_ (_22511_, _06938_, _22494_);
  or _73250_ (_22512_, _22511_, _06102_);
  or _73251_ (_22513_, _22512_, _22509_);
  and _73252_ (_22514_, _22513_, _06848_);
  and _73253_ (_22515_, _22514_, _22506_);
  nor _73254_ (_22516_, _22502_, _06848_);
  or _73255_ (_22517_, _22516_, _22515_);
  nand _73256_ (_22518_, _22517_, _06220_);
  or _73257_ (_22519_, _22508_, _06220_);
  and _73258_ (_22520_, _22519_, _09817_);
  nand _73259_ (_22522_, _22520_, _22518_);
  and _73260_ (_22523_, _22522_, _22503_);
  and _73261_ (_22524_, _22523_, _22500_);
  or _73262_ (_22525_, _22524_, _09833_);
  and _73263_ (_22526_, _14778_, _07659_);
  or _73264_ (_22527_, _22526_, _22497_);
  or _73265_ (_22528_, _22527_, _05669_);
  and _73266_ (_22529_, _22528_, _06020_);
  and _73267_ (_22530_, _22529_, _22525_);
  and _73268_ (_22531_, _07659_, _08662_);
  or _73269_ (_22533_, _22531_, _22497_);
  and _73270_ (_22534_, _22533_, _06019_);
  or _73271_ (_22535_, _22534_, _06112_);
  or _73272_ (_22536_, _22535_, _22530_);
  and _73273_ (_22537_, _14793_, _07659_);
  or _73274_ (_22538_, _22537_, _22497_);
  or _73275_ (_22539_, _22538_, _08751_);
  and _73276_ (_22540_, _22539_, _08756_);
  and _73277_ (_22541_, _22540_, _22536_);
  and _73278_ (_22542_, _12299_, _07659_);
  or _73279_ (_22544_, _22542_, _22497_);
  and _73280_ (_22545_, _22544_, _06284_);
  or _73281_ (_22546_, _22545_, _22541_);
  and _73282_ (_22547_, _22546_, _07032_);
  or _73283_ (_22548_, _22497_, _08029_);
  and _73284_ (_22549_, _22533_, _06108_);
  and _73285_ (_22550_, _22549_, _22548_);
  or _73286_ (_22551_, _22550_, _22547_);
  and _73287_ (_22552_, _22551_, _06278_);
  nor _73288_ (_22553_, _22508_, _06278_);
  and _73289_ (_22555_, _22553_, _22548_);
  or _73290_ (_22556_, _22555_, _06130_);
  or _73291_ (_22557_, _22556_, _22552_);
  and _73292_ (_22558_, _14792_, _07659_);
  or _73293_ (_22559_, _22497_, _08777_);
  or _73294_ (_22560_, _22559_, _22558_);
  and _73295_ (_22561_, _22560_, _08782_);
  and _73296_ (_22562_, _22561_, _22557_);
  nor _73297_ (_22563_, _10988_, _11528_);
  or _73298_ (_22564_, _22563_, _22497_);
  and _73299_ (_22566_, _22564_, _06292_);
  or _73300_ (_22567_, _22566_, _22562_);
  and _73301_ (_22568_, _22567_, _06718_);
  and _73302_ (_22569_, _22505_, _06316_);
  or _73303_ (_22570_, _22569_, _06047_);
  or _73304_ (_22571_, _22570_, _22568_);
  and _73305_ (_22572_, _14849_, _07659_);
  or _73306_ (_22573_, _22497_, _06048_);
  or _73307_ (_22574_, _22573_, _22572_);
  and _73308_ (_22575_, _22574_, _01336_);
  and _73309_ (_22577_, _22575_, _22571_);
  or _73310_ (_22578_, _22577_, _22495_);
  and _73311_ (_43386_, _22578_, _42882_);
  and _73312_ (_22579_, _01340_, \oc8051_golden_model_1.TL0 [4]);
  and _73313_ (_22580_, _11528_, \oc8051_golden_model_1.TL0 [4]);
  or _73314_ (_22581_, _22580_, _08273_);
  and _73315_ (_22582_, _08665_, _07659_);
  or _73316_ (_22583_, _22582_, _22580_);
  and _73317_ (_22584_, _22583_, _06108_);
  and _73318_ (_22585_, _22584_, _22581_);
  or _73319_ (_22587_, _22583_, _06020_);
  and _73320_ (_22588_, _14887_, _07659_);
  or _73321_ (_22589_, _22588_, _22580_);
  or _73322_ (_22590_, _22589_, _06954_);
  and _73323_ (_22591_, _07659_, \oc8051_golden_model_1.ACC [4]);
  or _73324_ (_22592_, _22591_, _22580_);
  and _73325_ (_22593_, _22592_, _06938_);
  and _73326_ (_22594_, _06939_, \oc8051_golden_model_1.TL0 [4]);
  or _73327_ (_22595_, _22594_, _06102_);
  or _73328_ (_22596_, _22595_, _22593_);
  and _73329_ (_22597_, _22596_, _06848_);
  and _73330_ (_22598_, _22597_, _22590_);
  nor _73331_ (_22599_, _08270_, _11528_);
  or _73332_ (_22600_, _22599_, _22580_);
  and _73333_ (_22601_, _22600_, _06239_);
  or _73334_ (_22602_, _22601_, _22598_);
  and _73335_ (_22603_, _22602_, _06220_);
  and _73336_ (_22604_, _22592_, _06219_);
  or _73337_ (_22605_, _22604_, _09818_);
  or _73338_ (_22606_, _22605_, _22603_);
  and _73339_ (_22609_, _09180_, _07659_);
  or _73340_ (_22610_, _22580_, _07012_);
  or _73341_ (_22611_, _22610_, _22609_);
  or _73342_ (_22612_, _22600_, _09827_);
  and _73343_ (_22613_, _22612_, _05669_);
  and _73344_ (_22614_, _22613_, _22611_);
  and _73345_ (_22615_, _22614_, _22606_);
  and _73346_ (_22616_, _14983_, _07659_);
  or _73347_ (_22617_, _22616_, _22580_);
  and _73348_ (_22618_, _22617_, _09833_);
  or _73349_ (_22620_, _22618_, _06019_);
  or _73350_ (_22621_, _22620_, _22615_);
  and _73351_ (_22622_, _22621_, _22587_);
  or _73352_ (_22623_, _22622_, _06112_);
  and _73353_ (_22624_, _14876_, _07659_);
  or _73354_ (_22625_, _22580_, _08751_);
  or _73355_ (_22626_, _22625_, _22624_);
  and _73356_ (_22627_, _22626_, _08756_);
  and _73357_ (_22628_, _22627_, _22623_);
  and _73358_ (_22629_, _10986_, _07659_);
  or _73359_ (_22631_, _22629_, _22580_);
  and _73360_ (_22632_, _22631_, _06284_);
  or _73361_ (_22633_, _22632_, _22628_);
  and _73362_ (_22634_, _22633_, _07032_);
  or _73363_ (_22635_, _22634_, _22585_);
  and _73364_ (_22636_, _22635_, _06278_);
  and _73365_ (_22637_, _22592_, _06277_);
  and _73366_ (_22638_, _22637_, _22581_);
  or _73367_ (_22639_, _22638_, _06130_);
  or _73368_ (_22640_, _22639_, _22636_);
  and _73369_ (_22642_, _14873_, _07659_);
  or _73370_ (_22643_, _22580_, _08777_);
  or _73371_ (_22644_, _22643_, _22642_);
  and _73372_ (_22645_, _22644_, _08782_);
  and _73373_ (_22646_, _22645_, _22640_);
  nor _73374_ (_22647_, _10985_, _11528_);
  or _73375_ (_22648_, _22647_, _22580_);
  and _73376_ (_22649_, _22648_, _06292_);
  or _73377_ (_22650_, _22649_, _22646_);
  and _73378_ (_22651_, _22650_, _06718_);
  and _73379_ (_22653_, _22589_, _06316_);
  or _73380_ (_22654_, _22653_, _06047_);
  or _73381_ (_22655_, _22654_, _22651_);
  and _73382_ (_22656_, _15055_, _07659_);
  or _73383_ (_22657_, _22580_, _06048_);
  or _73384_ (_22658_, _22657_, _22656_);
  and _73385_ (_22659_, _22658_, _01336_);
  and _73386_ (_22660_, _22659_, _22655_);
  or _73387_ (_22661_, _22660_, _22579_);
  and _73388_ (_43387_, _22661_, _42882_);
  and _73389_ (_22663_, _01340_, \oc8051_golden_model_1.TL0 [5]);
  and _73390_ (_22664_, _11528_, \oc8051_golden_model_1.TL0 [5]);
  or _73391_ (_22665_, _22664_, _07980_);
  and _73392_ (_22666_, _08652_, _07659_);
  or _73393_ (_22667_, _22666_, _22664_);
  and _73394_ (_22668_, _22667_, _06108_);
  and _73395_ (_22669_, _22668_, _22665_);
  or _73396_ (_22670_, _22667_, _06020_);
  and _73397_ (_22671_, _15093_, _07659_);
  or _73398_ (_22672_, _22671_, _22664_);
  or _73399_ (_22674_, _22672_, _06954_);
  and _73400_ (_22675_, _07659_, \oc8051_golden_model_1.ACC [5]);
  or _73401_ (_22676_, _22675_, _22664_);
  and _73402_ (_22677_, _22676_, _06938_);
  and _73403_ (_22678_, _06939_, \oc8051_golden_model_1.TL0 [5]);
  or _73404_ (_22679_, _22678_, _06102_);
  or _73405_ (_22680_, _22679_, _22677_);
  and _73406_ (_22681_, _22680_, _06848_);
  and _73407_ (_22682_, _22681_, _22674_);
  nor _73408_ (_22683_, _07977_, _11528_);
  or _73409_ (_22685_, _22683_, _22664_);
  and _73410_ (_22686_, _22685_, _06239_);
  or _73411_ (_22687_, _22686_, _22682_);
  and _73412_ (_22688_, _22687_, _06220_);
  and _73413_ (_22689_, _22676_, _06219_);
  or _73414_ (_22690_, _22689_, _09818_);
  or _73415_ (_22691_, _22690_, _22688_);
  and _73416_ (_22692_, _09179_, _07659_);
  or _73417_ (_22693_, _22664_, _07012_);
  or _73418_ (_22694_, _22693_, _22692_);
  or _73419_ (_22696_, _22685_, _09827_);
  and _73420_ (_22697_, _22696_, _05669_);
  and _73421_ (_22698_, _22697_, _22694_);
  and _73422_ (_22699_, _22698_, _22691_);
  and _73423_ (_22700_, _15179_, _07659_);
  or _73424_ (_22701_, _22700_, _22664_);
  and _73425_ (_22702_, _22701_, _09833_);
  or _73426_ (_22703_, _22702_, _06019_);
  or _73427_ (_22704_, _22703_, _22699_);
  and _73428_ (_22705_, _22704_, _22670_);
  or _73429_ (_22706_, _22705_, _06112_);
  and _73430_ (_22707_, _15195_, _07659_);
  or _73431_ (_22708_, _22707_, _22664_);
  or _73432_ (_22709_, _22708_, _08751_);
  and _73433_ (_22710_, _22709_, _08756_);
  and _73434_ (_22711_, _22710_, _22706_);
  and _73435_ (_22712_, _12306_, _07659_);
  or _73436_ (_22713_, _22712_, _22664_);
  and _73437_ (_22714_, _22713_, _06284_);
  or _73438_ (_22715_, _22714_, _22711_);
  and _73439_ (_22718_, _22715_, _07032_);
  or _73440_ (_22719_, _22718_, _22669_);
  and _73441_ (_22720_, _22719_, _06278_);
  and _73442_ (_22721_, _22676_, _06277_);
  and _73443_ (_22722_, _22721_, _22665_);
  or _73444_ (_22723_, _22722_, _06130_);
  or _73445_ (_22724_, _22723_, _22720_);
  and _73446_ (_22725_, _15194_, _07659_);
  or _73447_ (_22726_, _22664_, _08777_);
  or _73448_ (_22727_, _22726_, _22725_);
  and _73449_ (_22729_, _22727_, _08782_);
  and _73450_ (_22730_, _22729_, _22724_);
  nor _73451_ (_22731_, _10982_, _11528_);
  or _73452_ (_22732_, _22731_, _22664_);
  and _73453_ (_22733_, _22732_, _06292_);
  or _73454_ (_22734_, _22733_, _22730_);
  and _73455_ (_22735_, _22734_, _06718_);
  and _73456_ (_22736_, _22672_, _06316_);
  or _73457_ (_22737_, _22736_, _06047_);
  or _73458_ (_22738_, _22737_, _22735_);
  and _73459_ (_22740_, _15253_, _07659_);
  or _73460_ (_22741_, _22664_, _06048_);
  or _73461_ (_22742_, _22741_, _22740_);
  and _73462_ (_22743_, _22742_, _01336_);
  and _73463_ (_22744_, _22743_, _22738_);
  or _73464_ (_22745_, _22744_, _22663_);
  and _73465_ (_43388_, _22745_, _42882_);
  and _73466_ (_22746_, _01340_, \oc8051_golden_model_1.TL0 [6]);
  and _73467_ (_22747_, _11528_, \oc8051_golden_model_1.TL0 [6]);
  or _73468_ (_22748_, _22747_, _07886_);
  and _73469_ (_22750_, _15389_, _07659_);
  or _73470_ (_22751_, _22750_, _22747_);
  and _73471_ (_22752_, _22751_, _06108_);
  and _73472_ (_22753_, _22752_, _22748_);
  or _73473_ (_22754_, _22751_, _06020_);
  and _73474_ (_22755_, _15293_, _07659_);
  or _73475_ (_22756_, _22755_, _22747_);
  or _73476_ (_22757_, _22756_, _06954_);
  and _73477_ (_22758_, _07659_, \oc8051_golden_model_1.ACC [6]);
  or _73478_ (_22759_, _22758_, _22747_);
  and _73479_ (_22761_, _22759_, _06938_);
  and _73480_ (_22762_, _06939_, \oc8051_golden_model_1.TL0 [6]);
  or _73481_ (_22763_, _22762_, _06102_);
  or _73482_ (_22764_, _22763_, _22761_);
  and _73483_ (_22765_, _22764_, _06848_);
  and _73484_ (_22766_, _22765_, _22757_);
  nor _73485_ (_22767_, _07883_, _11528_);
  or _73486_ (_22768_, _22767_, _22747_);
  and _73487_ (_22769_, _22768_, _06239_);
  or _73488_ (_22770_, _22769_, _22766_);
  and _73489_ (_22772_, _22770_, _06220_);
  and _73490_ (_22773_, _22759_, _06219_);
  or _73491_ (_22774_, _22773_, _09818_);
  or _73492_ (_22775_, _22774_, _22772_);
  and _73493_ (_22776_, _09178_, _07659_);
  or _73494_ (_22777_, _22747_, _07012_);
  or _73495_ (_22778_, _22777_, _22776_);
  or _73496_ (_22779_, _22768_, _09827_);
  and _73497_ (_22780_, _22779_, _05669_);
  and _73498_ (_22781_, _22780_, _22778_);
  and _73499_ (_22783_, _22781_, _22775_);
  and _73500_ (_22784_, _15382_, _07659_);
  or _73501_ (_22785_, _22784_, _22747_);
  and _73502_ (_22786_, _22785_, _09833_);
  or _73503_ (_22787_, _22786_, _06019_);
  or _73504_ (_22788_, _22787_, _22783_);
  and _73505_ (_22789_, _22788_, _22754_);
  or _73506_ (_22790_, _22789_, _06112_);
  and _73507_ (_22791_, _15399_, _07659_);
  or _73508_ (_22792_, _22747_, _08751_);
  or _73509_ (_22794_, _22792_, _22791_);
  and _73510_ (_22795_, _22794_, _08756_);
  and _73511_ (_22796_, _22795_, _22790_);
  and _73512_ (_22797_, _10980_, _07659_);
  or _73513_ (_22798_, _22797_, _22747_);
  and _73514_ (_22799_, _22798_, _06284_);
  or _73515_ (_22800_, _22799_, _22796_);
  and _73516_ (_22801_, _22800_, _07032_);
  or _73517_ (_22802_, _22801_, _22753_);
  and _73518_ (_22803_, _22802_, _06278_);
  and _73519_ (_22805_, _22759_, _06277_);
  and _73520_ (_22806_, _22805_, _22748_);
  or _73521_ (_22807_, _22806_, _06130_);
  or _73522_ (_22808_, _22807_, _22803_);
  and _73523_ (_22809_, _15396_, _07659_);
  or _73524_ (_22810_, _22747_, _08777_);
  or _73525_ (_22811_, _22810_, _22809_);
  and _73526_ (_22812_, _22811_, _08782_);
  and _73527_ (_22813_, _22812_, _22808_);
  nor _73528_ (_22814_, _10979_, _11528_);
  or _73529_ (_22816_, _22814_, _22747_);
  and _73530_ (_22817_, _22816_, _06292_);
  or _73531_ (_22818_, _22817_, _22813_);
  and _73532_ (_22819_, _22818_, _06718_);
  and _73533_ (_22820_, _22756_, _06316_);
  or _73534_ (_22821_, _22820_, _06047_);
  or _73535_ (_22822_, _22821_, _22819_);
  and _73536_ (_22823_, _15451_, _07659_);
  or _73537_ (_22824_, _22747_, _06048_);
  or _73538_ (_22825_, _22824_, _22823_);
  and _73539_ (_22827_, _22825_, _01336_);
  and _73540_ (_22828_, _22827_, _22822_);
  or _73541_ (_22829_, _22828_, _22746_);
  and _73542_ (_43389_, _22829_, _42882_);
  not _73543_ (_22830_, \oc8051_golden_model_1.TCON [0]);
  nor _73544_ (_22831_, _01336_, _22830_);
  nand _73545_ (_22832_, _10995_, _07648_);
  nor _73546_ (_22833_, _07648_, _22830_);
  nor _73547_ (_22834_, _22833_, _06278_);
  nand _73548_ (_22835_, _22834_, _22832_);
  and _73549_ (_22837_, _07648_, _08672_);
  or _73550_ (_22838_, _22837_, _22833_);
  or _73551_ (_22839_, _22838_, _06020_);
  and _73552_ (_22840_, _09120_, _07648_);
  or _73553_ (_22841_, _22833_, _07012_);
  or _73554_ (_22842_, _22841_, _22840_);
  nor _73555_ (_22843_, _08127_, _11605_);
  or _73556_ (_22844_, _22843_, _22833_);
  or _73557_ (_22845_, _22844_, _06954_);
  and _73558_ (_22846_, _07648_, \oc8051_golden_model_1.ACC [0]);
  or _73559_ (_22848_, _22846_, _22833_);
  and _73560_ (_22849_, _22848_, _06938_);
  nor _73561_ (_22850_, _06938_, _22830_);
  or _73562_ (_22851_, _22850_, _06102_);
  or _73563_ (_22852_, _22851_, _22849_);
  and _73564_ (_22853_, _22852_, _06044_);
  and _73565_ (_22854_, _22853_, _22845_);
  nor _73566_ (_22855_, _08341_, _22830_);
  and _73567_ (_22856_, _14102_, _08341_);
  or _73568_ (_22857_, _22856_, _22855_);
  and _73569_ (_22859_, _22857_, _06043_);
  or _73570_ (_22860_, _22859_, _22854_);
  and _73571_ (_22861_, _22860_, _06848_);
  and _73572_ (_22862_, _07648_, _06931_);
  or _73573_ (_22863_, _22862_, _22833_);
  and _73574_ (_22864_, _22863_, _06239_);
  or _73575_ (_22865_, _22864_, _06219_);
  or _73576_ (_22866_, _22865_, _22861_);
  or _73577_ (_22867_, _22848_, _06220_);
  and _73578_ (_22868_, _22867_, _06040_);
  and _73579_ (_22870_, _22868_, _22866_);
  and _73580_ (_22871_, _22833_, _06039_);
  or _73581_ (_22872_, _22871_, _06032_);
  or _73582_ (_22873_, _22872_, _22870_);
  or _73583_ (_22874_, _22844_, _06033_);
  and _73584_ (_22875_, _22874_, _06027_);
  and _73585_ (_22876_, _22875_, _22873_);
  or _73586_ (_22877_, _22855_, _14131_);
  and _73587_ (_22878_, _22877_, _06026_);
  and _73588_ (_22879_, _22878_, _22857_);
  or _73589_ (_22881_, _22879_, _09818_);
  or _73590_ (_22882_, _22881_, _22876_);
  or _73591_ (_22883_, _22863_, _09827_);
  and _73592_ (_22884_, _22883_, _05669_);
  and _73593_ (_22885_, _22884_, _22882_);
  and _73594_ (_22886_, _22885_, _22842_);
  and _73595_ (_22887_, _14186_, _07648_);
  or _73596_ (_22888_, _22887_, _22833_);
  and _73597_ (_22889_, _22888_, _09833_);
  or _73598_ (_22890_, _22889_, _06019_);
  or _73599_ (_22892_, _22890_, _22886_);
  and _73600_ (_22893_, _22892_, _22839_);
  or _73601_ (_22894_, _22893_, _06112_);
  and _73602_ (_22895_, _14086_, _07648_);
  or _73603_ (_22896_, _22833_, _08751_);
  or _73604_ (_22897_, _22896_, _22895_);
  and _73605_ (_22898_, _22897_, _08756_);
  and _73606_ (_22899_, _22898_, _22894_);
  nor _73607_ (_22900_, _12302_, _11605_);
  or _73608_ (_22901_, _22900_, _22833_);
  and _73609_ (_22903_, _22832_, _06284_);
  and _73610_ (_22904_, _22903_, _22901_);
  or _73611_ (_22905_, _22904_, _22899_);
  and _73612_ (_22906_, _22905_, _07032_);
  nand _73613_ (_22907_, _22838_, _06108_);
  nor _73614_ (_22908_, _22907_, _22843_);
  or _73615_ (_22909_, _22908_, _06277_);
  or _73616_ (_22910_, _22909_, _22906_);
  and _73617_ (_22911_, _22910_, _22835_);
  or _73618_ (_22912_, _22911_, _06130_);
  and _73619_ (_22914_, _14083_, _07648_);
  or _73620_ (_22915_, _22833_, _08777_);
  or _73621_ (_22916_, _22915_, _22914_);
  and _73622_ (_22917_, _22916_, _08782_);
  and _73623_ (_22918_, _22917_, _22912_);
  and _73624_ (_22919_, _22901_, _06292_);
  or _73625_ (_22920_, _22919_, _06316_);
  or _73626_ (_22921_, _22920_, _22918_);
  or _73627_ (_22922_, _22844_, _06718_);
  and _73628_ (_22923_, _22922_, _22921_);
  or _73629_ (_22924_, _22923_, _05652_);
  or _73630_ (_22925_, _22833_, _05653_);
  and _73631_ (_22926_, _22925_, _22924_);
  or _73632_ (_22927_, _22926_, _06047_);
  or _73633_ (_22928_, _22844_, _06048_);
  and _73634_ (_22929_, _22928_, _01336_);
  and _73635_ (_22930_, _22929_, _22927_);
  or _73636_ (_22931_, _22930_, _22831_);
  and _73637_ (_43391_, _22931_, _42882_);
  and _73638_ (_22932_, _01340_, \oc8051_golden_model_1.TCON [1]);
  and _73639_ (_22935_, _11605_, \oc8051_golden_model_1.TCON [1]);
  nor _73640_ (_22936_, _10993_, _11605_);
  or _73641_ (_22937_, _22936_, _22935_);
  or _73642_ (_22938_, _22937_, _08782_);
  or _73643_ (_22939_, _14367_, _11605_);
  or _73644_ (_22940_, _07648_, \oc8051_golden_model_1.TCON [1]);
  and _73645_ (_22941_, _22940_, _09833_);
  and _73646_ (_22942_, _22941_, _22939_);
  nor _73647_ (_22943_, _11605_, _07132_);
  or _73648_ (_22944_, _22943_, _22935_);
  or _73649_ (_22946_, _22944_, _06848_);
  and _73650_ (_22947_, _14284_, _07648_);
  not _73651_ (_22948_, _22947_);
  and _73652_ (_22949_, _22948_, _22940_);
  or _73653_ (_22950_, _22949_, _06954_);
  and _73654_ (_22951_, _07648_, \oc8051_golden_model_1.ACC [1]);
  or _73655_ (_22952_, _22951_, _22935_);
  and _73656_ (_22953_, _22952_, _06938_);
  and _73657_ (_22954_, _06939_, \oc8051_golden_model_1.TCON [1]);
  or _73658_ (_22955_, _22954_, _06102_);
  or _73659_ (_22957_, _22955_, _22953_);
  and _73660_ (_22958_, _22957_, _06044_);
  and _73661_ (_22959_, _22958_, _22950_);
  and _73662_ (_22960_, _11624_, \oc8051_golden_model_1.TCON [1]);
  and _73663_ (_22961_, _14266_, _08341_);
  or _73664_ (_22962_, _22961_, _22960_);
  and _73665_ (_22963_, _22962_, _06043_);
  or _73666_ (_22964_, _22963_, _06239_);
  or _73667_ (_22965_, _22964_, _22959_);
  and _73668_ (_22966_, _22965_, _22946_);
  or _73669_ (_22968_, _22966_, _06219_);
  or _73670_ (_22969_, _22952_, _06220_);
  and _73671_ (_22970_, _22969_, _06040_);
  and _73672_ (_22971_, _22970_, _22968_);
  and _73673_ (_22972_, _14273_, _08341_);
  or _73674_ (_22973_, _22972_, _22960_);
  and _73675_ (_22974_, _22973_, _06039_);
  or _73676_ (_22975_, _22974_, _06032_);
  or _73677_ (_22976_, _22975_, _22971_);
  and _73678_ (_22977_, _22961_, _14302_);
  or _73679_ (_22979_, _22960_, _06033_);
  or _73680_ (_22980_, _22979_, _22977_);
  and _73681_ (_22981_, _22980_, _06027_);
  and _73682_ (_22982_, _22981_, _22976_);
  or _73683_ (_22983_, _22960_, _14267_);
  and _73684_ (_22984_, _22983_, _06026_);
  and _73685_ (_22985_, _22984_, _22962_);
  or _73686_ (_22986_, _22985_, _09818_);
  or _73687_ (_22987_, _22986_, _22982_);
  and _73688_ (_22988_, _09075_, _07648_);
  or _73689_ (_22990_, _22935_, _07012_);
  or _73690_ (_22991_, _22990_, _22988_);
  or _73691_ (_22992_, _22944_, _09827_);
  and _73692_ (_22993_, _22992_, _05669_);
  and _73693_ (_22994_, _22993_, _22991_);
  and _73694_ (_22995_, _22994_, _22987_);
  or _73695_ (_22996_, _22995_, _22942_);
  and _73696_ (_22997_, _22996_, _06020_);
  nand _73697_ (_22998_, _07648_, _06832_);
  and _73698_ (_22999_, _22940_, _06019_);
  and _73699_ (_23001_, _22999_, _22998_);
  or _73700_ (_23002_, _23001_, _22997_);
  and _73701_ (_23003_, _23002_, _08751_);
  or _73702_ (_23004_, _14263_, _11605_);
  and _73703_ (_23005_, _22940_, _06112_);
  and _73704_ (_23006_, _23005_, _23004_);
  or _73705_ (_23007_, _23006_, _06284_);
  or _73706_ (_23008_, _23007_, _23003_);
  and _73707_ (_23009_, _10994_, _07648_);
  or _73708_ (_23010_, _23009_, _22935_);
  or _73709_ (_23012_, _23010_, _08756_);
  and _73710_ (_23013_, _23012_, _07032_);
  and _73711_ (_23014_, _23013_, _23008_);
  or _73712_ (_23015_, _14261_, _11605_);
  and _73713_ (_23016_, _22940_, _06108_);
  and _73714_ (_23017_, _23016_, _23015_);
  or _73715_ (_23018_, _23017_, _06277_);
  or _73716_ (_23019_, _23018_, _23014_);
  and _73717_ (_23020_, _22951_, _08078_);
  or _73718_ (_23021_, _22935_, _06278_);
  or _73719_ (_23023_, _23021_, _23020_);
  and _73720_ (_23024_, _23023_, _08777_);
  and _73721_ (_23025_, _23024_, _23019_);
  or _73722_ (_23026_, _22998_, _08078_);
  and _73723_ (_23027_, _22940_, _06130_);
  and _73724_ (_23028_, _23027_, _23026_);
  or _73725_ (_23029_, _23028_, _06292_);
  or _73726_ (_23030_, _23029_, _23025_);
  and _73727_ (_23031_, _23030_, _22938_);
  or _73728_ (_23032_, _23031_, _06316_);
  or _73729_ (_23034_, _22949_, _06718_);
  and _73730_ (_23035_, _23034_, _05653_);
  and _73731_ (_23036_, _23035_, _23032_);
  and _73732_ (_23037_, _22973_, _05652_);
  or _73733_ (_23038_, _23037_, _06047_);
  or _73734_ (_23039_, _23038_, _23036_);
  or _73735_ (_23040_, _22935_, _06048_);
  or _73736_ (_23041_, _23040_, _22947_);
  and _73737_ (_23042_, _23041_, _01336_);
  and _73738_ (_23043_, _23042_, _23039_);
  or _73739_ (_23044_, _23043_, _22932_);
  and _73740_ (_43392_, _23044_, _42882_);
  and _73741_ (_23045_, _01340_, \oc8051_golden_model_1.TCON [2]);
  and _73742_ (_23046_, _11605_, \oc8051_golden_model_1.TCON [2]);
  and _73743_ (_23047_, _07648_, _08730_);
  or _73744_ (_23048_, _23047_, _23046_);
  or _73745_ (_23049_, _23048_, _06020_);
  nor _73746_ (_23050_, _11605_, _07530_);
  or _73747_ (_23051_, _23050_, _23046_);
  and _73748_ (_23052_, _23051_, _06239_);
  and _73749_ (_23054_, _11624_, \oc8051_golden_model_1.TCON [2]);
  and _73750_ (_23055_, _14497_, _08341_);
  or _73751_ (_23056_, _23055_, _23054_);
  or _73752_ (_23057_, _23056_, _06044_);
  and _73753_ (_23058_, _14493_, _07648_);
  or _73754_ (_23059_, _23058_, _23046_);
  and _73755_ (_23060_, _23059_, _06102_);
  and _73756_ (_23061_, _06939_, \oc8051_golden_model_1.TCON [2]);
  and _73757_ (_23062_, _07648_, \oc8051_golden_model_1.ACC [2]);
  or _73758_ (_23063_, _23062_, _23046_);
  and _73759_ (_23065_, _23063_, _06938_);
  or _73760_ (_23066_, _23065_, _23061_);
  and _73761_ (_23067_, _23066_, _06954_);
  or _73762_ (_23068_, _23067_, _06043_);
  or _73763_ (_23069_, _23068_, _23060_);
  and _73764_ (_23070_, _23069_, _23057_);
  and _73765_ (_23071_, _23070_, _06848_);
  or _73766_ (_23072_, _23071_, _23052_);
  or _73767_ (_23073_, _23072_, _06219_);
  or _73768_ (_23074_, _23063_, _06220_);
  and _73769_ (_23076_, _23074_, _06040_);
  and _73770_ (_23077_, _23076_, _23073_);
  and _73771_ (_23078_, _14479_, _08341_);
  or _73772_ (_23079_, _23078_, _23054_);
  and _73773_ (_23080_, _23079_, _06039_);
  or _73774_ (_23081_, _23080_, _06032_);
  or _73775_ (_23082_, _23081_, _23077_);
  or _73776_ (_23083_, _23054_, _14512_);
  and _73777_ (_23084_, _23083_, _23056_);
  or _73778_ (_23085_, _23084_, _06033_);
  and _73779_ (_23086_, _23085_, _06027_);
  and _73780_ (_23087_, _23086_, _23082_);
  or _73781_ (_23088_, _23054_, _14525_);
  and _73782_ (_23089_, _23088_, _06026_);
  and _73783_ (_23090_, _23089_, _23056_);
  or _73784_ (_23091_, _23090_, _09818_);
  or _73785_ (_23092_, _23091_, _23087_);
  and _73786_ (_23093_, _09182_, _07648_);
  or _73787_ (_23094_, _23046_, _07012_);
  or _73788_ (_23095_, _23094_, _23093_);
  or _73789_ (_23097_, _23051_, _09827_);
  and _73790_ (_23098_, _23097_, _05669_);
  and _73791_ (_23099_, _23098_, _23095_);
  and _73792_ (_23100_, _23099_, _23092_);
  and _73793_ (_23101_, _14580_, _07648_);
  or _73794_ (_23102_, _23101_, _23046_);
  and _73795_ (_23103_, _23102_, _09833_);
  or _73796_ (_23104_, _23103_, _06019_);
  or _73797_ (_23105_, _23104_, _23100_);
  and _73798_ (_23106_, _23105_, _23049_);
  or _73799_ (_23107_, _23106_, _06112_);
  and _73800_ (_23108_, _14596_, _07648_);
  or _73801_ (_23109_, _23108_, _23046_);
  or _73802_ (_23110_, _23109_, _08751_);
  and _73803_ (_23111_, _23110_, _08756_);
  and _73804_ (_23112_, _23111_, _23107_);
  and _73805_ (_23113_, _10991_, _07648_);
  or _73806_ (_23114_, _23113_, _23046_);
  and _73807_ (_23115_, _23114_, _06284_);
  or _73808_ (_23116_, _23115_, _23112_);
  and _73809_ (_23118_, _23116_, _07032_);
  or _73810_ (_23119_, _23046_, _08177_);
  and _73811_ (_23120_, _23048_, _06108_);
  and _73812_ (_23121_, _23120_, _23119_);
  or _73813_ (_23122_, _23121_, _23118_);
  and _73814_ (_23123_, _23122_, _06278_);
  and _73815_ (_23124_, _23063_, _06277_);
  and _73816_ (_23125_, _23124_, _23119_);
  or _73817_ (_23126_, _23125_, _06130_);
  or _73818_ (_23127_, _23126_, _23123_);
  and _73819_ (_23129_, _14593_, _07648_);
  or _73820_ (_23130_, _23046_, _08777_);
  or _73821_ (_23131_, _23130_, _23129_);
  and _73822_ (_23132_, _23131_, _08782_);
  and _73823_ (_23133_, _23132_, _23127_);
  nor _73824_ (_23134_, _10990_, _11605_);
  or _73825_ (_23135_, _23134_, _23046_);
  and _73826_ (_23136_, _23135_, _06292_);
  or _73827_ (_23137_, _23136_, _06316_);
  or _73828_ (_23138_, _23137_, _23133_);
  or _73829_ (_23139_, _23059_, _06718_);
  and _73830_ (_23140_, _23139_, _05653_);
  and _73831_ (_23141_, _23140_, _23138_);
  and _73832_ (_23142_, _23079_, _05652_);
  or _73833_ (_23143_, _23142_, _06047_);
  or _73834_ (_23144_, _23143_, _23141_);
  and _73835_ (_23145_, _14657_, _07648_);
  or _73836_ (_23146_, _23046_, _06048_);
  or _73837_ (_23147_, _23146_, _23145_);
  and _73838_ (_23148_, _23147_, _01336_);
  and _73839_ (_23150_, _23148_, _23144_);
  or _73840_ (_23151_, _23150_, _23045_);
  and _73841_ (_43393_, _23151_, _42882_);
  and _73842_ (_23152_, _01340_, \oc8051_golden_model_1.TCON [3]);
  and _73843_ (_23153_, _11605_, \oc8051_golden_model_1.TCON [3]);
  and _73844_ (_23154_, _07648_, _08662_);
  or _73845_ (_23155_, _23154_, _23153_);
  or _73846_ (_23156_, _23155_, _06020_);
  and _73847_ (_23157_, _14672_, _07648_);
  or _73848_ (_23158_, _23157_, _23153_);
  or _73849_ (_23160_, _23158_, _06954_);
  and _73850_ (_23161_, _07648_, \oc8051_golden_model_1.ACC [3]);
  or _73851_ (_23162_, _23161_, _23153_);
  and _73852_ (_23163_, _23162_, _06938_);
  and _73853_ (_23164_, _06939_, \oc8051_golden_model_1.TCON [3]);
  or _73854_ (_23165_, _23164_, _06102_);
  or _73855_ (_23166_, _23165_, _23163_);
  and _73856_ (_23167_, _23166_, _06044_);
  and _73857_ (_23168_, _23167_, _23160_);
  and _73858_ (_23169_, _11624_, \oc8051_golden_model_1.TCON [3]);
  and _73859_ (_23170_, _14683_, _08341_);
  or _73860_ (_23171_, _23170_, _23169_);
  and _73861_ (_23172_, _23171_, _06043_);
  or _73862_ (_23173_, _23172_, _06239_);
  or _73863_ (_23174_, _23173_, _23168_);
  nor _73864_ (_23175_, _11605_, _07353_);
  or _73865_ (_23176_, _23175_, _23153_);
  or _73866_ (_23177_, _23176_, _06848_);
  and _73867_ (_23178_, _23177_, _23174_);
  or _73868_ (_23179_, _23178_, _06219_);
  or _73869_ (_23180_, _23162_, _06220_);
  and _73870_ (_23181_, _23180_, _06040_);
  and _73871_ (_23182_, _23181_, _23179_);
  and _73872_ (_23183_, _14681_, _08341_);
  or _73873_ (_23184_, _23183_, _23169_);
  and _73874_ (_23185_, _23184_, _06039_);
  or _73875_ (_23186_, _23185_, _06032_);
  or _73876_ (_23187_, _23186_, _23182_);
  or _73877_ (_23188_, _23169_, _14708_);
  and _73878_ (_23189_, _23188_, _23171_);
  or _73879_ (_23192_, _23189_, _06033_);
  and _73880_ (_23193_, _23192_, _06027_);
  and _73881_ (_23194_, _23193_, _23187_);
  and _73882_ (_23195_, _14724_, _08341_);
  or _73883_ (_23196_, _23195_, _23169_);
  and _73884_ (_23197_, _23196_, _06026_);
  or _73885_ (_23198_, _23197_, _09818_);
  or _73886_ (_23199_, _23198_, _23194_);
  and _73887_ (_23200_, _09181_, _07648_);
  or _73888_ (_23201_, _23153_, _07012_);
  or _73889_ (_23202_, _23201_, _23200_);
  or _73890_ (_23203_, _23176_, _09827_);
  and _73891_ (_23204_, _23203_, _05669_);
  and _73892_ (_23205_, _23204_, _23202_);
  and _73893_ (_23206_, _23205_, _23199_);
  and _73894_ (_23207_, _14778_, _07648_);
  or _73895_ (_23208_, _23207_, _23153_);
  and _73896_ (_23209_, _23208_, _09833_);
  or _73897_ (_23210_, _23209_, _06019_);
  or _73898_ (_23211_, _23210_, _23206_);
  and _73899_ (_23213_, _23211_, _23156_);
  or _73900_ (_23214_, _23213_, _06112_);
  and _73901_ (_23215_, _14793_, _07648_);
  or _73902_ (_23216_, _23153_, _08751_);
  or _73903_ (_23217_, _23216_, _23215_);
  and _73904_ (_23218_, _23217_, _08756_);
  and _73905_ (_23219_, _23218_, _23214_);
  and _73906_ (_23220_, _12299_, _07648_);
  or _73907_ (_23221_, _23220_, _23153_);
  and _73908_ (_23222_, _23221_, _06284_);
  or _73909_ (_23224_, _23222_, _23219_);
  and _73910_ (_23225_, _23224_, _07032_);
  or _73911_ (_23226_, _23153_, _08029_);
  and _73912_ (_23227_, _23155_, _06108_);
  and _73913_ (_23228_, _23227_, _23226_);
  or _73914_ (_23229_, _23228_, _23225_);
  and _73915_ (_23230_, _23229_, _06278_);
  and _73916_ (_23231_, _23162_, _06277_);
  and _73917_ (_23232_, _23231_, _23226_);
  or _73918_ (_23233_, _23232_, _06130_);
  or _73919_ (_23234_, _23233_, _23230_);
  and _73920_ (_23235_, _14792_, _07648_);
  or _73921_ (_23236_, _23153_, _08777_);
  or _73922_ (_23237_, _23236_, _23235_);
  and _73923_ (_23238_, _23237_, _08782_);
  and _73924_ (_23239_, _23238_, _23234_);
  nor _73925_ (_23240_, _10988_, _11605_);
  or _73926_ (_23241_, _23240_, _23153_);
  and _73927_ (_23242_, _23241_, _06292_);
  or _73928_ (_23243_, _23242_, _06316_);
  or _73929_ (_23245_, _23243_, _23239_);
  or _73930_ (_23246_, _23158_, _06718_);
  and _73931_ (_23247_, _23246_, _05653_);
  and _73932_ (_23248_, _23247_, _23245_);
  and _73933_ (_23249_, _23184_, _05652_);
  or _73934_ (_23250_, _23249_, _06047_);
  or _73935_ (_23251_, _23250_, _23248_);
  and _73936_ (_23252_, _14849_, _07648_);
  or _73937_ (_23253_, _23153_, _06048_);
  or _73938_ (_23254_, _23253_, _23252_);
  and _73939_ (_23256_, _23254_, _01336_);
  and _73940_ (_23257_, _23256_, _23251_);
  or _73941_ (_23258_, _23257_, _23152_);
  and _73942_ (_43394_, _23258_, _42882_);
  and _73943_ (_23259_, _01340_, \oc8051_golden_model_1.TCON [4]);
  and _73944_ (_23260_, _11605_, \oc8051_golden_model_1.TCON [4]);
  and _73945_ (_23261_, _08665_, _07648_);
  or _73946_ (_23262_, _23261_, _23260_);
  or _73947_ (_23263_, _23262_, _06020_);
  and _73948_ (_23264_, _14887_, _07648_);
  or _73949_ (_23265_, _23264_, _23260_);
  or _73950_ (_23266_, _23265_, _06954_);
  and _73951_ (_23267_, _07648_, \oc8051_golden_model_1.ACC [4]);
  or _73952_ (_23268_, _23267_, _23260_);
  and _73953_ (_23269_, _23268_, _06938_);
  and _73954_ (_23270_, _06939_, \oc8051_golden_model_1.TCON [4]);
  or _73955_ (_23271_, _23270_, _06102_);
  or _73956_ (_23272_, _23271_, _23269_);
  and _73957_ (_23273_, _23272_, _06044_);
  and _73958_ (_23274_, _23273_, _23266_);
  and _73959_ (_23276_, _11624_, \oc8051_golden_model_1.TCON [4]);
  and _73960_ (_23277_, _14878_, _08341_);
  or _73961_ (_23278_, _23277_, _23276_);
  and _73962_ (_23279_, _23278_, _06043_);
  or _73963_ (_23280_, _23279_, _06239_);
  or _73964_ (_23281_, _23280_, _23274_);
  nor _73965_ (_23282_, _08270_, _11605_);
  or _73966_ (_23283_, _23282_, _23260_);
  or _73967_ (_23284_, _23283_, _06848_);
  and _73968_ (_23285_, _23284_, _23281_);
  or _73969_ (_23287_, _23285_, _06219_);
  or _73970_ (_23288_, _23268_, _06220_);
  and _73971_ (_23289_, _23288_, _06040_);
  and _73972_ (_23290_, _23289_, _23287_);
  and _73973_ (_23291_, _14882_, _08341_);
  or _73974_ (_23292_, _23291_, _23276_);
  and _73975_ (_23293_, _23292_, _06039_);
  or _73976_ (_23294_, _23293_, _06032_);
  or _73977_ (_23295_, _23294_, _23290_);
  or _73978_ (_23296_, _23276_, _14914_);
  and _73979_ (_23297_, _23296_, _23278_);
  or _73980_ (_23298_, _23297_, _06033_);
  and _73981_ (_23299_, _23298_, _06027_);
  and _73982_ (_23300_, _23299_, _23295_);
  or _73983_ (_23301_, _23276_, _14879_);
  and _73984_ (_23302_, _23301_, _06026_);
  and _73985_ (_23303_, _23302_, _23278_);
  or _73986_ (_23304_, _23303_, _09818_);
  or _73987_ (_23305_, _23304_, _23300_);
  and _73988_ (_23306_, _09180_, _07648_);
  or _73989_ (_23308_, _23260_, _07012_);
  or _73990_ (_23309_, _23308_, _23306_);
  or _73991_ (_23310_, _23283_, _09827_);
  and _73992_ (_23311_, _23310_, _05669_);
  and _73993_ (_23312_, _23311_, _23309_);
  and _73994_ (_23313_, _23312_, _23305_);
  and _73995_ (_23314_, _14983_, _07648_);
  or _73996_ (_23315_, _23314_, _23260_);
  and _73997_ (_23316_, _23315_, _09833_);
  or _73998_ (_23317_, _23316_, _06019_);
  or _73999_ (_23319_, _23317_, _23313_);
  and _74000_ (_23320_, _23319_, _23263_);
  or _74001_ (_23321_, _23320_, _06112_);
  and _74002_ (_23322_, _14876_, _07648_);
  or _74003_ (_23323_, _23260_, _08751_);
  or _74004_ (_23324_, _23323_, _23322_);
  and _74005_ (_23325_, _23324_, _08756_);
  and _74006_ (_23326_, _23325_, _23321_);
  and _74007_ (_23327_, _10986_, _07648_);
  or _74008_ (_23328_, _23327_, _23260_);
  and _74009_ (_23329_, _23328_, _06284_);
  or _74010_ (_23330_, _23329_, _23326_);
  and _74011_ (_23331_, _23330_, _07032_);
  or _74012_ (_23332_, _23260_, _08273_);
  and _74013_ (_23333_, _23262_, _06108_);
  and _74014_ (_23334_, _23333_, _23332_);
  or _74015_ (_23335_, _23334_, _23331_);
  and _74016_ (_23336_, _23335_, _06278_);
  and _74017_ (_23337_, _23268_, _06277_);
  and _74018_ (_23338_, _23337_, _23332_);
  or _74019_ (_23340_, _23338_, _06130_);
  or _74020_ (_23341_, _23340_, _23336_);
  and _74021_ (_23342_, _14873_, _07648_);
  or _74022_ (_23343_, _23260_, _08777_);
  or _74023_ (_23344_, _23343_, _23342_);
  and _74024_ (_23345_, _23344_, _08782_);
  and _74025_ (_23346_, _23345_, _23341_);
  nor _74026_ (_23347_, _10985_, _11605_);
  or _74027_ (_23348_, _23347_, _23260_);
  and _74028_ (_23349_, _23348_, _06292_);
  or _74029_ (_23351_, _23349_, _06316_);
  or _74030_ (_23352_, _23351_, _23346_);
  or _74031_ (_23353_, _23265_, _06718_);
  and _74032_ (_23354_, _23353_, _05653_);
  and _74033_ (_23355_, _23354_, _23352_);
  and _74034_ (_23356_, _23292_, _05652_);
  or _74035_ (_23357_, _23356_, _06047_);
  or _74036_ (_23358_, _23357_, _23355_);
  and _74037_ (_23359_, _15055_, _07648_);
  or _74038_ (_23360_, _23260_, _06048_);
  or _74039_ (_23361_, _23360_, _23359_);
  and _74040_ (_23362_, _23361_, _01336_);
  and _74041_ (_23363_, _23362_, _23358_);
  or _74042_ (_23364_, _23363_, _23259_);
  and _74043_ (_43395_, _23364_, _42882_);
  and _74044_ (_23365_, _01340_, \oc8051_golden_model_1.TCON [5]);
  and _74045_ (_23366_, _11605_, \oc8051_golden_model_1.TCON [5]);
  and _74046_ (_23367_, _08652_, _07648_);
  or _74047_ (_23368_, _23367_, _23366_);
  or _74048_ (_23369_, _23368_, _06020_);
  and _74049_ (_23371_, _15093_, _07648_);
  or _74050_ (_23372_, _23371_, _23366_);
  or _74051_ (_23373_, _23372_, _06954_);
  and _74052_ (_23374_, _07648_, \oc8051_golden_model_1.ACC [5]);
  or _74053_ (_23375_, _23374_, _23366_);
  and _74054_ (_23376_, _23375_, _06938_);
  and _74055_ (_23377_, _06939_, \oc8051_golden_model_1.TCON [5]);
  or _74056_ (_23378_, _23377_, _06102_);
  or _74057_ (_23379_, _23378_, _23376_);
  and _74058_ (_23380_, _23379_, _06044_);
  and _74059_ (_23382_, _23380_, _23373_);
  and _74060_ (_23383_, _11624_, \oc8051_golden_model_1.TCON [5]);
  and _74061_ (_23384_, _15073_, _08341_);
  or _74062_ (_23385_, _23384_, _23383_);
  and _74063_ (_23386_, _23385_, _06043_);
  or _74064_ (_23387_, _23386_, _06239_);
  or _74065_ (_23388_, _23387_, _23382_);
  nor _74066_ (_23389_, _07977_, _11605_);
  or _74067_ (_23390_, _23389_, _23366_);
  or _74068_ (_23391_, _23390_, _06848_);
  and _74069_ (_23392_, _23391_, _23388_);
  or _74070_ (_23393_, _23392_, _06219_);
  or _74071_ (_23394_, _23375_, _06220_);
  and _74072_ (_23395_, _23394_, _06040_);
  and _74073_ (_23396_, _23395_, _23393_);
  and _74074_ (_23397_, _15077_, _08341_);
  or _74075_ (_23398_, _23397_, _23383_);
  and _74076_ (_23399_, _23398_, _06039_);
  or _74077_ (_23400_, _23399_, _06032_);
  or _74078_ (_23401_, _23400_, _23396_);
  or _74079_ (_23403_, _23383_, _15110_);
  and _74080_ (_23404_, _23403_, _23385_);
  or _74081_ (_23405_, _23404_, _06033_);
  and _74082_ (_23406_, _23405_, _06027_);
  and _74083_ (_23407_, _23406_, _23401_);
  or _74084_ (_23408_, _23383_, _15074_);
  and _74085_ (_23409_, _23408_, _06026_);
  and _74086_ (_23410_, _23409_, _23385_);
  or _74087_ (_23411_, _23410_, _09818_);
  or _74088_ (_23412_, _23411_, _23407_);
  and _74089_ (_23414_, _09179_, _07648_);
  or _74090_ (_23415_, _23366_, _07012_);
  or _74091_ (_23416_, _23415_, _23414_);
  or _74092_ (_23417_, _23390_, _09827_);
  and _74093_ (_23418_, _23417_, _05669_);
  and _74094_ (_23419_, _23418_, _23416_);
  and _74095_ (_23420_, _23419_, _23412_);
  and _74096_ (_23421_, _15179_, _07648_);
  or _74097_ (_23422_, _23421_, _23366_);
  and _74098_ (_23423_, _23422_, _09833_);
  or _74099_ (_23424_, _23423_, _06019_);
  or _74100_ (_23425_, _23424_, _23420_);
  and _74101_ (_23426_, _23425_, _23369_);
  or _74102_ (_23427_, _23426_, _06112_);
  and _74103_ (_23428_, _15195_, _07648_);
  or _74104_ (_23429_, _23428_, _23366_);
  or _74105_ (_23430_, _23429_, _08751_);
  and _74106_ (_23431_, _23430_, _08756_);
  and _74107_ (_23432_, _23431_, _23427_);
  and _74108_ (_23433_, _12306_, _07648_);
  or _74109_ (_23435_, _23433_, _23366_);
  and _74110_ (_23436_, _23435_, _06284_);
  or _74111_ (_23437_, _23436_, _23432_);
  and _74112_ (_23438_, _23437_, _07032_);
  or _74113_ (_23439_, _23366_, _07980_);
  and _74114_ (_23440_, _23368_, _06108_);
  and _74115_ (_23441_, _23440_, _23439_);
  or _74116_ (_23442_, _23441_, _23438_);
  and _74117_ (_23443_, _23442_, _06278_);
  and _74118_ (_23444_, _23375_, _06277_);
  and _74119_ (_23446_, _23444_, _23439_);
  or _74120_ (_23447_, _23446_, _06130_);
  or _74121_ (_23448_, _23447_, _23443_);
  and _74122_ (_23449_, _15194_, _07648_);
  or _74123_ (_23450_, _23366_, _08777_);
  or _74124_ (_23451_, _23450_, _23449_);
  and _74125_ (_23452_, _23451_, _08782_);
  and _74126_ (_23453_, _23452_, _23448_);
  nor _74127_ (_23454_, _10982_, _11605_);
  or _74128_ (_23455_, _23454_, _23366_);
  and _74129_ (_23456_, _23455_, _06292_);
  or _74130_ (_23457_, _23456_, _06316_);
  or _74131_ (_23458_, _23457_, _23453_);
  or _74132_ (_23459_, _23372_, _06718_);
  and _74133_ (_23460_, _23459_, _05653_);
  and _74134_ (_23461_, _23460_, _23458_);
  and _74135_ (_23462_, _23398_, _05652_);
  or _74136_ (_23463_, _23462_, _06047_);
  or _74137_ (_23464_, _23463_, _23461_);
  and _74138_ (_23465_, _15253_, _07648_);
  or _74139_ (_23467_, _23366_, _06048_);
  or _74140_ (_23468_, _23467_, _23465_);
  and _74141_ (_23469_, _23468_, _01336_);
  and _74142_ (_23470_, _23469_, _23464_);
  or _74143_ (_23471_, _23470_, _23365_);
  and _74144_ (_43396_, _23471_, _42882_);
  and _74145_ (_23472_, _01340_, \oc8051_golden_model_1.TCON [6]);
  and _74146_ (_23473_, _11605_, \oc8051_golden_model_1.TCON [6]);
  and _74147_ (_23474_, _15389_, _07648_);
  or _74148_ (_23475_, _23474_, _23473_);
  or _74149_ (_23477_, _23475_, _06020_);
  and _74150_ (_23478_, _15293_, _07648_);
  or _74151_ (_23479_, _23478_, _23473_);
  or _74152_ (_23480_, _23479_, _06954_);
  and _74153_ (_23481_, _07648_, \oc8051_golden_model_1.ACC [6]);
  or _74154_ (_23482_, _23481_, _23473_);
  and _74155_ (_23483_, _23482_, _06938_);
  and _74156_ (_23484_, _06939_, \oc8051_golden_model_1.TCON [6]);
  or _74157_ (_23485_, _23484_, _06102_);
  or _74158_ (_23486_, _23485_, _23483_);
  and _74159_ (_23488_, _23486_, _06044_);
  and _74160_ (_23489_, _23488_, _23480_);
  and _74161_ (_23490_, _11624_, \oc8051_golden_model_1.TCON [6]);
  and _74162_ (_23491_, _15280_, _08341_);
  or _74163_ (_23492_, _23491_, _23490_);
  and _74164_ (_23493_, _23492_, _06043_);
  or _74165_ (_23494_, _23493_, _06239_);
  or _74166_ (_23495_, _23494_, _23489_);
  nor _74167_ (_23496_, _07883_, _11605_);
  or _74168_ (_23497_, _23496_, _23473_);
  or _74169_ (_23498_, _23497_, _06848_);
  and _74170_ (_23499_, _23498_, _23495_);
  or _74171_ (_23500_, _23499_, _06219_);
  or _74172_ (_23501_, _23482_, _06220_);
  and _74173_ (_23502_, _23501_, _06040_);
  and _74174_ (_23503_, _23502_, _23500_);
  and _74175_ (_23504_, _15278_, _08341_);
  or _74176_ (_23505_, _23504_, _23490_);
  and _74177_ (_23506_, _23505_, _06039_);
  or _74178_ (_23507_, _23506_, _06032_);
  or _74179_ (_23509_, _23507_, _23503_);
  or _74180_ (_23510_, _23490_, _15310_);
  and _74181_ (_23511_, _23510_, _23492_);
  or _74182_ (_23512_, _23511_, _06033_);
  and _74183_ (_23513_, _23512_, _06027_);
  and _74184_ (_23514_, _23513_, _23509_);
  or _74185_ (_23515_, _23490_, _15326_);
  and _74186_ (_23516_, _23515_, _06026_);
  and _74187_ (_23517_, _23516_, _23492_);
  or _74188_ (_23518_, _23517_, _09818_);
  or _74189_ (_23520_, _23518_, _23514_);
  and _74190_ (_23521_, _09178_, _07648_);
  or _74191_ (_23522_, _23473_, _07012_);
  or _74192_ (_23523_, _23522_, _23521_);
  or _74193_ (_23524_, _23497_, _09827_);
  and _74194_ (_23525_, _23524_, _05669_);
  and _74195_ (_23526_, _23525_, _23523_);
  and _74196_ (_23527_, _23526_, _23520_);
  and _74197_ (_23528_, _15382_, _07648_);
  or _74198_ (_23529_, _23528_, _23473_);
  and _74199_ (_23531_, _23529_, _09833_);
  or _74200_ (_23532_, _23531_, _06019_);
  or _74201_ (_23533_, _23532_, _23527_);
  and _74202_ (_23534_, _23533_, _23477_);
  or _74203_ (_23535_, _23534_, _06112_);
  and _74204_ (_23536_, _15399_, _07648_);
  or _74205_ (_23537_, _23473_, _08751_);
  or _74206_ (_23538_, _23537_, _23536_);
  and _74207_ (_23539_, _23538_, _08756_);
  and _74208_ (_23540_, _23539_, _23535_);
  and _74209_ (_23541_, _10980_, _07648_);
  or _74210_ (_23542_, _23541_, _23473_);
  and _74211_ (_23543_, _23542_, _06284_);
  or _74212_ (_23544_, _23543_, _23540_);
  and _74213_ (_23545_, _23544_, _07032_);
  or _74214_ (_23546_, _23473_, _07886_);
  and _74215_ (_23547_, _23475_, _06108_);
  and _74216_ (_23548_, _23547_, _23546_);
  or _74217_ (_23549_, _23548_, _23545_);
  and _74218_ (_23550_, _23549_, _06278_);
  and _74219_ (_23552_, _23482_, _06277_);
  and _74220_ (_23553_, _23552_, _23546_);
  or _74221_ (_23554_, _23553_, _06130_);
  or _74222_ (_23555_, _23554_, _23550_);
  and _74223_ (_23556_, _15396_, _07648_);
  or _74224_ (_23557_, _23473_, _08777_);
  or _74225_ (_23558_, _23557_, _23556_);
  and _74226_ (_23559_, _23558_, _08782_);
  and _74227_ (_23560_, _23559_, _23555_);
  nor _74228_ (_23561_, _10979_, _11605_);
  or _74229_ (_23563_, _23561_, _23473_);
  and _74230_ (_23564_, _23563_, _06292_);
  or _74231_ (_23565_, _23564_, _06316_);
  or _74232_ (_23566_, _23565_, _23560_);
  or _74233_ (_23567_, _23479_, _06718_);
  and _74234_ (_23568_, _23567_, _05653_);
  and _74235_ (_23569_, _23568_, _23566_);
  and _74236_ (_23570_, _23505_, _05652_);
  or _74237_ (_23571_, _23570_, _06047_);
  or _74238_ (_23572_, _23571_, _23569_);
  and _74239_ (_23573_, _15451_, _07648_);
  or _74240_ (_23574_, _23473_, _06048_);
  or _74241_ (_23575_, _23574_, _23573_);
  and _74242_ (_23576_, _23575_, _01336_);
  and _74243_ (_23577_, _23576_, _23572_);
  or _74244_ (_23578_, _23577_, _23472_);
  and _74245_ (_43397_, _23578_, _42882_);
  not _74246_ (_23579_, \oc8051_golden_model_1.TH1 [0]);
  nor _74247_ (_23580_, _01336_, _23579_);
  nand _74248_ (_23581_, _10995_, _07670_);
  nor _74249_ (_23583_, _07670_, _23579_);
  nor _74250_ (_23584_, _23583_, _06278_);
  nand _74251_ (_23585_, _23584_, _23581_);
  and _74252_ (_23586_, _09120_, _07670_);
  or _74253_ (_23587_, _23583_, _07012_);
  or _74254_ (_23588_, _23587_, _23586_);
  and _74255_ (_23589_, _07670_, _06931_);
  nor _74256_ (_23590_, _23589_, _23583_);
  nand _74257_ (_23591_, _23590_, _09815_);
  nor _74258_ (_23592_, _08127_, _11707_);
  or _74259_ (_23594_, _23592_, _23583_);
  or _74260_ (_23595_, _23594_, _06954_);
  and _74261_ (_23596_, _07670_, \oc8051_golden_model_1.ACC [0]);
  nor _74262_ (_23597_, _23596_, _23583_);
  nor _74263_ (_23598_, _23597_, _06939_);
  nor _74264_ (_23599_, _06938_, _23579_);
  or _74265_ (_23600_, _23599_, _06102_);
  or _74266_ (_23601_, _23600_, _23598_);
  and _74267_ (_23602_, _23601_, _06848_);
  and _74268_ (_23603_, _23602_, _23595_);
  nor _74269_ (_23605_, _23590_, _06848_);
  or _74270_ (_23606_, _23605_, _23603_);
  nand _74271_ (_23607_, _23606_, _06220_);
  or _74272_ (_23608_, _23597_, _06220_);
  and _74273_ (_23609_, _23608_, _09817_);
  nand _74274_ (_23610_, _23609_, _23607_);
  and _74275_ (_23611_, _23610_, _23591_);
  and _74276_ (_23612_, _23611_, _23588_);
  or _74277_ (_23613_, _23612_, _09833_);
  and _74278_ (_23614_, _14186_, _07670_);
  or _74279_ (_23616_, _23614_, _23583_);
  or _74280_ (_23617_, _23616_, _05669_);
  and _74281_ (_23618_, _23617_, _06020_);
  and _74282_ (_23619_, _23618_, _23613_);
  and _74283_ (_23620_, _07670_, _08672_);
  or _74284_ (_23621_, _23620_, _23583_);
  and _74285_ (_23622_, _23621_, _06019_);
  or _74286_ (_23623_, _23622_, _06112_);
  or _74287_ (_23624_, _23623_, _23619_);
  and _74288_ (_23625_, _14086_, _07670_);
  or _74289_ (_23627_, _23583_, _08751_);
  or _74290_ (_23628_, _23627_, _23625_);
  and _74291_ (_23629_, _23628_, _08756_);
  and _74292_ (_23630_, _23629_, _23624_);
  nor _74293_ (_23631_, _12302_, _11707_);
  or _74294_ (_23632_, _23631_, _23583_);
  and _74295_ (_23633_, _23581_, _06284_);
  and _74296_ (_23634_, _23633_, _23632_);
  or _74297_ (_23635_, _23634_, _23630_);
  and _74298_ (_23636_, _23635_, _07032_);
  nand _74299_ (_23638_, _23621_, _06108_);
  nor _74300_ (_23639_, _23638_, _23592_);
  or _74301_ (_23640_, _23639_, _06277_);
  or _74302_ (_23641_, _23640_, _23636_);
  and _74303_ (_23642_, _23641_, _23585_);
  or _74304_ (_23643_, _23642_, _06130_);
  and _74305_ (_23644_, _14083_, _07670_);
  or _74306_ (_23645_, _23583_, _08777_);
  or _74307_ (_23646_, _23645_, _23644_);
  and _74308_ (_23647_, _23646_, _08782_);
  and _74309_ (_23649_, _23647_, _23643_);
  and _74310_ (_23650_, _23632_, _06292_);
  or _74311_ (_23651_, _23650_, _19256_);
  or _74312_ (_23652_, _23651_, _23649_);
  or _74313_ (_23653_, _23594_, _06408_);
  and _74314_ (_23654_, _23653_, _01336_);
  and _74315_ (_23655_, _23654_, _23652_);
  or _74316_ (_23656_, _23655_, _23580_);
  and _74317_ (_43399_, _23656_, _42882_);
  not _74318_ (_23657_, \oc8051_golden_model_1.TH1 [1]);
  nor _74319_ (_23659_, _01336_, _23657_);
  or _74320_ (_23660_, _14367_, _11707_);
  or _74321_ (_23661_, _07670_, \oc8051_golden_model_1.TH1 [1]);
  and _74322_ (_23662_, _23661_, _09833_);
  and _74323_ (_23663_, _23662_, _23660_);
  and _74324_ (_23664_, _09075_, _07670_);
  nor _74325_ (_23665_, _07670_, _23657_);
  or _74326_ (_23666_, _23665_, _07012_);
  or _74327_ (_23667_, _23666_, _23664_);
  and _74328_ (_23668_, _14284_, _07670_);
  not _74329_ (_23670_, _23668_);
  and _74330_ (_23671_, _23670_, _23661_);
  or _74331_ (_23672_, _23671_, _06954_);
  and _74332_ (_23673_, _07670_, \oc8051_golden_model_1.ACC [1]);
  or _74333_ (_23674_, _23673_, _23665_);
  and _74334_ (_23675_, _23674_, _06938_);
  nor _74335_ (_23676_, _06938_, _23657_);
  or _74336_ (_23677_, _23676_, _06102_);
  or _74337_ (_23678_, _23677_, _23675_);
  and _74338_ (_23679_, _23678_, _06848_);
  and _74339_ (_23680_, _23679_, _23672_);
  nor _74340_ (_23681_, _11707_, _07132_);
  or _74341_ (_23682_, _23681_, _23665_);
  and _74342_ (_23683_, _23682_, _06239_);
  or _74343_ (_23684_, _23683_, _23680_);
  and _74344_ (_23685_, _23684_, _06220_);
  and _74345_ (_23686_, _23674_, _06219_);
  or _74346_ (_23687_, _23686_, _09818_);
  or _74347_ (_23688_, _23687_, _23685_);
  or _74348_ (_23689_, _23682_, _09827_);
  and _74349_ (_23690_, _23689_, _05669_);
  and _74350_ (_23691_, _23690_, _23688_);
  and _74351_ (_23692_, _23691_, _23667_);
  or _74352_ (_23693_, _23692_, _23663_);
  and _74353_ (_23694_, _23693_, _06020_);
  nand _74354_ (_23695_, _07670_, _06832_);
  and _74355_ (_23696_, _23661_, _06019_);
  and _74356_ (_23697_, _23696_, _23695_);
  or _74357_ (_23698_, _23697_, _23694_);
  and _74358_ (_23699_, _23698_, _08751_);
  or _74359_ (_23701_, _14263_, _11707_);
  and _74360_ (_23702_, _23661_, _06112_);
  and _74361_ (_23703_, _23702_, _23701_);
  or _74362_ (_23704_, _23703_, _06284_);
  or _74363_ (_23705_, _23704_, _23699_);
  nor _74364_ (_23706_, _10993_, _11707_);
  or _74365_ (_23707_, _23706_, _23665_);
  nand _74366_ (_23708_, _10992_, _07670_);
  and _74367_ (_23709_, _23708_, _23707_);
  or _74368_ (_23710_, _23709_, _08756_);
  and _74369_ (_23712_, _23710_, _07032_);
  and _74370_ (_23713_, _23712_, _23705_);
  or _74371_ (_23714_, _14261_, _11707_);
  and _74372_ (_23715_, _23661_, _06108_);
  and _74373_ (_23716_, _23715_, _23714_);
  or _74374_ (_23717_, _23716_, _06277_);
  or _74375_ (_23718_, _23717_, _23713_);
  nor _74376_ (_23719_, _23665_, _06278_);
  nand _74377_ (_23720_, _23719_, _23708_);
  and _74378_ (_23721_, _23720_, _08777_);
  and _74379_ (_23723_, _23721_, _23718_);
  or _74380_ (_23724_, _23695_, _08078_);
  and _74381_ (_23725_, _23661_, _06130_);
  and _74382_ (_23726_, _23725_, _23724_);
  or _74383_ (_23727_, _23726_, _06292_);
  or _74384_ (_23728_, _23727_, _23723_);
  or _74385_ (_23729_, _23707_, _08782_);
  and _74386_ (_23730_, _23729_, _06718_);
  and _74387_ (_23731_, _23730_, _23728_);
  and _74388_ (_23732_, _23671_, _06316_);
  or _74389_ (_23734_, _23732_, _06047_);
  or _74390_ (_23735_, _23734_, _23731_);
  or _74391_ (_23736_, _23665_, _06048_);
  or _74392_ (_23737_, _23736_, _23668_);
  and _74393_ (_23738_, _23737_, _01336_);
  and _74394_ (_23739_, _23738_, _23735_);
  or _74395_ (_23740_, _23739_, _23659_);
  and _74396_ (_43400_, _23740_, _42882_);
  not _74397_ (_23741_, \oc8051_golden_model_1.TH1 [2]);
  nor _74398_ (_23742_, _01336_, _23741_);
  and _74399_ (_23744_, _09182_, _07670_);
  nor _74400_ (_23745_, _07670_, _23741_);
  or _74401_ (_23746_, _23745_, _07012_);
  or _74402_ (_23747_, _23746_, _23744_);
  nor _74403_ (_23748_, _11707_, _07530_);
  nor _74404_ (_23749_, _23748_, _23745_);
  nand _74405_ (_23750_, _23749_, _09815_);
  and _74406_ (_23751_, _14493_, _07670_);
  or _74407_ (_23752_, _23751_, _23745_);
  or _74408_ (_23753_, _23752_, _06954_);
  and _74409_ (_23755_, _07670_, \oc8051_golden_model_1.ACC [2]);
  nor _74410_ (_23756_, _23755_, _23745_);
  nor _74411_ (_23757_, _23756_, _06939_);
  nor _74412_ (_23758_, _06938_, _23741_);
  or _74413_ (_23759_, _23758_, _06102_);
  or _74414_ (_23760_, _23759_, _23757_);
  and _74415_ (_23761_, _23760_, _06848_);
  and _74416_ (_23762_, _23761_, _23753_);
  nor _74417_ (_23763_, _23749_, _06848_);
  or _74418_ (_23764_, _23763_, _23762_);
  nand _74419_ (_23766_, _23764_, _06220_);
  or _74420_ (_23767_, _23756_, _06220_);
  and _74421_ (_23768_, _23767_, _09817_);
  nand _74422_ (_23769_, _23768_, _23766_);
  and _74423_ (_23770_, _23769_, _23750_);
  and _74424_ (_23771_, _23770_, _23747_);
  or _74425_ (_23772_, _23771_, _09833_);
  and _74426_ (_23773_, _14580_, _07670_);
  or _74427_ (_23774_, _23745_, _05669_);
  or _74428_ (_23775_, _23774_, _23773_);
  and _74429_ (_23777_, _23775_, _06020_);
  and _74430_ (_23778_, _23777_, _23772_);
  and _74431_ (_23779_, _07670_, _08730_);
  or _74432_ (_23780_, _23779_, _23745_);
  and _74433_ (_23781_, _23780_, _06019_);
  or _74434_ (_23782_, _23781_, _06112_);
  or _74435_ (_23783_, _23782_, _23778_);
  and _74436_ (_23784_, _14596_, _07670_);
  or _74437_ (_23785_, _23784_, _23745_);
  or _74438_ (_23786_, _23785_, _08751_);
  and _74439_ (_23788_, _23786_, _08756_);
  and _74440_ (_23789_, _23788_, _23783_);
  and _74441_ (_23790_, _10991_, _07670_);
  or _74442_ (_23791_, _23790_, _23745_);
  and _74443_ (_23792_, _23791_, _06284_);
  or _74444_ (_23793_, _23792_, _23789_);
  and _74445_ (_23794_, _23793_, _07032_);
  or _74446_ (_23795_, _23745_, _08177_);
  and _74447_ (_23796_, _23780_, _06108_);
  and _74448_ (_23797_, _23796_, _23795_);
  or _74449_ (_23799_, _23797_, _23794_);
  and _74450_ (_23800_, _23799_, _06278_);
  nor _74451_ (_23801_, _23756_, _06278_);
  and _74452_ (_23802_, _23801_, _23795_);
  or _74453_ (_23803_, _23802_, _06130_);
  or _74454_ (_23804_, _23803_, _23800_);
  and _74455_ (_23805_, _14593_, _07670_);
  or _74456_ (_23806_, _23745_, _08777_);
  or _74457_ (_23807_, _23806_, _23805_);
  and _74458_ (_23808_, _23807_, _08782_);
  and _74459_ (_23810_, _23808_, _23804_);
  nor _74460_ (_23811_, _10990_, _11707_);
  or _74461_ (_23812_, _23811_, _23745_);
  and _74462_ (_23813_, _23812_, _06292_);
  or _74463_ (_23814_, _23813_, _23810_);
  and _74464_ (_23815_, _23814_, _06718_);
  and _74465_ (_23816_, _23752_, _06316_);
  or _74466_ (_23817_, _23816_, _06047_);
  or _74467_ (_23818_, _23817_, _23815_);
  and _74468_ (_23819_, _14657_, _07670_);
  or _74469_ (_23821_, _23745_, _06048_);
  or _74470_ (_23822_, _23821_, _23819_);
  and _74471_ (_23823_, _23822_, _01336_);
  and _74472_ (_23824_, _23823_, _23818_);
  or _74473_ (_23825_, _23824_, _23742_);
  and _74474_ (_43401_, _23825_, _42882_);
  not _74475_ (_23826_, \oc8051_golden_model_1.TH1 [3]);
  nor _74476_ (_23827_, _01336_, _23826_);
  nor _74477_ (_23828_, _07670_, _23826_);
  or _74478_ (_23829_, _23828_, _08029_);
  and _74479_ (_23831_, _07670_, _08662_);
  or _74480_ (_23832_, _23831_, _23828_);
  and _74481_ (_23833_, _23832_, _06108_);
  and _74482_ (_23834_, _23833_, _23829_);
  and _74483_ (_23835_, _09181_, _07670_);
  or _74484_ (_23836_, _23828_, _07012_);
  or _74485_ (_23837_, _23836_, _23835_);
  nor _74486_ (_23838_, _11707_, _07353_);
  nor _74487_ (_23839_, _23838_, _23828_);
  nand _74488_ (_23840_, _23839_, _09815_);
  and _74489_ (_23842_, _14672_, _07670_);
  or _74490_ (_23843_, _23842_, _23828_);
  or _74491_ (_23844_, _23843_, _06954_);
  and _74492_ (_23845_, _07670_, \oc8051_golden_model_1.ACC [3]);
  nor _74493_ (_23846_, _23845_, _23828_);
  nor _74494_ (_23847_, _23846_, _06939_);
  nor _74495_ (_23848_, _06938_, _23826_);
  or _74496_ (_23849_, _23848_, _06102_);
  or _74497_ (_23850_, _23849_, _23847_);
  and _74498_ (_23851_, _23850_, _06848_);
  and _74499_ (_23853_, _23851_, _23844_);
  nor _74500_ (_23854_, _23839_, _06848_);
  or _74501_ (_23855_, _23854_, _23853_);
  nand _74502_ (_23856_, _23855_, _06220_);
  or _74503_ (_23857_, _23846_, _06220_);
  and _74504_ (_23858_, _23857_, _09817_);
  nand _74505_ (_23859_, _23858_, _23856_);
  and _74506_ (_23860_, _23859_, _23840_);
  and _74507_ (_23861_, _23860_, _23837_);
  or _74508_ (_23862_, _23861_, _09833_);
  and _74509_ (_23864_, _14778_, _07670_);
  or _74510_ (_23865_, _23864_, _23828_);
  or _74511_ (_23866_, _23865_, _05669_);
  and _74512_ (_23867_, _23866_, _06020_);
  and _74513_ (_23868_, _23867_, _23862_);
  and _74514_ (_23869_, _23832_, _06019_);
  or _74515_ (_23870_, _23869_, _06112_);
  or _74516_ (_23871_, _23870_, _23868_);
  and _74517_ (_23872_, _14793_, _07670_);
  or _74518_ (_23873_, _23828_, _08751_);
  or _74519_ (_23875_, _23873_, _23872_);
  and _74520_ (_23876_, _23875_, _08756_);
  and _74521_ (_23877_, _23876_, _23871_);
  and _74522_ (_23878_, _12299_, _07670_);
  or _74523_ (_23879_, _23878_, _23828_);
  and _74524_ (_23880_, _23879_, _06284_);
  or _74525_ (_23881_, _23880_, _23877_);
  and _74526_ (_23882_, _23881_, _07032_);
  or _74527_ (_23883_, _23882_, _23834_);
  and _74528_ (_23884_, _23883_, _06278_);
  nor _74529_ (_23885_, _23846_, _06278_);
  and _74530_ (_23886_, _23885_, _23829_);
  or _74531_ (_23887_, _23886_, _06130_);
  or _74532_ (_23888_, _23887_, _23884_);
  and _74533_ (_23889_, _14792_, _07670_);
  or _74534_ (_23890_, _23828_, _08777_);
  or _74535_ (_23891_, _23890_, _23889_);
  and _74536_ (_23892_, _23891_, _08782_);
  and _74537_ (_23893_, _23892_, _23888_);
  nor _74538_ (_23894_, _10988_, _11707_);
  or _74539_ (_23897_, _23894_, _23828_);
  and _74540_ (_23898_, _23897_, _06292_);
  or _74541_ (_23899_, _23898_, _23893_);
  and _74542_ (_23900_, _23899_, _06718_);
  and _74543_ (_23901_, _23843_, _06316_);
  or _74544_ (_23902_, _23901_, _06047_);
  or _74545_ (_23903_, _23902_, _23900_);
  and _74546_ (_23904_, _14849_, _07670_);
  or _74547_ (_23905_, _23828_, _06048_);
  or _74548_ (_23906_, _23905_, _23904_);
  and _74549_ (_23908_, _23906_, _01336_);
  and _74550_ (_23909_, _23908_, _23903_);
  or _74551_ (_23910_, _23909_, _23827_);
  and _74552_ (_43403_, _23910_, _42882_);
  and _74553_ (_23911_, _01340_, \oc8051_golden_model_1.TH1 [4]);
  and _74554_ (_23912_, _11707_, \oc8051_golden_model_1.TH1 [4]);
  or _74555_ (_23913_, _23912_, _08273_);
  and _74556_ (_23914_, _08665_, _07670_);
  or _74557_ (_23915_, _23914_, _23912_);
  and _74558_ (_23916_, _23915_, _06108_);
  and _74559_ (_23918_, _23916_, _23913_);
  or _74560_ (_23919_, _23915_, _06020_);
  and _74561_ (_23920_, _14887_, _07670_);
  or _74562_ (_23921_, _23920_, _23912_);
  or _74563_ (_23922_, _23921_, _06954_);
  and _74564_ (_23923_, _07670_, \oc8051_golden_model_1.ACC [4]);
  or _74565_ (_23924_, _23923_, _23912_);
  and _74566_ (_23925_, _23924_, _06938_);
  and _74567_ (_23926_, _06939_, \oc8051_golden_model_1.TH1 [4]);
  or _74568_ (_23927_, _23926_, _06102_);
  or _74569_ (_23929_, _23927_, _23925_);
  and _74570_ (_23930_, _23929_, _06848_);
  and _74571_ (_23931_, _23930_, _23922_);
  nor _74572_ (_23932_, _08270_, _11707_);
  or _74573_ (_23933_, _23932_, _23912_);
  and _74574_ (_23934_, _23933_, _06239_);
  or _74575_ (_23935_, _23934_, _23931_);
  and _74576_ (_23936_, _23935_, _06220_);
  and _74577_ (_23937_, _23924_, _06219_);
  or _74578_ (_23938_, _23937_, _09818_);
  or _74579_ (_23940_, _23938_, _23936_);
  and _74580_ (_23941_, _09180_, _07670_);
  or _74581_ (_23942_, _23912_, _07012_);
  or _74582_ (_23943_, _23942_, _23941_);
  or _74583_ (_23944_, _23933_, _09827_);
  and _74584_ (_23945_, _23944_, _05669_);
  and _74585_ (_23946_, _23945_, _23943_);
  and _74586_ (_23947_, _23946_, _23940_);
  and _74587_ (_23948_, _14983_, _07670_);
  or _74588_ (_23949_, _23948_, _23912_);
  and _74589_ (_23951_, _23949_, _09833_);
  or _74590_ (_23952_, _23951_, _06019_);
  or _74591_ (_23953_, _23952_, _23947_);
  and _74592_ (_23954_, _23953_, _23919_);
  or _74593_ (_23955_, _23954_, _06112_);
  and _74594_ (_23956_, _14876_, _07670_);
  or _74595_ (_23957_, _23912_, _08751_);
  or _74596_ (_23958_, _23957_, _23956_);
  and _74597_ (_23959_, _23958_, _08756_);
  and _74598_ (_23960_, _23959_, _23955_);
  and _74599_ (_23962_, _10986_, _07670_);
  or _74600_ (_23963_, _23962_, _23912_);
  and _74601_ (_23964_, _23963_, _06284_);
  or _74602_ (_23965_, _23964_, _23960_);
  and _74603_ (_23966_, _23965_, _07032_);
  or _74604_ (_23967_, _23966_, _23918_);
  and _74605_ (_23968_, _23967_, _06278_);
  and _74606_ (_23969_, _23924_, _06277_);
  and _74607_ (_23970_, _23969_, _23913_);
  or _74608_ (_23971_, _23970_, _06130_);
  or _74609_ (_23973_, _23971_, _23968_);
  and _74610_ (_23974_, _14873_, _07670_);
  or _74611_ (_23975_, _23912_, _08777_);
  or _74612_ (_23976_, _23975_, _23974_);
  and _74613_ (_23977_, _23976_, _08782_);
  and _74614_ (_23978_, _23977_, _23973_);
  nor _74615_ (_23979_, _10985_, _11707_);
  or _74616_ (_23980_, _23979_, _23912_);
  and _74617_ (_23981_, _23980_, _06292_);
  or _74618_ (_23982_, _23981_, _23978_);
  and _74619_ (_23984_, _23982_, _06718_);
  and _74620_ (_23985_, _23921_, _06316_);
  or _74621_ (_23986_, _23985_, _06047_);
  or _74622_ (_23987_, _23986_, _23984_);
  and _74623_ (_23988_, _15055_, _07670_);
  or _74624_ (_23989_, _23912_, _06048_);
  or _74625_ (_23990_, _23989_, _23988_);
  and _74626_ (_23991_, _23990_, _01336_);
  and _74627_ (_23992_, _23991_, _23987_);
  or _74628_ (_23993_, _23992_, _23911_);
  and _74629_ (_43404_, _23993_, _42882_);
  and _74630_ (_23995_, _01340_, \oc8051_golden_model_1.TH1 [5]);
  and _74631_ (_23996_, _11707_, \oc8051_golden_model_1.TH1 [5]);
  or _74632_ (_23997_, _23996_, _07980_);
  and _74633_ (_23998_, _08652_, _07670_);
  or _74634_ (_23999_, _23998_, _23996_);
  and _74635_ (_24000_, _23999_, _06108_);
  and _74636_ (_24001_, _24000_, _23997_);
  or _74637_ (_24002_, _23999_, _06020_);
  and _74638_ (_24003_, _15093_, _07670_);
  or _74639_ (_24005_, _24003_, _23996_);
  or _74640_ (_24006_, _24005_, _06954_);
  and _74641_ (_24007_, _07670_, \oc8051_golden_model_1.ACC [5]);
  or _74642_ (_24008_, _24007_, _23996_);
  and _74643_ (_24009_, _24008_, _06938_);
  and _74644_ (_24010_, _06939_, \oc8051_golden_model_1.TH1 [5]);
  or _74645_ (_24011_, _24010_, _06102_);
  or _74646_ (_24012_, _24011_, _24009_);
  and _74647_ (_24013_, _24012_, _06848_);
  and _74648_ (_24014_, _24013_, _24006_);
  nor _74649_ (_24016_, _07977_, _11707_);
  or _74650_ (_24017_, _24016_, _23996_);
  and _74651_ (_24018_, _24017_, _06239_);
  or _74652_ (_24019_, _24018_, _24014_);
  and _74653_ (_24020_, _24019_, _06220_);
  and _74654_ (_24021_, _24008_, _06219_);
  or _74655_ (_24022_, _24021_, _09818_);
  or _74656_ (_24023_, _24022_, _24020_);
  and _74657_ (_24024_, _09179_, _07670_);
  or _74658_ (_24025_, _23996_, _07012_);
  or _74659_ (_24027_, _24025_, _24024_);
  or _74660_ (_24028_, _24017_, _09827_);
  and _74661_ (_24029_, _24028_, _05669_);
  and _74662_ (_24030_, _24029_, _24027_);
  and _74663_ (_24031_, _24030_, _24023_);
  and _74664_ (_24032_, _15179_, _07670_);
  or _74665_ (_24033_, _24032_, _23996_);
  and _74666_ (_24034_, _24033_, _09833_);
  or _74667_ (_24035_, _24034_, _06019_);
  or _74668_ (_24036_, _24035_, _24031_);
  and _74669_ (_24038_, _24036_, _24002_);
  or _74670_ (_24039_, _24038_, _06112_);
  and _74671_ (_24040_, _15195_, _07670_);
  or _74672_ (_24041_, _23996_, _08751_);
  or _74673_ (_24042_, _24041_, _24040_);
  and _74674_ (_24043_, _24042_, _08756_);
  and _74675_ (_24044_, _24043_, _24039_);
  and _74676_ (_24045_, _12306_, _07670_);
  or _74677_ (_24046_, _24045_, _23996_);
  and _74678_ (_24047_, _24046_, _06284_);
  or _74679_ (_24049_, _24047_, _24044_);
  and _74680_ (_24050_, _24049_, _07032_);
  or _74681_ (_24051_, _24050_, _24001_);
  and _74682_ (_24052_, _24051_, _06278_);
  and _74683_ (_24053_, _24008_, _06277_);
  and _74684_ (_24054_, _24053_, _23997_);
  or _74685_ (_24055_, _24054_, _06130_);
  or _74686_ (_24056_, _24055_, _24052_);
  and _74687_ (_24057_, _15194_, _07670_);
  or _74688_ (_24058_, _23996_, _08777_);
  or _74689_ (_24060_, _24058_, _24057_);
  and _74690_ (_24061_, _24060_, _08782_);
  and _74691_ (_24062_, _24061_, _24056_);
  nor _74692_ (_24063_, _10982_, _11707_);
  or _74693_ (_24064_, _24063_, _23996_);
  and _74694_ (_24065_, _24064_, _06292_);
  or _74695_ (_24066_, _24065_, _24062_);
  and _74696_ (_24067_, _24066_, _06718_);
  and _74697_ (_24068_, _24005_, _06316_);
  or _74698_ (_24069_, _24068_, _06047_);
  or _74699_ (_24070_, _24069_, _24067_);
  and _74700_ (_24071_, _15253_, _07670_);
  or _74701_ (_24072_, _23996_, _06048_);
  or _74702_ (_24073_, _24072_, _24071_);
  and _74703_ (_24074_, _24073_, _01336_);
  and _74704_ (_24075_, _24074_, _24070_);
  or _74705_ (_24076_, _24075_, _23995_);
  and _74706_ (_43405_, _24076_, _42882_);
  and _74707_ (_24077_, _01340_, \oc8051_golden_model_1.TH1 [6]);
  and _74708_ (_24078_, _11707_, \oc8051_golden_model_1.TH1 [6]);
  or _74709_ (_24081_, _24078_, _07886_);
  and _74710_ (_24082_, _15389_, _07670_);
  or _74711_ (_24083_, _24082_, _24078_);
  and _74712_ (_24084_, _24083_, _06108_);
  and _74713_ (_24085_, _24084_, _24081_);
  or _74714_ (_24086_, _24083_, _06020_);
  and _74715_ (_24087_, _15293_, _07670_);
  or _74716_ (_24088_, _24087_, _24078_);
  or _74717_ (_24089_, _24088_, _06954_);
  and _74718_ (_24090_, _07670_, \oc8051_golden_model_1.ACC [6]);
  or _74719_ (_24092_, _24090_, _24078_);
  and _74720_ (_24093_, _24092_, _06938_);
  and _74721_ (_24094_, _06939_, \oc8051_golden_model_1.TH1 [6]);
  or _74722_ (_24095_, _24094_, _06102_);
  or _74723_ (_24096_, _24095_, _24093_);
  and _74724_ (_24097_, _24096_, _06848_);
  and _74725_ (_24098_, _24097_, _24089_);
  nor _74726_ (_24099_, _07883_, _11707_);
  or _74727_ (_24100_, _24099_, _24078_);
  and _74728_ (_24101_, _24100_, _06239_);
  or _74729_ (_24103_, _24101_, _24098_);
  and _74730_ (_24104_, _24103_, _06220_);
  and _74731_ (_24105_, _24092_, _06219_);
  or _74732_ (_24106_, _24105_, _09818_);
  or _74733_ (_24107_, _24106_, _24104_);
  and _74734_ (_24108_, _09178_, _07670_);
  or _74735_ (_24109_, _24078_, _07012_);
  or _74736_ (_24110_, _24109_, _24108_);
  or _74737_ (_24111_, _24100_, _09827_);
  and _74738_ (_24112_, _24111_, _05669_);
  and _74739_ (_24114_, _24112_, _24110_);
  and _74740_ (_24115_, _24114_, _24107_);
  and _74741_ (_24116_, _15382_, _07670_);
  or _74742_ (_24117_, _24116_, _24078_);
  and _74743_ (_24118_, _24117_, _09833_);
  or _74744_ (_24119_, _24118_, _06019_);
  or _74745_ (_24120_, _24119_, _24115_);
  and _74746_ (_24121_, _24120_, _24086_);
  or _74747_ (_24122_, _24121_, _06112_);
  and _74748_ (_24123_, _15399_, _07670_);
  or _74749_ (_24125_, _24123_, _24078_);
  or _74750_ (_24126_, _24125_, _08751_);
  and _74751_ (_24127_, _24126_, _08756_);
  and _74752_ (_24128_, _24127_, _24122_);
  and _74753_ (_24129_, _10980_, _07670_);
  or _74754_ (_24130_, _24129_, _24078_);
  and _74755_ (_24131_, _24130_, _06284_);
  or _74756_ (_24132_, _24131_, _24128_);
  and _74757_ (_24133_, _24132_, _07032_);
  or _74758_ (_24134_, _24133_, _24085_);
  and _74759_ (_24136_, _24134_, _06278_);
  and _74760_ (_24137_, _24092_, _06277_);
  and _74761_ (_24138_, _24137_, _24081_);
  or _74762_ (_24139_, _24138_, _06130_);
  or _74763_ (_24140_, _24139_, _24136_);
  and _74764_ (_24141_, _15396_, _07670_);
  or _74765_ (_24142_, _24078_, _08777_);
  or _74766_ (_24143_, _24142_, _24141_);
  and _74767_ (_24144_, _24143_, _08782_);
  and _74768_ (_24145_, _24144_, _24140_);
  nor _74769_ (_24147_, _10979_, _11707_);
  or _74770_ (_24148_, _24147_, _24078_);
  and _74771_ (_24149_, _24148_, _06292_);
  or _74772_ (_24150_, _24149_, _24145_);
  and _74773_ (_24151_, _24150_, _06718_);
  and _74774_ (_24152_, _24088_, _06316_);
  or _74775_ (_24153_, _24152_, _06047_);
  or _74776_ (_24154_, _24153_, _24151_);
  and _74777_ (_24155_, _15451_, _07670_);
  or _74778_ (_24156_, _24078_, _06048_);
  or _74779_ (_24158_, _24156_, _24155_);
  and _74780_ (_24159_, _24158_, _01336_);
  and _74781_ (_24160_, _24159_, _24154_);
  or _74782_ (_24161_, _24160_, _24077_);
  and _74783_ (_43406_, _24161_, _42882_);
  not _74784_ (_24162_, \oc8051_golden_model_1.TH0 [0]);
  nor _74785_ (_24163_, _01336_, _24162_);
  nand _74786_ (_24164_, _10995_, _07663_);
  nor _74787_ (_24165_, _07663_, _24162_);
  nor _74788_ (_24166_, _24165_, _06278_);
  nand _74789_ (_24168_, _24166_, _24164_);
  and _74790_ (_24169_, _09120_, _07663_);
  or _74791_ (_24170_, _24165_, _07012_);
  or _74792_ (_24171_, _24170_, _24169_);
  and _74793_ (_24172_, _07663_, _06931_);
  nor _74794_ (_24173_, _24172_, _24165_);
  nand _74795_ (_24174_, _24173_, _09815_);
  nor _74796_ (_24175_, _08127_, _11784_);
  or _74797_ (_24176_, _24175_, _24165_);
  and _74798_ (_24177_, _24176_, _06102_);
  nor _74799_ (_24179_, _06938_, _24162_);
  and _74800_ (_24180_, _07663_, \oc8051_golden_model_1.ACC [0]);
  nor _74801_ (_24181_, _24180_, _24165_);
  nor _74802_ (_24182_, _24181_, _06939_);
  or _74803_ (_24183_, _24182_, _24179_);
  and _74804_ (_24184_, _24183_, _06954_);
  or _74805_ (_24185_, _24184_, _06239_);
  or _74806_ (_24186_, _24185_, _24177_);
  nand _74807_ (_24187_, _24173_, _06239_);
  and _74808_ (_24188_, _24187_, _06220_);
  nand _74809_ (_24190_, _24188_, _24186_);
  or _74810_ (_24191_, _24181_, _06220_);
  and _74811_ (_24192_, _24191_, _09817_);
  nand _74812_ (_24193_, _24192_, _24190_);
  and _74813_ (_24194_, _24193_, _24174_);
  and _74814_ (_24195_, _24194_, _24171_);
  or _74815_ (_24196_, _24195_, _09833_);
  and _74816_ (_24197_, _14186_, _07663_);
  or _74817_ (_24198_, _24165_, _05669_);
  or _74818_ (_24199_, _24198_, _24197_);
  and _74819_ (_24201_, _24199_, _06020_);
  and _74820_ (_24202_, _24201_, _24196_);
  and _74821_ (_24203_, _07663_, _08672_);
  or _74822_ (_24204_, _24203_, _24165_);
  and _74823_ (_24205_, _24204_, _06019_);
  or _74824_ (_24206_, _24205_, _06112_);
  or _74825_ (_24207_, _24206_, _24202_);
  and _74826_ (_24208_, _14086_, _07663_);
  or _74827_ (_24209_, _24165_, _08751_);
  or _74828_ (_24210_, _24209_, _24208_);
  and _74829_ (_24212_, _24210_, _08756_);
  and _74830_ (_24213_, _24212_, _24207_);
  nor _74831_ (_24214_, _12302_, _11784_);
  or _74832_ (_24215_, _24214_, _24165_);
  and _74833_ (_24216_, _24164_, _06284_);
  and _74834_ (_24217_, _24216_, _24215_);
  or _74835_ (_24218_, _24217_, _24213_);
  and _74836_ (_24219_, _24218_, _07032_);
  nand _74837_ (_24220_, _24204_, _06108_);
  nor _74838_ (_24221_, _24220_, _24175_);
  or _74839_ (_24223_, _24221_, _06277_);
  or _74840_ (_24224_, _24223_, _24219_);
  and _74841_ (_24225_, _24224_, _24168_);
  or _74842_ (_24226_, _24225_, _06130_);
  and _74843_ (_24227_, _14083_, _07663_);
  or _74844_ (_24228_, _24165_, _08777_);
  or _74845_ (_24229_, _24228_, _24227_);
  and _74846_ (_24230_, _24229_, _08782_);
  and _74847_ (_24231_, _24230_, _24226_);
  and _74848_ (_24232_, _24215_, _06292_);
  or _74849_ (_24234_, _24232_, _19256_);
  or _74850_ (_24235_, _24234_, _24231_);
  or _74851_ (_24236_, _24176_, _06408_);
  and _74852_ (_24237_, _24236_, _01336_);
  and _74853_ (_24238_, _24237_, _24235_);
  or _74854_ (_24239_, _24238_, _24163_);
  and _74855_ (_43408_, _24239_, _42882_);
  not _74856_ (_24240_, \oc8051_golden_model_1.TH0 [1]);
  nor _74857_ (_24241_, _01336_, _24240_);
  or _74858_ (_24242_, _14367_, _11784_);
  or _74859_ (_24244_, _07663_, \oc8051_golden_model_1.TH0 [1]);
  and _74860_ (_24245_, _24244_, _09833_);
  and _74861_ (_24246_, _24245_, _24242_);
  and _74862_ (_24247_, _09075_, _07663_);
  nor _74863_ (_24248_, _07663_, _24240_);
  or _74864_ (_24249_, _24248_, _07012_);
  or _74865_ (_24250_, _24249_, _24247_);
  and _74866_ (_24251_, _14284_, _07663_);
  not _74867_ (_24252_, _24251_);
  and _74868_ (_24253_, _24252_, _24244_);
  or _74869_ (_24255_, _24253_, _06954_);
  and _74870_ (_24256_, _07663_, \oc8051_golden_model_1.ACC [1]);
  or _74871_ (_24257_, _24256_, _24248_);
  and _74872_ (_24258_, _24257_, _06938_);
  nor _74873_ (_24259_, _06938_, _24240_);
  or _74874_ (_24260_, _24259_, _06102_);
  or _74875_ (_24261_, _24260_, _24258_);
  and _74876_ (_24262_, _24261_, _06848_);
  and _74877_ (_24263_, _24262_, _24255_);
  nor _74878_ (_24264_, _11784_, _07132_);
  or _74879_ (_24266_, _24264_, _24248_);
  and _74880_ (_24267_, _24266_, _06239_);
  or _74881_ (_24268_, _24267_, _24263_);
  and _74882_ (_24269_, _24268_, _06220_);
  and _74883_ (_24270_, _24257_, _06219_);
  or _74884_ (_24271_, _24270_, _09818_);
  or _74885_ (_24272_, _24271_, _24269_);
  or _74886_ (_24273_, _24266_, _09827_);
  and _74887_ (_24274_, _24273_, _05669_);
  and _74888_ (_24275_, _24274_, _24272_);
  and _74889_ (_24277_, _24275_, _24250_);
  or _74890_ (_24278_, _24277_, _24246_);
  and _74891_ (_24279_, _24278_, _06020_);
  nand _74892_ (_24280_, _07663_, _06832_);
  and _74893_ (_24281_, _24244_, _06019_);
  and _74894_ (_24282_, _24281_, _24280_);
  or _74895_ (_24283_, _24282_, _24279_);
  and _74896_ (_24284_, _24283_, _08751_);
  or _74897_ (_24285_, _14263_, _11784_);
  and _74898_ (_24286_, _24244_, _06112_);
  and _74899_ (_24288_, _24286_, _24285_);
  or _74900_ (_24289_, _24288_, _06284_);
  or _74901_ (_24290_, _24289_, _24284_);
  nor _74902_ (_24291_, _10993_, _11784_);
  or _74903_ (_24292_, _24291_, _24248_);
  nand _74904_ (_24293_, _10992_, _07663_);
  and _74905_ (_24294_, _24293_, _24292_);
  or _74906_ (_24295_, _24294_, _08756_);
  and _74907_ (_24296_, _24295_, _07032_);
  and _74908_ (_24297_, _24296_, _24290_);
  or _74909_ (_24299_, _14261_, _11784_);
  and _74910_ (_24300_, _24244_, _06108_);
  and _74911_ (_24301_, _24300_, _24299_);
  or _74912_ (_24302_, _24301_, _06277_);
  or _74913_ (_24303_, _24302_, _24297_);
  nor _74914_ (_24304_, _24248_, _06278_);
  nand _74915_ (_24305_, _24304_, _24293_);
  and _74916_ (_24306_, _24305_, _08777_);
  and _74917_ (_24307_, _24306_, _24303_);
  or _74918_ (_24308_, _24280_, _08078_);
  and _74919_ (_24310_, _24244_, _06130_);
  and _74920_ (_24311_, _24310_, _24308_);
  or _74921_ (_24312_, _24311_, _06292_);
  or _74922_ (_24313_, _24312_, _24307_);
  or _74923_ (_24314_, _24292_, _08782_);
  and _74924_ (_24315_, _24314_, _06718_);
  and _74925_ (_24316_, _24315_, _24313_);
  and _74926_ (_24317_, _24253_, _06316_);
  or _74927_ (_24318_, _24317_, _06047_);
  or _74928_ (_24319_, _24318_, _24316_);
  or _74929_ (_24321_, _24248_, _06048_);
  or _74930_ (_24322_, _24321_, _24251_);
  and _74931_ (_24323_, _24322_, _01336_);
  and _74932_ (_24324_, _24323_, _24319_);
  or _74933_ (_24325_, _24324_, _24241_);
  and _74934_ (_43409_, _24325_, _42882_);
  not _74935_ (_24326_, \oc8051_golden_model_1.TH0 [2]);
  nor _74936_ (_24327_, _01336_, _24326_);
  and _74937_ (_24328_, _09182_, _07663_);
  nor _74938_ (_24329_, _07663_, _24326_);
  or _74939_ (_24331_, _24329_, _07012_);
  or _74940_ (_24332_, _24331_, _24328_);
  nor _74941_ (_24333_, _11784_, _07530_);
  nor _74942_ (_24334_, _24333_, _24329_);
  nand _74943_ (_24335_, _24334_, _09815_);
  and _74944_ (_24336_, _14493_, _07663_);
  or _74945_ (_24337_, _24336_, _24329_);
  or _74946_ (_24338_, _24337_, _06954_);
  and _74947_ (_24339_, _07663_, \oc8051_golden_model_1.ACC [2]);
  nor _74948_ (_24340_, _24339_, _24329_);
  nor _74949_ (_24342_, _24340_, _06939_);
  nor _74950_ (_24343_, _06938_, _24326_);
  or _74951_ (_24344_, _24343_, _06102_);
  or _74952_ (_24345_, _24344_, _24342_);
  and _74953_ (_24346_, _24345_, _06848_);
  and _74954_ (_24347_, _24346_, _24338_);
  nor _74955_ (_24348_, _24334_, _06848_);
  or _74956_ (_24349_, _24348_, _24347_);
  nand _74957_ (_24350_, _24349_, _06220_);
  or _74958_ (_24351_, _24340_, _06220_);
  and _74959_ (_24353_, _24351_, _09817_);
  nand _74960_ (_24354_, _24353_, _24350_);
  and _74961_ (_24355_, _24354_, _24335_);
  and _74962_ (_24356_, _24355_, _24332_);
  or _74963_ (_24357_, _24356_, _09833_);
  and _74964_ (_24358_, _14580_, _07663_);
  or _74965_ (_24359_, _24358_, _24329_);
  or _74966_ (_24360_, _24359_, _05669_);
  and _74967_ (_24361_, _24360_, _06020_);
  and _74968_ (_24362_, _24361_, _24357_);
  and _74969_ (_24364_, _07663_, _08730_);
  or _74970_ (_24365_, _24364_, _24329_);
  and _74971_ (_24366_, _24365_, _06019_);
  or _74972_ (_24367_, _24366_, _06112_);
  or _74973_ (_24368_, _24367_, _24362_);
  and _74974_ (_24369_, _14596_, _07663_);
  or _74975_ (_24370_, _24369_, _24329_);
  or _74976_ (_24371_, _24370_, _08751_);
  and _74977_ (_24372_, _24371_, _08756_);
  and _74978_ (_24373_, _24372_, _24368_);
  and _74979_ (_24376_, _10991_, _07663_);
  or _74980_ (_24377_, _24376_, _24329_);
  and _74981_ (_24378_, _24377_, _06284_);
  or _74982_ (_24379_, _24378_, _24373_);
  and _74983_ (_24380_, _24379_, _07032_);
  or _74984_ (_24381_, _24329_, _08177_);
  and _74985_ (_24382_, _24365_, _06108_);
  and _74986_ (_24383_, _24382_, _24381_);
  or _74987_ (_24384_, _24383_, _24380_);
  and _74988_ (_24385_, _24384_, _06278_);
  nor _74989_ (_24387_, _24340_, _06278_);
  and _74990_ (_24388_, _24387_, _24381_);
  or _74991_ (_24389_, _24388_, _06130_);
  or _74992_ (_24390_, _24389_, _24385_);
  and _74993_ (_24391_, _14593_, _07663_);
  or _74994_ (_24392_, _24329_, _08777_);
  or _74995_ (_24393_, _24392_, _24391_);
  and _74996_ (_24394_, _24393_, _08782_);
  and _74997_ (_24395_, _24394_, _24390_);
  nor _74998_ (_24396_, _10990_, _11784_);
  or _74999_ (_24398_, _24396_, _24329_);
  and _75000_ (_24399_, _24398_, _06292_);
  or _75001_ (_24400_, _24399_, _24395_);
  and _75002_ (_24401_, _24400_, _06718_);
  and _75003_ (_24402_, _24337_, _06316_);
  or _75004_ (_24403_, _24402_, _06047_);
  or _75005_ (_24404_, _24403_, _24401_);
  and _75006_ (_24405_, _14657_, _07663_);
  or _75007_ (_24406_, _24329_, _06048_);
  or _75008_ (_24407_, _24406_, _24405_);
  and _75009_ (_24409_, _24407_, _01336_);
  and _75010_ (_24410_, _24409_, _24404_);
  or _75011_ (_24411_, _24410_, _24327_);
  and _75012_ (_43410_, _24411_, _42882_);
  not _75013_ (_24412_, \oc8051_golden_model_1.TH0 [3]);
  nor _75014_ (_24413_, _01336_, _24412_);
  nor _75015_ (_24414_, _07663_, _24412_);
  or _75016_ (_24415_, _24414_, _08029_);
  and _75017_ (_24416_, _07663_, _08662_);
  or _75018_ (_24417_, _24416_, _24414_);
  and _75019_ (_24419_, _24417_, _06108_);
  and _75020_ (_24420_, _24419_, _24415_);
  and _75021_ (_24421_, _09181_, _07663_);
  or _75022_ (_24422_, _24414_, _07012_);
  or _75023_ (_24423_, _24422_, _24421_);
  nor _75024_ (_24424_, _11784_, _07353_);
  nor _75025_ (_24425_, _24424_, _24414_);
  nand _75026_ (_24426_, _24425_, _09815_);
  and _75027_ (_24427_, _14672_, _07663_);
  or _75028_ (_24428_, _24427_, _24414_);
  or _75029_ (_24430_, _24428_, _06954_);
  and _75030_ (_24431_, _07663_, \oc8051_golden_model_1.ACC [3]);
  nor _75031_ (_24432_, _24431_, _24414_);
  nor _75032_ (_24433_, _24432_, _06939_);
  nor _75033_ (_24434_, _06938_, _24412_);
  or _75034_ (_24435_, _24434_, _06102_);
  or _75035_ (_24436_, _24435_, _24433_);
  and _75036_ (_24437_, _24436_, _06848_);
  and _75037_ (_24438_, _24437_, _24430_);
  nor _75038_ (_24439_, _24425_, _06848_);
  or _75039_ (_24441_, _24439_, _24438_);
  nand _75040_ (_24442_, _24441_, _06220_);
  or _75041_ (_24443_, _24432_, _06220_);
  and _75042_ (_24444_, _24443_, _09817_);
  nand _75043_ (_24445_, _24444_, _24442_);
  and _75044_ (_24446_, _24445_, _24426_);
  and _75045_ (_24447_, _24446_, _24423_);
  or _75046_ (_24448_, _24447_, _09833_);
  and _75047_ (_24449_, _14778_, _07663_);
  or _75048_ (_24450_, _24414_, _05669_);
  or _75049_ (_24452_, _24450_, _24449_);
  and _75050_ (_24453_, _24452_, _06020_);
  and _75051_ (_24454_, _24453_, _24448_);
  and _75052_ (_24455_, _24417_, _06019_);
  or _75053_ (_24456_, _24455_, _06112_);
  or _75054_ (_24457_, _24456_, _24454_);
  and _75055_ (_24458_, _14793_, _07663_);
  or _75056_ (_24459_, _24414_, _08751_);
  or _75057_ (_24460_, _24459_, _24458_);
  and _75058_ (_24461_, _24460_, _08756_);
  and _75059_ (_24463_, _24461_, _24457_);
  and _75060_ (_24464_, _12299_, _07663_);
  or _75061_ (_24465_, _24464_, _24414_);
  and _75062_ (_24466_, _24465_, _06284_);
  or _75063_ (_24467_, _24466_, _24463_);
  and _75064_ (_24468_, _24467_, _07032_);
  or _75065_ (_24469_, _24468_, _24420_);
  and _75066_ (_24470_, _24469_, _06278_);
  nor _75067_ (_24471_, _24432_, _06278_);
  and _75068_ (_24472_, _24471_, _24415_);
  or _75069_ (_24474_, _24472_, _06130_);
  or _75070_ (_24475_, _24474_, _24470_);
  and _75071_ (_24476_, _14792_, _07663_);
  or _75072_ (_24477_, _24414_, _08777_);
  or _75073_ (_24478_, _24477_, _24476_);
  and _75074_ (_24479_, _24478_, _08782_);
  and _75075_ (_24480_, _24479_, _24475_);
  nor _75076_ (_24481_, _10988_, _11784_);
  or _75077_ (_24482_, _24481_, _24414_);
  and _75078_ (_24483_, _24482_, _06292_);
  or _75079_ (_24485_, _24483_, _24480_);
  and _75080_ (_24486_, _24485_, _06718_);
  and _75081_ (_24487_, _24428_, _06316_);
  or _75082_ (_24488_, _24487_, _06047_);
  or _75083_ (_24489_, _24488_, _24486_);
  and _75084_ (_24490_, _14849_, _07663_);
  or _75085_ (_24491_, _24414_, _06048_);
  or _75086_ (_24492_, _24491_, _24490_);
  and _75087_ (_24493_, _24492_, _01336_);
  and _75088_ (_24494_, _24493_, _24489_);
  or _75089_ (_24496_, _24494_, _24413_);
  and _75090_ (_43411_, _24496_, _42882_);
  and _75091_ (_24497_, _01340_, \oc8051_golden_model_1.TH0 [4]);
  and _75092_ (_24498_, _11784_, \oc8051_golden_model_1.TH0 [4]);
  or _75093_ (_24499_, _24498_, _08273_);
  and _75094_ (_24500_, _08665_, _07663_);
  or _75095_ (_24501_, _24500_, _24498_);
  and _75096_ (_24502_, _24501_, _06108_);
  and _75097_ (_24503_, _24502_, _24499_);
  or _75098_ (_24504_, _24501_, _06020_);
  and _75099_ (_24506_, _14887_, _07663_);
  or _75100_ (_24507_, _24506_, _24498_);
  or _75101_ (_24508_, _24507_, _06954_);
  and _75102_ (_24509_, _07663_, \oc8051_golden_model_1.ACC [4]);
  or _75103_ (_24510_, _24509_, _24498_);
  and _75104_ (_24511_, _24510_, _06938_);
  and _75105_ (_24512_, _06939_, \oc8051_golden_model_1.TH0 [4]);
  or _75106_ (_24513_, _24512_, _06102_);
  or _75107_ (_24514_, _24513_, _24511_);
  and _75108_ (_24515_, _24514_, _06848_);
  and _75109_ (_24517_, _24515_, _24508_);
  nor _75110_ (_24518_, _08270_, _11784_);
  or _75111_ (_24519_, _24518_, _24498_);
  and _75112_ (_24520_, _24519_, _06239_);
  or _75113_ (_24521_, _24520_, _24517_);
  and _75114_ (_24522_, _24521_, _06220_);
  and _75115_ (_24523_, _24510_, _06219_);
  or _75116_ (_24524_, _24523_, _09818_);
  or _75117_ (_24525_, _24524_, _24522_);
  and _75118_ (_24526_, _09180_, _07663_);
  or _75119_ (_24528_, _24498_, _07012_);
  or _75120_ (_24529_, _24528_, _24526_);
  or _75121_ (_24530_, _24519_, _09827_);
  and _75122_ (_24531_, _24530_, _05669_);
  and _75123_ (_24532_, _24531_, _24529_);
  and _75124_ (_24533_, _24532_, _24525_);
  and _75125_ (_24534_, _14983_, _07663_);
  or _75126_ (_24535_, _24534_, _24498_);
  and _75127_ (_24536_, _24535_, _09833_);
  or _75128_ (_24537_, _24536_, _06019_);
  or _75129_ (_24539_, _24537_, _24533_);
  and _75130_ (_24540_, _24539_, _24504_);
  or _75131_ (_24541_, _24540_, _06112_);
  and _75132_ (_24542_, _14876_, _07663_);
  or _75133_ (_24543_, _24542_, _24498_);
  or _75134_ (_24544_, _24543_, _08751_);
  and _75135_ (_24545_, _24544_, _08756_);
  and _75136_ (_24546_, _24545_, _24541_);
  and _75137_ (_24547_, _10986_, _07663_);
  or _75138_ (_24548_, _24547_, _24498_);
  and _75139_ (_24550_, _24548_, _06284_);
  or _75140_ (_24551_, _24550_, _24546_);
  and _75141_ (_24552_, _24551_, _07032_);
  or _75142_ (_24553_, _24552_, _24503_);
  and _75143_ (_24554_, _24553_, _06278_);
  and _75144_ (_24555_, _24510_, _06277_);
  and _75145_ (_24556_, _24555_, _24499_);
  or _75146_ (_24557_, _24556_, _06130_);
  or _75147_ (_24558_, _24557_, _24554_);
  and _75148_ (_24559_, _14873_, _07663_);
  or _75149_ (_24561_, _24498_, _08777_);
  or _75150_ (_24562_, _24561_, _24559_);
  and _75151_ (_24563_, _24562_, _08782_);
  and _75152_ (_24564_, _24563_, _24558_);
  nor _75153_ (_24565_, _10985_, _11784_);
  or _75154_ (_24566_, _24565_, _24498_);
  and _75155_ (_24567_, _24566_, _06292_);
  or _75156_ (_24568_, _24567_, _24564_);
  and _75157_ (_24569_, _24568_, _06718_);
  and _75158_ (_24570_, _24507_, _06316_);
  or _75159_ (_24572_, _24570_, _06047_);
  or _75160_ (_24573_, _24572_, _24569_);
  and _75161_ (_24574_, _15055_, _07663_);
  or _75162_ (_24575_, _24498_, _06048_);
  or _75163_ (_24576_, _24575_, _24574_);
  and _75164_ (_24577_, _24576_, _01336_);
  and _75165_ (_24578_, _24577_, _24573_);
  or _75166_ (_24579_, _24578_, _24497_);
  and _75167_ (_43412_, _24579_, _42882_);
  and _75168_ (_24580_, _01340_, \oc8051_golden_model_1.TH0 [5]);
  and _75169_ (_24582_, _11784_, \oc8051_golden_model_1.TH0 [5]);
  or _75170_ (_24583_, _24582_, _07980_);
  and _75171_ (_24584_, _08652_, _07663_);
  or _75172_ (_24585_, _24584_, _24582_);
  and _75173_ (_24586_, _24585_, _06108_);
  and _75174_ (_24587_, _24586_, _24583_);
  or _75175_ (_24588_, _24585_, _06020_);
  and _75176_ (_24589_, _15093_, _07663_);
  or _75177_ (_24590_, _24589_, _24582_);
  or _75178_ (_24591_, _24590_, _06954_);
  and _75179_ (_24593_, _07663_, \oc8051_golden_model_1.ACC [5]);
  or _75180_ (_24594_, _24593_, _24582_);
  and _75181_ (_24595_, _24594_, _06938_);
  and _75182_ (_24596_, _06939_, \oc8051_golden_model_1.TH0 [5]);
  or _75183_ (_24597_, _24596_, _06102_);
  or _75184_ (_24598_, _24597_, _24595_);
  and _75185_ (_24599_, _24598_, _06848_);
  and _75186_ (_24600_, _24599_, _24591_);
  nor _75187_ (_24601_, _07977_, _11784_);
  or _75188_ (_24602_, _24601_, _24582_);
  and _75189_ (_24603_, _24602_, _06239_);
  or _75190_ (_24604_, _24603_, _24600_);
  and _75191_ (_24605_, _24604_, _06220_);
  and _75192_ (_24606_, _24594_, _06219_);
  or _75193_ (_24607_, _24606_, _09818_);
  or _75194_ (_24608_, _24607_, _24605_);
  and _75195_ (_24609_, _09179_, _07663_);
  or _75196_ (_24610_, _24582_, _07012_);
  or _75197_ (_24611_, _24610_, _24609_);
  or _75198_ (_24612_, _24602_, _09827_);
  and _75199_ (_24615_, _24612_, _05669_);
  and _75200_ (_24616_, _24615_, _24611_);
  and _75201_ (_24617_, _24616_, _24608_);
  and _75202_ (_24618_, _15179_, _07663_);
  or _75203_ (_24619_, _24618_, _24582_);
  and _75204_ (_24620_, _24619_, _09833_);
  or _75205_ (_24621_, _24620_, _06019_);
  or _75206_ (_24622_, _24621_, _24617_);
  and _75207_ (_24623_, _24622_, _24588_);
  or _75208_ (_24624_, _24623_, _06112_);
  and _75209_ (_24626_, _15195_, _07663_);
  or _75210_ (_24627_, _24582_, _08751_);
  or _75211_ (_24628_, _24627_, _24626_);
  and _75212_ (_24629_, _24628_, _08756_);
  and _75213_ (_24630_, _24629_, _24624_);
  and _75214_ (_24631_, _12306_, _07663_);
  or _75215_ (_24632_, _24631_, _24582_);
  and _75216_ (_24633_, _24632_, _06284_);
  or _75217_ (_24634_, _24633_, _24630_);
  and _75218_ (_24635_, _24634_, _07032_);
  or _75219_ (_24637_, _24635_, _24587_);
  and _75220_ (_24638_, _24637_, _06278_);
  and _75221_ (_24639_, _24594_, _06277_);
  and _75222_ (_24640_, _24639_, _24583_);
  or _75223_ (_24641_, _24640_, _06130_);
  or _75224_ (_24642_, _24641_, _24638_);
  and _75225_ (_24643_, _15194_, _07663_);
  or _75226_ (_24644_, _24582_, _08777_);
  or _75227_ (_24645_, _24644_, _24643_);
  and _75228_ (_24646_, _24645_, _08782_);
  and _75229_ (_24648_, _24646_, _24642_);
  nor _75230_ (_24649_, _10982_, _11784_);
  or _75231_ (_24650_, _24649_, _24582_);
  and _75232_ (_24651_, _24650_, _06292_);
  or _75233_ (_24652_, _24651_, _24648_);
  and _75234_ (_24653_, _24652_, _06718_);
  and _75235_ (_24654_, _24590_, _06316_);
  or _75236_ (_24655_, _24654_, _06047_);
  or _75237_ (_24656_, _24655_, _24653_);
  and _75238_ (_24657_, _15253_, _07663_);
  or _75239_ (_24659_, _24582_, _06048_);
  or _75240_ (_24660_, _24659_, _24657_);
  and _75241_ (_24661_, _24660_, _01336_);
  and _75242_ (_24662_, _24661_, _24656_);
  or _75243_ (_24663_, _24662_, _24580_);
  and _75244_ (_43413_, _24663_, _42882_);
  and _75245_ (_24664_, _01340_, \oc8051_golden_model_1.TH0 [6]);
  and _75246_ (_24665_, _11784_, \oc8051_golden_model_1.TH0 [6]);
  or _75247_ (_24666_, _24665_, _07886_);
  and _75248_ (_24667_, _15389_, _07663_);
  or _75249_ (_24669_, _24667_, _24665_);
  and _75250_ (_24670_, _24669_, _06108_);
  and _75251_ (_24671_, _24670_, _24666_);
  or _75252_ (_24672_, _24669_, _06020_);
  and _75253_ (_24673_, _15293_, _07663_);
  or _75254_ (_24674_, _24673_, _24665_);
  or _75255_ (_24675_, _24674_, _06954_);
  and _75256_ (_24676_, _07663_, \oc8051_golden_model_1.ACC [6]);
  or _75257_ (_24677_, _24676_, _24665_);
  and _75258_ (_24678_, _24677_, _06938_);
  and _75259_ (_24680_, _06939_, \oc8051_golden_model_1.TH0 [6]);
  or _75260_ (_24681_, _24680_, _06102_);
  or _75261_ (_24682_, _24681_, _24678_);
  and _75262_ (_24683_, _24682_, _06848_);
  and _75263_ (_24684_, _24683_, _24675_);
  nor _75264_ (_24685_, _07883_, _11784_);
  or _75265_ (_24686_, _24685_, _24665_);
  and _75266_ (_24687_, _24686_, _06239_);
  or _75267_ (_24688_, _24687_, _24684_);
  and _75268_ (_24689_, _24688_, _06220_);
  and _75269_ (_24691_, _24677_, _06219_);
  or _75270_ (_24692_, _24691_, _09818_);
  or _75271_ (_24693_, _24692_, _24689_);
  and _75272_ (_24694_, _09178_, _07663_);
  or _75273_ (_24695_, _24665_, _07012_);
  or _75274_ (_24696_, _24695_, _24694_);
  or _75275_ (_24697_, _24686_, _09827_);
  and _75276_ (_24698_, _24697_, _05669_);
  and _75277_ (_24699_, _24698_, _24696_);
  and _75278_ (_24700_, _24699_, _24693_);
  and _75279_ (_24702_, _15382_, _07663_);
  or _75280_ (_24703_, _24702_, _24665_);
  and _75281_ (_24704_, _24703_, _09833_);
  or _75282_ (_24705_, _24704_, _06019_);
  or _75283_ (_24706_, _24705_, _24700_);
  and _75284_ (_24707_, _24706_, _24672_);
  or _75285_ (_24708_, _24707_, _06112_);
  and _75286_ (_24709_, _15399_, _07663_);
  or _75287_ (_24710_, _24665_, _08751_);
  or _75288_ (_24711_, _24710_, _24709_);
  and _75289_ (_24713_, _24711_, _08756_);
  and _75290_ (_24714_, _24713_, _24708_);
  and _75291_ (_24715_, _10980_, _07663_);
  or _75292_ (_24716_, _24715_, _24665_);
  and _75293_ (_24717_, _24716_, _06284_);
  or _75294_ (_24718_, _24717_, _24714_);
  and _75295_ (_24719_, _24718_, _07032_);
  or _75296_ (_24720_, _24719_, _24671_);
  and _75297_ (_24721_, _24720_, _06278_);
  and _75298_ (_24722_, _24677_, _06277_);
  and _75299_ (_24724_, _24722_, _24666_);
  or _75300_ (_24725_, _24724_, _06130_);
  or _75301_ (_24726_, _24725_, _24721_);
  and _75302_ (_24727_, _15396_, _07663_);
  or _75303_ (_24728_, _24665_, _08777_);
  or _75304_ (_24729_, _24728_, _24727_);
  and _75305_ (_24730_, _24729_, _08782_);
  and _75306_ (_24731_, _24730_, _24726_);
  nor _75307_ (_24732_, _10979_, _11784_);
  or _75308_ (_24733_, _24732_, _24665_);
  and _75309_ (_24735_, _24733_, _06292_);
  or _75310_ (_24736_, _24735_, _24731_);
  and _75311_ (_24737_, _24736_, _06718_);
  and _75312_ (_24738_, _24674_, _06316_);
  or _75313_ (_24739_, _24738_, _06047_);
  or _75314_ (_24740_, _24739_, _24737_);
  and _75315_ (_24741_, _15451_, _07663_);
  or _75316_ (_24742_, _24665_, _06048_);
  or _75317_ (_24743_, _24742_, _24741_);
  and _75318_ (_24744_, _24743_, _01336_);
  and _75319_ (_24746_, _24744_, _24740_);
  or _75320_ (_24747_, _24746_, _24664_);
  and _75321_ (_43414_, _24747_, _42882_);
  nor _75322_ (_24748_, _06119_, _05751_);
  not _75323_ (_24749_, _24748_);
  and _75324_ (_24750_, _24749_, _06633_);
  and _75325_ (_24751_, _12779_, _12771_);
  nor _75326_ (_24752_, _24751_, _05346_);
  and _75327_ (_24753_, _12749_, _12756_);
  nor _75328_ (_24754_, _24753_, _05346_);
  and _75329_ (_24756_, _11872_, _11016_);
  nor _75330_ (_24757_, _24756_, _05346_);
  and _75331_ (_24758_, _12523_, _10855_);
  not _75332_ (_24759_, _05740_);
  nor _75333_ (_24760_, _06633_, _24759_);
  nor _75334_ (_24761_, _10612_, _05346_);
  and _75335_ (_24762_, _10612_, _05346_);
  nor _75336_ (_24763_, _24762_, _24761_);
  nor _75337_ (_24764_, _24763_, _12498_);
  not _75338_ (_24765_, _05736_);
  and _75339_ (_24767_, _12002_, _07032_);
  nor _75340_ (_24768_, _24767_, _05346_);
  not _75341_ (_24769_, _05727_);
  nor _75342_ (_24770_, _12006_, _06112_);
  nor _75343_ (_24771_, _24770_, _05346_);
  and _75344_ (_24772_, _06019_, _05346_);
  nor _75345_ (_24773_, _06110_, _09833_);
  and _75346_ (_24774_, _24773_, _12389_);
  nor _75347_ (_24775_, _24774_, _05346_);
  nor _75348_ (_24776_, _06633_, _05694_);
  and _75349_ (_24778_, _12239_, _12231_);
  nor _75350_ (_24779_, _24778_, _05346_);
  and _75351_ (_24780_, _06633_, _06943_);
  nor _75352_ (_24781_, _12205_, _05346_);
  nor _75353_ (_24782_, _12214_, _05346_);
  and _75354_ (_24783_, _12214_, _05346_);
  nor _75355_ (_24784_, _24783_, _24782_);
  and _75356_ (_24785_, _12205_, _07233_);
  not _75357_ (_24786_, _24785_);
  nor _75358_ (_24787_, _24786_, _24784_);
  nor _75359_ (_24789_, _24787_, _24781_);
  not _75360_ (_24790_, _24789_);
  nor _75361_ (_24791_, _24790_, _24780_);
  nor _75362_ (_24792_, _24791_, _08384_);
  and _75363_ (_24793_, _12197_, \oc8051_golden_model_1.PC [0]);
  and _75364_ (_24794_, _06016_, _05346_);
  nor _75365_ (_24795_, _24794_, _11928_);
  and _75366_ (_24796_, _24795_, _12199_);
  or _75367_ (_24797_, _24796_, _24793_);
  nor _75368_ (_24798_, _24797_, _08383_);
  nor _75369_ (_24800_, _24798_, _24792_);
  nor _75370_ (_24801_, _24800_, _06948_);
  and _75371_ (_24802_, _06948_, \oc8051_golden_model_1.PC [0]);
  nor _75372_ (_24803_, _24802_, _24801_);
  and _75373_ (_24804_, _24803_, _06954_);
  not _75374_ (_24805_, _12182_);
  and _75375_ (_24806_, _06633_, \oc8051_golden_model_1.PC [0]);
  nor _75376_ (_24807_, _24806_, _12088_);
  not _75377_ (_24808_, _24807_);
  and _75378_ (_24809_, _24808_, _12187_);
  and _75379_ (_24811_, _12189_, \oc8051_golden_model_1.PC [0]);
  or _75380_ (_24812_, _24811_, _06954_);
  nor _75381_ (_24813_, _24812_, _24809_);
  nor _75382_ (_24814_, _24813_, _24805_);
  not _75383_ (_24815_, _24814_);
  nor _75384_ (_24816_, _24815_, _24804_);
  nor _75385_ (_24817_, _12182_, _05346_);
  nor _75386_ (_24818_, _24817_, _07272_);
  not _75387_ (_24819_, _24818_);
  nor _75388_ (_24820_, _24819_, _24816_);
  nor _75389_ (_24822_, _06633_, _05690_);
  not _75390_ (_24823_, _24778_);
  nor _75391_ (_24824_, _24823_, _24822_);
  not _75392_ (_24825_, _24824_);
  nor _75393_ (_24826_, _24825_, _24820_);
  or _75394_ (_24827_, _24826_, _12243_);
  nor _75395_ (_24828_, _24827_, _24779_);
  nor _75396_ (_24829_, _24828_, _24776_);
  or _75397_ (_24830_, _24829_, _12256_);
  and _75398_ (_24831_, _12289_, \oc8051_golden_model_1.PC [0]);
  nor _75399_ (_24833_, _24807_, _12289_);
  or _75400_ (_24834_, _24833_, _12255_);
  or _75401_ (_24835_, _24834_, _24831_);
  and _75402_ (_24836_, _24835_, _12258_);
  and _75403_ (_24837_, _24836_, _24830_);
  nor _75404_ (_24838_, _24837_, _06121_);
  and _75405_ (_24839_, _12172_, _05346_);
  and _75406_ (_24840_, _24807_, _12174_);
  or _75407_ (_24841_, _24840_, _12258_);
  or _75408_ (_24842_, _24841_, _24839_);
  and _75409_ (_24844_, _24842_, _24838_);
  and _75410_ (_24845_, _12310_, _05346_);
  nor _75411_ (_24846_, _24808_, _12310_);
  nor _75412_ (_24847_, _24846_, _24845_);
  nor _75413_ (_24848_, _24847_, _06509_);
  nor _75414_ (_24849_, _24848_, _24844_);
  nor _75415_ (_24850_, _24849_, _06115_);
  and _75416_ (_24851_, _12329_, _05346_);
  nor _75417_ (_24852_, _24808_, _12329_);
  or _75418_ (_24853_, _24852_, _24851_);
  and _75419_ (_24855_, _24853_, _06115_);
  or _75420_ (_24856_, _24855_, _24850_);
  and _75421_ (_24857_, _24856_, _12013_);
  and _75422_ (_24858_, _12012_, _05346_);
  or _75423_ (_24859_, _24858_, _24857_);
  and _75424_ (_24860_, _24859_, _05686_);
  nor _75425_ (_24861_, _06633_, _05686_);
  nor _75426_ (_24862_, _24861_, _12355_);
  not _75427_ (_24863_, _24862_);
  nor _75428_ (_24864_, _24863_, _24860_);
  not _75429_ (_24866_, _05702_);
  nor _75430_ (_24867_, _12351_, _05346_);
  nor _75431_ (_24868_, _24867_, _24866_);
  not _75432_ (_24869_, _24868_);
  nor _75433_ (_24870_, _24869_, _24864_);
  nor _75434_ (_24871_, _06633_, _05702_);
  and _75435_ (_24872_, _12362_, _05675_);
  not _75436_ (_24873_, _24872_);
  nor _75437_ (_24874_, _24873_, _24871_);
  not _75438_ (_24875_, _24874_);
  nor _75439_ (_24877_, _24875_, _24870_);
  nor _75440_ (_24878_, _24872_, _05346_);
  nor _75441_ (_24879_, _24878_, _06023_);
  not _75442_ (_24880_, _24879_);
  nor _75443_ (_24881_, _24880_, _24877_);
  not _75444_ (_24882_, _24774_);
  nor _75445_ (_24883_, _06633_, _05673_);
  nor _75446_ (_24884_, _24883_, _24882_);
  not _75447_ (_24885_, _24884_);
  nor _75448_ (_24886_, _24885_, _24881_);
  nor _75449_ (_24888_, _24886_, _24775_);
  and _75450_ (_24889_, _24888_, _05720_);
  nor _75451_ (_24890_, _06633_, _05720_);
  or _75452_ (_24891_, _24890_, _24889_);
  and _75453_ (_24892_, _24891_, _12398_);
  and _75454_ (_24893_, _24795_, _12397_);
  or _75455_ (_24894_, _24893_, _24892_);
  and _75456_ (_24895_, _24894_, _06020_);
  or _75457_ (_24896_, _24895_, _24772_);
  and _75458_ (_24897_, _24896_, _12413_);
  and _75459_ (_24899_, _12412_, _05681_);
  or _75460_ (_24900_, _24899_, _24897_);
  and _75461_ (_24901_, _24900_, _13587_);
  nor _75462_ (_24902_, _06633_, _13587_);
  or _75463_ (_24903_, _24902_, _24901_);
  and _75464_ (_24904_, _24903_, _12454_);
  not _75465_ (_24905_, _24770_);
  nor _75466_ (_24906_, _24795_, _11071_);
  and _75467_ (_24907_, _11071_, _05346_);
  nor _75468_ (_24908_, _24907_, _12454_);
  not _75469_ (_24910_, _24908_);
  nor _75470_ (_24911_, _24910_, _24906_);
  nor _75471_ (_24912_, _24911_, _24905_);
  not _75472_ (_24913_, _24912_);
  nor _75473_ (_24914_, _24913_, _24904_);
  nor _75474_ (_24915_, _24914_, _24771_);
  and _75475_ (_24916_, _24915_, _24769_);
  nor _75476_ (_24917_, _06633_, _24769_);
  or _75477_ (_24918_, _24917_, _24916_);
  and _75478_ (_24919_, _24918_, _12477_);
  not _75479_ (_24921_, _24767_);
  nor _75480_ (_24922_, _24795_, _12459_);
  nor _75481_ (_24923_, _11071_, \oc8051_golden_model_1.PC [0]);
  nor _75482_ (_24924_, _24923_, _12477_);
  not _75483_ (_24925_, _24924_);
  nor _75484_ (_24926_, _24925_, _24922_);
  nor _75485_ (_24927_, _24926_, _24921_);
  not _75486_ (_24928_, _24927_);
  nor _75487_ (_24929_, _24928_, _24919_);
  nor _75488_ (_24930_, _24929_, _24768_);
  and _75489_ (_24932_, _24930_, _24765_);
  nor _75490_ (_24933_, _06633_, _24765_);
  or _75491_ (_24934_, _24933_, _24932_);
  and _75492_ (_24935_, _24934_, _12498_);
  and _75493_ (_24936_, _11993_, _08777_);
  not _75494_ (_24937_, _24936_);
  or _75495_ (_24938_, _24937_, _24935_);
  nor _75496_ (_24939_, _24938_, _24764_);
  nor _75497_ (_24940_, _24936_, _05346_);
  nor _75498_ (_24941_, _24940_, _05740_);
  not _75499_ (_24943_, _24941_);
  nor _75500_ (_24944_, _24943_, _24939_);
  nor _75501_ (_24945_, _24944_, _24760_);
  nor _75502_ (_24946_, _24945_, _11982_);
  nor _75503_ (_24947_, _10607_, _05346_);
  and _75504_ (_24948_, _10607_, _05346_);
  nor _75505_ (_24949_, _24948_, _24947_);
  nor _75506_ (_24950_, _24949_, _12518_);
  nor _75507_ (_24951_, _24950_, _24946_);
  and _75508_ (_24952_, _24951_, _24758_);
  nor _75509_ (_24954_, _24758_, _05346_);
  nor _75510_ (_24955_, _24954_, _06298_);
  not _75511_ (_24956_, _24955_);
  nor _75512_ (_24957_, _24956_, _24952_);
  and _75513_ (_24958_, _09120_, _06298_);
  or _75514_ (_24959_, _24958_, _24957_);
  and _75515_ (_24960_, _24959_, _05734_);
  nor _75516_ (_24961_, _06633_, _05734_);
  or _75517_ (_24962_, _24961_, _24960_);
  and _75518_ (_24963_, _24962_, _06306_);
  and _75519_ (_24965_, _24808_, _12722_);
  nor _75520_ (_24966_, _12722_, _05346_);
  or _75521_ (_24967_, _24966_, _06306_);
  or _75522_ (_24968_, _24967_, _24965_);
  and _75523_ (_24969_, _24968_, _24756_);
  not _75524_ (_24970_, _24969_);
  nor _75525_ (_24971_, _24970_, _24963_);
  nor _75526_ (_24972_, _24971_, _24757_);
  and _75527_ (_24973_, _24972_, _06050_);
  and _75528_ (_24974_, _09120_, _06049_);
  or _75529_ (_24976_, _24974_, _24973_);
  and _75530_ (_24977_, _24976_, _05748_);
  nor _75531_ (_24978_, _06633_, _05748_);
  nor _75532_ (_24979_, _24978_, _24977_);
  nor _75533_ (_24980_, _24979_, _06126_);
  not _75534_ (_24981_, _24753_);
  and _75535_ (_24982_, _12722_, \oc8051_golden_model_1.PC [0]);
  nor _75536_ (_24983_, _24807_, _12722_);
  nor _75537_ (_24984_, _24983_, _24982_);
  and _75538_ (_24985_, _24984_, _06126_);
  nor _75539_ (_24987_, _24985_, _24981_);
  not _75540_ (_24988_, _24987_);
  nor _75541_ (_24989_, _24988_, _24980_);
  nor _75542_ (_24990_, _24989_, _24754_);
  nor _75543_ (_24991_, _24990_, _07458_);
  and _75544_ (_24992_, _07458_, _06633_);
  nor _75545_ (_24993_, _24992_, _05652_);
  not _75546_ (_24994_, _24993_);
  nor _75547_ (_24995_, _24994_, _24991_);
  not _75548_ (_24996_, _24751_);
  and _75549_ (_24998_, _24984_, _05652_);
  nor _75550_ (_24999_, _24998_, _24996_);
  not _75551_ (_25000_, _24999_);
  nor _75552_ (_25001_, _25000_, _24995_);
  nor _75553_ (_25002_, _25001_, _24752_);
  nor _75554_ (_25003_, _24749_, _25002_);
  or _75555_ (_25004_, _25003_, _12789_);
  nor _75556_ (_25005_, _25004_, _24750_);
  and _75557_ (_25006_, _12789_, _05346_);
  or _75558_ (_25007_, _25006_, _25005_);
  or _75559_ (_25009_, _25007_, _01340_);
  or _75560_ (_25010_, _01336_, \oc8051_golden_model_1.PC [0]);
  and _75561_ (_25011_, _25010_, _42882_);
  and _75562_ (_43417_, _25011_, _25009_);
  and _75563_ (_25012_, _12789_, _12086_);
  and _75564_ (_25013_, _06047_, _05312_);
  nor _75565_ (_25014_, _12756_, _12086_);
  nor _75566_ (_25015_, _08286_, _12086_);
  nor _75567_ (_25016_, _11872_, _12086_);
  nor _75568_ (_25017_, _12523_, _12086_);
  and _75569_ (_25019_, _11989_, _05777_);
  nor _75570_ (_25020_, _12002_, _12086_);
  and _75571_ (_25021_, _12006_, _05777_);
  nor _75572_ (_25022_, _08742_, _05312_);
  not _75573_ (_25023_, _06089_);
  nor _75574_ (_25024_, _12389_, _12086_);
  nor _75575_ (_25025_, _12362_, _12086_);
  and _75576_ (_25026_, _12172_, _05777_);
  nor _75577_ (_25027_, _12090_, _12088_);
  nor _75578_ (_25028_, _25027_, _12091_);
  and _75579_ (_25030_, _25028_, _12174_);
  nor _75580_ (_25031_, _25030_, _25026_);
  nand _75581_ (_25032_, _25031_, _06104_);
  and _75582_ (_25033_, _06948_, _12086_);
  or _75583_ (_25034_, _12199_, \oc8051_golden_model_1.PC [1]);
  nor _75584_ (_25035_, _11930_, _11928_);
  nor _75585_ (_25036_, _25035_, _11931_);
  nand _75586_ (_25037_, _25036_, _12199_);
  and _75587_ (_25038_, _25037_, _25034_);
  nand _75588_ (_25039_, _25038_, _08384_);
  and _75589_ (_25041_, _06832_, _06943_);
  nor _75590_ (_25042_, _12205_, _12086_);
  and _75591_ (_25043_, _07250_, \oc8051_golden_model_1.PC [0]);
  nand _75592_ (_25044_, _06450_, _06523_);
  and _75593_ (_25045_, _06530_, _05346_);
  nor _75594_ (_25046_, _25045_, _25044_);
  nor _75595_ (_25047_, _25046_, _25043_);
  nor _75596_ (_25048_, _25047_, _05312_);
  and _75597_ (_25049_, _25047_, _05312_);
  nor _75598_ (_25050_, _25049_, _25048_);
  nor _75599_ (_25052_, _25050_, _24786_);
  nor _75600_ (_25053_, _25052_, _25042_);
  not _75601_ (_25054_, _25053_);
  nor _75602_ (_25055_, _25054_, _25041_);
  nor _75603_ (_25056_, _25055_, _08384_);
  nor _75604_ (_25057_, _25056_, _06948_);
  and _75605_ (_25058_, _25057_, _25039_);
  or _75606_ (_25059_, _25058_, _25033_);
  nand _75607_ (_25060_, _25059_, _06954_);
  or _75608_ (_25061_, _12187_, _12086_);
  not _75609_ (_25063_, _25028_);
  or _75610_ (_25064_, _25063_, _12189_);
  nand _75611_ (_25065_, _25064_, _25061_);
  nand _75612_ (_25066_, _25065_, _06102_);
  and _75613_ (_25067_, _25066_, _12182_);
  nand _75614_ (_25068_, _25067_, _25060_);
  nor _75615_ (_25069_, _12182_, _12086_);
  nor _75616_ (_25070_, _25069_, _06043_);
  nand _75617_ (_25071_, _25070_, _25068_);
  and _75618_ (_25072_, _06043_, _05312_);
  nor _75619_ (_25074_, _25072_, _07272_);
  nand _75620_ (_25075_, _25074_, _25071_);
  and _75621_ (_25076_, _06832_, _07272_);
  nor _75622_ (_25077_, _25076_, _06239_);
  nand _75623_ (_25078_, _25077_, _25075_);
  and _75624_ (_25079_, _06239_, _05312_);
  nor _75625_ (_25080_, _25079_, _12232_);
  nand _75626_ (_25081_, _25080_, _25078_);
  nor _75627_ (_25082_, _12231_, _12086_);
  nor _75628_ (_25083_, _25082_, _06219_);
  nand _75629_ (_25085_, _25083_, _25081_);
  and _75630_ (_25086_, _06219_, _05312_);
  nor _75631_ (_25087_, _25086_, _12241_);
  nand _75632_ (_25088_, _25087_, _25085_);
  nor _75633_ (_25089_, _12239_, _12086_);
  nor _75634_ (_25090_, _25089_, _06039_);
  nand _75635_ (_25091_, _25090_, _25088_);
  and _75636_ (_25092_, _06039_, _05312_);
  nor _75637_ (_25093_, _25092_, _12243_);
  nand _75638_ (_25094_, _25093_, _25091_);
  and _75639_ (_25096_, _06832_, _12243_);
  nor _75640_ (_25097_, _25096_, _06038_);
  nand _75641_ (_25098_, _25097_, _25094_);
  and _75642_ (_25099_, _06038_, _05312_);
  nor _75643_ (_25100_, _25099_, _12256_);
  and _75644_ (_25101_, _25100_, _25098_);
  and _75645_ (_25102_, _12289_, _05777_);
  nor _75646_ (_25103_, _25063_, _12289_);
  or _75647_ (_25104_, _25103_, _25102_);
  nor _75648_ (_25105_, _25104_, _12255_);
  or _75649_ (_25107_, _25105_, _25101_);
  nand _75650_ (_25108_, _25107_, _12258_);
  nand _75651_ (_25109_, _25108_, _25032_);
  nand _75652_ (_25110_, _25109_, _06509_);
  nor _75653_ (_25111_, _25063_, _12310_);
  not _75654_ (_25112_, _25111_);
  and _75655_ (_25113_, _12310_, _05777_);
  nor _75656_ (_25114_, _25113_, _06509_);
  and _75657_ (_25115_, _25114_, _25112_);
  nor _75658_ (_25116_, _25115_, _06115_);
  nand _75659_ (_25118_, _25116_, _25110_);
  and _75660_ (_25119_, _12329_, _12086_);
  not _75661_ (_25120_, _25119_);
  nor _75662_ (_25121_, _25028_, _12329_);
  nor _75663_ (_25122_, _25121_, _12298_);
  and _75664_ (_25123_, _25122_, _25120_);
  nor _75665_ (_25124_, _25123_, _12012_);
  nand _75666_ (_25125_, _25124_, _25118_);
  and _75667_ (_25126_, _12012_, _05777_);
  not _75668_ (_25127_, _25126_);
  and _75669_ (_25129_, _25127_, _12337_);
  nand _75670_ (_25130_, _25129_, _25125_);
  and _75671_ (_25131_, _06032_, _05312_);
  not _75672_ (_25132_, _25131_);
  not _75673_ (_25133_, _12344_);
  nor _75674_ (_25134_, _06832_, _05686_);
  nor _75675_ (_25135_, _25134_, _25133_);
  and _75676_ (_25136_, _25135_, _25132_);
  nand _75677_ (_25137_, _25136_, _25130_);
  nor _75678_ (_25138_, _12344_, _05312_);
  nor _75679_ (_25140_, _25138_, _12348_);
  nand _75680_ (_25141_, _25140_, _25137_);
  and _75681_ (_25142_, _12350_, _05777_);
  or _75682_ (_25143_, _25142_, _12351_);
  nand _75683_ (_25144_, _25143_, _25141_);
  nor _75684_ (_25145_, _12350_, _12086_);
  nor _75685_ (_25146_, _25145_, _06251_);
  nand _75686_ (_25147_, _25146_, _25144_);
  and _75687_ (_25148_, _06251_, _05312_);
  nor _75688_ (_25149_, _25148_, _24866_);
  nand _75689_ (_25150_, _25149_, _25147_);
  and _75690_ (_25151_, _06832_, _24866_);
  nor _75691_ (_25152_, _25151_, _06250_);
  nand _75692_ (_25153_, _25152_, _25150_);
  and _75693_ (_25154_, _06250_, _05312_);
  nor _75694_ (_25155_, _25154_, _12368_);
  and _75695_ (_25156_, _25155_, _25153_);
  or _75696_ (_25157_, _25156_, _25025_);
  nand _75697_ (_25158_, _25157_, _12366_);
  nor _75698_ (_25159_, _12366_, _05312_);
  nor _75699_ (_25162_, _25159_, _05676_);
  nand _75700_ (_25163_, _25162_, _25158_);
  nor _75701_ (_25164_, _05777_, _05675_);
  nor _75702_ (_25165_, _25164_, _06026_);
  and _75703_ (_25166_, _25165_, _25163_);
  and _75704_ (_25167_, _06026_, \oc8051_golden_model_1.PC [1]);
  or _75705_ (_25168_, _25167_, _25166_);
  nand _75706_ (_25169_, _25168_, _05673_);
  and _75707_ (_25170_, _06832_, _06023_);
  nor _75708_ (_25171_, _25170_, _06110_);
  nand _75709_ (_25173_, _25171_, _25169_);
  and _75710_ (_25174_, _06110_, _05777_);
  nor _75711_ (_25175_, _25174_, _09818_);
  nand _75712_ (_25176_, _25175_, _25173_);
  nor _75713_ (_25177_, _09817_, _05312_);
  nor _75714_ (_25178_, _25177_, _09833_);
  nand _75715_ (_25179_, _25178_, _25176_);
  nor _75716_ (_25180_, _12086_, _05669_);
  nor _75717_ (_25181_, _25180_, _12393_);
  and _75718_ (_25182_, _25181_, _25179_);
  or _75719_ (_25184_, _25182_, _25024_);
  nand _75720_ (_25185_, _25184_, _25023_);
  and _75721_ (_25186_, _06089_, \oc8051_golden_model_1.PC [1]);
  nor _75722_ (_25187_, _25186_, _05719_);
  and _75723_ (_25188_, _25187_, _25185_);
  nor _75724_ (_25189_, _06832_, _05720_);
  or _75725_ (_25190_, _25189_, _25188_);
  nand _75726_ (_25191_, _25190_, _12398_);
  and _75727_ (_25192_, _25036_, _12397_);
  nor _75728_ (_25193_, _25192_, _08743_);
  and _75729_ (_25195_, _25193_, _25191_);
  or _75730_ (_25196_, _25195_, _25022_);
  nand _75731_ (_25197_, _25196_, _06020_);
  and _75732_ (_25198_, _06019_, _12086_);
  nor _75733_ (_25199_, _25198_, _10661_);
  nand _75734_ (_25200_, _25199_, _25197_);
  and _75735_ (_25201_, _10661_, _05312_);
  nor _75736_ (_25202_, _25201_, _12412_);
  nand _75737_ (_25203_, _25202_, _25200_);
  nor _75738_ (_25204_, _12413_, _05775_);
  nor _75739_ (_25206_, _25204_, _06088_);
  nand _75740_ (_25207_, _25206_, _25203_);
  and _75741_ (_25208_, _06088_, _05312_);
  nor _75742_ (_25209_, _25208_, _05724_);
  nand _75743_ (_25210_, _25209_, _25207_);
  and _75744_ (_25211_, _06832_, _05724_);
  nor _75745_ (_25212_, _25211_, _12453_);
  nand _75746_ (_25213_, _25212_, _25210_);
  nor _75747_ (_25214_, _25036_, _11071_);
  and _75748_ (_25215_, _11071_, \oc8051_golden_model_1.PC [1]);
  nor _75749_ (_25217_, _25215_, _12454_);
  not _75750_ (_25218_, _25217_);
  nor _75751_ (_25219_, _25218_, _25214_);
  nor _75752_ (_25220_, _25219_, _12006_);
  and _75753_ (_25221_, _25220_, _25213_);
  or _75754_ (_25222_, _25221_, _25021_);
  nand _75755_ (_25223_, _25222_, _12466_);
  nor _75756_ (_25224_, _12466_, _05312_);
  nor _75757_ (_25225_, _25224_, _06112_);
  nand _75758_ (_25226_, _25225_, _25223_);
  and _75759_ (_25228_, _06112_, _05777_);
  nor _75760_ (_25229_, _25228_, _06284_);
  and _75761_ (_25230_, _25229_, _25226_);
  and _75762_ (_25231_, _06284_, \oc8051_golden_model_1.PC [1]);
  or _75763_ (_25232_, _25231_, _25230_);
  nand _75764_ (_25233_, _25232_, _24769_);
  and _75765_ (_25234_, _06832_, _05727_);
  nor _75766_ (_25235_, _25234_, _12476_);
  nand _75767_ (_25236_, _25235_, _25233_);
  nor _75768_ (_25237_, _25036_, _12459_);
  nor _75769_ (_25239_, _11071_, _05312_);
  nor _75770_ (_25240_, _25239_, _12477_);
  not _75771_ (_25241_, _25240_);
  nor _75772_ (_25242_, _25241_, _25237_);
  nor _75773_ (_25243_, _25242_, _12481_);
  and _75774_ (_25244_, _25243_, _25236_);
  or _75775_ (_25245_, _25244_, _25020_);
  nand _75776_ (_25246_, _25245_, _10742_);
  nor _75777_ (_25247_, _10742_, _05312_);
  nor _75778_ (_25248_, _25247_, _06108_);
  nand _75779_ (_25250_, _25248_, _25246_);
  and _75780_ (_25251_, _06108_, _05777_);
  nor _75781_ (_25252_, _25251_, _06277_);
  and _75782_ (_25253_, _25252_, _25250_);
  and _75783_ (_25254_, _06277_, \oc8051_golden_model_1.PC [1]);
  or _75784_ (_25255_, _25254_, _25253_);
  nand _75785_ (_25256_, _25255_, _24765_);
  and _75786_ (_25257_, _06832_, _05736_);
  nor _75787_ (_25258_, _25257_, _12497_);
  nand _75788_ (_25259_, _25258_, _25256_);
  and _75789_ (_25261_, \oc8051_golden_model_1.PSW [7], _05312_);
  and _75790_ (_25262_, _25036_, _10606_);
  or _75791_ (_25263_, _25262_, _25261_);
  and _75792_ (_25264_, _25263_, _12497_);
  nor _75793_ (_25265_, _25264_, _11989_);
  and _75794_ (_25266_, _25265_, _25259_);
  nor _75795_ (_25267_, _25266_, _25019_);
  nor _75796_ (_25268_, _07002_, _10394_);
  nor _75797_ (_25269_, _25268_, _10757_);
  or _75798_ (_25270_, _25269_, _25267_);
  and _75799_ (_25272_, _25269_, _05777_);
  nor _75800_ (_25273_, _25272_, _06669_);
  nand _75801_ (_25274_, _25273_, _25270_);
  and _75802_ (_25275_, _06669_, _12086_);
  nor _75803_ (_25276_, _25275_, _11987_);
  nand _75804_ (_25277_, _25276_, _25274_);
  nor _75805_ (_25278_, _11986_, _05312_);
  nor _75806_ (_25279_, _25278_, _06130_);
  and _75807_ (_25280_, _25279_, _25277_);
  and _75808_ (_25281_, _06130_, _05777_);
  or _75809_ (_25283_, _25281_, _06292_);
  nor _75810_ (_25284_, _25283_, _25280_);
  and _75811_ (_25285_, _06292_, \oc8051_golden_model_1.PC [1]);
  or _75812_ (_25286_, _25285_, _25284_);
  nand _75813_ (_25287_, _25286_, _24759_);
  and _75814_ (_25288_, _06832_, _05740_);
  nor _75815_ (_25289_, _25288_, _11982_);
  nand _75816_ (_25290_, _25289_, _25287_);
  nor _75817_ (_25291_, _25036_, _10606_);
  and _75818_ (_25292_, _10606_, \oc8051_golden_model_1.PC [1]);
  nor _75819_ (_25294_, _25292_, _12518_);
  not _75820_ (_25295_, _25294_);
  nor _75821_ (_25296_, _25295_, _25291_);
  nor _75822_ (_25297_, _25296_, _12525_);
  and _75823_ (_25298_, _25297_, _25290_);
  or _75824_ (_25299_, _25298_, _25017_);
  nand _75825_ (_25300_, _25299_, _10825_);
  nor _75826_ (_25301_, _10825_, _05312_);
  nor _75827_ (_25302_, _25301_, _10854_);
  nand _75828_ (_25303_, _25302_, _25300_);
  and _75829_ (_25305_, _10854_, _12086_);
  nor _75830_ (_25306_, _25305_, _06298_);
  and _75831_ (_25307_, _25306_, _25303_);
  and _75832_ (_25308_, _12150_, _06298_);
  or _75833_ (_25309_, _25308_, _25307_);
  nand _75834_ (_25310_, _25309_, _05734_);
  and _75835_ (_25311_, _06832_, _05732_);
  nor _75836_ (_25312_, _25311_, _06129_);
  nand _75837_ (_25313_, _25312_, _25310_);
  nor _75838_ (_25314_, _12722_, _05777_);
  not _75839_ (_25316_, _25314_);
  and _75840_ (_25317_, _25063_, _12722_);
  nor _75841_ (_25318_, _25317_, _06306_);
  and _75842_ (_25319_, _25318_, _25316_);
  nor _75843_ (_25320_, _25319_, _12541_);
  and _75844_ (_25321_, _25320_, _25313_);
  or _75845_ (_25322_, _25321_, _25016_);
  nand _75846_ (_25323_, _25322_, _10975_);
  nor _75847_ (_25324_, _10975_, _05312_);
  nor _75848_ (_25325_, _25324_, _11015_);
  nand _75849_ (_25327_, _25325_, _25323_);
  and _75850_ (_25328_, _11015_, _12086_);
  nor _75851_ (_25329_, _25328_, _06049_);
  and _75852_ (_25330_, _25329_, _25327_);
  and _75853_ (_25331_, _12150_, _06049_);
  or _75854_ (_25332_, _25331_, _25330_);
  nand _75855_ (_25333_, _25332_, _05748_);
  and _75856_ (_25334_, _06832_, _05747_);
  nor _75857_ (_25335_, _25334_, _06126_);
  nand _75858_ (_25336_, _25335_, _25333_);
  not _75859_ (_25338_, _08286_);
  nor _75860_ (_25339_, _25028_, _12722_);
  and _75861_ (_25340_, _12722_, _12086_);
  nor _75862_ (_25341_, _25340_, _25339_);
  and _75863_ (_25342_, _25341_, _06126_);
  nor _75864_ (_25343_, _25342_, _25338_);
  and _75865_ (_25344_, _25343_, _25336_);
  nor _75866_ (_25345_, _25344_, _25015_);
  not _75867_ (_25346_, _05495_);
  nor _75868_ (_25347_, _07248_, _25346_);
  or _75869_ (_25349_, _25347_, _25345_);
  and _75870_ (_25350_, _25347_, _05777_);
  nor _75871_ (_25351_, _25350_, _06316_);
  nand _75872_ (_25352_, _25351_, _25349_);
  not _75873_ (_25353_, _12756_);
  and _75874_ (_25354_, _06316_, _05312_);
  nor _75875_ (_25355_, _25354_, _25353_);
  and _75876_ (_25356_, _25355_, _25352_);
  or _75877_ (_25357_, _25356_, _25014_);
  nand _75878_ (_25358_, _25357_, _07059_);
  and _75879_ (_25360_, _07458_, _06832_);
  nor _75880_ (_25361_, _25360_, _05652_);
  nand _75881_ (_25362_, _25361_, _25358_);
  and _75882_ (_25363_, _25341_, _05652_);
  nor _75883_ (_25364_, _25363_, _12772_);
  nand _75884_ (_25365_, _25364_, _25362_);
  nor _75885_ (_25366_, _12771_, _12086_);
  nor _75886_ (_25367_, _25366_, _06047_);
  and _75887_ (_25368_, _25367_, _25365_);
  or _75888_ (_25369_, _25368_, _25013_);
  nand _75889_ (_25371_, _25369_, _12779_);
  nor _75890_ (_25372_, _12779_, _05777_);
  nor _75891_ (_25373_, _25372_, _24749_);
  nand _75892_ (_25374_, _25373_, _25371_);
  and _75893_ (_25375_, _24749_, _06832_);
  nor _75894_ (_25376_, _25375_, _12789_);
  and _75895_ (_25377_, _25376_, _25374_);
  or _75896_ (_25378_, _25377_, _25012_);
  or _75897_ (_25379_, _25378_, _01340_);
  or _75898_ (_25380_, _01336_, \oc8051_golden_model_1.PC [1]);
  and _75899_ (_25382_, _25380_, _42882_);
  and _75900_ (_43418_, _25382_, _25379_);
  and _75901_ (_25383_, _06047_, _05803_);
  and _75902_ (_25384_, _06316_, _05803_);
  nor _75903_ (_25385_, _11872_, _05823_);
  nor _75904_ (_25386_, _12523_, _05823_);
  nor _75905_ (_25387_, _11993_, _05823_);
  nor _75906_ (_25388_, _12002_, _05823_);
  and _75907_ (_25389_, _12006_, _05824_);
  nor _75908_ (_25390_, _08741_, _05803_);
  nor _75909_ (_25392_, _12344_, _05803_);
  and _75910_ (_25393_, _12012_, _05824_);
  or _75911_ (_25394_, _12174_, _12083_);
  and _75912_ (_25395_, _12095_, _12092_);
  nor _75913_ (_25396_, _25395_, _12096_);
  or _75914_ (_25397_, _25396_, _12172_);
  nand _75915_ (_25398_, _25397_, _25394_);
  nand _75916_ (_25399_, _25398_, _06104_);
  and _75917_ (_25400_, _06943_, _06445_);
  nor _75918_ (_25401_, _12205_, _05823_);
  nor _75919_ (_25403_, _12214_, _05823_);
  and _75920_ (_25404_, _06938_, _05804_);
  nor _75921_ (_25405_, _06938_, \oc8051_golden_model_1.PC [2]);
  and _75922_ (_25406_, _25405_, _07251_);
  nor _75923_ (_25407_, _25406_, _25404_);
  nor _75924_ (_25408_, _25407_, _06530_);
  nor _75925_ (_25409_, _25408_, _25403_);
  nor _75926_ (_25410_, _25409_, _24786_);
  or _75927_ (_25411_, _25410_, _25401_);
  nor _75928_ (_25412_, _25411_, _25400_);
  nor _75929_ (_25413_, _25412_, _08384_);
  and _75930_ (_25414_, _11935_, _11932_);
  nor _75931_ (_25415_, _25414_, _11936_);
  nand _75932_ (_25416_, _25415_, _12199_);
  or _75933_ (_25417_, _12199_, _05804_);
  and _75934_ (_25418_, _25417_, _08384_);
  and _75935_ (_25419_, _25418_, _25416_);
  or _75936_ (_25420_, _25419_, _25413_);
  nand _75937_ (_25421_, _25420_, _06949_);
  and _75938_ (_25422_, _06948_, _05824_);
  nor _75939_ (_25425_, _25422_, _06102_);
  nand _75940_ (_25426_, _25425_, _25421_);
  or _75941_ (_25427_, _25396_, _12189_);
  or _75942_ (_25428_, _12187_, _12083_);
  and _75943_ (_25429_, _25428_, _06102_);
  nand _75944_ (_25430_, _25429_, _25427_);
  and _75945_ (_25431_, _25430_, _12182_);
  nand _75946_ (_25432_, _25431_, _25426_);
  nor _75947_ (_25433_, _12182_, _05823_);
  nor _75948_ (_25434_, _25433_, _06043_);
  nand _75949_ (_25436_, _25434_, _25432_);
  and _75950_ (_25437_, _06043_, _05803_);
  nor _75951_ (_25438_, _25437_, _07272_);
  nand _75952_ (_25439_, _25438_, _25436_);
  and _75953_ (_25440_, _06445_, _07272_);
  nor _75954_ (_25441_, _25440_, _06239_);
  nand _75955_ (_25442_, _25441_, _25439_);
  and _75956_ (_25443_, _06239_, _05803_);
  nor _75957_ (_25444_, _25443_, _12232_);
  nand _75958_ (_25445_, _25444_, _25442_);
  nor _75959_ (_25447_, _12231_, _05823_);
  nor _75960_ (_25448_, _25447_, _06219_);
  nand _75961_ (_25449_, _25448_, _25445_);
  and _75962_ (_25450_, _06219_, _05803_);
  nor _75963_ (_25451_, _25450_, _12241_);
  nand _75964_ (_25452_, _25451_, _25449_);
  nor _75965_ (_25453_, _12239_, _05823_);
  nor _75966_ (_25454_, _25453_, _06039_);
  nand _75967_ (_25455_, _25454_, _25452_);
  and _75968_ (_25456_, _06039_, _05803_);
  nor _75969_ (_25458_, _25456_, _12243_);
  nand _75970_ (_25459_, _25458_, _25455_);
  and _75971_ (_25460_, _06445_, _12243_);
  nor _75972_ (_25461_, _25460_, _06038_);
  nand _75973_ (_25462_, _25461_, _25459_);
  and _75974_ (_25463_, _06038_, _05803_);
  nor _75975_ (_25464_, _25463_, _12256_);
  and _75976_ (_25465_, _25464_, _25462_);
  and _75977_ (_25466_, _12289_, _12083_);
  not _75978_ (_25467_, _25466_);
  not _75979_ (_25469_, _25396_);
  nor _75980_ (_25470_, _25469_, _12289_);
  nor _75981_ (_25471_, _25470_, _12255_);
  and _75982_ (_25472_, _25471_, _25467_);
  or _75983_ (_25473_, _25472_, _25465_);
  nand _75984_ (_25474_, _25473_, _12258_);
  nand _75985_ (_25475_, _25474_, _25399_);
  nand _75986_ (_25476_, _25475_, _06509_);
  nor _75987_ (_25477_, _25469_, _12310_);
  not _75988_ (_25478_, _25477_);
  and _75989_ (_25480_, _12310_, _12083_);
  nor _75990_ (_25481_, _25480_, _06509_);
  and _75991_ (_25482_, _25481_, _25478_);
  nor _75992_ (_25483_, _25482_, _06115_);
  nand _75993_ (_25484_, _25483_, _25476_);
  and _75994_ (_25485_, _12329_, _12084_);
  nor _75995_ (_25486_, _25396_, _12329_);
  or _75996_ (_25487_, _25486_, _12298_);
  or _75997_ (_25488_, _25487_, _25485_);
  and _75998_ (_25489_, _25488_, _12013_);
  and _75999_ (_25491_, _25489_, _25484_);
  or _76000_ (_25492_, _25491_, _25393_);
  nand _76001_ (_25493_, _25492_, _06033_);
  and _76002_ (_25494_, _06032_, _05804_);
  nor _76003_ (_25495_, _25494_, _07355_);
  nand _76004_ (_25496_, _25495_, _25493_);
  nor _76005_ (_25497_, _06445_, _05686_);
  nor _76006_ (_25498_, _25497_, _25133_);
  and _76007_ (_25499_, _25498_, _25496_);
  or _76008_ (_25500_, _25499_, _25392_);
  nand _76009_ (_25502_, _25500_, _12351_);
  nor _76010_ (_25503_, _12351_, _05823_);
  nor _76011_ (_25504_, _25503_, _06251_);
  nand _76012_ (_25505_, _25504_, _25502_);
  and _76013_ (_25506_, _06251_, _05803_);
  nor _76014_ (_25507_, _25506_, _24866_);
  nand _76015_ (_25508_, _25507_, _25505_);
  and _76016_ (_25509_, _06445_, _24866_);
  nor _76017_ (_25510_, _25509_, _06250_);
  nand _76018_ (_25511_, _25510_, _25508_);
  and _76019_ (_25513_, _06250_, _05803_);
  nor _76020_ (_25514_, _25513_, _12368_);
  and _76021_ (_25515_, _25514_, _25511_);
  nor _76022_ (_25516_, _12362_, _05823_);
  or _76023_ (_25517_, _25516_, _25515_);
  nand _76024_ (_25518_, _25517_, _12366_);
  nor _76025_ (_25519_, _12366_, _05803_);
  nor _76026_ (_25520_, _25519_, _05676_);
  nand _76027_ (_25521_, _25520_, _25518_);
  nor _76028_ (_25522_, _05824_, _05675_);
  nor _76029_ (_25524_, _25522_, _06026_);
  and _76030_ (_25525_, _25524_, _25521_);
  and _76031_ (_25526_, _06026_, _05804_);
  or _76032_ (_25527_, _25526_, _25525_);
  nand _76033_ (_25528_, _25527_, _05673_);
  and _76034_ (_25529_, _06445_, _06023_);
  nor _76035_ (_25530_, _25529_, _06110_);
  nand _76036_ (_25531_, _25530_, _25528_);
  and _76037_ (_25532_, _12083_, _06110_);
  nor _76038_ (_25533_, _25532_, _07011_);
  and _76039_ (_25535_, _25533_, _09827_);
  nand _76040_ (_25536_, _25535_, _25531_);
  nor _76041_ (_25537_, _09817_, _05803_);
  nor _76042_ (_25538_, _25537_, _09833_);
  nand _76043_ (_25539_, _25538_, _25536_);
  nor _76044_ (_25540_, _12084_, _05669_);
  nor _76045_ (_25541_, _25540_, _12393_);
  nand _76046_ (_25542_, _25541_, _25539_);
  nor _76047_ (_25543_, _12389_, _05823_);
  nor _76048_ (_25544_, _25543_, _06089_);
  and _76049_ (_25546_, _25544_, _25542_);
  and _76050_ (_25547_, _06089_, _05803_);
  or _76051_ (_25548_, _25547_, _05719_);
  nor _76052_ (_25549_, _25548_, _25546_);
  and _76053_ (_25550_, _06445_, _05719_);
  or _76054_ (_25551_, _25550_, _25549_);
  nand _76055_ (_25552_, _25551_, _12398_);
  not _76056_ (_25553_, _08740_);
  nor _76057_ (_25554_, _25415_, _12398_);
  nor _76058_ (_25555_, _25554_, _25553_);
  nand _76059_ (_25557_, _25555_, _25552_);
  not _76060_ (_25558_, _08741_);
  nor _76061_ (_25559_, _08740_, _05804_);
  nor _76062_ (_25560_, _25559_, _25558_);
  and _76063_ (_25561_, _25560_, _25557_);
  or _76064_ (_25562_, _25561_, _25390_);
  nand _76065_ (_25563_, _25562_, _06020_);
  and _76066_ (_25564_, _12084_, _06019_);
  nor _76067_ (_25565_, _25564_, _10661_);
  nand _76068_ (_25566_, _25565_, _25563_);
  and _76069_ (_25568_, _10661_, _05803_);
  nor _76070_ (_25569_, _25568_, _12412_);
  nand _76071_ (_25570_, _25569_, _25566_);
  and _76072_ (_25571_, _12412_, _05818_);
  nor _76073_ (_25572_, _25571_, _06088_);
  nand _76074_ (_25573_, _25572_, _25570_);
  and _76075_ (_25574_, _06088_, _05803_);
  nor _76076_ (_25575_, _25574_, _05724_);
  nand _76077_ (_25576_, _25575_, _25573_);
  and _76078_ (_25577_, _06445_, _05724_);
  nor _76079_ (_25579_, _25577_, _12453_);
  nand _76080_ (_25580_, _25579_, _25576_);
  nor _76081_ (_25581_, _25415_, _11071_);
  and _76082_ (_25582_, _11071_, _05804_);
  nor _76083_ (_25583_, _25582_, _12454_);
  not _76084_ (_25584_, _25583_);
  nor _76085_ (_25585_, _25584_, _25581_);
  nor _76086_ (_25586_, _25585_, _12006_);
  and _76087_ (_25587_, _25586_, _25580_);
  or _76088_ (_25588_, _25587_, _25389_);
  nand _76089_ (_25590_, _25588_, _12466_);
  nor _76090_ (_25591_, _12466_, _05803_);
  nor _76091_ (_25592_, _25591_, _06112_);
  nand _76092_ (_25593_, _25592_, _25590_);
  and _76093_ (_25594_, _12083_, _06112_);
  nor _76094_ (_25595_, _25594_, _06284_);
  and _76095_ (_25596_, _25595_, _25593_);
  and _76096_ (_25597_, _06284_, _05804_);
  or _76097_ (_25598_, _25597_, _25596_);
  nand _76098_ (_25599_, _25598_, _24769_);
  and _76099_ (_25601_, _06445_, _05727_);
  nor _76100_ (_25602_, _25601_, _12476_);
  nand _76101_ (_25603_, _25602_, _25599_);
  nor _76102_ (_25604_, _25415_, _12459_);
  nor _76103_ (_25605_, _11071_, _05803_);
  nor _76104_ (_25606_, _25605_, _12477_);
  not _76105_ (_25607_, _25606_);
  nor _76106_ (_25608_, _25607_, _25604_);
  nor _76107_ (_25609_, _25608_, _12481_);
  and _76108_ (_25610_, _25609_, _25603_);
  or _76109_ (_25612_, _25610_, _25388_);
  nand _76110_ (_25613_, _25612_, _10742_);
  nor _76111_ (_25614_, _10742_, _05803_);
  nor _76112_ (_25615_, _25614_, _06108_);
  nand _76113_ (_25616_, _25615_, _25613_);
  and _76114_ (_25617_, _12083_, _06108_);
  nor _76115_ (_25618_, _25617_, _06277_);
  and _76116_ (_25619_, _25618_, _25616_);
  and _76117_ (_25620_, _06277_, _05804_);
  or _76118_ (_25621_, _25620_, _25619_);
  nand _76119_ (_25623_, _25621_, _24765_);
  and _76120_ (_25624_, _06445_, _05736_);
  nor _76121_ (_25625_, _25624_, _12497_);
  nand _76122_ (_25626_, _25625_, _25623_);
  nor _76123_ (_25627_, _25415_, \oc8051_golden_model_1.PSW [7]);
  nor _76124_ (_25628_, _05803_, _10606_);
  nor _76125_ (_25629_, _25628_, _12498_);
  not _76126_ (_25630_, _25629_);
  nor _76127_ (_25631_, _25630_, _25627_);
  nor _76128_ (_25632_, _25631_, _12502_);
  and _76129_ (_25634_, _25632_, _25626_);
  or _76130_ (_25635_, _25634_, _25387_);
  nand _76131_ (_25636_, _25635_, _11986_);
  nor _76132_ (_25637_, _11986_, _05803_);
  nor _76133_ (_25638_, _25637_, _06130_);
  and _76134_ (_25639_, _25638_, _25636_);
  and _76135_ (_25640_, _12083_, _06130_);
  or _76136_ (_25641_, _25640_, _06292_);
  nor _76137_ (_25642_, _25641_, _25639_);
  and _76138_ (_25643_, _06292_, _05804_);
  or _76139_ (_25645_, _25643_, _25642_);
  nand _76140_ (_25646_, _25645_, _24759_);
  and _76141_ (_25647_, _06445_, _05740_);
  nor _76142_ (_25648_, _25647_, _11982_);
  nand _76143_ (_25649_, _25648_, _25646_);
  or _76144_ (_25650_, _25415_, _10606_);
  or _76145_ (_25651_, _05803_, \oc8051_golden_model_1.PSW [7]);
  and _76146_ (_25652_, _25651_, _11982_);
  and _76147_ (_25653_, _25652_, _25650_);
  nor _76148_ (_25654_, _25653_, _12525_);
  and _76149_ (_25656_, _25654_, _25649_);
  or _76150_ (_25657_, _25656_, _25386_);
  nand _76151_ (_25658_, _25657_, _10825_);
  nor _76152_ (_25659_, _10825_, _05803_);
  nor _76153_ (_25660_, _25659_, _10854_);
  nand _76154_ (_25661_, _25660_, _25658_);
  and _76155_ (_25662_, _10854_, _05823_);
  nor _76156_ (_25663_, _25662_, _06298_);
  and _76157_ (_25664_, _25663_, _25661_);
  and _76158_ (_25665_, _09030_, _06298_);
  or _76159_ (_25667_, _25665_, _25664_);
  nand _76160_ (_25668_, _25667_, _05734_);
  and _76161_ (_25669_, _06445_, _05732_);
  nor _76162_ (_25670_, _25669_, _06129_);
  nand _76163_ (_25671_, _25670_, _25668_);
  nor _76164_ (_25672_, _12083_, _12722_);
  and _76165_ (_25673_, _25469_, _12722_);
  or _76166_ (_25674_, _25673_, _06306_);
  nor _76167_ (_25675_, _25674_, _25672_);
  nor _76168_ (_25676_, _25675_, _12541_);
  and _76169_ (_25678_, _25676_, _25671_);
  or _76170_ (_25679_, _25678_, _25385_);
  nand _76171_ (_25680_, _25679_, _10975_);
  nor _76172_ (_25681_, _10975_, _05803_);
  nor _76173_ (_25682_, _25681_, _11015_);
  nand _76174_ (_25683_, _25682_, _25680_);
  and _76175_ (_25684_, _11015_, _05823_);
  nor _76176_ (_25685_, _25684_, _06049_);
  and _76177_ (_25686_, _25685_, _25683_);
  and _76178_ (_25687_, _09030_, _06049_);
  or _76179_ (_25689_, _25687_, _25686_);
  nand _76180_ (_25690_, _25689_, _05748_);
  and _76181_ (_25691_, _06445_, _05747_);
  nor _76182_ (_25692_, _25691_, _06126_);
  nand _76183_ (_25693_, _25692_, _25690_);
  nor _76184_ (_25694_, _25396_, _12722_);
  and _76185_ (_25695_, _12084_, _12722_);
  nor _76186_ (_25696_, _25695_, _25694_);
  and _76187_ (_25697_, _25696_, _06126_);
  nor _76188_ (_25698_, _25697_, _12750_);
  nand _76189_ (_25700_, _25698_, _25693_);
  nor _76190_ (_25701_, _12749_, _05823_);
  nor _76191_ (_25702_, _25701_, _06316_);
  and _76192_ (_25703_, _25702_, _25700_);
  or _76193_ (_25704_, _25703_, _25384_);
  nand _76194_ (_25705_, _25704_, _12756_);
  nor _76195_ (_25706_, _12756_, _05824_);
  nor _76196_ (_25707_, _25706_, _07458_);
  nand _76197_ (_25708_, _25707_, _25705_);
  and _76198_ (_25709_, _07458_, _06445_);
  nor _76199_ (_25711_, _25709_, _05652_);
  nand _76200_ (_25712_, _25711_, _25708_);
  and _76201_ (_25713_, _25696_, _05652_);
  nor _76202_ (_25714_, _25713_, _12772_);
  nand _76203_ (_25715_, _25714_, _25712_);
  nor _76204_ (_25716_, _12771_, _05823_);
  nor _76205_ (_25717_, _25716_, _06047_);
  and _76206_ (_25718_, _25717_, _25715_);
  or _76207_ (_25719_, _25718_, _25383_);
  nand _76208_ (_25720_, _25719_, _12779_);
  nor _76209_ (_25721_, _12779_, _05824_);
  nor _76210_ (_25722_, _25721_, _24749_);
  nand _76211_ (_25723_, _25722_, _25720_);
  and _76212_ (_25724_, _24749_, _06445_);
  nor _76213_ (_25725_, _25724_, _12789_);
  and _76214_ (_25726_, _25725_, _25723_);
  and _76215_ (_25727_, _12789_, _05823_);
  or _76216_ (_25728_, _25727_, _25726_);
  or _76217_ (_25729_, _25728_, _01340_);
  or _76218_ (_25730_, _01336_, \oc8051_golden_model_1.PC [2]);
  and _76219_ (_25733_, _25730_, _42882_);
  and _76220_ (_43419_, _25733_, _25729_);
  and _76221_ (_25734_, _06047_, _05853_);
  nor _76222_ (_25735_, _11872_, _06150_);
  nor _76223_ (_25736_, _12523_, _06150_);
  or _76224_ (_25737_, _11993_, _06150_);
  or _76225_ (_25738_, _12002_, _06150_);
  nand _76226_ (_25739_, _12006_, _05870_);
  or _76227_ (_25740_, _08742_, _05853_);
  nand _76228_ (_25741_, _12012_, _05870_);
  and _76229_ (_25743_, _12172_, _12078_);
  or _76230_ (_25744_, _12081_, _12080_);
  and _76231_ (_25745_, _25744_, _12097_);
  nor _76232_ (_25746_, _25744_, _12097_);
  nor _76233_ (_25747_, _25746_, _25745_);
  and _76234_ (_25748_, _25747_, _12174_);
  or _76235_ (_25749_, _25748_, _25743_);
  or _76236_ (_25750_, _25749_, _12258_);
  and _76237_ (_25751_, _12289_, _12078_);
  not _76238_ (_25752_, _25747_);
  nor _76239_ (_25754_, _25752_, _12289_);
  or _76240_ (_25755_, _25754_, _25751_);
  or _76241_ (_25756_, _25755_, _12255_);
  nor _76242_ (_25757_, _07233_, _06215_);
  not _76243_ (_25758_, _06530_);
  nand _76244_ (_25759_, _06938_, _06148_);
  and _76245_ (_25760_, _25759_, _25758_);
  nor _76246_ (_25761_, _07250_, _05307_);
  or _76247_ (_25762_, _25761_, _06938_);
  and _76248_ (_25763_, _25762_, _25760_);
  or _76249_ (_25765_, _12214_, _05870_);
  nand _76250_ (_25766_, _25765_, _12205_);
  or _76251_ (_25767_, _25766_, _25763_);
  and _76252_ (_25768_, _25767_, _07233_);
  or _76253_ (_25769_, _25768_, _25757_);
  or _76254_ (_25770_, _12205_, _06150_);
  and _76255_ (_25771_, _25770_, _25769_);
  or _76256_ (_25772_, _25771_, _08384_);
  or _76257_ (_25773_, _11925_, _11924_);
  and _76258_ (_25774_, _25773_, _11937_);
  nor _76259_ (_25776_, _25773_, _11937_);
  nor _76260_ (_25777_, _25776_, _25774_);
  and _76261_ (_25778_, _25777_, _12199_);
  and _76262_ (_25779_, _12197_, _05853_);
  or _76263_ (_25780_, _25779_, _08383_);
  or _76264_ (_25781_, _25780_, _25778_);
  and _76265_ (_25782_, _25781_, _25772_);
  or _76266_ (_25783_, _25782_, _06948_);
  nand _76267_ (_25784_, _06948_, _05870_);
  and _76268_ (_25785_, _25784_, _06954_);
  and _76269_ (_25787_, _25785_, _25783_);
  or _76270_ (_25788_, _12187_, _12078_);
  or _76271_ (_25789_, _25747_, _12189_);
  and _76272_ (_25790_, _25789_, _06102_);
  and _76273_ (_25791_, _25790_, _25788_);
  or _76274_ (_25792_, _25791_, _24805_);
  or _76275_ (_25793_, _25792_, _25787_);
  or _76276_ (_25794_, _12182_, _06150_);
  and _76277_ (_25795_, _25794_, _06044_);
  and _76278_ (_25796_, _25795_, _25793_);
  and _76279_ (_25798_, _06043_, _05853_);
  or _76280_ (_25799_, _25798_, _07272_);
  or _76281_ (_25800_, _25799_, _25796_);
  nand _76282_ (_25801_, _06215_, _07272_);
  and _76283_ (_25802_, _25801_, _06848_);
  and _76284_ (_25803_, _25802_, _25800_);
  nand _76285_ (_25804_, _06239_, _05853_);
  nand _76286_ (_25805_, _25804_, _12231_);
  or _76287_ (_25806_, _25805_, _25803_);
  or _76288_ (_25807_, _12231_, _06150_);
  and _76289_ (_25809_, _25807_, _06220_);
  and _76290_ (_25810_, _25809_, _25806_);
  nand _76291_ (_25811_, _06219_, _05853_);
  nand _76292_ (_25812_, _25811_, _12239_);
  or _76293_ (_25813_, _25812_, _25810_);
  or _76294_ (_25814_, _12239_, _06150_);
  and _76295_ (_25815_, _25814_, _06040_);
  and _76296_ (_25816_, _25815_, _25813_);
  and _76297_ (_25817_, _06039_, _05853_);
  or _76298_ (_25818_, _25817_, _12243_);
  or _76299_ (_25820_, _25818_, _25816_);
  nand _76300_ (_25821_, _06215_, _12243_);
  and _76301_ (_25822_, _25821_, _07364_);
  and _76302_ (_25823_, _25822_, _25820_);
  nand _76303_ (_25824_, _06038_, _05853_);
  nand _76304_ (_25825_, _25824_, _12255_);
  or _76305_ (_25826_, _25825_, _25823_);
  and _76306_ (_25827_, _25826_, _25756_);
  or _76307_ (_25828_, _25827_, _13850_);
  and _76308_ (_25829_, _25828_, _25750_);
  or _76309_ (_25831_, _25829_, _06121_);
  nor _76310_ (_25832_, _25752_, _12310_);
  and _76311_ (_25833_, _12310_, _12078_);
  or _76312_ (_25834_, _25833_, _06509_);
  or _76313_ (_25835_, _25834_, _25832_);
  and _76314_ (_25836_, _25835_, _12298_);
  and _76315_ (_25837_, _25836_, _25831_);
  nand _76316_ (_25838_, _12329_, _12079_);
  or _76317_ (_25839_, _25747_, _12329_);
  and _76318_ (_25840_, _25839_, _06115_);
  and _76319_ (_25842_, _25840_, _25838_);
  or _76320_ (_25843_, _25842_, _12012_);
  or _76321_ (_25844_, _25843_, _25837_);
  and _76322_ (_25845_, _25844_, _25741_);
  or _76323_ (_25846_, _25845_, _06032_);
  nand _76324_ (_25847_, _06032_, _06148_);
  and _76325_ (_25848_, _25847_, _05686_);
  and _76326_ (_25849_, _25848_, _25846_);
  nor _76327_ (_25850_, _06215_, _05686_);
  or _76328_ (_25851_, _25850_, _25133_);
  or _76329_ (_25853_, _25851_, _25849_);
  or _76330_ (_25854_, _12344_, _05853_);
  and _76331_ (_25855_, _25854_, _25853_);
  or _76332_ (_25856_, _25855_, _12355_);
  or _76333_ (_25857_, _12351_, _06150_);
  and _76334_ (_25858_, _25857_, _13765_);
  and _76335_ (_25859_, _25858_, _25856_);
  and _76336_ (_25860_, _06251_, _05853_);
  or _76337_ (_25861_, _25860_, _24866_);
  or _76338_ (_25862_, _25861_, _25859_);
  nand _76339_ (_25864_, _06215_, _24866_);
  and _76340_ (_25865_, _25864_, _13764_);
  and _76341_ (_25866_, _25865_, _25862_);
  nand _76342_ (_25867_, _06250_, _05853_);
  nand _76343_ (_25868_, _25867_, _12362_);
  or _76344_ (_25869_, _25868_, _25866_);
  or _76345_ (_25870_, _12362_, _06150_);
  and _76346_ (_25871_, _25870_, _25869_);
  or _76347_ (_25872_, _25871_, _12367_);
  or _76348_ (_25873_, _12366_, _05853_);
  and _76349_ (_25875_, _25873_, _05675_);
  and _76350_ (_25876_, _25875_, _25872_);
  nor _76351_ (_25877_, _05675_, _05870_);
  or _76352_ (_25878_, _25877_, _06026_);
  or _76353_ (_25879_, _25878_, _25876_);
  nand _76354_ (_25880_, _06026_, _06148_);
  and _76355_ (_25881_, _25880_, _25879_);
  or _76356_ (_25882_, _25881_, _06023_);
  nand _76357_ (_25883_, _06215_, _06023_);
  and _76358_ (_25884_, _25883_, _06111_);
  and _76359_ (_25886_, _25884_, _25882_);
  nand _76360_ (_25887_, _12078_, _06110_);
  nand _76361_ (_25888_, _25887_, _09817_);
  or _76362_ (_25889_, _25888_, _25886_);
  or _76363_ (_25890_, _09817_, _05853_);
  and _76364_ (_25891_, _25890_, _05669_);
  and _76365_ (_25892_, _25891_, _25889_);
  or _76366_ (_25893_, _12079_, _05669_);
  nand _76367_ (_25894_, _25893_, _12389_);
  or _76368_ (_25895_, _25894_, _25892_);
  or _76369_ (_25896_, _12389_, _06150_);
  and _76370_ (_25897_, _25896_, _25023_);
  and _76371_ (_25898_, _25897_, _25895_);
  and _76372_ (_25899_, _06089_, _05853_);
  or _76373_ (_25900_, _25899_, _05719_);
  or _76374_ (_25901_, _25900_, _25898_);
  nand _76375_ (_25902_, _06215_, _05719_);
  and _76376_ (_25903_, _25902_, _12398_);
  and _76377_ (_25904_, _25903_, _25901_);
  and _76378_ (_25905_, _25777_, _12397_);
  or _76379_ (_25907_, _25905_, _08743_);
  or _76380_ (_25908_, _25907_, _25904_);
  and _76381_ (_25909_, _25908_, _25740_);
  or _76382_ (_25910_, _25909_, _06019_);
  nand _76383_ (_25911_, _12079_, _06019_);
  and _76384_ (_25912_, _25911_, _10662_);
  and _76385_ (_25913_, _25912_, _25910_);
  and _76386_ (_25914_, _10661_, _05853_);
  or _76387_ (_25915_, _25914_, _12412_);
  or _76388_ (_25916_, _25915_, _25913_);
  or _76389_ (_25918_, _12413_, _05865_);
  and _76390_ (_25919_, _25918_, _06636_);
  and _76391_ (_25920_, _25919_, _25916_);
  and _76392_ (_25921_, _06088_, _05853_);
  or _76393_ (_25922_, _25921_, _05724_);
  or _76394_ (_25923_, _25922_, _25920_);
  nand _76395_ (_25924_, _06215_, _05724_);
  and _76396_ (_25925_, _25924_, _12454_);
  and _76397_ (_25926_, _25925_, _25923_);
  or _76398_ (_25927_, _25777_, _11071_);
  nand _76399_ (_25928_, _11071_, _06148_);
  and _76400_ (_25929_, _25928_, _12453_);
  and _76401_ (_25930_, _25929_, _25927_);
  or _76402_ (_25931_, _25930_, _12006_);
  or _76403_ (_25932_, _25931_, _25926_);
  and _76404_ (_25933_, _25932_, _25739_);
  or _76405_ (_25934_, _25933_, _12467_);
  or _76406_ (_25935_, _12466_, _05853_);
  and _76407_ (_25936_, _25935_, _08751_);
  and _76408_ (_25937_, _25936_, _25934_);
  and _76409_ (_25938_, _12078_, _06112_);
  or _76410_ (_25939_, _25938_, _06284_);
  or _76411_ (_25940_, _25939_, _25937_);
  nand _76412_ (_25941_, _06284_, _06148_);
  and _76413_ (_25942_, _25941_, _25940_);
  or _76414_ (_25943_, _25942_, _05727_);
  nand _76415_ (_25944_, _06215_, _05727_);
  and _76416_ (_25945_, _25944_, _12477_);
  and _76417_ (_25946_, _25945_, _25943_);
  or _76418_ (_25947_, _25777_, _12459_);
  or _76419_ (_25948_, _11071_, _05853_);
  and _76420_ (_25949_, _25948_, _12476_);
  and _76421_ (_25950_, _25949_, _25947_);
  or _76422_ (_25951_, _25950_, _12481_);
  or _76423_ (_25952_, _25951_, _25946_);
  and _76424_ (_25953_, _25952_, _25738_);
  or _76425_ (_25954_, _25953_, _10743_);
  or _76426_ (_25955_, _10742_, _05853_);
  and _76427_ (_25956_, _25955_, _07032_);
  and _76428_ (_25957_, _25956_, _25954_);
  and _76429_ (_25958_, _12078_, _06108_);
  or _76430_ (_25959_, _25958_, _06277_);
  or _76431_ (_25960_, _25959_, _25957_);
  nand _76432_ (_25961_, _06277_, _06148_);
  and _76433_ (_25962_, _25961_, _25960_);
  or _76434_ (_25963_, _25962_, _05736_);
  nand _76435_ (_25964_, _06215_, _05736_);
  and _76436_ (_25965_, _25964_, _12498_);
  and _76437_ (_25966_, _25965_, _25963_);
  or _76438_ (_25967_, _25777_, \oc8051_golden_model_1.PSW [7]);
  or _76439_ (_25968_, _05853_, _10606_);
  and _76440_ (_25969_, _25968_, _12497_);
  and _76441_ (_25970_, _25969_, _25967_);
  or _76442_ (_25971_, _25970_, _12502_);
  or _76443_ (_25972_, _25971_, _25966_);
  nand _76444_ (_25973_, _25972_, _25737_);
  nand _76445_ (_25974_, _25973_, _11986_);
  nor _76446_ (_25975_, _11986_, _05853_);
  nor _76447_ (_25976_, _25975_, _06130_);
  and _76448_ (_25977_, _25976_, _25974_);
  and _76449_ (_25979_, _12078_, _06130_);
  or _76450_ (_25980_, _25979_, _06292_);
  nor _76451_ (_25981_, _25980_, _25977_);
  and _76452_ (_25982_, _06292_, _06148_);
  or _76453_ (_25983_, _25982_, _25981_);
  nand _76454_ (_25984_, _25983_, _24759_);
  and _76455_ (_25985_, _06215_, _05740_);
  nor _76456_ (_25986_, _25985_, _11982_);
  nand _76457_ (_25987_, _25986_, _25984_);
  and _76458_ (_25988_, _05853_, _10606_);
  and _76459_ (_25990_, _25777_, \oc8051_golden_model_1.PSW [7]);
  or _76460_ (_25991_, _25990_, _25988_);
  and _76461_ (_25992_, _25991_, _11982_);
  nor _76462_ (_25993_, _25992_, _12525_);
  and _76463_ (_25994_, _25993_, _25987_);
  or _76464_ (_25995_, _25994_, _25736_);
  nand _76465_ (_25996_, _25995_, _10825_);
  nor _76466_ (_25997_, _10825_, _05853_);
  nor _76467_ (_25998_, _25997_, _10854_);
  nand _76468_ (_25999_, _25998_, _25996_);
  and _76469_ (_26000_, _10854_, _06150_);
  nor _76470_ (_26001_, _26000_, _06298_);
  and _76471_ (_26002_, _26001_, _25999_);
  and _76472_ (_26003_, _08985_, _06298_);
  or _76473_ (_26004_, _26003_, _26002_);
  nand _76474_ (_26005_, _26004_, _05734_);
  and _76475_ (_26006_, _06215_, _05732_);
  nor _76476_ (_26007_, _26006_, _06129_);
  nand _76477_ (_26008_, _26007_, _26005_);
  and _76478_ (_26009_, _25752_, _12722_);
  nor _76479_ (_26011_, _12078_, _12722_);
  or _76480_ (_26012_, _26011_, _06306_);
  nor _76481_ (_26013_, _26012_, _26009_);
  nor _76482_ (_26014_, _26013_, _12541_);
  and _76483_ (_26015_, _26014_, _26008_);
  or _76484_ (_26016_, _26015_, _25735_);
  nand _76485_ (_26017_, _26016_, _10975_);
  nor _76486_ (_26018_, _10975_, _05853_);
  nor _76487_ (_26019_, _26018_, _11015_);
  nand _76488_ (_26020_, _26019_, _26017_);
  and _76489_ (_26022_, _11015_, _06150_);
  nor _76490_ (_26023_, _26022_, _06049_);
  and _76491_ (_26024_, _26023_, _26020_);
  and _76492_ (_26025_, _08985_, _06049_);
  or _76493_ (_26026_, _26025_, _26024_);
  nand _76494_ (_26027_, _26026_, _05748_);
  and _76495_ (_26028_, _06215_, _05747_);
  nor _76496_ (_26029_, _26028_, _06126_);
  nand _76497_ (_26030_, _26029_, _26027_);
  nor _76498_ (_26031_, _25747_, _12722_);
  and _76499_ (_26033_, _12079_, _12722_);
  nor _76500_ (_26034_, _26033_, _26031_);
  and _76501_ (_26035_, _26034_, _06126_);
  nor _76502_ (_26036_, _26035_, _12750_);
  nand _76503_ (_26037_, _26036_, _26030_);
  nor _76504_ (_26038_, _12749_, _06150_);
  nor _76505_ (_26039_, _26038_, _06316_);
  nand _76506_ (_26040_, _26039_, _26037_);
  and _76507_ (_26041_, _06316_, _05853_);
  nor _76508_ (_26042_, _26041_, _25353_);
  and _76509_ (_26043_, _26042_, _26040_);
  nor _76510_ (_26044_, _12756_, _06150_);
  or _76511_ (_26045_, _26044_, _26043_);
  nand _76512_ (_26046_, _26045_, _07059_);
  and _76513_ (_26047_, _07458_, _06215_);
  nor _76514_ (_26048_, _26047_, _05652_);
  nand _76515_ (_26049_, _26048_, _26046_);
  and _76516_ (_26050_, _26034_, _05652_);
  nor _76517_ (_26051_, _26050_, _12772_);
  nand _76518_ (_26052_, _26051_, _26049_);
  nor _76519_ (_26055_, _12771_, _06150_);
  nor _76520_ (_26056_, _26055_, _06047_);
  and _76521_ (_26057_, _26056_, _26052_);
  or _76522_ (_26058_, _26057_, _25734_);
  nand _76523_ (_26059_, _26058_, _12779_);
  nor _76524_ (_26060_, _12779_, _05870_);
  nor _76525_ (_26061_, _26060_, _24749_);
  nand _76526_ (_26062_, _26061_, _26059_);
  and _76527_ (_26063_, _24749_, _06215_);
  nor _76528_ (_26064_, _26063_, _12789_);
  and _76529_ (_26065_, _26064_, _26062_);
  and _76530_ (_26066_, _12789_, _06150_);
  or _76531_ (_26067_, _26066_, _26065_);
  or _76532_ (_26068_, _26067_, _01340_);
  or _76533_ (_26069_, _01336_, \oc8051_golden_model_1.PC [3]);
  and _76534_ (_26070_, _26069_, _42882_);
  and _76535_ (_43420_, _26070_, _26068_);
  and _76536_ (_26071_, _08581_, _07458_);
  nor _76537_ (_26072_, _11921_, _08742_);
  nor _76538_ (_26073_, _12344_, _11921_);
  not _76539_ (_26075_, \oc8051_golden_model_1.PC [4]);
  nor _76540_ (_26076_, _05331_, _26075_);
  and _76541_ (_26077_, _05331_, _26075_);
  nor _76542_ (_26078_, _26077_, _26076_);
  not _76543_ (_26079_, _26078_);
  and _76544_ (_26080_, _26079_, _12012_);
  or _76545_ (_26081_, _12174_, _12074_);
  and _76546_ (_26082_, _12102_, _12099_);
  nor _76547_ (_26083_, _26082_, _12103_);
  not _76548_ (_26084_, _26083_);
  nand _76549_ (_26086_, _26084_, _12174_);
  nand _76550_ (_26087_, _26086_, _26081_);
  nand _76551_ (_26088_, _26087_, _06104_);
  and _76552_ (_26089_, _11922_, _06039_);
  and _76553_ (_26090_, _08581_, _06943_);
  not _76554_ (_26091_, _12205_);
  and _76555_ (_26092_, _11922_, _06938_);
  nor _76556_ (_26093_, _26092_, _06530_);
  nor _76557_ (_26094_, _07250_, _26075_);
  or _76558_ (_26095_, _26094_, _06938_);
  and _76559_ (_26097_, _26095_, _26093_);
  nor _76560_ (_26098_, _26079_, _12214_);
  or _76561_ (_26099_, _26098_, _06943_);
  nor _76562_ (_26100_, _26099_, _26097_);
  nor _76563_ (_26101_, _26100_, _26091_);
  not _76564_ (_26102_, _26101_);
  nor _76565_ (_26103_, _26102_, _26090_);
  nor _76566_ (_26104_, _26079_, _12205_);
  nor _76567_ (_26105_, _26104_, _08384_);
  not _76568_ (_26106_, _26105_);
  nor _76569_ (_26108_, _26106_, _26103_);
  and _76570_ (_26109_, _11942_, _11939_);
  nor _76571_ (_26110_, _26109_, _11943_);
  nand _76572_ (_26111_, _26110_, _12199_);
  or _76573_ (_26112_, _12199_, _11922_);
  and _76574_ (_26113_, _26112_, _26111_);
  and _76575_ (_26114_, _26113_, _08384_);
  or _76576_ (_26115_, _26114_, _26108_);
  nand _76577_ (_26116_, _26115_, _06949_);
  and _76578_ (_26117_, _26079_, _06948_);
  nor _76579_ (_26119_, _26117_, _06102_);
  nand _76580_ (_26120_, _26119_, _26116_);
  or _76581_ (_26121_, _12187_, _12074_);
  or _76582_ (_26122_, _26083_, _12189_);
  and _76583_ (_26123_, _26122_, _06102_);
  nand _76584_ (_26124_, _26123_, _26121_);
  nand _76585_ (_26125_, _26124_, _26120_);
  nand _76586_ (_26126_, _26125_, _12182_);
  nor _76587_ (_26127_, _26079_, _12182_);
  nor _76588_ (_26128_, _26127_, _06043_);
  nand _76589_ (_26129_, _26128_, _26126_);
  and _76590_ (_26130_, _11922_, _06043_);
  nor _76591_ (_26131_, _26130_, _07272_);
  nand _76592_ (_26132_, _26131_, _26129_);
  nor _76593_ (_26133_, _08581_, _05690_);
  nor _76594_ (_26134_, _26133_, _06239_);
  nand _76595_ (_26135_, _26134_, _26132_);
  and _76596_ (_26136_, _11922_, _06239_);
  nor _76597_ (_26137_, _26136_, _12232_);
  nand _76598_ (_26138_, _26137_, _26135_);
  nor _76599_ (_26140_, _26079_, _12231_);
  nor _76600_ (_26141_, _26140_, _06219_);
  nand _76601_ (_26142_, _26141_, _26138_);
  and _76602_ (_26143_, _11922_, _06219_);
  nor _76603_ (_26144_, _26143_, _12241_);
  nand _76604_ (_26145_, _26144_, _26142_);
  nor _76605_ (_26146_, _26079_, _12239_);
  nor _76606_ (_26147_, _26146_, _06039_);
  and _76607_ (_26148_, _26147_, _26145_);
  or _76608_ (_26149_, _26148_, _26089_);
  nand _76609_ (_26151_, _26149_, _05694_);
  and _76610_ (_26152_, _08581_, _12243_);
  nor _76611_ (_26153_, _26152_, _06038_);
  nand _76612_ (_26154_, _26153_, _26151_);
  and _76613_ (_26155_, _11921_, _06038_);
  nor _76614_ (_26156_, _26155_, _12256_);
  and _76615_ (_26157_, _26156_, _26154_);
  and _76616_ (_26158_, _12289_, _12074_);
  nor _76617_ (_26159_, _26084_, _12289_);
  or _76618_ (_26160_, _26159_, _12255_);
  nor _76619_ (_26162_, _26160_, _26158_);
  or _76620_ (_26163_, _26162_, _26157_);
  nand _76621_ (_26164_, _26163_, _12258_);
  nand _76622_ (_26165_, _26164_, _26088_);
  nand _76623_ (_26166_, _26165_, _06509_);
  nor _76624_ (_26167_, _26084_, _12310_);
  not _76625_ (_26168_, _26167_);
  and _76626_ (_26169_, _12310_, _12074_);
  nor _76627_ (_26170_, _26169_, _06509_);
  and _76628_ (_26171_, _26170_, _26168_);
  nor _76629_ (_26173_, _26171_, _06115_);
  nand _76630_ (_26174_, _26173_, _26166_);
  nor _76631_ (_26175_, _26083_, _12329_);
  and _76632_ (_26176_, _12329_, _12075_);
  nor _76633_ (_26177_, _26176_, _12298_);
  not _76634_ (_26178_, _26177_);
  nor _76635_ (_26179_, _26178_, _26175_);
  nor _76636_ (_26180_, _26179_, _12012_);
  and _76637_ (_26181_, _26180_, _26174_);
  or _76638_ (_26182_, _26181_, _26080_);
  nand _76639_ (_26184_, _26182_, _06033_);
  and _76640_ (_26185_, _11922_, _06032_);
  nor _76641_ (_26186_, _26185_, _07355_);
  nand _76642_ (_26187_, _26186_, _26184_);
  nor _76643_ (_26188_, _08581_, _05686_);
  nor _76644_ (_26189_, _26188_, _25133_);
  and _76645_ (_26190_, _26189_, _26187_);
  or _76646_ (_26191_, _26190_, _26073_);
  nand _76647_ (_26192_, _26191_, _12351_);
  nor _76648_ (_26193_, _26078_, _12351_);
  nor _76649_ (_26194_, _26193_, _06251_);
  nand _76650_ (_26195_, _26194_, _26192_);
  and _76651_ (_26196_, _11921_, _06251_);
  nor _76652_ (_26197_, _26196_, _24866_);
  nand _76653_ (_26198_, _26197_, _26195_);
  and _76654_ (_26199_, _08581_, _24866_);
  nor _76655_ (_26200_, _26199_, _06250_);
  and _76656_ (_26201_, _26200_, _26198_);
  and _76657_ (_26202_, _11921_, _06250_);
  or _76658_ (_26203_, _26202_, _26201_);
  nand _76659_ (_26205_, _26203_, _12362_);
  nor _76660_ (_26206_, _26079_, _12362_);
  nor _76661_ (_26207_, _26206_, _12367_);
  nand _76662_ (_26208_, _26207_, _26205_);
  nor _76663_ (_26209_, _11921_, _12366_);
  nor _76664_ (_26210_, _26209_, _05676_);
  nand _76665_ (_26211_, _26210_, _26208_);
  nor _76666_ (_26212_, _26079_, _05675_);
  nor _76667_ (_26213_, _26212_, _06026_);
  and _76668_ (_26214_, _26213_, _26211_);
  and _76669_ (_26216_, _11922_, _06026_);
  or _76670_ (_26217_, _26216_, _26214_);
  nand _76671_ (_26218_, _26217_, _05673_);
  and _76672_ (_26219_, _08581_, _06023_);
  nor _76673_ (_26220_, _26219_, _06110_);
  nand _76674_ (_26221_, _26220_, _26218_);
  and _76675_ (_26222_, _12074_, _06110_);
  nor _76676_ (_26223_, _26222_, _09818_);
  nand _76677_ (_26224_, _26223_, _26221_);
  nor _76678_ (_26225_, _11921_, _09817_);
  nor _76679_ (_26227_, _26225_, _09833_);
  nand _76680_ (_26228_, _26227_, _26224_);
  nor _76681_ (_26229_, _12075_, _05669_);
  nor _76682_ (_26230_, _26229_, _12393_);
  nand _76683_ (_26231_, _26230_, _26228_);
  nor _76684_ (_26232_, _26078_, _12389_);
  nor _76685_ (_26233_, _26232_, _06089_);
  nand _76686_ (_26234_, _26233_, _26231_);
  and _76687_ (_26235_, _11921_, _06089_);
  nor _76688_ (_26236_, _26235_, _05719_);
  nand _76689_ (_26238_, _26236_, _26234_);
  and _76690_ (_26239_, _08581_, _05719_);
  nor _76691_ (_26240_, _26239_, _12397_);
  nand _76692_ (_26241_, _26240_, _26238_);
  and _76693_ (_26242_, _26110_, _12397_);
  nor _76694_ (_26243_, _26242_, _08743_);
  and _76695_ (_26244_, _26243_, _26241_);
  or _76696_ (_26245_, _26244_, _26072_);
  nand _76697_ (_26246_, _26245_, _06020_);
  and _76698_ (_26247_, _12075_, _06019_);
  nor _76699_ (_26249_, _26247_, _10661_);
  and _76700_ (_26250_, _26249_, _26246_);
  and _76701_ (_26251_, _11921_, _10661_);
  or _76702_ (_26252_, _26251_, _26250_);
  nand _76703_ (_26253_, _26252_, _12413_);
  and _76704_ (_26254_, _12431_, _12428_);
  nor _76705_ (_26255_, _26254_, _12432_);
  and _76706_ (_26256_, _26255_, _12412_);
  nor _76707_ (_26257_, _26256_, _06088_);
  and _76708_ (_26258_, _26257_, _26253_);
  and _76709_ (_26259_, _11922_, _06088_);
  or _76710_ (_26260_, _26259_, _26258_);
  nand _76711_ (_26261_, _26260_, _13587_);
  and _76712_ (_26262_, _08581_, _05724_);
  nor _76713_ (_26263_, _26262_, _12453_);
  and _76714_ (_26264_, _26263_, _26261_);
  and _76715_ (_26265_, _11921_, _11071_);
  and _76716_ (_26266_, _26110_, _12459_);
  or _76717_ (_26267_, _26266_, _26265_);
  and _76718_ (_26268_, _26267_, _12453_);
  or _76719_ (_26270_, _26268_, _26264_);
  nand _76720_ (_26271_, _26270_, _12007_);
  and _76721_ (_26272_, _26078_, _12006_);
  nor _76722_ (_26273_, _26272_, _12467_);
  nand _76723_ (_26274_, _26273_, _26271_);
  nor _76724_ (_26275_, _12466_, _11921_);
  nor _76725_ (_26276_, _26275_, _06112_);
  nand _76726_ (_26277_, _26276_, _26274_);
  and _76727_ (_26278_, _12074_, _06112_);
  nor _76728_ (_26279_, _26278_, _06284_);
  and _76729_ (_26281_, _26279_, _26277_);
  and _76730_ (_26282_, _11922_, _06284_);
  or _76731_ (_26283_, _26282_, _26281_);
  nand _76732_ (_26284_, _26283_, _24769_);
  and _76733_ (_26285_, _08581_, _05727_);
  nor _76734_ (_26286_, _26285_, _12476_);
  and _76735_ (_26287_, _26286_, _26284_);
  nor _76736_ (_26288_, _11922_, _11071_);
  and _76737_ (_26289_, _26110_, _11071_);
  or _76738_ (_26290_, _26289_, _26288_);
  and _76739_ (_26292_, _26290_, _12476_);
  or _76740_ (_26293_, _26292_, _26287_);
  nand _76741_ (_26294_, _26293_, _12002_);
  nor _76742_ (_26295_, _26079_, _12002_);
  nor _76743_ (_26296_, _26295_, _10743_);
  nand _76744_ (_26297_, _26296_, _26294_);
  nor _76745_ (_26298_, _11921_, _10742_);
  nor _76746_ (_26299_, _26298_, _06108_);
  nand _76747_ (_26300_, _26299_, _26297_);
  and _76748_ (_26301_, _12074_, _06108_);
  nor _76749_ (_26303_, _26301_, _06277_);
  and _76750_ (_26304_, _26303_, _26300_);
  and _76751_ (_26305_, _11922_, _06277_);
  or _76752_ (_26306_, _26305_, _26304_);
  nand _76753_ (_26307_, _26306_, _24765_);
  and _76754_ (_26308_, _08581_, _05736_);
  nor _76755_ (_26309_, _26308_, _12497_);
  and _76756_ (_26310_, _26309_, _26307_);
  and _76757_ (_26311_, _11921_, \oc8051_golden_model_1.PSW [7]);
  and _76758_ (_26312_, _26110_, _10606_);
  or _76759_ (_26314_, _26312_, _26311_);
  and _76760_ (_26315_, _26314_, _12497_);
  or _76761_ (_26316_, _26315_, _26310_);
  nand _76762_ (_26317_, _26316_, _11993_);
  nor _76763_ (_26318_, _26079_, _11993_);
  nor _76764_ (_26319_, _26318_, _11987_);
  nand _76765_ (_26320_, _26319_, _26317_);
  nor _76766_ (_26321_, _11921_, _11986_);
  nor _76767_ (_26322_, _26321_, _06130_);
  nand _76768_ (_26323_, _26322_, _26320_);
  and _76769_ (_26324_, _12074_, _06130_);
  nor _76770_ (_26325_, _26324_, _06292_);
  and _76771_ (_26326_, _26325_, _26323_);
  and _76772_ (_26327_, _11922_, _06292_);
  or _76773_ (_26328_, _26327_, _26326_);
  nand _76774_ (_26329_, _26328_, _24759_);
  and _76775_ (_26330_, _08581_, _05740_);
  nor _76776_ (_26331_, _26330_, _11982_);
  and _76777_ (_26332_, _26331_, _26329_);
  and _76778_ (_26333_, _11921_, _10606_);
  and _76779_ (_26335_, _26110_, \oc8051_golden_model_1.PSW [7]);
  or _76780_ (_26336_, _26335_, _26333_);
  and _76781_ (_26337_, _26336_, _11982_);
  or _76782_ (_26338_, _26337_, _26332_);
  nand _76783_ (_26339_, _26338_, _12523_);
  nor _76784_ (_26340_, _26079_, _12523_);
  nor _76785_ (_26341_, _26340_, _10826_);
  nand _76786_ (_26342_, _26341_, _26339_);
  nor _76787_ (_26343_, _11921_, _10825_);
  nor _76788_ (_26344_, _26343_, _10854_);
  nand _76789_ (_26346_, _26344_, _26342_);
  and _76790_ (_26347_, _26078_, _10854_);
  nor _76791_ (_26348_, _26347_, _06298_);
  and _76792_ (_26349_, _26348_, _26346_);
  and _76793_ (_26350_, _08937_, _06298_);
  or _76794_ (_26351_, _26350_, _26349_);
  nand _76795_ (_26352_, _26351_, _05734_);
  and _76796_ (_26353_, _08581_, _05732_);
  nor _76797_ (_26354_, _26353_, _06129_);
  and _76798_ (_26355_, _26354_, _26352_);
  nor _76799_ (_26357_, _12075_, _12722_);
  and _76800_ (_26358_, _26083_, _12722_);
  nor _76801_ (_26359_, _26358_, _26357_);
  nor _76802_ (_26360_, _26359_, _06306_);
  or _76803_ (_26361_, _26360_, _26355_);
  nand _76804_ (_26362_, _26361_, _11872_);
  nor _76805_ (_26363_, _26079_, _11872_);
  nor _76806_ (_26364_, _26363_, _10976_);
  nand _76807_ (_26365_, _26364_, _26362_);
  nor _76808_ (_26366_, _11921_, _10975_);
  nor _76809_ (_26368_, _26366_, _11015_);
  nand _76810_ (_26369_, _26368_, _26365_);
  and _76811_ (_26370_, _26078_, _11015_);
  nor _76812_ (_26371_, _26370_, _06049_);
  nand _76813_ (_26372_, _26371_, _26369_);
  and _76814_ (_26373_, _08937_, _06049_);
  nor _76815_ (_26374_, _26373_, _05747_);
  nand _76816_ (_26375_, _26374_, _26372_);
  nor _76817_ (_26376_, _08581_, _05748_);
  nor _76818_ (_26377_, _26376_, _06126_);
  nand _76819_ (_26379_, _26377_, _26375_);
  nor _76820_ (_26380_, _26083_, _12722_);
  and _76821_ (_26381_, _12075_, _12722_);
  nor _76822_ (_26382_, _26381_, _26380_);
  nor _76823_ (_26383_, _26382_, _06704_);
  nor _76824_ (_26384_, _26383_, _12750_);
  nand _76825_ (_26385_, _26384_, _26379_);
  nor _76826_ (_26386_, _26079_, _12749_);
  nor _76827_ (_26387_, _26386_, _06316_);
  nand _76828_ (_26388_, _26387_, _26385_);
  and _76829_ (_26390_, _11922_, _06316_);
  nor _76830_ (_26391_, _26390_, _25353_);
  nand _76831_ (_26392_, _26391_, _26388_);
  nor _76832_ (_26393_, _26079_, _12756_);
  nor _76833_ (_26394_, _26393_, _07458_);
  and _76834_ (_26395_, _26394_, _26392_);
  or _76835_ (_26396_, _26395_, _26071_);
  nand _76836_ (_26397_, _26396_, _05653_);
  nor _76837_ (_26398_, _26382_, _05653_);
  nor _76838_ (_26399_, _26398_, _12772_);
  nand _76839_ (_26401_, _26399_, _26397_);
  nor _76840_ (_26402_, _26079_, _12771_);
  nor _76841_ (_26403_, _26402_, _06047_);
  nand _76842_ (_26404_, _26403_, _26401_);
  not _76843_ (_26405_, _12779_);
  and _76844_ (_26406_, _11922_, _06047_);
  nor _76845_ (_26407_, _26406_, _26405_);
  nand _76846_ (_26408_, _26407_, _26404_);
  nor _76847_ (_26409_, _26079_, _12779_);
  nor _76848_ (_26410_, _26409_, _24749_);
  nand _76849_ (_26411_, _26410_, _26408_);
  and _76850_ (_26412_, _24749_, _08581_);
  nor _76851_ (_26413_, _26412_, _12789_);
  and _76852_ (_26414_, _26413_, _26411_);
  and _76853_ (_26415_, _26078_, _12789_);
  or _76854_ (_26416_, _26415_, _26414_);
  or _76855_ (_26417_, _26416_, _01340_);
  or _76856_ (_26418_, _01336_, \oc8051_golden_model_1.PC [4]);
  and _76857_ (_26419_, _26418_, _42882_);
  and _76858_ (_43421_, _26419_, _26417_);
  nor _76859_ (_26421_, \oc8051_golden_model_1.PC [5], \oc8051_golden_model_1.PC [0]);
  nor _76860_ (_26422_, _11916_, _05346_);
  nor _76861_ (_26423_, _26422_, _26421_);
  and _76862_ (_26424_, _26423_, _12789_);
  and _76863_ (_26425_, _11916_, _06047_);
  nor _76864_ (_26426_, _26423_, _11872_);
  nor _76865_ (_26427_, _26423_, _12523_);
  nor _76866_ (_26428_, _26423_, _11993_);
  nor _76867_ (_26429_, _26423_, _12002_);
  not _76868_ (_26430_, _26423_);
  and _76869_ (_26432_, _26430_, _12006_);
  nor _76870_ (_26433_, _11916_, _08742_);
  and _76871_ (_26434_, _26430_, _12012_);
  and _76872_ (_26435_, _12172_, _12069_);
  or _76873_ (_26436_, _12071_, _12072_);
  and _76874_ (_26437_, _26436_, _12104_);
  nor _76875_ (_26438_, _26436_, _12104_);
  nor _76876_ (_26439_, _26438_, _26437_);
  and _76877_ (_26440_, _26439_, _12174_);
  nor _76878_ (_26441_, _26440_, _26435_);
  nand _76879_ (_26443_, _26441_, _06104_);
  nor _76880_ (_26444_, _08612_, _07233_);
  nand _76881_ (_26445_, _11917_, _06938_);
  and _76882_ (_26446_, _26445_, _25758_);
  and _76883_ (_26447_, _07251_, \oc8051_golden_model_1.PC [5]);
  or _76884_ (_26448_, _26447_, _06938_);
  and _76885_ (_26449_, _26448_, _26446_);
  or _76886_ (_26450_, _26430_, _12214_);
  nand _76887_ (_26451_, _26450_, _12205_);
  or _76888_ (_26452_, _26451_, _26449_);
  and _76889_ (_26454_, _26452_, _07233_);
  or _76890_ (_26455_, _26454_, _26444_);
  or _76891_ (_26456_, _26423_, _12205_);
  and _76892_ (_26457_, _26456_, _26455_);
  nor _76893_ (_26458_, _26457_, _08384_);
  or _76894_ (_26459_, _11919_, _11918_);
  and _76895_ (_26460_, _26459_, _11944_);
  nor _76896_ (_26461_, _26459_, _11944_);
  or _76897_ (_26462_, _26461_, _26460_);
  or _76898_ (_26463_, _26462_, _12197_);
  or _76899_ (_26465_, _12199_, _11917_);
  and _76900_ (_26466_, _26465_, _08384_);
  and _76901_ (_26467_, _26466_, _26463_);
  or _76902_ (_26468_, _26467_, _26458_);
  nand _76903_ (_26469_, _26468_, _06949_);
  and _76904_ (_26470_, _26430_, _06948_);
  nor _76905_ (_26471_, _26470_, _06102_);
  nand _76906_ (_26472_, _26471_, _26469_);
  or _76907_ (_26473_, _12187_, _12069_);
  or _76908_ (_26474_, _26439_, _12189_);
  and _76909_ (_26475_, _26474_, _06102_);
  nand _76910_ (_26476_, _26475_, _26473_);
  and _76911_ (_26477_, _26476_, _12182_);
  nand _76912_ (_26478_, _26477_, _26472_);
  nor _76913_ (_26479_, _26423_, _12182_);
  nor _76914_ (_26480_, _26479_, _06043_);
  nand _76915_ (_26481_, _26480_, _26478_);
  and _76916_ (_26482_, _11916_, _06043_);
  nor _76917_ (_26483_, _26482_, _07272_);
  nand _76918_ (_26484_, _26483_, _26481_);
  and _76919_ (_26486_, _08612_, _07272_);
  nor _76920_ (_26487_, _26486_, _06239_);
  nand _76921_ (_26488_, _26487_, _26484_);
  and _76922_ (_26489_, _11916_, _06239_);
  nor _76923_ (_26490_, _26489_, _12232_);
  nand _76924_ (_26491_, _26490_, _26488_);
  nor _76925_ (_26492_, _26423_, _12231_);
  nor _76926_ (_26493_, _26492_, _06219_);
  nand _76927_ (_26494_, _26493_, _26491_);
  and _76928_ (_26495_, _11916_, _06219_);
  nor _76929_ (_26497_, _26495_, _12241_);
  nand _76930_ (_26498_, _26497_, _26494_);
  nor _76931_ (_26499_, _26423_, _12239_);
  nor _76932_ (_26500_, _26499_, _06039_);
  nand _76933_ (_26501_, _26500_, _26498_);
  and _76934_ (_26502_, _11916_, _06039_);
  nor _76935_ (_26503_, _26502_, _12243_);
  nand _76936_ (_26504_, _26503_, _26501_);
  and _76937_ (_26505_, _08612_, _12243_);
  nor _76938_ (_26506_, _26505_, _06038_);
  nand _76939_ (_26508_, _26506_, _26504_);
  and _76940_ (_26509_, _11916_, _06038_);
  nor _76941_ (_26510_, _26509_, _12256_);
  and _76942_ (_26511_, _26510_, _26508_);
  and _76943_ (_26512_, _12289_, _12069_);
  not _76944_ (_26513_, _26439_);
  nor _76945_ (_26514_, _26513_, _12289_);
  or _76946_ (_26515_, _26514_, _26512_);
  nor _76947_ (_26516_, _26515_, _12255_);
  or _76948_ (_26517_, _26516_, _26511_);
  nand _76949_ (_26518_, _26517_, _12258_);
  nand _76950_ (_26519_, _26518_, _26443_);
  nand _76951_ (_26520_, _26519_, _06509_);
  nor _76952_ (_26521_, _26513_, _12310_);
  not _76953_ (_26522_, _26521_);
  and _76954_ (_26523_, _12310_, _12069_);
  nor _76955_ (_26524_, _26523_, _06509_);
  and _76956_ (_26525_, _26524_, _26522_);
  nor _76957_ (_26526_, _26525_, _06115_);
  nand _76958_ (_26527_, _26526_, _26520_);
  nor _76959_ (_26530_, _26439_, _12329_);
  and _76960_ (_26531_, _12329_, _12070_);
  nor _76961_ (_26532_, _26531_, _12298_);
  not _76962_ (_26533_, _26532_);
  nor _76963_ (_26534_, _26533_, _26530_);
  nor _76964_ (_26535_, _26534_, _12012_);
  and _76965_ (_26536_, _26535_, _26527_);
  or _76966_ (_26537_, _26536_, _26434_);
  nand _76967_ (_26538_, _26537_, _06033_);
  and _76968_ (_26539_, _11917_, _06032_);
  nor _76969_ (_26541_, _26539_, _07355_);
  nand _76970_ (_26542_, _26541_, _26538_);
  nor _76971_ (_26543_, _08612_, _05686_);
  nor _76972_ (_26544_, _26543_, _25133_);
  and _76973_ (_26545_, _26544_, _26542_);
  nor _76974_ (_26546_, _12344_, _11916_);
  or _76975_ (_26547_, _26546_, _26545_);
  nand _76976_ (_26548_, _26547_, _12351_);
  nor _76977_ (_26549_, _26423_, _12351_);
  nor _76978_ (_26550_, _26549_, _06251_);
  nand _76979_ (_26552_, _26550_, _26548_);
  and _76980_ (_26553_, _11916_, _06251_);
  nor _76981_ (_26554_, _26553_, _24866_);
  nand _76982_ (_26555_, _26554_, _26552_);
  and _76983_ (_26556_, _08612_, _24866_);
  nor _76984_ (_26557_, _26556_, _06250_);
  nand _76985_ (_26558_, _26557_, _26555_);
  and _76986_ (_26559_, _11916_, _06250_);
  nor _76987_ (_26560_, _26559_, _12368_);
  and _76988_ (_26561_, _26560_, _26558_);
  nor _76989_ (_26563_, _26423_, _12362_);
  or _76990_ (_26564_, _26563_, _26561_);
  nand _76991_ (_26565_, _26564_, _12366_);
  nor _76992_ (_26566_, _11916_, _12366_);
  nor _76993_ (_26567_, _26566_, _05676_);
  nand _76994_ (_26568_, _26567_, _26565_);
  nor _76995_ (_26569_, _26430_, _05675_);
  nor _76996_ (_26570_, _26569_, _06026_);
  and _76997_ (_26571_, _26570_, _26568_);
  and _76998_ (_26572_, _11917_, _06026_);
  or _76999_ (_26574_, _26572_, _26571_);
  nand _77000_ (_26575_, _26574_, _05673_);
  and _77001_ (_26576_, _08612_, _06023_);
  nor _77002_ (_26577_, _26576_, _06110_);
  nand _77003_ (_26578_, _26577_, _26575_);
  and _77004_ (_26579_, _12069_, _06110_);
  nor _77005_ (_26580_, _26579_, _09818_);
  nand _77006_ (_26581_, _26580_, _26578_);
  nor _77007_ (_26582_, _11916_, _09817_);
  nor _77008_ (_26583_, _26582_, _09833_);
  nand _77009_ (_26585_, _26583_, _26581_);
  nor _77010_ (_26586_, _12070_, _05669_);
  nor _77011_ (_26587_, _26586_, _12393_);
  nand _77012_ (_26588_, _26587_, _26585_);
  nor _77013_ (_26589_, _26423_, _12389_);
  nor _77014_ (_26590_, _26589_, _06089_);
  nand _77015_ (_26591_, _26590_, _26588_);
  and _77016_ (_26592_, _11916_, _06089_);
  nor _77017_ (_26593_, _26592_, _05719_);
  nand _77018_ (_26594_, _26593_, _26591_);
  and _77019_ (_26596_, _08612_, _05719_);
  nor _77020_ (_26597_, _26596_, _12397_);
  nand _77021_ (_26598_, _26597_, _26594_);
  nor _77022_ (_26599_, _26462_, _12398_);
  nor _77023_ (_26600_, _26599_, _08743_);
  and _77024_ (_26601_, _26600_, _26598_);
  or _77025_ (_26602_, _26601_, _26433_);
  nand _77026_ (_26603_, _26602_, _06020_);
  and _77027_ (_26604_, _12070_, _06019_);
  nor _77028_ (_26605_, _26604_, _10661_);
  and _77029_ (_26607_, _26605_, _26603_);
  and _77030_ (_26608_, _11916_, _10661_);
  or _77031_ (_26609_, _26608_, _26607_);
  nand _77032_ (_26610_, _26609_, _12413_);
  and _77033_ (_26611_, _12433_, _12426_);
  nor _77034_ (_26612_, _26611_, _12434_);
  and _77035_ (_26613_, _26612_, _12412_);
  nor _77036_ (_26614_, _26613_, _06088_);
  and _77037_ (_26615_, _26614_, _26610_);
  and _77038_ (_26616_, _11917_, _06088_);
  or _77039_ (_26618_, _26616_, _26615_);
  nand _77040_ (_26619_, _26618_, _13587_);
  and _77041_ (_26620_, _08612_, _05724_);
  nor _77042_ (_26621_, _26620_, _12453_);
  nand _77043_ (_26622_, _26621_, _26619_);
  and _77044_ (_26623_, _11916_, _11071_);
  nor _77045_ (_26624_, _26462_, _11071_);
  or _77046_ (_26625_, _26624_, _26623_);
  and _77047_ (_26626_, _26625_, _12453_);
  nor _77048_ (_26627_, _26626_, _12006_);
  and _77049_ (_26629_, _26627_, _26622_);
  or _77050_ (_26630_, _26629_, _26432_);
  nand _77051_ (_26631_, _26630_, _12466_);
  nor _77052_ (_26632_, _12466_, _11916_);
  nor _77053_ (_26633_, _26632_, _06112_);
  nand _77054_ (_26634_, _26633_, _26631_);
  and _77055_ (_26635_, _12069_, _06112_);
  nor _77056_ (_26636_, _26635_, _06284_);
  and _77057_ (_26637_, _26636_, _26634_);
  and _77058_ (_26638_, _11917_, _06284_);
  or _77059_ (_26640_, _26638_, _26637_);
  nand _77060_ (_26641_, _26640_, _24769_);
  and _77061_ (_26642_, _08612_, _05727_);
  nor _77062_ (_26643_, _26642_, _12476_);
  nand _77063_ (_26644_, _26643_, _26641_);
  and _77064_ (_26645_, _26462_, _11071_);
  nor _77065_ (_26646_, _11916_, _11071_);
  nor _77066_ (_26647_, _26646_, _12477_);
  not _77067_ (_26648_, _26647_);
  nor _77068_ (_26649_, _26648_, _26645_);
  nor _77069_ (_26651_, _26649_, _12481_);
  and _77070_ (_26652_, _26651_, _26644_);
  or _77071_ (_26653_, _26652_, _26429_);
  nand _77072_ (_26654_, _26653_, _10742_);
  nor _77073_ (_26655_, _11916_, _10742_);
  nor _77074_ (_26656_, _26655_, _06108_);
  nand _77075_ (_26657_, _26656_, _26654_);
  and _77076_ (_26658_, _12069_, _06108_);
  nor _77077_ (_26659_, _26658_, _06277_);
  and _77078_ (_26660_, _26659_, _26657_);
  and _77079_ (_26662_, _11917_, _06277_);
  or _77080_ (_26663_, _26662_, _26660_);
  nand _77081_ (_26664_, _26663_, _24765_);
  and _77082_ (_26665_, _08612_, _05736_);
  nor _77083_ (_26666_, _26665_, _12497_);
  nand _77084_ (_26667_, _26666_, _26664_);
  and _77085_ (_26668_, _11916_, \oc8051_golden_model_1.PSW [7]);
  nor _77086_ (_26669_, _26462_, \oc8051_golden_model_1.PSW [7]);
  or _77087_ (_26670_, _26669_, _26668_);
  and _77088_ (_26671_, _26670_, _12497_);
  nor _77089_ (_26673_, _26671_, _12502_);
  and _77090_ (_26674_, _26673_, _26667_);
  or _77091_ (_26675_, _26674_, _26428_);
  nand _77092_ (_26676_, _26675_, _11986_);
  nor _77093_ (_26677_, _11916_, _11986_);
  nor _77094_ (_26678_, _26677_, _06130_);
  nand _77095_ (_26679_, _26678_, _26676_);
  and _77096_ (_26680_, _12069_, _06130_);
  nor _77097_ (_26681_, _26680_, _06292_);
  and _77098_ (_26682_, _26681_, _26679_);
  and _77099_ (_26684_, _11917_, _06292_);
  or _77100_ (_26685_, _26684_, _26682_);
  nand _77101_ (_26686_, _26685_, _24759_);
  and _77102_ (_26687_, _08612_, _05740_);
  nor _77103_ (_26688_, _26687_, _11982_);
  nand _77104_ (_26689_, _26688_, _26686_);
  nand _77105_ (_26690_, _26462_, \oc8051_golden_model_1.PSW [7]);
  or _77106_ (_26691_, _11916_, \oc8051_golden_model_1.PSW [7]);
  and _77107_ (_26692_, _26691_, _11982_);
  and _77108_ (_26693_, _26692_, _26690_);
  nor _77109_ (_26695_, _26693_, _12525_);
  and _77110_ (_26696_, _26695_, _26689_);
  or _77111_ (_26697_, _26696_, _26427_);
  nand _77112_ (_26698_, _26697_, _10825_);
  nor _77113_ (_26699_, _11916_, _10825_);
  nor _77114_ (_26700_, _26699_, _10854_);
  nand _77115_ (_26701_, _26700_, _26698_);
  and _77116_ (_26702_, _26423_, _10854_);
  nor _77117_ (_26703_, _26702_, _06298_);
  and _77118_ (_26704_, _26703_, _26701_);
  and _77119_ (_26706_, _08888_, _06298_);
  or _77120_ (_26707_, _26706_, _26704_);
  nand _77121_ (_26708_, _26707_, _05734_);
  and _77122_ (_26709_, _08612_, _05732_);
  nor _77123_ (_26710_, _26709_, _06129_);
  nand _77124_ (_26711_, _26710_, _26708_);
  and _77125_ (_26712_, _26513_, _12722_);
  nor _77126_ (_26713_, _12069_, _12722_);
  or _77127_ (_26714_, _26713_, _06306_);
  or _77128_ (_26715_, _26714_, _26712_);
  and _77129_ (_26717_, _26715_, _11872_);
  and _77130_ (_26718_, _26717_, _26711_);
  or _77131_ (_26719_, _26718_, _26426_);
  nand _77132_ (_26720_, _26719_, _10975_);
  nor _77133_ (_26721_, _11916_, _10975_);
  nor _77134_ (_26722_, _26721_, _11015_);
  nand _77135_ (_26723_, _26722_, _26720_);
  and _77136_ (_26724_, _26423_, _11015_);
  nor _77137_ (_26725_, _26724_, _06049_);
  and _77138_ (_26726_, _26725_, _26723_);
  and _77139_ (_26728_, _08888_, _06049_);
  or _77140_ (_26729_, _26728_, _26726_);
  nand _77141_ (_26730_, _26729_, _05748_);
  and _77142_ (_26731_, _08612_, _05747_);
  nor _77143_ (_26732_, _26731_, _06126_);
  nand _77144_ (_26733_, _26732_, _26730_);
  and _77145_ (_26734_, _12070_, _12722_);
  nor _77146_ (_26735_, _26439_, _12722_);
  nor _77147_ (_26736_, _26735_, _26734_);
  and _77148_ (_26737_, _26736_, _06126_);
  nor _77149_ (_26739_, _26737_, _12750_);
  nand _77150_ (_26740_, _26739_, _26733_);
  nor _77151_ (_26741_, _26423_, _12749_);
  nor _77152_ (_26742_, _26741_, _06316_);
  nand _77153_ (_26743_, _26742_, _26740_);
  and _77154_ (_26744_, _11916_, _06316_);
  nor _77155_ (_26745_, _26744_, _25353_);
  and _77156_ (_26746_, _26745_, _26743_);
  nor _77157_ (_26747_, _26423_, _12756_);
  or _77158_ (_26748_, _26747_, _26746_);
  nand _77159_ (_26749_, _26748_, _07059_);
  and _77160_ (_26750_, _08612_, _07458_);
  nor _77161_ (_26751_, _26750_, _05652_);
  nand _77162_ (_26752_, _26751_, _26749_);
  and _77163_ (_26753_, _26736_, _05652_);
  nor _77164_ (_26754_, _26753_, _12772_);
  nand _77165_ (_26755_, _26754_, _26752_);
  nor _77166_ (_26756_, _26423_, _12771_);
  nor _77167_ (_26757_, _26756_, _06047_);
  and _77168_ (_26758_, _26757_, _26755_);
  or _77169_ (_26761_, _26758_, _26425_);
  nand _77170_ (_26762_, _26761_, _12779_);
  nor _77171_ (_26763_, _26430_, _12779_);
  nor _77172_ (_26764_, _26763_, _24749_);
  nand _77173_ (_26765_, _26764_, _26762_);
  and _77174_ (_26766_, _24749_, _08612_);
  nor _77175_ (_26767_, _26766_, _12789_);
  and _77176_ (_26768_, _26767_, _26765_);
  or _77177_ (_26769_, _26768_, _26424_);
  or _77178_ (_26770_, _26769_, _01340_);
  or _77179_ (_26772_, _01336_, \oc8051_golden_model_1.PC [5]);
  and _77180_ (_26773_, _26772_, _42882_);
  and _77181_ (_43422_, _26773_, _26770_);
  and _77182_ (_26774_, _08647_, _07458_);
  and _77183_ (_26775_, _08386_, _11860_);
  nor _77184_ (_26776_, _26775_, \oc8051_golden_model_1.PC [6]);
  nor _77185_ (_26777_, _26776_, _11861_);
  not _77186_ (_26778_, _26777_);
  and _77187_ (_26779_, _26778_, _11015_);
  and _77188_ (_26780_, _12063_, _06130_);
  and _77189_ (_26782_, _12063_, _06108_);
  and _77190_ (_26783_, _12063_, _06112_);
  and _77191_ (_26784_, _11909_, _06088_);
  nor _77192_ (_26785_, _12344_, _11908_);
  and _77193_ (_26786_, _26778_, _12012_);
  nor _77194_ (_26787_, _12106_, _12066_);
  nor _77195_ (_26788_, _26787_, _12107_);
  or _77196_ (_26789_, _26788_, _12172_);
  or _77197_ (_26790_, _12174_, _12062_);
  nand _77198_ (_26791_, _26790_, _26789_);
  nand _77199_ (_26793_, _26791_, _06104_);
  and _77200_ (_26794_, _11909_, _06039_);
  or _77201_ (_26795_, _26788_, _12189_);
  or _77202_ (_26796_, _12187_, _12062_);
  and _77203_ (_26797_, _26796_, _06102_);
  nand _77204_ (_26798_, _26797_, _26795_);
  and _77205_ (_26799_, _11946_, _11913_);
  nor _77206_ (_26800_, _26799_, _11947_);
  nand _77207_ (_26801_, _26800_, _12199_);
  or _77208_ (_26802_, _12199_, _11909_);
  and _77209_ (_26804_, _26802_, _08384_);
  nand _77210_ (_26805_, _26804_, _26801_);
  not _77211_ (_26806_, _12219_);
  and _77212_ (_26807_, _08647_, _06943_);
  and _77213_ (_26808_, _11909_, _06938_);
  nor _77214_ (_26809_, _26808_, _06530_);
  and _77215_ (_26810_, _07251_, \oc8051_golden_model_1.PC [6]);
  or _77216_ (_26811_, _26810_, _06938_);
  and _77217_ (_26812_, _26811_, _26809_);
  nor _77218_ (_26813_, _26778_, _12214_);
  or _77219_ (_26815_, _26813_, _06943_);
  nor _77220_ (_26816_, _26815_, _26812_);
  nor _77221_ (_26817_, _26816_, _26091_);
  not _77222_ (_26818_, _26817_);
  nor _77223_ (_26819_, _26818_, _26807_);
  nor _77224_ (_26820_, _26778_, _12205_);
  nor _77225_ (_26821_, _26820_, _08384_);
  not _77226_ (_26822_, _26821_);
  nor _77227_ (_26823_, _26822_, _26819_);
  nor _77228_ (_26824_, _26823_, _26806_);
  nand _77229_ (_26826_, _26824_, _26805_);
  nand _77230_ (_26827_, _26826_, _26798_);
  nand _77231_ (_26828_, _26827_, _12182_);
  nor _77232_ (_26829_, _26778_, _12225_);
  nor _77233_ (_26830_, _26829_, _06043_);
  nand _77234_ (_26831_, _26830_, _26828_);
  and _77235_ (_26832_, _11909_, _06043_);
  nor _77236_ (_26833_, _26832_, _07272_);
  nand _77237_ (_26834_, _26833_, _26831_);
  nor _77238_ (_26835_, _08647_, _05690_);
  nor _77239_ (_26837_, _26835_, _06239_);
  nand _77240_ (_26838_, _26837_, _26834_);
  and _77241_ (_26839_, _11909_, _06239_);
  nor _77242_ (_26840_, _26839_, _12232_);
  nand _77243_ (_26841_, _26840_, _26838_);
  nor _77244_ (_26842_, _26778_, _12231_);
  nor _77245_ (_26843_, _26842_, _06219_);
  nand _77246_ (_26844_, _26843_, _26841_);
  and _77247_ (_26845_, _11909_, _06219_);
  nor _77248_ (_26846_, _26845_, _12241_);
  nand _77249_ (_26848_, _26846_, _26844_);
  nor _77250_ (_26849_, _26778_, _12239_);
  nor _77251_ (_26850_, _26849_, _06039_);
  and _77252_ (_26851_, _26850_, _26848_);
  or _77253_ (_26852_, _26851_, _26794_);
  nand _77254_ (_26853_, _26852_, _05694_);
  and _77255_ (_26854_, _08647_, _12243_);
  nor _77256_ (_26855_, _26854_, _06038_);
  nand _77257_ (_26856_, _26855_, _26853_);
  and _77258_ (_26857_, _11908_, _06038_);
  nor _77259_ (_26859_, _26857_, _12256_);
  and _77260_ (_26860_, _26859_, _26856_);
  and _77261_ (_26861_, _12289_, _12062_);
  not _77262_ (_26862_, _26861_);
  not _77263_ (_26863_, _26788_);
  nor _77264_ (_26864_, _26863_, _12289_);
  nor _77265_ (_26865_, _26864_, _12255_);
  and _77266_ (_26866_, _26865_, _26862_);
  or _77267_ (_26867_, _26866_, _26860_);
  nand _77268_ (_26868_, _26867_, _12258_);
  nand _77269_ (_26870_, _26868_, _26793_);
  nand _77270_ (_26871_, _26870_, _06509_);
  nor _77271_ (_26872_, _26863_, _12310_);
  not _77272_ (_26873_, _26872_);
  and _77273_ (_26874_, _12310_, _12062_);
  nor _77274_ (_26875_, _26874_, _06509_);
  and _77275_ (_26876_, _26875_, _26873_);
  nor _77276_ (_26877_, _26876_, _06115_);
  nand _77277_ (_26878_, _26877_, _26871_);
  and _77278_ (_26879_, _12329_, _12062_);
  not _77279_ (_26881_, _12329_);
  and _77280_ (_26882_, _26788_, _26881_);
  nor _77281_ (_26883_, _26882_, _26879_);
  nor _77282_ (_26884_, _26883_, _12298_);
  nor _77283_ (_26885_, _26884_, _12012_);
  and _77284_ (_26886_, _26885_, _26878_);
  or _77285_ (_26887_, _26886_, _26786_);
  nand _77286_ (_26888_, _26887_, _06033_);
  and _77287_ (_26889_, _11909_, _06032_);
  nor _77288_ (_26890_, _26889_, _07355_);
  nand _77289_ (_26892_, _26890_, _26888_);
  nor _77290_ (_26893_, _08647_, _05686_);
  nor _77291_ (_26894_, _26893_, _25133_);
  and _77292_ (_26895_, _26894_, _26892_);
  or _77293_ (_26896_, _26895_, _26785_);
  nand _77294_ (_26897_, _26896_, _12351_);
  nor _77295_ (_26898_, _26777_, _12351_);
  nor _77296_ (_26899_, _26898_, _06251_);
  nand _77297_ (_26900_, _26899_, _26897_);
  and _77298_ (_26901_, _11908_, _06251_);
  nor _77299_ (_26903_, _26901_, _24866_);
  nand _77300_ (_26904_, _26903_, _26900_);
  and _77301_ (_26905_, _08647_, _24866_);
  nor _77302_ (_26906_, _26905_, _06250_);
  nand _77303_ (_26907_, _26906_, _26904_);
  and _77304_ (_26908_, _11908_, _06250_);
  nor _77305_ (_26909_, _26908_, _12368_);
  nand _77306_ (_26910_, _26909_, _26907_);
  nor _77307_ (_26911_, _26777_, _12362_);
  nor _77308_ (_26912_, _26911_, _12367_);
  nand _77309_ (_26914_, _26912_, _26910_);
  nor _77310_ (_26915_, _11909_, _12366_);
  nor _77311_ (_26916_, _26915_, _05676_);
  and _77312_ (_26917_, _26916_, _26914_);
  nor _77313_ (_26918_, _26777_, _05675_);
  or _77314_ (_26919_, _26918_, _26917_);
  nand _77315_ (_26920_, _26919_, _06027_);
  and _77316_ (_26921_, _11909_, _06026_);
  nor _77317_ (_26922_, _26921_, _06023_);
  nand _77318_ (_26923_, _26922_, _26920_);
  nor _77319_ (_26925_, _08647_, _05673_);
  nor _77320_ (_26926_, _26925_, _06110_);
  nand _77321_ (_26927_, _26926_, _26923_);
  and _77322_ (_26928_, _12063_, _06110_);
  nor _77323_ (_26929_, _26928_, _09818_);
  nand _77324_ (_26930_, _26929_, _26927_);
  nor _77325_ (_26931_, _11909_, _09817_);
  nor _77326_ (_26932_, _26931_, _09833_);
  nand _77327_ (_26933_, _26932_, _26930_);
  nor _77328_ (_26934_, _12062_, _05669_);
  nor _77329_ (_26936_, _26934_, _12393_);
  nand _77330_ (_26937_, _26936_, _26933_);
  nor _77331_ (_26938_, _26778_, _12389_);
  nor _77332_ (_26939_, _26938_, _06089_);
  nand _77333_ (_26940_, _26939_, _26937_);
  and _77334_ (_26941_, _11909_, _06089_);
  nor _77335_ (_26942_, _26941_, _05719_);
  nand _77336_ (_26943_, _26942_, _26940_);
  nor _77337_ (_26944_, _08647_, _05720_);
  nor _77338_ (_26945_, _26944_, _12397_);
  nand _77339_ (_26947_, _26945_, _26943_);
  nor _77340_ (_26948_, _26800_, _12398_);
  nor _77341_ (_26949_, _26948_, _08743_);
  nand _77342_ (_26950_, _26949_, _26947_);
  nor _77343_ (_26951_, _11909_, _08742_);
  nor _77344_ (_26952_, _26951_, _06019_);
  nand _77345_ (_26953_, _26952_, _26950_);
  and _77346_ (_26954_, _12063_, _06019_);
  nor _77347_ (_26955_, _26954_, _10661_);
  nand _77348_ (_26956_, _26955_, _26953_);
  and _77349_ (_26958_, _11908_, _10661_);
  nor _77350_ (_26959_, _26958_, _12412_);
  and _77351_ (_26960_, _26959_, _26956_);
  and _77352_ (_26961_, _12435_, _12422_);
  nor _77353_ (_26962_, _26961_, _12436_);
  nor _77354_ (_26963_, _26962_, _12413_);
  or _77355_ (_26964_, _26963_, _26960_);
  and _77356_ (_26965_, _26964_, _06636_);
  or _77357_ (_26966_, _26965_, _26784_);
  nand _77358_ (_26967_, _26966_, _13587_);
  and _77359_ (_26969_, _08647_, _05724_);
  nor _77360_ (_26970_, _26969_, _12453_);
  nand _77361_ (_26971_, _26970_, _26967_);
  and _77362_ (_26972_, _11908_, _11071_);
  and _77363_ (_26973_, _26800_, _12459_);
  or _77364_ (_26974_, _26973_, _26972_);
  and _77365_ (_26975_, _26974_, _12453_);
  nor _77366_ (_26976_, _26975_, _12006_);
  nand _77367_ (_26977_, _26976_, _26971_);
  and _77368_ (_26978_, _26778_, _12006_);
  nor _77369_ (_26980_, _26978_, _12467_);
  nand _77370_ (_26981_, _26980_, _26977_);
  nor _77371_ (_26982_, _12466_, _11909_);
  nor _77372_ (_26983_, _26982_, _06112_);
  and _77373_ (_26984_, _26983_, _26981_);
  or _77374_ (_26985_, _26984_, _26783_);
  nand _77375_ (_26986_, _26985_, _08756_);
  and _77376_ (_26987_, _11909_, _06284_);
  nor _77377_ (_26988_, _26987_, _05727_);
  and _77378_ (_26989_, _26988_, _26986_);
  nor _77379_ (_26991_, _08647_, _24769_);
  or _77380_ (_26992_, _26991_, _26989_);
  nand _77381_ (_26993_, _26992_, _12477_);
  nor _77382_ (_26994_, _11909_, _11071_);
  and _77383_ (_26995_, _26800_, _11071_);
  or _77384_ (_26996_, _26995_, _26994_);
  and _77385_ (_26997_, _26996_, _12476_);
  nor _77386_ (_26998_, _26997_, _12481_);
  nand _77387_ (_26999_, _26998_, _26993_);
  nor _77388_ (_27000_, _26777_, _12002_);
  nor _77389_ (_27002_, _27000_, _10743_);
  nand _77390_ (_27003_, _27002_, _26999_);
  nor _77391_ (_27004_, _11909_, _10742_);
  nor _77392_ (_27005_, _27004_, _06108_);
  and _77393_ (_27006_, _27005_, _27003_);
  or _77394_ (_27007_, _27006_, _26782_);
  nand _77395_ (_27008_, _27007_, _06278_);
  and _77396_ (_27009_, _11909_, _06277_);
  nor _77397_ (_27010_, _27009_, _05736_);
  and _77398_ (_27011_, _27010_, _27008_);
  nor _77399_ (_27013_, _08647_, _24765_);
  or _77400_ (_27014_, _27013_, _27011_);
  nand _77401_ (_27015_, _27014_, _12498_);
  and _77402_ (_27016_, _11908_, \oc8051_golden_model_1.PSW [7]);
  and _77403_ (_27017_, _26800_, _10606_);
  or _77404_ (_27018_, _27017_, _27016_);
  and _77405_ (_27019_, _27018_, _12497_);
  nor _77406_ (_27020_, _27019_, _12502_);
  nand _77407_ (_27021_, _27020_, _27015_);
  nor _77408_ (_27022_, _26777_, _11993_);
  nor _77409_ (_27024_, _27022_, _11987_);
  nand _77410_ (_27025_, _27024_, _27021_);
  nor _77411_ (_27026_, _11909_, _11986_);
  nor _77412_ (_27027_, _27026_, _06130_);
  and _77413_ (_27028_, _27027_, _27025_);
  or _77414_ (_27029_, _27028_, _26780_);
  nand _77415_ (_27030_, _27029_, _08782_);
  and _77416_ (_27031_, _11909_, _06292_);
  nor _77417_ (_27032_, _27031_, _05740_);
  and _77418_ (_27033_, _27032_, _27030_);
  nor _77419_ (_27035_, _08647_, _24759_);
  or _77420_ (_27036_, _27035_, _27033_);
  nand _77421_ (_27037_, _27036_, _12518_);
  or _77422_ (_27038_, _26800_, _10606_);
  or _77423_ (_27039_, _11908_, \oc8051_golden_model_1.PSW [7]);
  and _77424_ (_27040_, _27039_, _11982_);
  and _77425_ (_27041_, _27040_, _27038_);
  nor _77426_ (_27042_, _27041_, _12525_);
  nand _77427_ (_27043_, _27042_, _27037_);
  nor _77428_ (_27044_, _26777_, _12523_);
  nor _77429_ (_27046_, _27044_, _10826_);
  nand _77430_ (_27047_, _27046_, _27043_);
  nor _77431_ (_27048_, _11909_, _10825_);
  nor _77432_ (_27049_, _27048_, _10854_);
  nand _77433_ (_27050_, _27049_, _27047_);
  and _77434_ (_27051_, _26778_, _10854_);
  nor _77435_ (_27052_, _27051_, _06298_);
  nand _77436_ (_27053_, _27052_, _27050_);
  and _77437_ (_27054_, _09178_, _06298_);
  nor _77438_ (_27055_, _27054_, _05732_);
  nand _77439_ (_27057_, _27055_, _27053_);
  and _77440_ (_27058_, _08647_, _05732_);
  nor _77441_ (_27059_, _27058_, _06129_);
  nand _77442_ (_27060_, _27059_, _27057_);
  and _77443_ (_27061_, _26863_, _12722_);
  nor _77444_ (_27062_, _12062_, _12722_);
  or _77445_ (_27063_, _27062_, _06306_);
  nor _77446_ (_27064_, _27063_, _27061_);
  nor _77447_ (_27065_, _27064_, _12541_);
  nand _77448_ (_27066_, _27065_, _27060_);
  nor _77449_ (_27068_, _26777_, _11872_);
  nor _77450_ (_27069_, _27068_, _10976_);
  nand _77451_ (_27070_, _27069_, _27066_);
  nor _77452_ (_27071_, _11909_, _10975_);
  nor _77453_ (_27072_, _27071_, _11015_);
  and _77454_ (_27073_, _27072_, _27070_);
  or _77455_ (_27074_, _27073_, _26779_);
  nand _77456_ (_27075_, _27074_, _06050_);
  and _77457_ (_27076_, _08843_, _06049_);
  nor _77458_ (_27077_, _27076_, _05747_);
  nand _77459_ (_27079_, _27077_, _27075_);
  nor _77460_ (_27080_, _08647_, _05748_);
  nor _77461_ (_27081_, _27080_, _06126_);
  and _77462_ (_27082_, _27081_, _27079_);
  nor _77463_ (_27083_, _26788_, _12722_);
  and _77464_ (_27084_, _12063_, _12722_);
  nor _77465_ (_27085_, _27084_, _27083_);
  nor _77466_ (_27086_, _27085_, _06704_);
  or _77467_ (_27087_, _27086_, _27082_);
  and _77468_ (_27088_, _27087_, _12749_);
  nor _77469_ (_27090_, _26777_, _12749_);
  or _77470_ (_27091_, _27090_, _27088_);
  nand _77471_ (_27092_, _27091_, _06718_);
  and _77472_ (_27093_, _11909_, _06316_);
  nor _77473_ (_27094_, _27093_, _25353_);
  nand _77474_ (_27095_, _27094_, _27092_);
  nor _77475_ (_27096_, _26778_, _12756_);
  nor _77476_ (_27097_, _27096_, _07458_);
  and _77477_ (_27098_, _27097_, _27095_);
  or _77478_ (_27099_, _27098_, _26774_);
  nand _77479_ (_27101_, _27099_, _05653_);
  nor _77480_ (_27102_, _27085_, _05653_);
  nor _77481_ (_27103_, _27102_, _12772_);
  nand _77482_ (_27104_, _27103_, _27101_);
  nor _77483_ (_27105_, _26778_, _12771_);
  nor _77484_ (_27106_, _27105_, _06047_);
  nand _77485_ (_27107_, _27106_, _27104_);
  and _77486_ (_27108_, _11909_, _06047_);
  nor _77487_ (_27109_, _27108_, _26405_);
  nand _77488_ (_27110_, _27109_, _27107_);
  nor _77489_ (_27112_, _26778_, _12779_);
  nor _77490_ (_27113_, _27112_, _24749_);
  nand _77491_ (_27114_, _27113_, _27110_);
  and _77492_ (_27115_, _24749_, _08647_);
  nor _77493_ (_27116_, _27115_, _12789_);
  and _77494_ (_27117_, _27116_, _27114_);
  and _77495_ (_27118_, _26777_, _12789_);
  or _77496_ (_27119_, _27118_, _27117_);
  or _77497_ (_27120_, _27119_, _01340_);
  or _77498_ (_27121_, _01336_, \oc8051_golden_model_1.PC [6]);
  and _77499_ (_27123_, _27121_, _42882_);
  and _77500_ (_43423_, _27123_, _27120_);
  and _77501_ (_27124_, _08391_, _06047_);
  and _77502_ (_27125_, _08391_, _06316_);
  nor _77503_ (_27126_, _11861_, \oc8051_golden_model_1.PC [7]);
  nor _77504_ (_27127_, _27126_, _11862_);
  nor _77505_ (_27128_, _27127_, _11872_);
  nor _77506_ (_27129_, _27127_, _12523_);
  nor _77507_ (_27130_, _27127_, _11993_);
  nor _77508_ (_27131_, _27127_, _12002_);
  not _77509_ (_27133_, _27127_);
  and _77510_ (_27134_, _27133_, _12006_);
  nor _77511_ (_27135_, _08742_, _08391_);
  nor _77512_ (_27136_, _12344_, _08391_);
  and _77513_ (_27137_, _27133_, _12012_);
  nor _77514_ (_27138_, _08332_, _07233_);
  nand _77515_ (_27139_, _08524_, _06938_);
  and _77516_ (_27140_, _27139_, _25758_);
  and _77517_ (_27141_, _07251_, \oc8051_golden_model_1.PC [7]);
  or _77518_ (_27142_, _27141_, _06938_);
  and _77519_ (_27144_, _27142_, _27140_);
  or _77520_ (_27145_, _27133_, _12214_);
  nand _77521_ (_27146_, _27145_, _12205_);
  or _77522_ (_27147_, _27146_, _27144_);
  and _77523_ (_27148_, _27147_, _07233_);
  or _77524_ (_27149_, _27148_, _27138_);
  or _77525_ (_27150_, _27127_, _12205_);
  and _77526_ (_27151_, _27150_, _27149_);
  nor _77527_ (_27152_, _27151_, _08384_);
  or _77528_ (_27153_, _11904_, _11905_);
  and _77529_ (_27155_, _27153_, _11948_);
  nor _77530_ (_27156_, _27153_, _11948_);
  nor _77531_ (_27157_, _27156_, _27155_);
  nand _77532_ (_27158_, _27157_, _12199_);
  or _77533_ (_27159_, _12199_, _08524_);
  and _77534_ (_27160_, _27159_, _08384_);
  and _77535_ (_27161_, _27160_, _27158_);
  or _77536_ (_27162_, _27161_, _27152_);
  nand _77537_ (_27163_, _27162_, _06949_);
  and _77538_ (_27164_, _27133_, _06948_);
  nor _77539_ (_27166_, _27164_, _06102_);
  nand _77540_ (_27167_, _27166_, _27163_);
  or _77541_ (_27168_, _12187_, _09141_);
  and _77542_ (_27169_, _12108_, _12059_);
  nor _77543_ (_27170_, _27169_, _12109_);
  or _77544_ (_27171_, _27170_, _12189_);
  and _77545_ (_27172_, _27171_, _06102_);
  nand _77546_ (_27173_, _27172_, _27168_);
  and _77547_ (_27174_, _27173_, _12182_);
  nand _77548_ (_27175_, _27174_, _27167_);
  nor _77549_ (_27177_, _27127_, _12182_);
  nor _77550_ (_27178_, _27177_, _06043_);
  nand _77551_ (_27179_, _27178_, _27175_);
  and _77552_ (_27180_, _08391_, _06043_);
  nor _77553_ (_27181_, _27180_, _07272_);
  nand _77554_ (_27182_, _27181_, _27179_);
  and _77555_ (_27183_, _08332_, _07272_);
  nor _77556_ (_27184_, _27183_, _06239_);
  nand _77557_ (_27185_, _27184_, _27182_);
  and _77558_ (_27186_, _08391_, _06239_);
  nor _77559_ (_27188_, _27186_, _12232_);
  nand _77560_ (_27189_, _27188_, _27185_);
  nor _77561_ (_27190_, _27127_, _12231_);
  nor _77562_ (_27191_, _27190_, _06219_);
  nand _77563_ (_27192_, _27191_, _27189_);
  and _77564_ (_27193_, _08391_, _06219_);
  nor _77565_ (_27194_, _27193_, _12241_);
  nand _77566_ (_27195_, _27194_, _27192_);
  nor _77567_ (_27196_, _27127_, _12239_);
  nor _77568_ (_27197_, _27196_, _06039_);
  nand _77569_ (_27199_, _27197_, _27195_);
  and _77570_ (_27200_, _08391_, _06039_);
  nor _77571_ (_27201_, _27200_, _12243_);
  nand _77572_ (_27202_, _27201_, _27199_);
  and _77573_ (_27203_, _08332_, _12243_);
  nor _77574_ (_27204_, _27203_, _06038_);
  nand _77575_ (_27205_, _27204_, _27202_);
  and _77576_ (_27206_, _08391_, _06038_);
  nor _77577_ (_27207_, _27206_, _12256_);
  nand _77578_ (_27208_, _27207_, _27205_);
  not _77579_ (_27210_, _27170_);
  nor _77580_ (_27211_, _27210_, _12289_);
  not _77581_ (_27212_, _27211_);
  and _77582_ (_27213_, _12289_, _09141_);
  nor _77583_ (_27214_, _27213_, _12255_);
  and _77584_ (_27215_, _27214_, _27212_);
  nor _77585_ (_27216_, _27215_, _06104_);
  nand _77586_ (_27217_, _27216_, _27208_);
  or _77587_ (_27218_, _12174_, _09141_);
  or _77588_ (_27219_, _27170_, _12172_);
  and _77589_ (_27221_, _27219_, _06104_);
  nand _77590_ (_27222_, _27221_, _27218_);
  and _77591_ (_27223_, _27222_, _06509_);
  nand _77592_ (_27224_, _27223_, _27217_);
  nor _77593_ (_27225_, _27210_, _12310_);
  not _77594_ (_27226_, _27225_);
  and _77595_ (_27227_, _12310_, _09141_);
  nor _77596_ (_27228_, _27227_, _06509_);
  and _77597_ (_27229_, _27228_, _27226_);
  nor _77598_ (_27230_, _27229_, _06115_);
  nand _77599_ (_27232_, _27230_, _27224_);
  nor _77600_ (_27233_, _27170_, _12329_);
  and _77601_ (_27234_, _12329_, _09142_);
  nor _77602_ (_27235_, _27234_, _12298_);
  not _77603_ (_27236_, _27235_);
  nor _77604_ (_27237_, _27236_, _27233_);
  nor _77605_ (_27238_, _27237_, _12012_);
  and _77606_ (_27239_, _27238_, _27232_);
  or _77607_ (_27240_, _27239_, _27137_);
  nand _77608_ (_27241_, _27240_, _06033_);
  and _77609_ (_27243_, _08524_, _06032_);
  nor _77610_ (_27244_, _27243_, _07355_);
  nand _77611_ (_27245_, _27244_, _27241_);
  nor _77612_ (_27246_, _08332_, _05686_);
  nor _77613_ (_27247_, _27246_, _25133_);
  and _77614_ (_27248_, _27247_, _27245_);
  or _77615_ (_27249_, _27248_, _27136_);
  nand _77616_ (_27250_, _27249_, _12351_);
  nor _77617_ (_27251_, _27127_, _12351_);
  nor _77618_ (_27252_, _27251_, _06251_);
  nand _77619_ (_27254_, _27252_, _27250_);
  and _77620_ (_27255_, _08391_, _06251_);
  nor _77621_ (_27256_, _27255_, _24866_);
  nand _77622_ (_27257_, _27256_, _27254_);
  and _77623_ (_27258_, _08332_, _24866_);
  nor _77624_ (_27259_, _27258_, _06250_);
  nand _77625_ (_27260_, _27259_, _27257_);
  and _77626_ (_27261_, _08391_, _06250_);
  nor _77627_ (_27262_, _27261_, _12368_);
  and _77628_ (_27263_, _27262_, _27260_);
  nor _77629_ (_27265_, _27127_, _12362_);
  or _77630_ (_27266_, _27265_, _27263_);
  nand _77631_ (_27267_, _27266_, _12366_);
  nor _77632_ (_27268_, _12366_, _08391_);
  nor _77633_ (_27269_, _27268_, _05676_);
  nand _77634_ (_27270_, _27269_, _27267_);
  nor _77635_ (_27271_, _27133_, _05675_);
  nor _77636_ (_27272_, _27271_, _06026_);
  and _77637_ (_27273_, _27272_, _27270_);
  and _77638_ (_27274_, _08524_, _06026_);
  or _77639_ (_27276_, _27274_, _27273_);
  nand _77640_ (_27277_, _27276_, _05673_);
  and _77641_ (_27278_, _08332_, _06023_);
  nor _77642_ (_27279_, _27278_, _06110_);
  nand _77643_ (_27280_, _27279_, _27277_);
  and _77644_ (_27281_, _09141_, _06110_);
  nor _77645_ (_27282_, _27281_, _09818_);
  nand _77646_ (_27283_, _27282_, _27280_);
  nor _77647_ (_27284_, _09817_, _08391_);
  nor _77648_ (_27285_, _27284_, _09833_);
  nand _77649_ (_27287_, _27285_, _27283_);
  nor _77650_ (_27288_, _09142_, _05669_);
  nor _77651_ (_27289_, _27288_, _12393_);
  nand _77652_ (_27290_, _27289_, _27287_);
  nor _77653_ (_27291_, _27127_, _12389_);
  nor _77654_ (_27292_, _27291_, _06089_);
  nand _77655_ (_27293_, _27292_, _27290_);
  and _77656_ (_27294_, _08391_, _06089_);
  nor _77657_ (_27295_, _27294_, _05719_);
  nand _77658_ (_27296_, _27295_, _27293_);
  and _77659_ (_27298_, _08332_, _05719_);
  nor _77660_ (_27299_, _27298_, _12397_);
  nand _77661_ (_27300_, _27299_, _27296_);
  and _77662_ (_27301_, _27157_, _12397_);
  nor _77663_ (_27302_, _27301_, _08743_);
  and _77664_ (_27303_, _27302_, _27300_);
  or _77665_ (_27304_, _27303_, _27135_);
  nand _77666_ (_27305_, _27304_, _06020_);
  and _77667_ (_27306_, _09142_, _06019_);
  nor _77668_ (_27307_, _27306_, _10661_);
  and _77669_ (_27309_, _27307_, _27305_);
  and _77670_ (_27310_, _10661_, _08391_);
  or _77671_ (_27311_, _27310_, _27309_);
  nand _77672_ (_27312_, _27311_, _12413_);
  or _77673_ (_27313_, _12417_, _12418_);
  nor _77674_ (_27314_, _27313_, _12437_);
  and _77675_ (_27315_, _27313_, _12437_);
  nor _77676_ (_27316_, _27315_, _27314_);
  and _77677_ (_27317_, _27316_, _12412_);
  nor _77678_ (_27318_, _27317_, _06088_);
  and _77679_ (_27320_, _27318_, _27312_);
  and _77680_ (_27321_, _08524_, _06088_);
  or _77681_ (_27322_, _27321_, _27320_);
  nand _77682_ (_27323_, _27322_, _13587_);
  and _77683_ (_27324_, _08332_, _05724_);
  nor _77684_ (_27325_, _27324_, _12453_);
  nand _77685_ (_27326_, _27325_, _27323_);
  and _77686_ (_27327_, _11071_, _08391_);
  and _77687_ (_27328_, _27157_, _12459_);
  or _77688_ (_27329_, _27328_, _27327_);
  and _77689_ (_27330_, _27329_, _12453_);
  nor _77690_ (_27331_, _27330_, _12006_);
  and _77691_ (_27332_, _27331_, _27326_);
  or _77692_ (_27333_, _27332_, _27134_);
  nand _77693_ (_27334_, _27333_, _12466_);
  nor _77694_ (_27335_, _12466_, _08391_);
  nor _77695_ (_27336_, _27335_, _06112_);
  nand _77696_ (_27337_, _27336_, _27334_);
  and _77697_ (_27338_, _09141_, _06112_);
  nor _77698_ (_27339_, _27338_, _06284_);
  and _77699_ (_27342_, _27339_, _27337_);
  and _77700_ (_27343_, _08524_, _06284_);
  or _77701_ (_27344_, _27343_, _27342_);
  nand _77702_ (_27345_, _27344_, _24769_);
  and _77703_ (_27346_, _08332_, _05727_);
  nor _77704_ (_27347_, _27346_, _12476_);
  nand _77705_ (_27348_, _27347_, _27345_);
  nor _77706_ (_27349_, _27157_, _12459_);
  nor _77707_ (_27350_, _11071_, _08391_);
  nor _77708_ (_27351_, _27350_, _12477_);
  not _77709_ (_27353_, _27351_);
  nor _77710_ (_27354_, _27353_, _27349_);
  nor _77711_ (_27355_, _27354_, _12481_);
  and _77712_ (_27356_, _27355_, _27348_);
  or _77713_ (_27357_, _27356_, _27131_);
  nand _77714_ (_27358_, _27357_, _10742_);
  nor _77715_ (_27359_, _10742_, _08391_);
  nor _77716_ (_27360_, _27359_, _06108_);
  nand _77717_ (_27361_, _27360_, _27358_);
  and _77718_ (_27362_, _09141_, _06108_);
  nor _77719_ (_27364_, _27362_, _06277_);
  and _77720_ (_27365_, _27364_, _27361_);
  and _77721_ (_27366_, _08524_, _06277_);
  or _77722_ (_27367_, _27366_, _27365_);
  nand _77723_ (_27368_, _27367_, _24765_);
  and _77724_ (_27369_, _08332_, _05736_);
  nor _77725_ (_27370_, _27369_, _12497_);
  nand _77726_ (_27371_, _27370_, _27368_);
  and _77727_ (_27372_, _08391_, \oc8051_golden_model_1.PSW [7]);
  and _77728_ (_27373_, _27157_, _10606_);
  or _77729_ (_27375_, _27373_, _27372_);
  and _77730_ (_27376_, _27375_, _12497_);
  nor _77731_ (_27377_, _27376_, _12502_);
  and _77732_ (_27378_, _27377_, _27371_);
  or _77733_ (_27379_, _27378_, _27130_);
  nand _77734_ (_27380_, _27379_, _11986_);
  nor _77735_ (_27381_, _11986_, _08391_);
  nor _77736_ (_27382_, _27381_, _06130_);
  nand _77737_ (_27383_, _27382_, _27380_);
  and _77738_ (_27384_, _09141_, _06130_);
  nor _77739_ (_27386_, _27384_, _06292_);
  and _77740_ (_27387_, _27386_, _27383_);
  and _77741_ (_27388_, _08524_, _06292_);
  or _77742_ (_27389_, _27388_, _27387_);
  nand _77743_ (_27390_, _27389_, _24759_);
  and _77744_ (_27391_, _08332_, _05740_);
  nor _77745_ (_27392_, _27391_, _11982_);
  nand _77746_ (_27393_, _27392_, _27390_);
  and _77747_ (_27394_, _08391_, _10606_);
  and _77748_ (_27395_, _27157_, \oc8051_golden_model_1.PSW [7]);
  or _77749_ (_27397_, _27395_, _27394_);
  and _77750_ (_27398_, _27397_, _11982_);
  nor _77751_ (_27399_, _27398_, _12525_);
  and _77752_ (_27400_, _27399_, _27393_);
  or _77753_ (_27401_, _27400_, _27129_);
  nand _77754_ (_27402_, _27401_, _10825_);
  nor _77755_ (_27403_, _10825_, _08391_);
  nor _77756_ (_27404_, _27403_, _10854_);
  nand _77757_ (_27405_, _27404_, _27402_);
  and _77758_ (_27406_, _27127_, _10854_);
  nor _77759_ (_27408_, _27406_, _06298_);
  and _77760_ (_27409_, _27408_, _27405_);
  and _77761_ (_27410_, _08798_, _06298_);
  or _77762_ (_27411_, _27410_, _27409_);
  nand _77763_ (_27412_, _27411_, _05734_);
  and _77764_ (_27413_, _08332_, _05732_);
  nor _77765_ (_27414_, _27413_, _06129_);
  nand _77766_ (_27415_, _27414_, _27412_);
  and _77767_ (_27416_, _27210_, _12722_);
  nor _77768_ (_27417_, _09141_, _12722_);
  or _77769_ (_27419_, _27417_, _06306_);
  nor _77770_ (_27420_, _27419_, _27416_);
  nor _77771_ (_27421_, _27420_, _12541_);
  and _77772_ (_27422_, _27421_, _27415_);
  or _77773_ (_27423_, _27422_, _27128_);
  nand _77774_ (_27424_, _27423_, _10975_);
  nor _77775_ (_27425_, _10975_, _08391_);
  nor _77776_ (_27426_, _27425_, _11015_);
  nand _77777_ (_27427_, _27426_, _27424_);
  and _77778_ (_27428_, _27127_, _11015_);
  nor _77779_ (_27430_, _27428_, _06049_);
  and _77780_ (_27431_, _27430_, _27427_);
  and _77781_ (_27432_, _08798_, _06049_);
  or _77782_ (_27433_, _27432_, _27431_);
  nand _77783_ (_27434_, _27433_, _05748_);
  and _77784_ (_27435_, _08332_, _05747_);
  nor _77785_ (_27436_, _27435_, _06126_);
  nand _77786_ (_27437_, _27436_, _27434_);
  and _77787_ (_27438_, _09142_, _12722_);
  nor _77788_ (_27439_, _27170_, _12722_);
  nor _77789_ (_27441_, _27439_, _27438_);
  and _77790_ (_27442_, _27441_, _06126_);
  nor _77791_ (_27443_, _27442_, _12750_);
  nand _77792_ (_27444_, _27443_, _27437_);
  nor _77793_ (_27445_, _27127_, _12749_);
  nor _77794_ (_27446_, _27445_, _06316_);
  and _77795_ (_27447_, _27446_, _27444_);
  or _77796_ (_27448_, _27447_, _27125_);
  nand _77797_ (_27449_, _27448_, _12756_);
  nor _77798_ (_27450_, _27133_, _12756_);
  nor _77799_ (_27452_, _27450_, _07458_);
  nand _77800_ (_27453_, _27452_, _27449_);
  and _77801_ (_27454_, _08332_, _07458_);
  nor _77802_ (_27455_, _27454_, _05652_);
  nand _77803_ (_27456_, _27455_, _27453_);
  and _77804_ (_27457_, _27441_, _05652_);
  nor _77805_ (_27458_, _27457_, _12772_);
  nand _77806_ (_27459_, _27458_, _27456_);
  nor _77807_ (_27460_, _27127_, _12771_);
  nor _77808_ (_27461_, _27460_, _06047_);
  and _77809_ (_27463_, _27461_, _27459_);
  or _77810_ (_27464_, _27463_, _27124_);
  nand _77811_ (_27465_, _27464_, _12779_);
  nor _77812_ (_27466_, _27133_, _12779_);
  nor _77813_ (_27467_, _27466_, _24749_);
  nand _77814_ (_27468_, _27467_, _27465_);
  and _77815_ (_27469_, _24749_, _08332_);
  nor _77816_ (_27470_, _27469_, _12789_);
  and _77817_ (_27471_, _27470_, _27468_);
  and _77818_ (_27472_, _27127_, _12789_);
  or _77819_ (_27474_, _27472_, _27471_);
  or _77820_ (_27475_, _27474_, _01340_);
  or _77821_ (_27476_, _01336_, \oc8051_golden_model_1.PC [7]);
  and _77822_ (_27477_, _27476_, _42882_);
  and _77823_ (_43425_, _27477_, _27475_);
  and _77824_ (_27478_, _11862_, \oc8051_golden_model_1.PC [8]);
  nor _77825_ (_27479_, _11862_, \oc8051_golden_model_1.PC [8]);
  nor _77826_ (_27480_, _27479_, _27478_);
  nor _77827_ (_27481_, _27480_, _12779_);
  nor _77828_ (_27482_, _09200_, _06016_);
  nor _77829_ (_27484_, _11982_, _05740_);
  nor _77830_ (_27485_, _11952_, _08742_);
  and _77831_ (_27486_, _11952_, _06089_);
  or _77832_ (_27487_, _27480_, _05675_);
  and _77833_ (_27488_, _11952_, _06039_);
  nor _77834_ (_27489_, _06239_, _07272_);
  and _77835_ (_27490_, _11952_, _06043_);
  and _77836_ (_27491_, _12205_, _07251_);
  or _77837_ (_27492_, _27491_, _27480_);
  nand _77838_ (_27493_, _14066_, _06938_);
  and _77839_ (_27495_, _27493_, _25758_);
  or _77840_ (_27496_, _06938_, \oc8051_golden_model_1.PC [8]);
  or _77841_ (_27497_, _27496_, _07250_);
  nand _77842_ (_27498_, _27497_, _27495_);
  nand _77843_ (_27499_, _27498_, _24785_);
  and _77844_ (_27500_, _27499_, _27492_);
  and _77845_ (_27501_, _27480_, _06530_);
  or _77846_ (_27502_, _27501_, _08384_);
  or _77847_ (_27503_, _27502_, _27500_);
  nor _77848_ (_27504_, _11955_, _11950_);
  nor _77849_ (_27506_, _27504_, _11956_);
  and _77850_ (_27507_, _27506_, _12199_);
  and _77851_ (_27508_, _12197_, _11952_);
  or _77852_ (_27509_, _27508_, _08383_);
  or _77853_ (_27510_, _27509_, _27507_);
  and _77854_ (_27511_, _27510_, _27503_);
  or _77855_ (_27512_, _27511_, _06948_);
  not _77856_ (_27513_, _27480_);
  nand _77857_ (_27514_, _27513_, _06948_);
  and _77858_ (_27515_, _27514_, _06954_);
  and _77859_ (_27517_, _27515_, _27512_);
  and _77860_ (_27518_, _12117_, _12110_);
  nor _77861_ (_27519_, _27518_, _12118_);
  or _77862_ (_27520_, _27519_, _12189_);
  or _77863_ (_27521_, _12187_, _12112_);
  and _77864_ (_27522_, _27521_, _06102_);
  and _77865_ (_27523_, _27522_, _27520_);
  or _77866_ (_27524_, _27523_, _24805_);
  or _77867_ (_27525_, _27524_, _27517_);
  or _77868_ (_27526_, _27480_, _12182_);
  and _77869_ (_27528_, _27526_, _06044_);
  and _77870_ (_27529_, _27528_, _27525_);
  or _77871_ (_27530_, _27529_, _27490_);
  and _77872_ (_27531_, _27530_, _27489_);
  nand _77873_ (_27532_, _11952_, _06239_);
  nand _77874_ (_27533_, _27532_, _12231_);
  or _77875_ (_27534_, _27533_, _27531_);
  or _77876_ (_27535_, _27480_, _12231_);
  and _77877_ (_27536_, _27535_, _06220_);
  and _77878_ (_27537_, _27536_, _27534_);
  nand _77879_ (_27539_, _11952_, _06219_);
  nand _77880_ (_27540_, _27539_, _12239_);
  or _77881_ (_27541_, _27540_, _27537_);
  or _77882_ (_27542_, _27480_, _12239_);
  and _77883_ (_27543_, _27542_, _06040_);
  and _77884_ (_27544_, _27543_, _27541_);
  or _77885_ (_27545_, _27544_, _27488_);
  and _77886_ (_27546_, _27545_, _12244_);
  nand _77887_ (_27547_, _11952_, _06038_);
  nand _77888_ (_27548_, _27547_, _12255_);
  or _77889_ (_27550_, _27548_, _27546_);
  not _77890_ (_27551_, _27519_);
  nor _77891_ (_27552_, _27551_, _12289_);
  and _77892_ (_27553_, _12289_, _12112_);
  or _77893_ (_27554_, _27553_, _12255_);
  or _77894_ (_27555_, _27554_, _27552_);
  and _77895_ (_27556_, _27555_, _12258_);
  and _77896_ (_27557_, _27556_, _27550_);
  and _77897_ (_27558_, _27519_, _12174_);
  and _77898_ (_27559_, _12172_, _12112_);
  or _77899_ (_27561_, _27559_, _27558_);
  and _77900_ (_27562_, _27561_, _06104_);
  or _77901_ (_27563_, _27562_, _06121_);
  or _77902_ (_27564_, _27563_, _27557_);
  nor _77903_ (_27565_, _27551_, _12310_);
  and _77904_ (_27566_, _12310_, _12112_);
  or _77905_ (_27567_, _27566_, _06509_);
  or _77906_ (_27568_, _27567_, _27565_);
  and _77907_ (_27569_, _27568_, _12298_);
  and _77908_ (_27570_, _27569_, _27564_);
  or _77909_ (_27572_, _27519_, _12329_);
  nand _77910_ (_27573_, _12329_, _12113_);
  and _77911_ (_27574_, _27573_, _06115_);
  and _77912_ (_27575_, _27574_, _27572_);
  or _77913_ (_27576_, _27575_, _12012_);
  or _77914_ (_27577_, _27576_, _27570_);
  nand _77915_ (_27578_, _27513_, _12012_);
  and _77916_ (_27579_, _27578_, _06033_);
  and _77917_ (_27580_, _27579_, _27577_);
  and _77918_ (_27581_, _11952_, _06032_);
  or _77919_ (_27583_, _27581_, _07355_);
  or _77920_ (_27584_, _27583_, _27580_);
  and _77921_ (_27585_, _27584_, _12344_);
  nor _77922_ (_27586_, _12344_, _14066_);
  or _77923_ (_27587_, _27586_, _12355_);
  or _77924_ (_27588_, _27587_, _27585_);
  or _77925_ (_27589_, _27480_, _12351_);
  and _77926_ (_27590_, _27589_, _13765_);
  and _77927_ (_27591_, _27590_, _27588_);
  and _77928_ (_27592_, _11952_, _06251_);
  or _77929_ (_27594_, _27592_, _24866_);
  or _77930_ (_27595_, _27594_, _27591_);
  and _77931_ (_27596_, _27595_, _13764_);
  nand _77932_ (_27597_, _11952_, _06250_);
  nand _77933_ (_27598_, _27597_, _12362_);
  or _77934_ (_27599_, _27598_, _27596_);
  or _77935_ (_27600_, _27480_, _12362_);
  and _77936_ (_27601_, _27600_, _12366_);
  and _77937_ (_27602_, _27601_, _27599_);
  nor _77938_ (_27603_, _14066_, _12366_);
  or _77939_ (_27605_, _27603_, _05676_);
  or _77940_ (_27606_, _27605_, _27602_);
  and _77941_ (_27607_, _27606_, _27487_);
  or _77942_ (_27608_, _27607_, _06026_);
  nand _77943_ (_27609_, _14066_, _06026_);
  nor _77944_ (_27610_, _06110_, _06023_);
  and _77945_ (_27611_, _27610_, _27609_);
  and _77946_ (_27612_, _27611_, _27608_);
  and _77947_ (_27613_, _12112_, _06110_);
  or _77948_ (_27614_, _27613_, _09818_);
  or _77949_ (_27616_, _27614_, _27612_);
  nor _77950_ (_27617_, _11952_, _09817_);
  nor _77951_ (_27618_, _27617_, _09833_);
  nand _77952_ (_27619_, _27618_, _27616_);
  nor _77953_ (_27620_, _12113_, _05669_);
  nor _77954_ (_27621_, _27620_, _12393_);
  nand _77955_ (_27622_, _27621_, _27619_);
  nor _77956_ (_27623_, _27480_, _12389_);
  nor _77957_ (_27624_, _27623_, _06089_);
  and _77958_ (_27625_, _27624_, _27622_);
  or _77959_ (_27627_, _27625_, _27486_);
  nor _77960_ (_27628_, _12397_, _05719_);
  nand _77961_ (_27629_, _27628_, _27627_);
  and _77962_ (_27630_, _27506_, _12397_);
  nor _77963_ (_27631_, _27630_, _08743_);
  and _77964_ (_27632_, _27631_, _27629_);
  or _77965_ (_27633_, _27632_, _27485_);
  nand _77966_ (_27634_, _27633_, _06020_);
  and _77967_ (_27635_, _12113_, _06019_);
  nor _77968_ (_27636_, _27635_, _10661_);
  nand _77969_ (_27638_, _27636_, _27634_);
  and _77970_ (_27639_, _11952_, _10661_);
  nor _77971_ (_27640_, _27639_, _12412_);
  nand _77972_ (_27641_, _27640_, _27638_);
  nor _77973_ (_27642_, _12439_, \oc8051_golden_model_1.DPH [0]);
  nor _77974_ (_27643_, _27642_, _12440_);
  nor _77975_ (_27644_, _27643_, _12413_);
  nor _77976_ (_27645_, _27644_, _06088_);
  nand _77977_ (_27646_, _27645_, _27641_);
  and _77978_ (_27647_, _11952_, _06088_);
  nor _77979_ (_27649_, _27647_, _05724_);
  nand _77980_ (_27650_, _27649_, _27646_);
  nand _77981_ (_27651_, _27650_, _12454_);
  and _77982_ (_27652_, _11952_, _11071_);
  and _77983_ (_27653_, _27506_, _12459_);
  or _77984_ (_27654_, _27653_, _27652_);
  and _77985_ (_27655_, _27654_, _12453_);
  nor _77986_ (_27656_, _27655_, _12006_);
  nand _77987_ (_27657_, _27656_, _27651_);
  and _77988_ (_27658_, _27513_, _12006_);
  nor _77989_ (_27660_, _27658_, _12467_);
  nand _77990_ (_27661_, _27660_, _27657_);
  nor _77991_ (_27662_, _12466_, _14066_);
  nor _77992_ (_27663_, _27662_, _06112_);
  nand _77993_ (_27664_, _27663_, _27661_);
  and _77994_ (_27665_, _12113_, _06112_);
  nor _77995_ (_27666_, _27665_, _06284_);
  nand _77996_ (_27667_, _27666_, _27664_);
  and _77997_ (_27668_, _11952_, _06284_);
  nor _77998_ (_27669_, _27668_, _05727_);
  nand _77999_ (_27671_, _27669_, _27667_);
  nand _78000_ (_27672_, _27671_, _12477_);
  nor _78001_ (_27673_, _27506_, _12459_);
  nor _78002_ (_27674_, _11952_, _11071_);
  nor _78003_ (_27675_, _27674_, _12477_);
  not _78004_ (_27676_, _27675_);
  nor _78005_ (_27677_, _27676_, _27673_);
  nor _78006_ (_27678_, _27677_, _12481_);
  nand _78007_ (_27679_, _27678_, _27672_);
  nor _78008_ (_27680_, _27480_, _12002_);
  nor _78009_ (_27682_, _27680_, _10743_);
  nand _78010_ (_27683_, _27682_, _27679_);
  nor _78011_ (_27684_, _14066_, _10742_);
  nor _78012_ (_27685_, _27684_, _06108_);
  and _78013_ (_27686_, _27685_, _27683_);
  and _78014_ (_27687_, _12113_, _06108_);
  or _78015_ (_27688_, _27687_, _27686_);
  nand _78016_ (_27689_, _27688_, _06278_);
  nor _78017_ (_27690_, _12497_, _05736_);
  and _78018_ (_27691_, _14066_, _06277_);
  not _78019_ (_27693_, _27691_);
  and _78020_ (_27694_, _27693_, _27690_);
  nand _78021_ (_27695_, _27694_, _27689_);
  and _78022_ (_27696_, _11952_, \oc8051_golden_model_1.PSW [7]);
  and _78023_ (_27697_, _27506_, _10606_);
  or _78024_ (_27698_, _27697_, _27696_);
  and _78025_ (_27699_, _27698_, _12497_);
  nor _78026_ (_27700_, _27699_, _12502_);
  nand _78027_ (_27701_, _27700_, _27695_);
  nor _78028_ (_27702_, _27480_, _11993_);
  nor _78029_ (_27704_, _27702_, _11987_);
  and _78030_ (_27705_, _27704_, _27701_);
  nor _78031_ (_27706_, _14066_, _11986_);
  or _78032_ (_27707_, _27706_, _06130_);
  or _78033_ (_27708_, _27707_, _27705_);
  and _78034_ (_27709_, _12113_, _06130_);
  nor _78035_ (_27710_, _27709_, _06292_);
  and _78036_ (_27711_, _27710_, _27708_);
  and _78037_ (_27712_, _11952_, _06292_);
  or _78038_ (_27713_, _27712_, _27711_);
  nand _78039_ (_27715_, _27713_, _27484_);
  and _78040_ (_27716_, _11952_, _10606_);
  and _78041_ (_27717_, _27506_, \oc8051_golden_model_1.PSW [7]);
  or _78042_ (_27718_, _27717_, _27716_);
  and _78043_ (_27719_, _27718_, _11982_);
  nor _78044_ (_27720_, _27719_, _12525_);
  nand _78045_ (_27721_, _27720_, _27715_);
  nor _78046_ (_27722_, _27480_, _12523_);
  nor _78047_ (_27723_, _27722_, _10826_);
  and _78048_ (_27724_, _27723_, _27721_);
  nor _78049_ (_27726_, _14066_, _10825_);
  or _78050_ (_27727_, _27726_, _10854_);
  or _78051_ (_27728_, _27727_, _27724_);
  and _78052_ (_27729_, _27513_, _10854_);
  nor _78053_ (_27730_, _27729_, _06298_);
  nand _78054_ (_27731_, _27730_, _27728_);
  and _78055_ (_27732_, _06931_, _06298_);
  nor _78056_ (_27733_, _27732_, _05732_);
  nand _78057_ (_27734_, _27733_, _27731_);
  nand _78058_ (_27735_, _27734_, _06306_);
  nor _78059_ (_27737_, _12112_, _12722_);
  and _78060_ (_27738_, _27551_, _12722_);
  or _78061_ (_27739_, _27738_, _06306_);
  nor _78062_ (_27740_, _27739_, _27737_);
  nor _78063_ (_27741_, _27740_, _12541_);
  nand _78064_ (_27742_, _27741_, _27735_);
  nor _78065_ (_27743_, _27480_, _11872_);
  nor _78066_ (_27744_, _27743_, _10976_);
  nand _78067_ (_27745_, _27744_, _27742_);
  nor _78068_ (_27746_, _14066_, _10975_);
  nor _78069_ (_27748_, _27746_, _11015_);
  nand _78070_ (_27749_, _27748_, _27745_);
  and _78071_ (_27750_, _27513_, _11015_);
  nor _78072_ (_27751_, _27750_, _06049_);
  nand _78073_ (_27752_, _27751_, _27749_);
  and _78074_ (_27753_, _06931_, _06049_);
  nor _78075_ (_27754_, _27753_, _05747_);
  nand _78076_ (_27755_, _27754_, _27752_);
  nand _78077_ (_27756_, _27755_, _06704_);
  and _78078_ (_27757_, _12113_, _12722_);
  nor _78079_ (_27759_, _27519_, _12722_);
  nor _78080_ (_27760_, _27759_, _27757_);
  and _78081_ (_27761_, _27760_, _06126_);
  nor _78082_ (_27762_, _27761_, _12750_);
  nand _78083_ (_27763_, _27762_, _27756_);
  nor _78084_ (_27764_, _27480_, _12749_);
  nor _78085_ (_27765_, _27764_, _06316_);
  nand _78086_ (_27766_, _27765_, _27763_);
  and _78087_ (_27767_, _11952_, _06316_);
  nor _78088_ (_27768_, _27767_, _25353_);
  nand _78089_ (_27770_, _27768_, _27766_);
  nor _78090_ (_27771_, _27480_, _12756_);
  nor _78091_ (_27772_, _27771_, _06127_);
  and _78092_ (_27773_, _27772_, _27770_);
  or _78093_ (_27774_, _27773_, _27482_);
  nor _78094_ (_27775_, _05752_, _05652_);
  nand _78095_ (_27776_, _27775_, _27774_);
  and _78096_ (_27777_, _27760_, _05652_);
  nor _78097_ (_27778_, _27777_, _12772_);
  nand _78098_ (_27779_, _27778_, _27776_);
  nor _78099_ (_27781_, _27480_, _12771_);
  nor _78100_ (_27782_, _27781_, _06047_);
  nand _78101_ (_27783_, _27782_, _27779_);
  and _78102_ (_27784_, _11952_, _06047_);
  nor _78103_ (_27785_, _27784_, _26405_);
  and _78104_ (_27786_, _27785_, _27783_);
  or _78105_ (_27787_, _27786_, _27481_);
  nand _78106_ (_27788_, _27787_, _12782_);
  nor _78107_ (_27789_, _12789_, _05751_);
  not _78108_ (_27790_, _27789_);
  and _78109_ (_27792_, _06119_, _06016_);
  nor _78110_ (_27793_, _27792_, _27790_);
  and _78111_ (_27794_, _27793_, _27788_);
  and _78112_ (_27795_, _27480_, _12789_);
  or _78113_ (_27796_, _27795_, _27794_);
  or _78114_ (_27797_, _27796_, _01340_);
  or _78115_ (_27798_, _01336_, \oc8051_golden_model_1.PC [8]);
  and _78116_ (_27799_, _27798_, _42882_);
  and _78117_ (_43426_, _27799_, _27797_);
  nor _78118_ (_27800_, _06799_, _09200_);
  nor _78119_ (_27802_, _27478_, \oc8051_golden_model_1.PC [9]);
  nor _78120_ (_27803_, _27802_, _11863_);
  nor _78121_ (_27804_, _27803_, _11872_);
  nor _78122_ (_27805_, _27803_, _12523_);
  and _78123_ (_27806_, _12051_, _06130_);
  nor _78124_ (_27807_, _27803_, _11993_);
  and _78125_ (_27808_, _12051_, _06108_);
  nor _78126_ (_27809_, _27803_, _12002_);
  and _78127_ (_27810_, _12051_, _06112_);
  not _78128_ (_27811_, _27803_);
  and _78129_ (_27813_, _27811_, _12006_);
  nor _78130_ (_27814_, _11900_, _08742_);
  and _78131_ (_27815_, _11900_, _06089_);
  and _78132_ (_27816_, _11900_, _06250_);
  nor _78133_ (_27817_, _27803_, _12351_);
  or _78134_ (_27818_, _12187_, _12051_);
  nor _78135_ (_27819_, _12118_, _12114_);
  and _78136_ (_27820_, _27819_, _12055_);
  nor _78137_ (_27821_, _27819_, _12055_);
  nor _78138_ (_27822_, _27821_, _27820_);
  not _78139_ (_27824_, _27822_);
  or _78140_ (_27825_, _27824_, _12189_);
  and _78141_ (_27826_, _27825_, _27818_);
  or _78142_ (_27827_, _27826_, _06954_);
  nor _78143_ (_27828_, _11956_, _11953_);
  and _78144_ (_27829_, _27828_, _11903_);
  nor _78145_ (_27830_, _27828_, _11903_);
  nor _78146_ (_27831_, _27830_, _27829_);
  or _78147_ (_27832_, _27831_, _12197_);
  or _78148_ (_27833_, _12199_, _14461_);
  and _78149_ (_27835_, _27833_, _08384_);
  nand _78150_ (_27836_, _27835_, _27832_);
  and _78151_ (_27837_, _27803_, _06530_);
  or _78152_ (_27838_, _27803_, _27491_);
  and _78153_ (_27839_, _14461_, _06938_);
  nor _78154_ (_27840_, _27839_, _06530_);
  or _78155_ (_27841_, _06938_, \oc8051_golden_model_1.PC [9]);
  or _78156_ (_27842_, _27841_, _07250_);
  nand _78157_ (_27843_, _27842_, _27840_);
  nand _78158_ (_27844_, _27843_, _24785_);
  and _78159_ (_27846_, _27844_, _27838_);
  or _78160_ (_27847_, _27846_, _08384_);
  nor _78161_ (_27848_, _27847_, _27837_);
  nor _78162_ (_27849_, _27848_, _06948_);
  and _78163_ (_27850_, _27849_, _27836_);
  and _78164_ (_27851_, _27803_, _06948_);
  or _78165_ (_27852_, _27851_, _06102_);
  or _78166_ (_27853_, _27852_, _27850_);
  nand _78167_ (_27854_, _27853_, _27827_);
  nand _78168_ (_27855_, _27854_, _12182_);
  nor _78169_ (_27857_, _27803_, _12182_);
  nor _78170_ (_27858_, _27857_, _06043_);
  nand _78171_ (_27859_, _27858_, _27855_);
  and _78172_ (_27860_, _11900_, _06043_);
  nor _78173_ (_27861_, _27860_, _07272_);
  nand _78174_ (_27862_, _27861_, _27859_);
  nand _78175_ (_27863_, _27862_, _06848_);
  and _78176_ (_27864_, _11900_, _06239_);
  nor _78177_ (_27865_, _27864_, _12232_);
  nand _78178_ (_27866_, _27865_, _27863_);
  nor _78179_ (_27868_, _27803_, _12231_);
  nor _78180_ (_27869_, _27868_, _06219_);
  nand _78181_ (_27870_, _27869_, _27866_);
  and _78182_ (_27871_, _11900_, _06219_);
  nor _78183_ (_27872_, _27871_, _12241_);
  nand _78184_ (_27873_, _27872_, _27870_);
  nor _78185_ (_27874_, _27803_, _12239_);
  nor _78186_ (_27875_, _27874_, _06039_);
  nand _78187_ (_27876_, _27875_, _27873_);
  and _78188_ (_27877_, _11900_, _06039_);
  nor _78189_ (_27879_, _27877_, _12243_);
  nand _78190_ (_27880_, _27879_, _27876_);
  nand _78191_ (_27881_, _27880_, _07364_);
  and _78192_ (_27882_, _11900_, _06038_);
  nor _78193_ (_27883_, _27882_, _12256_);
  and _78194_ (_27884_, _27883_, _27881_);
  and _78195_ (_27885_, _12289_, _12051_);
  nor _78196_ (_27886_, _27822_, _12289_);
  or _78197_ (_27887_, _27886_, _27885_);
  nor _78198_ (_27888_, _27887_, _12255_);
  or _78199_ (_27890_, _27888_, _27884_);
  and _78200_ (_27891_, _27890_, _13849_);
  and _78201_ (_27892_, _12172_, _12051_);
  and _78202_ (_27893_, _27824_, _12174_);
  or _78203_ (_27894_, _27893_, _27892_);
  nor _78204_ (_27895_, _27894_, _12258_);
  or _78205_ (_27896_, _27895_, _27891_);
  or _78206_ (_27897_, _27896_, _06121_);
  and _78207_ (_27898_, _12310_, _12051_);
  nor _78208_ (_27899_, _27822_, _12310_);
  nor _78209_ (_27901_, _27899_, _27898_);
  or _78210_ (_27902_, _27901_, _06509_);
  and _78211_ (_27903_, _27902_, _27897_);
  or _78212_ (_27904_, _27903_, _06115_);
  nand _78213_ (_27905_, _12329_, _12051_);
  or _78214_ (_27906_, _27822_, _12329_);
  and _78215_ (_27907_, _27906_, _27905_);
  or _78216_ (_27908_, _27907_, _12298_);
  and _78217_ (_27909_, _27908_, _27904_);
  or _78218_ (_27910_, _27909_, _12012_);
  nand _78219_ (_27912_, _27803_, _12012_);
  and _78220_ (_27913_, _27912_, _27910_);
  nand _78221_ (_27914_, _27913_, _06033_);
  and _78222_ (_27915_, _14461_, _06032_);
  not _78223_ (_27916_, _27915_);
  and _78224_ (_27917_, _12344_, _05686_);
  and _78225_ (_27918_, _27917_, _27916_);
  nand _78226_ (_27919_, _27918_, _27914_);
  nor _78227_ (_27920_, _12344_, _14461_);
  nor _78228_ (_27921_, _27920_, _12355_);
  and _78229_ (_27923_, _27921_, _27919_);
  nor _78230_ (_27924_, _27923_, _27817_);
  or _78231_ (_27925_, _27924_, _06251_);
  nor _78232_ (_27926_, _06250_, _24866_);
  nand _78233_ (_27927_, _14461_, _06251_);
  and _78234_ (_27928_, _27927_, _27926_);
  and _78235_ (_27929_, _27928_, _27925_);
  or _78236_ (_27930_, _27929_, _27816_);
  nand _78237_ (_27931_, _27930_, _12362_);
  nor _78238_ (_27932_, _27811_, _12362_);
  nor _78239_ (_27934_, _27932_, _12367_);
  nand _78240_ (_27935_, _27934_, _27931_);
  nor _78241_ (_27936_, _11900_, _12366_);
  nor _78242_ (_27937_, _27936_, _05676_);
  nand _78243_ (_27938_, _27937_, _27935_);
  nor _78244_ (_27939_, _27811_, _05675_);
  nor _78245_ (_27940_, _27939_, _06026_);
  nand _78246_ (_27941_, _27940_, _27938_);
  not _78247_ (_27942_, _27610_);
  and _78248_ (_27943_, _14461_, _06026_);
  nor _78249_ (_27945_, _27943_, _27942_);
  nand _78250_ (_27946_, _27945_, _27941_);
  and _78251_ (_27947_, _12051_, _06110_);
  nor _78252_ (_27948_, _27947_, _09818_);
  nand _78253_ (_27949_, _27948_, _27946_);
  nor _78254_ (_27950_, _11900_, _09817_);
  nor _78255_ (_27951_, _27950_, _09833_);
  nand _78256_ (_27952_, _27951_, _27949_);
  nor _78257_ (_27953_, _12052_, _05669_);
  nor _78258_ (_27954_, _27953_, _12393_);
  nand _78259_ (_27956_, _27954_, _27952_);
  nor _78260_ (_27957_, _27803_, _12389_);
  nor _78261_ (_27958_, _27957_, _06089_);
  and _78262_ (_27959_, _27958_, _27956_);
  or _78263_ (_27960_, _27959_, _27815_);
  nand _78264_ (_27961_, _27960_, _27628_);
  nor _78265_ (_27962_, _27831_, _12398_);
  nor _78266_ (_27963_, _27962_, _08743_);
  and _78267_ (_27964_, _27963_, _27961_);
  or _78268_ (_27965_, _27964_, _27814_);
  nand _78269_ (_27966_, _27965_, _06020_);
  and _78270_ (_27967_, _12052_, _06019_);
  nor _78271_ (_27968_, _27967_, _10661_);
  nand _78272_ (_27969_, _27968_, _27966_);
  and _78273_ (_27970_, _11900_, _10661_);
  nor _78274_ (_27971_, _27970_, _12412_);
  nand _78275_ (_27972_, _27971_, _27969_);
  nor _78276_ (_27973_, _12440_, \oc8051_golden_model_1.DPH [1]);
  nor _78277_ (_27974_, _27973_, _12441_);
  nor _78278_ (_27975_, _27974_, _12413_);
  nor _78279_ (_27978_, _27975_, _06088_);
  nand _78280_ (_27979_, _27978_, _27972_);
  and _78281_ (_27980_, _11900_, _06088_);
  nor _78282_ (_27981_, _27980_, _05724_);
  nand _78283_ (_27982_, _27981_, _27979_);
  nand _78284_ (_27983_, _27982_, _12454_);
  and _78285_ (_27984_, _11900_, _11071_);
  nor _78286_ (_27985_, _27831_, _11071_);
  or _78287_ (_27986_, _27985_, _27984_);
  and _78288_ (_27987_, _27986_, _12453_);
  nor _78289_ (_27989_, _27987_, _12006_);
  and _78290_ (_27990_, _27989_, _27983_);
  or _78291_ (_27991_, _27990_, _27813_);
  nand _78292_ (_27992_, _27991_, _12466_);
  nor _78293_ (_27993_, _12466_, _11900_);
  nor _78294_ (_27994_, _27993_, _06112_);
  and _78295_ (_27995_, _27994_, _27992_);
  or _78296_ (_27996_, _27995_, _27810_);
  nand _78297_ (_27997_, _27996_, _08756_);
  and _78298_ (_27998_, _11900_, _06284_);
  nor _78299_ (_28000_, _27998_, _05727_);
  nand _78300_ (_28001_, _28000_, _27997_);
  nand _78301_ (_28002_, _28001_, _12477_);
  and _78302_ (_28003_, _11900_, _12459_);
  nor _78303_ (_28004_, _27831_, _12459_);
  or _78304_ (_28005_, _28004_, _28003_);
  and _78305_ (_28006_, _28005_, _12476_);
  nor _78306_ (_28007_, _28006_, _12481_);
  and _78307_ (_28008_, _28007_, _28002_);
  or _78308_ (_28009_, _28008_, _27809_);
  nand _78309_ (_28011_, _28009_, _10742_);
  nor _78310_ (_28012_, _11900_, _10742_);
  nor _78311_ (_28013_, _28012_, _06108_);
  and _78312_ (_28014_, _28013_, _28011_);
  or _78313_ (_28015_, _28014_, _27808_);
  nand _78314_ (_28016_, _28015_, _06278_);
  and _78315_ (_28017_, _11900_, _06277_);
  nor _78316_ (_28018_, _28017_, _05736_);
  nand _78317_ (_28019_, _28018_, _28016_);
  nand _78318_ (_28020_, _28019_, _12498_);
  and _78319_ (_28022_, _11900_, \oc8051_golden_model_1.PSW [7]);
  nor _78320_ (_28023_, _27831_, \oc8051_golden_model_1.PSW [7]);
  or _78321_ (_28024_, _28023_, _28022_);
  and _78322_ (_28025_, _28024_, _12497_);
  nor _78323_ (_28026_, _28025_, _12502_);
  and _78324_ (_28027_, _28026_, _28020_);
  or _78325_ (_28028_, _28027_, _27807_);
  nand _78326_ (_28029_, _28028_, _11986_);
  nor _78327_ (_28030_, _11900_, _11986_);
  nor _78328_ (_28031_, _28030_, _06130_);
  and _78329_ (_28033_, _28031_, _28029_);
  or _78330_ (_28034_, _28033_, _27806_);
  nand _78331_ (_28035_, _28034_, _08782_);
  and _78332_ (_28036_, _11900_, _06292_);
  nor _78333_ (_28037_, _28036_, _05740_);
  nand _78334_ (_28038_, _28037_, _28035_);
  nand _78335_ (_28039_, _28038_, _12518_);
  nand _78336_ (_28040_, _27831_, \oc8051_golden_model_1.PSW [7]);
  or _78337_ (_28041_, _11900_, \oc8051_golden_model_1.PSW [7]);
  and _78338_ (_28042_, _28041_, _11982_);
  and _78339_ (_28044_, _28042_, _28040_);
  nor _78340_ (_28045_, _28044_, _12525_);
  and _78341_ (_28046_, _28045_, _28039_);
  or _78342_ (_28047_, _28046_, _27805_);
  nand _78343_ (_28048_, _28047_, _10825_);
  nor _78344_ (_28049_, _11900_, _10825_);
  nor _78345_ (_28050_, _28049_, _10854_);
  nand _78346_ (_28051_, _28050_, _28048_);
  and _78347_ (_28052_, _27803_, _10854_);
  nor _78348_ (_28053_, _28052_, _06298_);
  nand _78349_ (_28055_, _28053_, _28051_);
  nor _78350_ (_28056_, _06129_, _05732_);
  not _78351_ (_28057_, _28056_);
  and _78352_ (_28058_, _07132_, _06298_);
  nor _78353_ (_28059_, _28058_, _28057_);
  nand _78354_ (_28060_, _28059_, _28055_);
  nor _78355_ (_28061_, _12051_, _12722_);
  and _78356_ (_28062_, _27822_, _12722_);
  or _78357_ (_28063_, _28062_, _06306_);
  nor _78358_ (_28064_, _28063_, _28061_);
  nor _78359_ (_28066_, _28064_, _12541_);
  and _78360_ (_28067_, _28066_, _28060_);
  or _78361_ (_28068_, _28067_, _27804_);
  nand _78362_ (_28069_, _28068_, _10975_);
  nor _78363_ (_28070_, _11900_, _10975_);
  nor _78364_ (_28071_, _28070_, _11015_);
  nand _78365_ (_28072_, _28071_, _28069_);
  and _78366_ (_28073_, _27803_, _11015_);
  nor _78367_ (_28074_, _28073_, _06049_);
  nand _78368_ (_28075_, _28074_, _28072_);
  nor _78369_ (_28077_, _06126_, _05747_);
  not _78370_ (_28078_, _28077_);
  and _78371_ (_28079_, _07132_, _06049_);
  nor _78372_ (_28080_, _28079_, _28078_);
  nand _78373_ (_28081_, _28080_, _28075_);
  and _78374_ (_28082_, _12052_, _12722_);
  nor _78375_ (_28083_, _27824_, _12722_);
  nor _78376_ (_28084_, _28083_, _28082_);
  and _78377_ (_28085_, _28084_, _06126_);
  nor _78378_ (_28086_, _28085_, _12750_);
  nand _78379_ (_28088_, _28086_, _28081_);
  nor _78380_ (_28089_, _27803_, _12749_);
  nor _78381_ (_28090_, _28089_, _06316_);
  nand _78382_ (_28091_, _28090_, _28088_);
  and _78383_ (_28092_, _11900_, _06316_);
  nor _78384_ (_28093_, _28092_, _25353_);
  nand _78385_ (_28094_, _28093_, _28091_);
  nor _78386_ (_28095_, _27803_, _12756_);
  nor _78387_ (_28096_, _28095_, _06127_);
  and _78388_ (_28097_, _28096_, _28094_);
  or _78389_ (_28099_, _28097_, _27800_);
  nand _78390_ (_28100_, _28099_, _27775_);
  and _78391_ (_28101_, _28084_, _05652_);
  nor _78392_ (_28102_, _28101_, _12772_);
  nand _78393_ (_28103_, _28102_, _28100_);
  nor _78394_ (_28104_, _27803_, _12771_);
  nor _78395_ (_28105_, _28104_, _06047_);
  nand _78396_ (_28106_, _28105_, _28103_);
  and _78397_ (_28107_, _11900_, _06047_);
  nor _78398_ (_28108_, _28107_, _26405_);
  nand _78399_ (_28110_, _28108_, _28106_);
  nor _78400_ (_28111_, _27803_, _12779_);
  nor _78401_ (_28112_, _28111_, _06119_);
  and _78402_ (_28113_, _28112_, _28110_);
  nor _78403_ (_28114_, _06799_, _12782_);
  or _78404_ (_28115_, _28114_, _28113_);
  and _78405_ (_28116_, _28115_, _27789_);
  and _78406_ (_28117_, _27803_, _12789_);
  or _78407_ (_28118_, _28117_, _28116_);
  or _78408_ (_28119_, _28118_, _01340_);
  or _78409_ (_28121_, _01336_, \oc8051_golden_model_1.PC [9]);
  and _78410_ (_28122_, _28121_, _42882_);
  and _78411_ (_43427_, _28122_, _28119_);
  nor _78412_ (_28123_, _11863_, \oc8051_golden_model_1.PC [10]);
  nor _78413_ (_28124_, _28123_, _11864_);
  and _78414_ (_28125_, _28124_, _12393_);
  or _78415_ (_28126_, _12344_, _11887_);
  or _78416_ (_28127_, _28124_, _12231_);
  nor _78417_ (_28128_, _12122_, _12119_);
  not _78418_ (_28129_, _28128_);
  and _78419_ (_28131_, _28129_, _12047_);
  nor _78420_ (_28132_, _28129_, _12047_);
  nor _78421_ (_28133_, _28132_, _28131_);
  and _78422_ (_28134_, _28133_, _12187_);
  and _78423_ (_28135_, _12189_, _12043_);
  or _78424_ (_28136_, _28135_, _06954_);
  or _78425_ (_28137_, _28136_, _28134_);
  nor _78426_ (_28138_, _11960_, _11957_);
  not _78427_ (_28139_, _28138_);
  and _78428_ (_28140_, _28139_, _11896_);
  nor _78429_ (_28142_, _28139_, _11896_);
  nor _78430_ (_28143_, _28142_, _28140_);
  or _78431_ (_28144_, _28143_, _12197_);
  or _78432_ (_28145_, _12199_, _11887_);
  and _78433_ (_28146_, _28145_, _28144_);
  or _78434_ (_28147_, _28146_, _08383_);
  and _78435_ (_28148_, _11887_, _06938_);
  nand _78436_ (_28149_, _06939_, \oc8051_golden_model_1.PC [10]);
  nor _78437_ (_28150_, _28149_, _07250_);
  or _78438_ (_28151_, _28150_, _28148_);
  and _78439_ (_28153_, _28151_, _25758_);
  or _78440_ (_28154_, _28153_, _06943_);
  and _78441_ (_28155_, _28154_, _12205_);
  not _78442_ (_28156_, _12215_);
  and _78443_ (_28157_, _28124_, _28156_);
  or _78444_ (_28158_, _28157_, _08384_);
  or _78445_ (_28159_, _28158_, _28155_);
  and _78446_ (_28160_, _28159_, _06949_);
  and _78447_ (_28161_, _28160_, _28147_);
  and _78448_ (_28162_, _28124_, _06948_);
  or _78449_ (_28164_, _28162_, _06102_);
  or _78450_ (_28165_, _28164_, _28161_);
  and _78451_ (_28166_, _28165_, _28137_);
  or _78452_ (_28167_, _28166_, _24805_);
  or _78453_ (_28168_, _28124_, _12182_);
  and _78454_ (_28169_, _28168_, _06044_);
  and _78455_ (_28170_, _28169_, _28167_);
  or _78456_ (_28171_, _28170_, _07272_);
  and _78457_ (_28172_, _28171_, _06848_);
  nor _78458_ (_28173_, _14664_, _06244_);
  or _78459_ (_28175_, _28173_, _12232_);
  or _78460_ (_28176_, _28175_, _28172_);
  and _78461_ (_28177_, _28176_, _28127_);
  or _78462_ (_28178_, _28177_, _06219_);
  nand _78463_ (_28179_, _14664_, _06219_);
  and _78464_ (_28180_, _28179_, _12239_);
  and _78465_ (_28181_, _28180_, _28178_);
  and _78466_ (_28182_, _28124_, _12241_);
  or _78467_ (_28183_, _28182_, _28181_);
  and _78468_ (_28184_, _28183_, _06040_);
  and _78469_ (_28186_, _11887_, _06039_);
  or _78470_ (_28187_, _28186_, _12243_);
  or _78471_ (_28188_, _28187_, _28184_);
  and _78472_ (_28189_, _28188_, _07364_);
  nand _78473_ (_28190_, _11887_, _06038_);
  nand _78474_ (_28191_, _28190_, _12255_);
  or _78475_ (_28192_, _28191_, _28189_);
  and _78476_ (_28193_, _28133_, _13828_);
  and _78477_ (_28194_, _12289_, _12043_);
  or _78478_ (_28195_, _28194_, _12255_);
  or _78479_ (_28197_, _28195_, _28193_);
  and _78480_ (_28198_, _28197_, _28192_);
  or _78481_ (_28199_, _28198_, _06104_);
  and _78482_ (_28200_, _28133_, _12174_);
  and _78483_ (_28201_, _12172_, _12043_);
  or _78484_ (_28202_, _28201_, _12258_);
  or _78485_ (_28203_, _28202_, _28200_);
  and _78486_ (_28204_, _28203_, _28199_);
  or _78487_ (_28205_, _28204_, _06121_);
  and _78488_ (_28206_, _28133_, _12312_);
  and _78489_ (_28208_, _12310_, _12043_);
  or _78490_ (_28209_, _28208_, _06509_);
  or _78491_ (_28210_, _28209_, _28206_);
  and _78492_ (_28211_, _28210_, _12298_);
  and _78493_ (_28212_, _28211_, _28205_);
  or _78494_ (_28213_, _28133_, _12329_);
  nand _78495_ (_28214_, _12329_, _12044_);
  and _78496_ (_28215_, _28214_, _06115_);
  and _78497_ (_28216_, _28215_, _28213_);
  or _78498_ (_28217_, _28216_, _12012_);
  or _78499_ (_28219_, _28217_, _28212_);
  or _78500_ (_28220_, _28124_, _12013_);
  and _78501_ (_28221_, _28220_, _06033_);
  and _78502_ (_28222_, _28221_, _28219_);
  and _78503_ (_28223_, _11887_, _06032_);
  nor _78504_ (_28224_, _28223_, _28222_);
  nand _78505_ (_28225_, _28224_, _27917_);
  and _78506_ (_28226_, _28225_, _28126_);
  or _78507_ (_28227_, _28226_, _12355_);
  or _78508_ (_28228_, _28124_, _12351_);
  and _78509_ (_28230_, _28228_, _13765_);
  and _78510_ (_28231_, _28230_, _28227_);
  or _78511_ (_28232_, _28231_, _24866_);
  and _78512_ (_28233_, _28232_, _13764_);
  nor _78513_ (_28234_, _14664_, _06252_);
  or _78514_ (_28235_, _28234_, _12368_);
  or _78515_ (_28236_, _28235_, _28233_);
  or _78516_ (_28237_, _28124_, _12362_);
  and _78517_ (_28238_, _28237_, _12366_);
  and _78518_ (_28239_, _28238_, _28236_);
  nor _78519_ (_28241_, _14664_, _12366_);
  or _78520_ (_28242_, _28241_, _05676_);
  or _78521_ (_28243_, _28242_, _28239_);
  or _78522_ (_28244_, _28124_, _05675_);
  and _78523_ (_28245_, _28244_, _06027_);
  and _78524_ (_28246_, _28245_, _28243_);
  nand _78525_ (_28247_, _11887_, _06026_);
  nand _78526_ (_28248_, _28247_, _27610_);
  or _78527_ (_28249_, _28248_, _28246_);
  nand _78528_ (_28250_, _12044_, _06110_);
  and _78529_ (_28252_, _28250_, _09817_);
  and _78530_ (_28253_, _28252_, _28249_);
  nor _78531_ (_28254_, _14664_, _09817_);
  or _78532_ (_28255_, _28254_, _09833_);
  or _78533_ (_28256_, _28255_, _28253_);
  or _78534_ (_28257_, _12043_, _05669_);
  and _78535_ (_28258_, _28257_, _12389_);
  and _78536_ (_28259_, _28258_, _28256_);
  or _78537_ (_28260_, _28259_, _28125_);
  and _78538_ (_28261_, _28260_, _25023_);
  nand _78539_ (_28263_, _11887_, _06089_);
  nand _78540_ (_28264_, _28263_, _27628_);
  or _78541_ (_28265_, _28264_, _28261_);
  or _78542_ (_28266_, _28143_, _12398_);
  and _78543_ (_28267_, _28266_, _08742_);
  and _78544_ (_28268_, _28267_, _28265_);
  nor _78545_ (_28269_, _14664_, _08742_);
  or _78546_ (_28270_, _28269_, _06019_);
  or _78547_ (_28271_, _28270_, _28268_);
  nand _78548_ (_28272_, _12044_, _06019_);
  and _78549_ (_28273_, _28272_, _10662_);
  and _78550_ (_28274_, _28273_, _28271_);
  and _78551_ (_28275_, _11887_, _10661_);
  or _78552_ (_28276_, _28275_, _12412_);
  or _78553_ (_28277_, _28276_, _28274_);
  nor _78554_ (_28278_, _12441_, \oc8051_golden_model_1.DPH [2]);
  nor _78555_ (_28279_, _28278_, _12442_);
  or _78556_ (_28280_, _28279_, _12413_);
  and _78557_ (_28281_, _28280_, _06636_);
  and _78558_ (_28282_, _28281_, _28277_);
  and _78559_ (_28285_, _11887_, _06088_);
  or _78560_ (_28286_, _28285_, _28282_);
  nand _78561_ (_28287_, _07187_, _05569_);
  and _78562_ (_28288_, _28287_, _28286_);
  or _78563_ (_28289_, _28143_, _11071_);
  or _78564_ (_28290_, _11887_, _12459_);
  and _78565_ (_28291_, _28290_, _12453_);
  and _78566_ (_28292_, _28291_, _28289_);
  or _78567_ (_28293_, _28292_, _12006_);
  or _78568_ (_28294_, _28293_, _28288_);
  or _78569_ (_28296_, _28124_, _12007_);
  and _78570_ (_28297_, _28296_, _12466_);
  and _78571_ (_28298_, _28297_, _28294_);
  nor _78572_ (_28299_, _12466_, _14664_);
  or _78573_ (_28300_, _28299_, _06112_);
  or _78574_ (_28301_, _28300_, _28298_);
  nand _78575_ (_28302_, _12044_, _06112_);
  and _78576_ (_28303_, _28302_, _28301_);
  or _78577_ (_28304_, _28303_, _06284_);
  nand _78578_ (_28305_, _14664_, _06284_);
  nor _78579_ (_28307_, _12476_, _05727_);
  and _78580_ (_28308_, _28307_, _28305_);
  and _78581_ (_28309_, _28308_, _28304_);
  or _78582_ (_28310_, _28143_, _12459_);
  or _78583_ (_28311_, _11887_, _11071_);
  and _78584_ (_28312_, _28311_, _12476_);
  and _78585_ (_28313_, _28312_, _28310_);
  or _78586_ (_28314_, _28313_, _12481_);
  or _78587_ (_28315_, _28314_, _28309_);
  or _78588_ (_28316_, _28124_, _12002_);
  and _78589_ (_28318_, _28316_, _10742_);
  and _78590_ (_28319_, _28318_, _28315_);
  nor _78591_ (_28320_, _14664_, _10742_);
  or _78592_ (_28321_, _28320_, _06108_);
  or _78593_ (_28322_, _28321_, _28319_);
  nand _78594_ (_28323_, _12044_, _06108_);
  and _78595_ (_28324_, _28323_, _28322_);
  or _78596_ (_28325_, _28324_, _06277_);
  nand _78597_ (_28326_, _14664_, _06277_);
  and _78598_ (_28327_, _28326_, _27690_);
  and _78599_ (_28329_, _28327_, _28325_);
  or _78600_ (_28330_, _28143_, \oc8051_golden_model_1.PSW [7]);
  or _78601_ (_28331_, _11887_, _10606_);
  and _78602_ (_28332_, _28331_, _12497_);
  and _78603_ (_28333_, _28332_, _28330_);
  or _78604_ (_28334_, _28333_, _12502_);
  or _78605_ (_28335_, _28334_, _28329_);
  or _78606_ (_28336_, _28124_, _11993_);
  and _78607_ (_28337_, _28336_, _11986_);
  and _78608_ (_28338_, _28337_, _28335_);
  nor _78609_ (_28340_, _14664_, _11986_);
  or _78610_ (_28341_, _28340_, _06130_);
  or _78611_ (_28342_, _28341_, _28338_);
  nand _78612_ (_28343_, _12044_, _06130_);
  and _78613_ (_28344_, _28343_, _28342_);
  or _78614_ (_28345_, _28344_, _06292_);
  nand _78615_ (_28346_, _14664_, _06292_);
  and _78616_ (_28347_, _28346_, _27484_);
  and _78617_ (_28348_, _28347_, _28345_);
  or _78618_ (_28349_, _28143_, _10606_);
  or _78619_ (_28351_, _11887_, \oc8051_golden_model_1.PSW [7]);
  and _78620_ (_28352_, _28351_, _11982_);
  and _78621_ (_28353_, _28352_, _28349_);
  or _78622_ (_28354_, _28353_, _12525_);
  or _78623_ (_28355_, _28354_, _28348_);
  or _78624_ (_28356_, _28124_, _12523_);
  and _78625_ (_28357_, _28356_, _10825_);
  and _78626_ (_28358_, _28357_, _28355_);
  nor _78627_ (_28359_, _14664_, _10825_);
  or _78628_ (_28360_, _28359_, _10854_);
  or _78629_ (_28362_, _28360_, _28358_);
  or _78630_ (_28363_, _28124_, _10855_);
  and _78631_ (_28364_, _28363_, _28362_);
  or _78632_ (_28365_, _28364_, _06298_);
  nand _78633_ (_28366_, _07530_, _06298_);
  and _78634_ (_28367_, _28366_, _28056_);
  and _78635_ (_28368_, _28367_, _28365_);
  or _78636_ (_28369_, _28133_, _12723_);
  or _78637_ (_28370_, _12043_, _12722_);
  and _78638_ (_28371_, _28370_, _06129_);
  and _78639_ (_28373_, _28371_, _28369_);
  or _78640_ (_28374_, _28373_, _12541_);
  or _78641_ (_28375_, _28374_, _28368_);
  or _78642_ (_28376_, _28124_, _11872_);
  and _78643_ (_28377_, _28376_, _10975_);
  and _78644_ (_28378_, _28377_, _28375_);
  nor _78645_ (_28379_, _14664_, _10975_);
  or _78646_ (_28380_, _28379_, _11015_);
  or _78647_ (_28381_, _28380_, _28378_);
  or _78648_ (_28382_, _28124_, _11016_);
  and _78649_ (_28384_, _28382_, _28381_);
  or _78650_ (_28385_, _28384_, _06049_);
  nand _78651_ (_28386_, _07530_, _06049_);
  and _78652_ (_28387_, _28386_, _28077_);
  and _78653_ (_28388_, _28387_, _28385_);
  or _78654_ (_28389_, _28133_, _12722_);
  nand _78655_ (_28390_, _12044_, _12722_);
  and _78656_ (_28391_, _28390_, _28389_);
  and _78657_ (_28392_, _28391_, _06126_);
  or _78658_ (_28393_, _28392_, _12750_);
  or _78659_ (_28395_, _28393_, _28388_);
  or _78660_ (_28396_, _28124_, _12749_);
  and _78661_ (_28397_, _28396_, _28395_);
  or _78662_ (_28398_, _28397_, _06316_);
  nand _78663_ (_28399_, _14664_, _06316_);
  and _78664_ (_28400_, _28399_, _12756_);
  and _78665_ (_28401_, _28400_, _28398_);
  and _78666_ (_28402_, _28124_, _25353_);
  or _78667_ (_28403_, _28402_, _06127_);
  or _78668_ (_28404_, _28403_, _28401_);
  nand _78669_ (_28406_, _06403_, _06127_);
  and _78670_ (_28407_, _28406_, _27775_);
  and _78671_ (_28408_, _28407_, _28404_);
  and _78672_ (_28409_, _28391_, _05652_);
  or _78673_ (_28410_, _28409_, _12772_);
  or _78674_ (_28411_, _28410_, _28408_);
  or _78675_ (_28412_, _28124_, _12771_);
  and _78676_ (_28413_, _28412_, _28411_);
  or _78677_ (_28414_, _28413_, _06047_);
  nand _78678_ (_28415_, _14664_, _06047_);
  and _78679_ (_28417_, _28415_, _12779_);
  and _78680_ (_28418_, _28417_, _28414_);
  and _78681_ (_28419_, _28124_, _26405_);
  or _78682_ (_28420_, _28419_, _06119_);
  or _78683_ (_28421_, _28420_, _28418_);
  nand _78684_ (_28422_, _06403_, _06119_);
  and _78685_ (_28423_, _28422_, _27789_);
  and _78686_ (_28424_, _28423_, _28421_);
  and _78687_ (_28425_, _28124_, _12789_);
  or _78688_ (_28426_, _28425_, _28424_);
  or _78689_ (_28428_, _28426_, _01340_);
  or _78690_ (_28429_, _01336_, \oc8051_golden_model_1.PC [10]);
  and _78691_ (_28430_, _28429_, _42882_);
  and _78692_ (_43428_, _28430_, _28428_);
  nor _78693_ (_28431_, _11864_, \oc8051_golden_model_1.PC [11]);
  nor _78694_ (_28432_, _28431_, _11865_);
  or _78695_ (_28433_, _28432_, _11872_);
  or _78696_ (_28434_, _28432_, _12523_);
  or _78697_ (_28435_, _28432_, _11993_);
  or _78698_ (_28436_, _28432_, _12007_);
  nor _78699_ (_28438_, _12037_, _05669_);
  nor _78700_ (_28439_, _28131_, _12045_);
  and _78701_ (_28440_, _28439_, _12040_);
  nor _78702_ (_28441_, _28439_, _12040_);
  or _78703_ (_28442_, _28441_, _28440_);
  or _78704_ (_28443_, _28442_, _12172_);
  or _78705_ (_28444_, _12174_, _12036_);
  and _78706_ (_28445_, _28444_, _06104_);
  and _78707_ (_28446_, _28445_, _28443_);
  and _78708_ (_28447_, _11891_, _06219_);
  or _78709_ (_28449_, _12179_, _11891_);
  or _78710_ (_28450_, _12187_, _12036_);
  or _78711_ (_28451_, _28442_, _12189_);
  and _78712_ (_28452_, _28451_, _06102_);
  and _78713_ (_28453_, _28452_, _28450_);
  nor _78714_ (_28454_, _28140_, _11888_);
  nor _78715_ (_28455_, _28454_, _11894_);
  and _78716_ (_28456_, _28454_, _11894_);
  or _78717_ (_28457_, _28456_, _28455_);
  and _78718_ (_28458_, _28457_, _12199_);
  and _78719_ (_28460_, _12197_, _11891_);
  or _78720_ (_28461_, _28460_, _08383_);
  or _78721_ (_28462_, _28461_, _28458_);
  or _78722_ (_28463_, _28432_, _12215_);
  or _78723_ (_28464_, _11891_, _07233_);
  or _78724_ (_28465_, _11891_, _06939_);
  or _78725_ (_28466_, _06938_, \oc8051_golden_model_1.PC [11]);
  or _78726_ (_28467_, _28466_, _07250_);
  and _78727_ (_28468_, _28467_, _28465_);
  nand _78728_ (_28469_, _24785_, _25758_);
  or _78729_ (_28471_, _28469_, _28468_);
  and _78730_ (_28472_, _28471_, _28464_);
  and _78731_ (_28473_, _28472_, _28463_);
  or _78732_ (_28474_, _28473_, _08384_);
  and _78733_ (_28475_, _28474_, _12219_);
  and _78734_ (_28476_, _28475_, _28462_);
  or _78735_ (_28477_, _28476_, _28453_);
  and _78736_ (_28478_, _28477_, _12182_);
  and _78737_ (_28479_, _28432_, _12226_);
  or _78738_ (_28480_, _28479_, _12224_);
  or _78739_ (_28482_, _28480_, _28478_);
  and _78740_ (_28483_, _28482_, _28449_);
  or _78741_ (_28484_, _28483_, _12232_);
  or _78742_ (_28485_, _28432_, _12231_);
  and _78743_ (_28486_, _28485_, _06220_);
  and _78744_ (_28487_, _28486_, _28484_);
  or _78745_ (_28488_, _28487_, _28447_);
  and _78746_ (_28489_, _28488_, _12239_);
  and _78747_ (_28490_, _28432_, _12241_);
  or _78748_ (_28491_, _28490_, _12246_);
  or _78749_ (_28493_, _28491_, _28489_);
  or _78750_ (_28494_, _12245_, _11891_);
  and _78751_ (_28495_, _28494_, _28493_);
  or _78752_ (_28496_, _28495_, _12256_);
  or _78753_ (_28497_, _28442_, _12289_);
  nand _78754_ (_28498_, _12289_, _12037_);
  and _78755_ (_28499_, _28498_, _28497_);
  or _78756_ (_28500_, _28499_, _12255_);
  and _78757_ (_28501_, _28500_, _12258_);
  and _78758_ (_28502_, _28501_, _28496_);
  or _78759_ (_28504_, _28502_, _06121_);
  or _78760_ (_28505_, _28504_, _28446_);
  and _78761_ (_28506_, _12310_, _12036_);
  and _78762_ (_28507_, _28442_, _12312_);
  or _78763_ (_28508_, _28507_, _06509_);
  or _78764_ (_28509_, _28508_, _28506_);
  and _78765_ (_28510_, _28509_, _12298_);
  and _78766_ (_28511_, _28510_, _28505_);
  or _78767_ (_28512_, _28442_, _12329_);
  nand _78768_ (_28513_, _12329_, _12037_);
  and _78769_ (_28515_, _28513_, _06115_);
  and _78770_ (_28516_, _28515_, _28512_);
  or _78771_ (_28517_, _28516_, _28511_);
  and _78772_ (_28518_, _28517_, _12013_);
  nand _78773_ (_28519_, _28432_, _12012_);
  nand _78774_ (_28520_, _28519_, _12345_);
  or _78775_ (_28521_, _28520_, _28518_);
  or _78776_ (_28522_, _12345_, _11891_);
  and _78777_ (_28523_, _28522_, _12351_);
  and _78778_ (_28524_, _28523_, _28521_);
  and _78779_ (_28526_, _28432_, _12355_);
  or _78780_ (_28527_, _28526_, _12358_);
  or _78781_ (_28528_, _28527_, _28524_);
  or _78782_ (_28529_, _12357_, _11891_);
  and _78783_ (_28530_, _28529_, _12362_);
  and _78784_ (_28531_, _28530_, _28528_);
  and _78785_ (_28532_, _28432_, _12368_);
  or _78786_ (_28533_, _28532_, _12367_);
  or _78787_ (_28534_, _28533_, _28531_);
  or _78788_ (_28535_, _11891_, _12366_);
  and _78789_ (_28537_, _28535_, _05675_);
  and _78790_ (_28538_, _28537_, _28534_);
  nand _78791_ (_28539_, _28432_, _05676_);
  nand _78792_ (_28540_, _28539_, _12376_);
  or _78793_ (_28541_, _28540_, _28538_);
  or _78794_ (_28542_, _12376_, _11891_);
  and _78795_ (_28543_, _28542_, _06111_);
  and _78796_ (_28544_, _28543_, _28541_);
  nand _78797_ (_28545_, _12036_, _06110_);
  nand _78798_ (_28546_, _28545_, _09817_);
  or _78799_ (_28548_, _28546_, _28544_);
  or _78800_ (_28549_, _11891_, _09817_);
  and _78801_ (_28550_, _28549_, _05669_);
  and _78802_ (_28551_, _28550_, _28548_);
  or _78803_ (_28552_, _28551_, _28438_);
  and _78804_ (_28553_, _28552_, _12389_);
  and _78805_ (_28554_, _28432_, _12393_);
  or _78806_ (_28555_, _28554_, _12392_);
  or _78807_ (_28556_, _28555_, _28553_);
  or _78808_ (_28557_, _12391_, _11891_);
  and _78809_ (_28559_, _28557_, _12398_);
  and _78810_ (_28560_, _28559_, _28556_);
  and _78811_ (_28561_, _28457_, _12397_);
  or _78812_ (_28562_, _28561_, _08743_);
  or _78813_ (_28563_, _28562_, _28560_);
  or _78814_ (_28564_, _11891_, _08742_);
  and _78815_ (_28565_, _28564_, _06020_);
  and _78816_ (_28566_, _28565_, _28563_);
  and _78817_ (_28567_, _12036_, _06019_);
  or _78818_ (_28568_, _28567_, _10661_);
  or _78819_ (_28570_, _28568_, _28566_);
  or _78820_ (_28571_, _11891_, _10662_);
  and _78821_ (_28572_, _28571_, _12413_);
  and _78822_ (_28573_, _28572_, _28570_);
  or _78823_ (_28574_, _12442_, \oc8051_golden_model_1.DPH [3]);
  nor _78824_ (_28575_, _12443_, _12413_);
  and _78825_ (_28576_, _28575_, _28574_);
  or _78826_ (_28577_, _28576_, _12416_);
  or _78827_ (_28578_, _28577_, _28573_);
  or _78828_ (_28579_, _12415_, _11891_);
  and _78829_ (_28581_, _28579_, _12454_);
  and _78830_ (_28582_, _28581_, _28578_);
  or _78831_ (_28583_, _28457_, _11071_);
  or _78832_ (_28584_, _11891_, _12459_);
  and _78833_ (_28585_, _28584_, _12453_);
  and _78834_ (_28586_, _28585_, _28583_);
  or _78835_ (_28587_, _28586_, _12006_);
  or _78836_ (_28588_, _28587_, _28582_);
  and _78837_ (_28589_, _28588_, _28436_);
  or _78838_ (_28590_, _28589_, _12467_);
  or _78839_ (_28592_, _12466_, _11891_);
  and _78840_ (_28593_, _28592_, _08751_);
  and _78841_ (_28594_, _28593_, _28590_);
  nand _78842_ (_28595_, _12036_, _06112_);
  nand _78843_ (_28596_, _28595_, _12473_);
  or _78844_ (_28597_, _28596_, _28594_);
  or _78845_ (_28598_, _12473_, _11891_);
  and _78846_ (_28599_, _28598_, _12477_);
  and _78847_ (_28600_, _28599_, _28597_);
  or _78848_ (_28601_, _28457_, _12459_);
  or _78849_ (_28603_, _11891_, _11071_);
  and _78850_ (_28604_, _28603_, _12476_);
  and _78851_ (_28605_, _28604_, _28601_);
  or _78852_ (_28606_, _28605_, _28600_);
  and _78853_ (_28607_, _28606_, _12002_);
  and _78854_ (_28608_, _28432_, _12481_);
  or _78855_ (_28609_, _28608_, _10743_);
  or _78856_ (_28610_, _28609_, _28607_);
  or _78857_ (_28611_, _11891_, _10742_);
  and _78858_ (_28612_, _28611_, _07032_);
  and _78859_ (_28614_, _28612_, _28610_);
  nand _78860_ (_28615_, _12036_, _06108_);
  nand _78861_ (_28616_, _28615_, _12494_);
  or _78862_ (_28617_, _28616_, _28614_);
  or _78863_ (_28618_, _12494_, _11891_);
  and _78864_ (_28619_, _28618_, _12498_);
  and _78865_ (_28620_, _28619_, _28617_);
  or _78866_ (_28621_, _28457_, \oc8051_golden_model_1.PSW [7]);
  or _78867_ (_28622_, _11891_, _10606_);
  and _78868_ (_28623_, _28622_, _12497_);
  and _78869_ (_28624_, _28623_, _28621_);
  or _78870_ (_28625_, _28624_, _12502_);
  or _78871_ (_28626_, _28625_, _28620_);
  and _78872_ (_28627_, _28626_, _28435_);
  or _78873_ (_28628_, _28627_, _11987_);
  or _78874_ (_28629_, _11891_, _11986_);
  and _78875_ (_28630_, _28629_, _08777_);
  and _78876_ (_28631_, _28630_, _28628_);
  nand _78877_ (_28632_, _12036_, _06130_);
  nand _78878_ (_28633_, _28632_, _12515_);
  or _78879_ (_28636_, _28633_, _28631_);
  or _78880_ (_28637_, _12515_, _11891_);
  and _78881_ (_28638_, _28637_, _12518_);
  and _78882_ (_28639_, _28638_, _28636_);
  or _78883_ (_28640_, _28457_, _10606_);
  or _78884_ (_28641_, _11891_, \oc8051_golden_model_1.PSW [7]);
  and _78885_ (_28642_, _28641_, _11982_);
  and _78886_ (_28643_, _28642_, _28640_);
  or _78887_ (_28644_, _28643_, _12525_);
  or _78888_ (_28645_, _28644_, _28639_);
  and _78889_ (_28647_, _28645_, _28434_);
  or _78890_ (_28648_, _28647_, _10826_);
  or _78891_ (_28649_, _11891_, _10825_);
  and _78892_ (_28650_, _28649_, _10855_);
  and _78893_ (_28651_, _28650_, _28648_);
  and _78894_ (_28652_, _28432_, _10854_);
  or _78895_ (_28653_, _28652_, _06298_);
  or _78896_ (_28654_, _28653_, _28651_);
  nand _78897_ (_28655_, _07353_, _06298_);
  and _78898_ (_28656_, _28655_, _28654_);
  or _78899_ (_28658_, _28656_, _05732_);
  or _78900_ (_28659_, _11891_, _05734_);
  and _78901_ (_28660_, _28659_, _06306_);
  and _78902_ (_28661_, _28660_, _28658_);
  or _78903_ (_28662_, _28442_, _12723_);
  or _78904_ (_28663_, _12036_, _12722_);
  and _78905_ (_28664_, _28663_, _06129_);
  and _78906_ (_28665_, _28664_, _28662_);
  or _78907_ (_28666_, _28665_, _12541_);
  or _78908_ (_28667_, _28666_, _28661_);
  and _78909_ (_28669_, _28667_, _28433_);
  or _78910_ (_28670_, _28669_, _10976_);
  or _78911_ (_28671_, _11891_, _10975_);
  and _78912_ (_28672_, _28671_, _11016_);
  and _78913_ (_28673_, _28672_, _28670_);
  and _78914_ (_28674_, _28432_, _11015_);
  or _78915_ (_28675_, _28674_, _06049_);
  or _78916_ (_28676_, _28675_, _28673_);
  nand _78917_ (_28677_, _07353_, _06049_);
  and _78918_ (_28678_, _28677_, _28676_);
  or _78919_ (_28680_, _28678_, _05747_);
  or _78920_ (_28681_, _11891_, _05748_);
  and _78921_ (_28682_, _28681_, _06704_);
  and _78922_ (_28683_, _28682_, _28680_);
  or _78923_ (_28684_, _28442_, _12722_);
  nand _78924_ (_28685_, _12037_, _12722_);
  and _78925_ (_28686_, _28685_, _28684_);
  and _78926_ (_28687_, _28686_, _06126_);
  or _78927_ (_28688_, _28687_, _12750_);
  or _78928_ (_28689_, _28688_, _28683_);
  or _78929_ (_28691_, _28432_, _12749_);
  and _78930_ (_28692_, _28691_, _06718_);
  and _78931_ (_28693_, _28692_, _28689_);
  nand _78932_ (_28694_, _11891_, _06316_);
  nand _78933_ (_28695_, _28694_, _12756_);
  or _78934_ (_28696_, _28695_, _28693_);
  or _78935_ (_28697_, _28432_, _12756_);
  and _78936_ (_28698_, _28697_, _09200_);
  and _78937_ (_28699_, _28698_, _28696_);
  nor _78938_ (_28700_, _09200_, _05983_);
  or _78939_ (_28702_, _28700_, _05752_);
  or _78940_ (_28703_, _28702_, _28699_);
  or _78941_ (_28704_, _11891_, _12766_);
  and _78942_ (_28705_, _28704_, _05653_);
  and _78943_ (_28706_, _28705_, _28703_);
  and _78944_ (_28707_, _28686_, _05652_);
  or _78945_ (_28708_, _28707_, _12772_);
  or _78946_ (_28709_, _28708_, _28706_);
  or _78947_ (_28710_, _28432_, _12771_);
  and _78948_ (_28711_, _28710_, _06048_);
  and _78949_ (_28713_, _28711_, _28709_);
  nand _78950_ (_28714_, _11891_, _06047_);
  nand _78951_ (_28715_, _28714_, _12779_);
  or _78952_ (_28716_, _28715_, _28713_);
  or _78953_ (_28717_, _28432_, _12779_);
  and _78954_ (_28718_, _28717_, _12782_);
  and _78955_ (_28719_, _28718_, _28716_);
  nor _78956_ (_28720_, _12782_, _05983_);
  or _78957_ (_28721_, _28720_, _05751_);
  or _78958_ (_28722_, _28721_, _28719_);
  or _78959_ (_28724_, _11891_, _12791_);
  and _78960_ (_28725_, _28724_, _12790_);
  and _78961_ (_28726_, _28725_, _28722_);
  and _78962_ (_28727_, _28432_, _12789_);
  or _78963_ (_28728_, _28727_, _28726_);
  or _78964_ (_28729_, _28728_, _01340_);
  or _78965_ (_28730_, _01336_, \oc8051_golden_model_1.PC [11]);
  and _78966_ (_28731_, _28730_, _42882_);
  and _78967_ (_43429_, _28731_, _28729_);
  and _78968_ (_28732_, _15062_, _05752_);
  and _78969_ (_28734_, _11884_, _10606_);
  and _78970_ (_28735_, _11967_, _11964_);
  nor _78971_ (_28736_, _28735_, _11968_);
  and _78972_ (_28737_, _28736_, \oc8051_golden_model_1.PSW [7]);
  or _78973_ (_28738_, _28737_, _28734_);
  and _78974_ (_28739_, _28738_, _11982_);
  nor _78975_ (_28740_, _11884_, _08742_);
  nor _78976_ (_28741_, _12033_, _05669_);
  and _78977_ (_28742_, _12129_, _12126_);
  nor _78978_ (_28743_, _28742_, _12130_);
  and _78979_ (_28745_, _28743_, _12174_);
  and _78980_ (_28746_, _12172_, _12032_);
  nor _78981_ (_28747_, _28746_, _28745_);
  nor _78982_ (_28748_, _28747_, _12258_);
  nand _78983_ (_28749_, _12289_, _12033_);
  or _78984_ (_28750_, _28743_, _12289_);
  and _78985_ (_28751_, _28750_, _12256_);
  and _78986_ (_28752_, _28751_, _28749_);
  and _78987_ (_28753_, _11862_, _09202_);
  and _78988_ (_28754_, _28753_, \oc8051_golden_model_1.PC [11]);
  and _78989_ (_28756_, _28754_, \oc8051_golden_model_1.PC [12]);
  nor _78990_ (_28757_, _28754_, \oc8051_golden_model_1.PC [12]);
  nor _78991_ (_28758_, _28757_, _28756_);
  nor _78992_ (_28759_, _28758_, _12225_);
  or _78993_ (_28760_, _12187_, _12033_);
  not _78994_ (_28761_, _28743_);
  or _78995_ (_28762_, _28761_, _12189_);
  and _78996_ (_28763_, _28762_, _06102_);
  and _78997_ (_28764_, _28763_, _28760_);
  nor _78998_ (_28765_, _12199_, _11884_);
  or _78999_ (_28767_, _28736_, _12197_);
  nand _79000_ (_28768_, _28767_, _08384_);
  or _79001_ (_28769_, _28768_, _28765_);
  nor _79002_ (_28770_, _28758_, _12215_);
  nor _79003_ (_28771_, _12206_, _11884_);
  or _79004_ (_28772_, _06938_, \oc8051_golden_model_1.PC [12]);
  or _79005_ (_28773_, _28772_, _12208_);
  nor _79006_ (_28774_, _28773_, _07250_);
  or _79007_ (_28775_, _28774_, _28771_);
  and _79008_ (_28776_, _28775_, _12205_);
  or _79009_ (_28778_, _28776_, _08384_);
  or _79010_ (_28779_, _28778_, _28770_);
  and _79011_ (_28780_, _28779_, _12219_);
  and _79012_ (_28781_, _28780_, _28769_);
  or _79013_ (_28782_, _28781_, _28764_);
  and _79014_ (_28783_, _28782_, _12182_);
  or _79015_ (_28784_, _28783_, _28759_);
  nand _79016_ (_28785_, _28784_, _12179_);
  nor _79017_ (_28786_, _12179_, _11884_);
  nor _79018_ (_28787_, _28786_, _12232_);
  nand _79019_ (_28789_, _28787_, _28785_);
  not _79020_ (_28790_, _28758_);
  nor _79021_ (_28791_, _28790_, _12231_);
  nor _79022_ (_28792_, _28791_, _06219_);
  nand _79023_ (_28793_, _28792_, _28789_);
  and _79024_ (_28794_, _15062_, _06219_);
  nor _79025_ (_28795_, _28794_, _12241_);
  nand _79026_ (_28796_, _28795_, _28793_);
  nor _79027_ (_28797_, _28790_, _12239_);
  nor _79028_ (_28798_, _28797_, _12246_);
  nand _79029_ (_28800_, _28798_, _28796_);
  nor _79030_ (_28801_, _12245_, _11884_);
  not _79031_ (_28802_, _28801_);
  and _79032_ (_28803_, _28802_, _12255_);
  and _79033_ (_28804_, _28803_, _28800_);
  or _79034_ (_28805_, _28804_, _28752_);
  and _79035_ (_28806_, _28805_, _12258_);
  or _79036_ (_28807_, _28806_, _28748_);
  and _79037_ (_28808_, _28807_, _06509_);
  and _79038_ (_28809_, _12310_, _12032_);
  nor _79039_ (_28811_, _28761_, _12310_);
  nor _79040_ (_28812_, _28811_, _28809_);
  nor _79041_ (_28813_, _28812_, _06509_);
  or _79042_ (_28814_, _28813_, _28808_);
  nand _79043_ (_28815_, _28814_, _12298_);
  nand _79044_ (_28816_, _12329_, _12032_);
  nand _79045_ (_28817_, _28743_, _26881_);
  and _79046_ (_28818_, _28817_, _28816_);
  or _79047_ (_28819_, _28818_, _12298_);
  nand _79048_ (_28820_, _28819_, _28815_);
  nand _79049_ (_28822_, _28820_, _12013_);
  and _79050_ (_28823_, _28758_, _12012_);
  not _79051_ (_28824_, _28823_);
  and _79052_ (_28825_, _28824_, _12345_);
  nand _79053_ (_28826_, _28825_, _28822_);
  nor _79054_ (_28827_, _12345_, _11884_);
  nor _79055_ (_28828_, _28827_, _12355_);
  nand _79056_ (_28829_, _28828_, _28826_);
  nor _79057_ (_28830_, _28790_, _12351_);
  nor _79058_ (_28831_, _28830_, _12358_);
  nand _79059_ (_28833_, _28831_, _28829_);
  nor _79060_ (_28834_, _12357_, _11884_);
  nor _79061_ (_28835_, _28834_, _12368_);
  nand _79062_ (_28836_, _28835_, _28833_);
  or _79063_ (_28837_, _28790_, _12362_);
  and _79064_ (_28838_, _28837_, _12366_);
  nand _79065_ (_28839_, _28838_, _28836_);
  nor _79066_ (_28840_, _11884_, _12366_);
  nor _79067_ (_28841_, _28840_, _05676_);
  nand _79068_ (_28842_, _28841_, _28839_);
  nor _79069_ (_28844_, _28790_, _05675_);
  not _79070_ (_28845_, _28844_);
  and _79071_ (_28846_, _28845_, _12376_);
  nand _79072_ (_28847_, _28846_, _28842_);
  nor _79073_ (_28848_, _12376_, _11884_);
  nor _79074_ (_28849_, _28848_, _06110_);
  nand _79075_ (_28850_, _28849_, _28847_);
  and _79076_ (_28851_, _12032_, _06110_);
  nor _79077_ (_28852_, _28851_, _09818_);
  nand _79078_ (_28853_, _28852_, _28850_);
  nor _79079_ (_28855_, _11884_, _09817_);
  nor _79080_ (_28856_, _28855_, _09833_);
  and _79081_ (_28857_, _28856_, _28853_);
  or _79082_ (_28858_, _28857_, _28741_);
  nand _79083_ (_28859_, _28858_, _12389_);
  nor _79084_ (_28860_, _28790_, _12389_);
  nor _79085_ (_28861_, _28860_, _12392_);
  nand _79086_ (_28862_, _28861_, _28859_);
  nor _79087_ (_28863_, _12391_, _11884_);
  nor _79088_ (_28864_, _28863_, _12397_);
  nand _79089_ (_28866_, _28864_, _28862_);
  and _79090_ (_28867_, _28736_, _12397_);
  nor _79091_ (_28868_, _28867_, _08743_);
  and _79092_ (_28869_, _28868_, _28866_);
  or _79093_ (_28870_, _28869_, _28740_);
  nand _79094_ (_28871_, _28870_, _06020_);
  and _79095_ (_28872_, _12033_, _06019_);
  nor _79096_ (_28873_, _28872_, _10661_);
  and _79097_ (_28874_, _28873_, _28871_);
  and _79098_ (_28875_, _11884_, _10661_);
  or _79099_ (_28877_, _28875_, _28874_);
  nand _79100_ (_28878_, _28877_, _12413_);
  nor _79101_ (_28879_, _12443_, \oc8051_golden_model_1.DPH [4]);
  nor _79102_ (_28880_, _28879_, _12444_);
  and _79103_ (_28881_, _28880_, _12412_);
  nor _79104_ (_28882_, _28881_, _12416_);
  nand _79105_ (_28883_, _28882_, _28878_);
  nor _79106_ (_28884_, _12415_, _11884_);
  nor _79107_ (_28885_, _28884_, _12453_);
  and _79108_ (_28886_, _28885_, _28883_);
  and _79109_ (_28888_, _11884_, _11071_);
  and _79110_ (_28889_, _28736_, _12459_);
  or _79111_ (_28890_, _28889_, _28888_);
  and _79112_ (_28891_, _28890_, _12453_);
  or _79113_ (_28892_, _28891_, _28886_);
  nand _79114_ (_28893_, _28892_, _12007_);
  and _79115_ (_28894_, _28758_, _12006_);
  nor _79116_ (_28895_, _28894_, _12467_);
  nand _79117_ (_28896_, _28895_, _28893_);
  nor _79118_ (_28897_, _12466_, _11884_);
  nor _79119_ (_28899_, _28897_, _06112_);
  nand _79120_ (_28900_, _28899_, _28896_);
  not _79121_ (_28901_, _12473_);
  and _79122_ (_28902_, _12032_, _06112_);
  nor _79123_ (_28903_, _28902_, _28901_);
  nand _79124_ (_28904_, _28903_, _28900_);
  nor _79125_ (_28905_, _12473_, _11884_);
  nor _79126_ (_28906_, _28905_, _12476_);
  and _79127_ (_28907_, _28906_, _28904_);
  and _79128_ (_28908_, _11884_, _12459_);
  and _79129_ (_28910_, _28736_, _11071_);
  or _79130_ (_28911_, _28910_, _28908_);
  and _79131_ (_28912_, _28911_, _12476_);
  or _79132_ (_28913_, _28912_, _28907_);
  nand _79133_ (_28914_, _28913_, _12002_);
  nor _79134_ (_28915_, _28790_, _12002_);
  nor _79135_ (_28916_, _28915_, _10743_);
  nand _79136_ (_28917_, _28916_, _28914_);
  nor _79137_ (_28918_, _11884_, _10742_);
  nor _79138_ (_28919_, _28918_, _06108_);
  nand _79139_ (_28921_, _28919_, _28917_);
  not _79140_ (_28922_, _12494_);
  and _79141_ (_28923_, _12032_, _06108_);
  nor _79142_ (_28924_, _28923_, _28922_);
  nand _79143_ (_28925_, _28924_, _28921_);
  nor _79144_ (_28926_, _12494_, _11884_);
  nor _79145_ (_28927_, _28926_, _12497_);
  and _79146_ (_28928_, _28927_, _28925_);
  and _79147_ (_28929_, _11884_, \oc8051_golden_model_1.PSW [7]);
  and _79148_ (_28930_, _28736_, _10606_);
  or _79149_ (_28932_, _28930_, _28929_);
  and _79150_ (_28933_, _28932_, _12497_);
  or _79151_ (_28934_, _28933_, _28928_);
  nand _79152_ (_28935_, _28934_, _11993_);
  nor _79153_ (_28936_, _28790_, _11993_);
  nor _79154_ (_28937_, _28936_, _11987_);
  nand _79155_ (_28938_, _28937_, _28935_);
  nor _79156_ (_28939_, _11884_, _11986_);
  nor _79157_ (_28940_, _28939_, _06130_);
  nand _79158_ (_28941_, _28940_, _28938_);
  not _79159_ (_28943_, _12515_);
  and _79160_ (_28944_, _12032_, _06130_);
  nor _79161_ (_28945_, _28944_, _28943_);
  nand _79162_ (_28946_, _28945_, _28941_);
  nor _79163_ (_28947_, _12515_, _11884_);
  nor _79164_ (_28948_, _28947_, _11982_);
  and _79165_ (_28949_, _28948_, _28946_);
  or _79166_ (_28950_, _28949_, _28739_);
  nand _79167_ (_28951_, _28950_, _12523_);
  nor _79168_ (_28952_, _28790_, _12523_);
  nor _79169_ (_28954_, _28952_, _10826_);
  nand _79170_ (_28955_, _28954_, _28951_);
  nor _79171_ (_28956_, _11884_, _10825_);
  nor _79172_ (_28957_, _28956_, _10854_);
  nand _79173_ (_28958_, _28957_, _28955_);
  and _79174_ (_28959_, _28758_, _10854_);
  nor _79175_ (_28960_, _28959_, _06298_);
  and _79176_ (_28961_, _28960_, _28958_);
  and _79177_ (_28962_, _08270_, _06298_);
  or _79178_ (_28963_, _28962_, _28961_);
  nand _79179_ (_28965_, _28963_, _05734_);
  and _79180_ (_28966_, _15062_, _05732_);
  nor _79181_ (_28967_, _28966_, _06129_);
  and _79182_ (_28968_, _28967_, _28965_);
  and _79183_ (_28969_, _28743_, _12722_);
  nor _79184_ (_28970_, _12033_, _12722_);
  nor _79185_ (_28971_, _28970_, _28969_);
  nor _79186_ (_28972_, _28971_, _06306_);
  or _79187_ (_28973_, _28972_, _28968_);
  nand _79188_ (_28974_, _28973_, _11872_);
  nor _79189_ (_28976_, _28790_, _11872_);
  nor _79190_ (_28977_, _28976_, _10976_);
  nand _79191_ (_28978_, _28977_, _28974_);
  nor _79192_ (_28979_, _11884_, _10975_);
  nor _79193_ (_28980_, _28979_, _11015_);
  nand _79194_ (_28981_, _28980_, _28978_);
  and _79195_ (_28982_, _28758_, _11015_);
  nor _79196_ (_28983_, _28982_, _06049_);
  nand _79197_ (_28984_, _28983_, _28981_);
  and _79198_ (_28985_, _08270_, _06049_);
  nor _79199_ (_28987_, _28985_, _05747_);
  and _79200_ (_28988_, _28987_, _28984_);
  and _79201_ (_28989_, _11884_, _05747_);
  or _79202_ (_28990_, _28989_, _06126_);
  or _79203_ (_28991_, _28990_, _28988_);
  nor _79204_ (_28992_, _28743_, _12722_);
  and _79205_ (_28993_, _12033_, _12722_);
  nor _79206_ (_28994_, _28993_, _28992_);
  nor _79207_ (_28995_, _28994_, _06704_);
  nor _79208_ (_28996_, _28995_, _12750_);
  nand _79209_ (_28997_, _28996_, _28991_);
  nor _79210_ (_28998_, _28790_, _12749_);
  nor _79211_ (_28999_, _28998_, _06316_);
  nand _79212_ (_29000_, _28999_, _28997_);
  and _79213_ (_29001_, _15062_, _06316_);
  nor _79214_ (_29002_, _29001_, _25353_);
  and _79215_ (_29003_, _29002_, _29000_);
  nor _79216_ (_29004_, _28790_, _12756_);
  or _79217_ (_29005_, _29004_, _06127_);
  nor _79218_ (_29006_, _29005_, _29003_);
  and _79219_ (_29009_, _06758_, _06127_);
  or _79220_ (_29010_, _29009_, _29006_);
  and _79221_ (_29011_, _29010_, _12766_);
  or _79222_ (_29012_, _29011_, _28732_);
  nand _79223_ (_29013_, _29012_, _05653_);
  nor _79224_ (_29014_, _28994_, _05653_);
  nor _79225_ (_29015_, _29014_, _12772_);
  nand _79226_ (_29016_, _29015_, _29013_);
  nor _79227_ (_29017_, _28790_, _12771_);
  nor _79228_ (_29018_, _29017_, _06047_);
  nand _79229_ (_29020_, _29018_, _29016_);
  and _79230_ (_29021_, _15062_, _06047_);
  nor _79231_ (_29022_, _29021_, _26405_);
  nand _79232_ (_29023_, _29022_, _29020_);
  nor _79233_ (_29024_, _28790_, _12779_);
  nor _79234_ (_29025_, _29024_, _06119_);
  nand _79235_ (_29026_, _29025_, _29023_);
  and _79236_ (_29027_, _06758_, _06119_);
  nor _79237_ (_29028_, _29027_, _05751_);
  nand _79238_ (_29029_, _29028_, _29026_);
  and _79239_ (_29031_, _11884_, _05751_);
  nor _79240_ (_29032_, _29031_, _12789_);
  and _79241_ (_29033_, _29032_, _29029_);
  and _79242_ (_29034_, _28790_, _12789_);
  nor _79243_ (_29035_, _29034_, _29033_);
  or _79244_ (_29036_, _29035_, _01340_);
  or _79245_ (_29037_, _01336_, \oc8051_golden_model_1.PC [12]);
  and _79246_ (_29038_, _29037_, _42882_);
  and _79247_ (_43430_, _29038_, _29036_);
  and _79248_ (_29039_, _28756_, \oc8051_golden_model_1.PC [13]);
  nor _79249_ (_29041_, _28756_, \oc8051_golden_model_1.PC [13]);
  nor _79250_ (_29042_, _29041_, _29039_);
  or _79251_ (_29043_, _29042_, _11872_);
  or _79252_ (_29044_, _29042_, _12523_);
  or _79253_ (_29045_, _29042_, _11993_);
  or _79254_ (_29046_, _11882_, _11881_);
  not _79255_ (_29047_, _29046_);
  nor _79256_ (_29048_, _29047_, _11969_);
  and _79257_ (_29049_, _29047_, _11969_);
  or _79258_ (_29050_, _29049_, _29048_);
  or _79259_ (_29052_, _29050_, _11071_);
  or _79260_ (_29053_, _11880_, _12459_);
  and _79261_ (_29054_, _29053_, _12453_);
  and _79262_ (_29055_, _29054_, _29052_);
  or _79263_ (_29056_, _11880_, _08742_);
  nor _79264_ (_29057_, _12028_, _05669_);
  or _79265_ (_29058_, _12030_, _12029_);
  not _79266_ (_29059_, _29058_);
  nor _79267_ (_29060_, _29059_, _12131_);
  and _79268_ (_29061_, _29059_, _12131_);
  or _79269_ (_29063_, _29061_, _29060_);
  or _79270_ (_29064_, _29063_, _12172_);
  nor _79271_ (_29065_, _12174_, _12027_);
  nor _79272_ (_29066_, _29065_, _12258_);
  and _79273_ (_29067_, _29066_, _29064_);
  and _79274_ (_29068_, _11880_, _06219_);
  or _79275_ (_29069_, _12179_, _11880_);
  or _79276_ (_29070_, _12187_, _12027_);
  or _79277_ (_29071_, _29063_, _12189_);
  and _79278_ (_29072_, _29071_, _06102_);
  and _79279_ (_29074_, _29072_, _29070_);
  and _79280_ (_29075_, _29050_, _12199_);
  and _79281_ (_29076_, _12197_, _11880_);
  or _79282_ (_29077_, _29076_, _08383_);
  or _79283_ (_29078_, _29077_, _29075_);
  or _79284_ (_29079_, _29042_, _12215_);
  or _79285_ (_29080_, _12206_, _11880_);
  or _79286_ (_29081_, _06530_, \oc8051_golden_model_1.PC [13]);
  or _79287_ (_29082_, _29081_, _06938_);
  nor _79288_ (_29083_, _29082_, _07250_);
  nand _79289_ (_29085_, _29083_, _24785_);
  and _79290_ (_29086_, _29085_, _29080_);
  and _79291_ (_29087_, _29086_, _29079_);
  or _79292_ (_29088_, _29087_, _08384_);
  and _79293_ (_29089_, _29088_, _12219_);
  and _79294_ (_29090_, _29089_, _29078_);
  or _79295_ (_29091_, _29090_, _29074_);
  and _79296_ (_29092_, _29091_, _12182_);
  not _79297_ (_29093_, _29042_);
  nor _79298_ (_29094_, _29093_, _12225_);
  or _79299_ (_29096_, _29094_, _12224_);
  or _79300_ (_29097_, _29096_, _29092_);
  and _79301_ (_29098_, _29097_, _29069_);
  or _79302_ (_29099_, _29098_, _12232_);
  or _79303_ (_29100_, _29042_, _12231_);
  and _79304_ (_29101_, _29100_, _06220_);
  and _79305_ (_29102_, _29101_, _29099_);
  or _79306_ (_29103_, _29102_, _29068_);
  and _79307_ (_29104_, _29103_, _12239_);
  or _79308_ (_29105_, _29093_, _12239_);
  nand _79309_ (_29107_, _29105_, _12245_);
  or _79310_ (_29108_, _29107_, _29104_);
  or _79311_ (_29109_, _12245_, _11880_);
  and _79312_ (_29110_, _29109_, _29108_);
  or _79313_ (_29111_, _29110_, _12256_);
  or _79314_ (_29112_, _29063_, _12289_);
  nand _79315_ (_29113_, _12289_, _12028_);
  and _79316_ (_29114_, _29113_, _29112_);
  or _79317_ (_29115_, _29114_, _12255_);
  and _79318_ (_29116_, _29115_, _12258_);
  and _79319_ (_29118_, _29116_, _29111_);
  or _79320_ (_29119_, _29118_, _06121_);
  or _79321_ (_29120_, _29119_, _29067_);
  and _79322_ (_29121_, _12310_, _12027_);
  and _79323_ (_29122_, _29063_, _12312_);
  or _79324_ (_29123_, _29122_, _06509_);
  or _79325_ (_29124_, _29123_, _29121_);
  and _79326_ (_29125_, _29124_, _12298_);
  and _79327_ (_29126_, _29125_, _29120_);
  or _79328_ (_29127_, _29063_, _12329_);
  nand _79329_ (_29129_, _12329_, _12028_);
  and _79330_ (_29130_, _29129_, _06115_);
  and _79331_ (_29131_, _29130_, _29127_);
  or _79332_ (_29132_, _29131_, _29126_);
  and _79333_ (_29133_, _29132_, _12013_);
  nand _79334_ (_29134_, _29042_, _12012_);
  nand _79335_ (_29135_, _29134_, _12345_);
  or _79336_ (_29136_, _29135_, _29133_);
  or _79337_ (_29137_, _12345_, _11880_);
  and _79338_ (_29138_, _29137_, _12351_);
  and _79339_ (_29140_, _29138_, _29136_);
  nor _79340_ (_29141_, _29093_, _12351_);
  or _79341_ (_29142_, _29141_, _12358_);
  or _79342_ (_29143_, _29142_, _29140_);
  or _79343_ (_29144_, _12357_, _11880_);
  and _79344_ (_29145_, _29144_, _12362_);
  and _79345_ (_29146_, _29145_, _29143_);
  or _79346_ (_29147_, _29093_, _12362_);
  nand _79347_ (_29148_, _29147_, _12366_);
  or _79348_ (_29149_, _29148_, _29146_);
  or _79349_ (_29151_, _11880_, _12366_);
  and _79350_ (_29152_, _29151_, _05675_);
  and _79351_ (_29153_, _29152_, _29149_);
  or _79352_ (_29154_, _29093_, _05675_);
  nand _79353_ (_29155_, _29154_, _12376_);
  or _79354_ (_29156_, _29155_, _29153_);
  or _79355_ (_29157_, _12376_, _11880_);
  and _79356_ (_29158_, _29157_, _06111_);
  and _79357_ (_29159_, _29158_, _29156_);
  nand _79358_ (_29160_, _12027_, _06110_);
  nand _79359_ (_29162_, _29160_, _09817_);
  or _79360_ (_29163_, _29162_, _29159_);
  or _79361_ (_29164_, _11880_, _09817_);
  and _79362_ (_29165_, _29164_, _05669_);
  and _79363_ (_29166_, _29165_, _29163_);
  or _79364_ (_29167_, _29166_, _29057_);
  and _79365_ (_29168_, _29167_, _12389_);
  nor _79366_ (_29169_, _29093_, _12389_);
  or _79367_ (_29170_, _29169_, _12392_);
  or _79368_ (_29171_, _29170_, _29168_);
  or _79369_ (_29173_, _12391_, _11880_);
  and _79370_ (_29174_, _29173_, _12398_);
  and _79371_ (_29175_, _29174_, _29171_);
  and _79372_ (_29176_, _29050_, _12397_);
  or _79373_ (_29177_, _29176_, _08743_);
  or _79374_ (_29178_, _29177_, _29175_);
  and _79375_ (_29179_, _29178_, _29056_);
  or _79376_ (_29180_, _29179_, _06019_);
  nand _79377_ (_29181_, _12028_, _06019_);
  and _79378_ (_29182_, _29181_, _10662_);
  and _79379_ (_29184_, _29182_, _29180_);
  and _79380_ (_29185_, _11880_, _10661_);
  or _79381_ (_29186_, _29185_, _29184_);
  and _79382_ (_29187_, _29186_, _12413_);
  or _79383_ (_29188_, _12444_, \oc8051_golden_model_1.DPH [5]);
  nor _79384_ (_29189_, _12445_, _12413_);
  and _79385_ (_29190_, _29189_, _29188_);
  or _79386_ (_29191_, _29190_, _12416_);
  or _79387_ (_29192_, _29191_, _29187_);
  or _79388_ (_29193_, _12415_, _11880_);
  and _79389_ (_29195_, _29193_, _12454_);
  and _79390_ (_29196_, _29195_, _29192_);
  or _79391_ (_29197_, _29196_, _29055_);
  and _79392_ (_29198_, _29197_, _12007_);
  and _79393_ (_29199_, _29042_, _12006_);
  or _79394_ (_29200_, _29199_, _12467_);
  or _79395_ (_29201_, _29200_, _29198_);
  or _79396_ (_29202_, _12466_, _11880_);
  and _79397_ (_29203_, _29202_, _08751_);
  and _79398_ (_29204_, _29203_, _29201_);
  nand _79399_ (_29206_, _12027_, _06112_);
  nand _79400_ (_29207_, _29206_, _12473_);
  or _79401_ (_29208_, _29207_, _29204_);
  or _79402_ (_29209_, _12473_, _11880_);
  and _79403_ (_29210_, _29209_, _12477_);
  and _79404_ (_29211_, _29210_, _29208_);
  or _79405_ (_29212_, _29050_, _12459_);
  or _79406_ (_29213_, _11880_, _11071_);
  and _79407_ (_29214_, _29213_, _12476_);
  and _79408_ (_29215_, _29214_, _29212_);
  or _79409_ (_29217_, _29215_, _29211_);
  and _79410_ (_29218_, _29217_, _12002_);
  nor _79411_ (_29219_, _29093_, _12002_);
  or _79412_ (_29220_, _29219_, _10743_);
  or _79413_ (_29221_, _29220_, _29218_);
  or _79414_ (_29222_, _11880_, _10742_);
  and _79415_ (_29223_, _29222_, _07032_);
  and _79416_ (_29224_, _29223_, _29221_);
  nand _79417_ (_29225_, _12027_, _06108_);
  nand _79418_ (_29226_, _29225_, _12494_);
  or _79419_ (_29228_, _29226_, _29224_);
  or _79420_ (_29229_, _12494_, _11880_);
  and _79421_ (_29230_, _29229_, _12498_);
  and _79422_ (_29231_, _29230_, _29228_);
  or _79423_ (_29232_, _29050_, \oc8051_golden_model_1.PSW [7]);
  or _79424_ (_29233_, _11880_, _10606_);
  and _79425_ (_29234_, _29233_, _12497_);
  and _79426_ (_29235_, _29234_, _29232_);
  or _79427_ (_29236_, _29235_, _12502_);
  or _79428_ (_29237_, _29236_, _29231_);
  and _79429_ (_29239_, _29237_, _29045_);
  or _79430_ (_29240_, _29239_, _11987_);
  or _79431_ (_29241_, _11880_, _11986_);
  and _79432_ (_29242_, _29241_, _08777_);
  and _79433_ (_29243_, _29242_, _29240_);
  nand _79434_ (_29244_, _12027_, _06130_);
  nand _79435_ (_29245_, _29244_, _12515_);
  or _79436_ (_29246_, _29245_, _29243_);
  or _79437_ (_29247_, _12515_, _11880_);
  and _79438_ (_29248_, _29247_, _12518_);
  and _79439_ (_29250_, _29248_, _29246_);
  or _79440_ (_29251_, _29050_, _10606_);
  or _79441_ (_29252_, _11880_, \oc8051_golden_model_1.PSW [7]);
  and _79442_ (_29253_, _29252_, _11982_);
  and _79443_ (_29254_, _29253_, _29251_);
  or _79444_ (_29255_, _29254_, _12525_);
  or _79445_ (_29256_, _29255_, _29250_);
  and _79446_ (_29257_, _29256_, _29044_);
  or _79447_ (_29258_, _29257_, _10826_);
  or _79448_ (_29259_, _11880_, _10825_);
  and _79449_ (_29261_, _29259_, _10855_);
  and _79450_ (_29262_, _29261_, _29258_);
  and _79451_ (_29263_, _29042_, _10854_);
  or _79452_ (_29264_, _29263_, _06298_);
  or _79453_ (_29265_, _29264_, _29262_);
  nand _79454_ (_29266_, _07977_, _06298_);
  and _79455_ (_29267_, _29266_, _29265_);
  or _79456_ (_29268_, _29267_, _05732_);
  nand _79457_ (_29269_, _15259_, _05732_);
  and _79458_ (_29270_, _29269_, _06306_);
  and _79459_ (_29272_, _29270_, _29268_);
  or _79460_ (_29273_, _29063_, _12723_);
  or _79461_ (_29274_, _12027_, _12722_);
  and _79462_ (_29275_, _29274_, _06129_);
  and _79463_ (_29276_, _29275_, _29273_);
  or _79464_ (_29277_, _29276_, _12541_);
  or _79465_ (_29278_, _29277_, _29272_);
  and _79466_ (_29279_, _29278_, _29043_);
  or _79467_ (_29280_, _29279_, _10976_);
  or _79468_ (_29281_, _11880_, _10975_);
  and _79469_ (_29283_, _29281_, _11016_);
  and _79470_ (_29284_, _29283_, _29280_);
  and _79471_ (_29285_, _29042_, _11015_);
  or _79472_ (_29286_, _29285_, _06049_);
  or _79473_ (_29287_, _29286_, _29284_);
  nand _79474_ (_29288_, _07977_, _06049_);
  and _79475_ (_29289_, _29288_, _29287_);
  or _79476_ (_29290_, _29289_, _05747_);
  nand _79477_ (_29291_, _15259_, _05747_);
  and _79478_ (_29292_, _29291_, _06704_);
  and _79479_ (_29294_, _29292_, _29290_);
  or _79480_ (_29295_, _29063_, _12722_);
  nand _79481_ (_29296_, _12028_, _12722_);
  and _79482_ (_29297_, _29296_, _29295_);
  and _79483_ (_29298_, _29297_, _06126_);
  or _79484_ (_29299_, _29298_, _12750_);
  or _79485_ (_29300_, _29299_, _29294_);
  or _79486_ (_29301_, _29042_, _12749_);
  and _79487_ (_29302_, _29301_, _06718_);
  and _79488_ (_29303_, _29302_, _29300_);
  nand _79489_ (_29305_, _11880_, _06316_);
  nand _79490_ (_29306_, _29305_, _12756_);
  or _79491_ (_29307_, _29306_, _29303_);
  or _79492_ (_29308_, _29042_, _12756_);
  and _79493_ (_29309_, _29308_, _09200_);
  and _79494_ (_29310_, _29309_, _29307_);
  nor _79495_ (_29311_, _06359_, _09200_);
  or _79496_ (_29312_, _29311_, _05752_);
  or _79497_ (_29313_, _29312_, _29310_);
  nand _79498_ (_29314_, _15259_, _05752_);
  and _79499_ (_29316_, _29314_, _05653_);
  and _79500_ (_29317_, _29316_, _29313_);
  and _79501_ (_29318_, _29297_, _05652_);
  or _79502_ (_29319_, _29318_, _12772_);
  or _79503_ (_29320_, _29319_, _29317_);
  or _79504_ (_29321_, _29042_, _12771_);
  and _79505_ (_29322_, _29321_, _06048_);
  and _79506_ (_29323_, _29322_, _29320_);
  nand _79507_ (_29324_, _11880_, _06047_);
  nand _79508_ (_29325_, _29324_, _12779_);
  or _79509_ (_29327_, _29325_, _29323_);
  or _79510_ (_29328_, _29042_, _12779_);
  and _79511_ (_29329_, _29328_, _12782_);
  and _79512_ (_29330_, _29329_, _29327_);
  nor _79513_ (_29331_, _06359_, _12782_);
  or _79514_ (_29332_, _29331_, _05751_);
  or _79515_ (_29333_, _29332_, _29330_);
  nand _79516_ (_29334_, _15259_, _05751_);
  and _79517_ (_29335_, _29334_, _12790_);
  and _79518_ (_29336_, _29335_, _29333_);
  and _79519_ (_29338_, _29042_, _12789_);
  or _79520_ (_29339_, _29338_, _29336_);
  or _79521_ (_29340_, _29339_, _01340_);
  or _79522_ (_29341_, _01336_, \oc8051_golden_model_1.PC [13]);
  and _79523_ (_29342_, _29341_, _42882_);
  and _79524_ (_43431_, _29342_, _29340_);
  and _79525_ (_29343_, _15457_, _06047_);
  nor _79526_ (_29344_, _29039_, \oc8051_golden_model_1.PC [14]);
  nor _79527_ (_29345_, _29344_, _11868_);
  not _79528_ (_29346_, _29345_);
  nand _79529_ (_29348_, _29346_, _11015_);
  nor _79530_ (_29349_, _12515_, _15457_);
  nor _79531_ (_29350_, _12494_, _15457_);
  nor _79532_ (_29351_, _12473_, _15457_);
  or _79533_ (_29352_, _29345_, _12231_);
  and _79534_ (_29353_, _29345_, _06948_);
  and _79535_ (_29354_, _12197_, _11875_);
  nor _79536_ (_29355_, _11972_, _11878_);
  nor _79537_ (_29356_, _29355_, _11973_);
  and _79538_ (_29357_, _29356_, _12199_);
  or _79539_ (_29359_, _29357_, _29354_);
  or _79540_ (_29360_, _29359_, _08383_);
  or _79541_ (_29361_, _29345_, _12205_);
  nand _79542_ (_29362_, _12205_, _15457_);
  and _79543_ (_29363_, _29362_, _29361_);
  or _79544_ (_29364_, _29363_, _24785_);
  nor _79545_ (_29365_, _29346_, _12215_);
  nand _79546_ (_29366_, _15457_, _06938_);
  and _79547_ (_29367_, _29366_, _25758_);
  and _79548_ (_29368_, _07251_, \oc8051_golden_model_1.PC [14]);
  or _79549_ (_29370_, _29368_, _06938_);
  and _79550_ (_29371_, _29370_, _29367_);
  or _79551_ (_29372_, _29371_, _06943_);
  or _79552_ (_29373_, _29372_, _29365_);
  and _79553_ (_29374_, _29373_, _29364_);
  or _79554_ (_29375_, _29374_, _08384_);
  and _79555_ (_29376_, _29375_, _06949_);
  and _79556_ (_29377_, _29376_, _29360_);
  or _79557_ (_29378_, _29377_, _29353_);
  or _79558_ (_29379_, _29378_, _06102_);
  or _79559_ (_29381_, _12187_, _12020_);
  and _79560_ (_29382_, _12133_, _12025_);
  nor _79561_ (_29383_, _29382_, _12134_);
  or _79562_ (_29384_, _29383_, _12189_);
  and _79563_ (_29385_, _29384_, _29381_);
  or _79564_ (_29386_, _29385_, _06954_);
  and _79565_ (_29387_, _29386_, _29379_);
  or _79566_ (_29388_, _29387_, _24805_);
  or _79567_ (_29389_, _29345_, _12182_);
  and _79568_ (_29390_, _29389_, _12179_);
  and _79569_ (_29392_, _29390_, _29388_);
  nor _79570_ (_29393_, _12179_, _15457_);
  or _79571_ (_29394_, _29393_, _12232_);
  or _79572_ (_29395_, _29394_, _29392_);
  and _79573_ (_29396_, _29395_, _29352_);
  or _79574_ (_29397_, _29396_, _06219_);
  nand _79575_ (_29398_, _15457_, _06219_);
  and _79576_ (_29399_, _29398_, _12239_);
  and _79577_ (_29400_, _29399_, _29397_);
  nor _79578_ (_29401_, _29346_, _12239_);
  or _79579_ (_29403_, _29401_, _29400_);
  and _79580_ (_29404_, _29403_, _12245_);
  or _79581_ (_29405_, _12245_, _15457_);
  nand _79582_ (_29406_, _29405_, _12255_);
  or _79583_ (_29407_, _29406_, _29404_);
  and _79584_ (_29408_, _12289_, _12020_);
  not _79585_ (_29409_, _29383_);
  nor _79586_ (_29410_, _29409_, _12289_);
  or _79587_ (_29411_, _29410_, _29408_);
  or _79588_ (_29412_, _29411_, _12255_);
  and _79589_ (_29414_, _29412_, _12258_);
  and _79590_ (_29415_, _29414_, _29407_);
  nand _79591_ (_29416_, _29409_, _12174_);
  or _79592_ (_29417_, _12174_, _12020_);
  and _79593_ (_29418_, _29417_, _06104_);
  and _79594_ (_29419_, _29418_, _29416_);
  or _79595_ (_29420_, _29419_, _06121_);
  or _79596_ (_29421_, _29420_, _29415_);
  and _79597_ (_29422_, _12310_, _12020_);
  nor _79598_ (_29423_, _29409_, _12310_);
  or _79599_ (_29425_, _29423_, _06509_);
  or _79600_ (_29426_, _29425_, _29422_);
  and _79601_ (_29427_, _29426_, _12298_);
  and _79602_ (_29428_, _29427_, _29421_);
  or _79603_ (_29429_, _29383_, _12329_);
  nand _79604_ (_29430_, _12329_, _12021_);
  and _79605_ (_29431_, _29430_, _06115_);
  and _79606_ (_29432_, _29431_, _29429_);
  or _79607_ (_29433_, _29432_, _12012_);
  or _79608_ (_29434_, _29433_, _29428_);
  or _79609_ (_29436_, _29345_, _12013_);
  and _79610_ (_29437_, _29436_, _12345_);
  and _79611_ (_29438_, _29437_, _29434_);
  nor _79612_ (_29439_, _12345_, _15457_);
  or _79613_ (_29440_, _29439_, _12355_);
  or _79614_ (_29441_, _29440_, _29438_);
  or _79615_ (_29442_, _29345_, _12351_);
  and _79616_ (_29443_, _29442_, _12357_);
  and _79617_ (_29444_, _29443_, _29441_);
  nor _79618_ (_29445_, _12357_, _15457_);
  or _79619_ (_29447_, _29445_, _12368_);
  or _79620_ (_29448_, _29447_, _29444_);
  or _79621_ (_29449_, _29345_, _12362_);
  and _79622_ (_29450_, _29449_, _12366_);
  and _79623_ (_29451_, _29450_, _29448_);
  nor _79624_ (_29452_, _15457_, _12366_);
  or _79625_ (_29453_, _29452_, _05676_);
  or _79626_ (_29454_, _29453_, _29451_);
  or _79627_ (_29455_, _29345_, _05675_);
  and _79628_ (_29456_, _29455_, _12376_);
  and _79629_ (_29458_, _29456_, _29454_);
  nor _79630_ (_29459_, _12376_, _15457_);
  or _79631_ (_29460_, _29459_, _06110_);
  or _79632_ (_29461_, _29460_, _29458_);
  nand _79633_ (_29462_, _12021_, _06110_);
  and _79634_ (_29463_, _29462_, _09817_);
  and _79635_ (_29464_, _29463_, _29461_);
  nor _79636_ (_29465_, _15457_, _09817_);
  or _79637_ (_29466_, _29465_, _09833_);
  or _79638_ (_29467_, _29466_, _29464_);
  or _79639_ (_29469_, _12020_, _05669_);
  and _79640_ (_29470_, _29469_, _12389_);
  and _79641_ (_29471_, _29470_, _29467_);
  nor _79642_ (_29472_, _29346_, _12389_);
  or _79643_ (_29473_, _29472_, _12392_);
  or _79644_ (_29474_, _29473_, _29471_);
  or _79645_ (_29475_, _12391_, _11875_);
  and _79646_ (_29476_, _29475_, _12398_);
  and _79647_ (_29477_, _29476_, _29474_);
  and _79648_ (_29478_, _29356_, _12397_);
  or _79649_ (_29480_, _29478_, _08743_);
  or _79650_ (_29481_, _29480_, _29477_);
  or _79651_ (_29482_, _11875_, _08742_);
  and _79652_ (_29483_, _29482_, _29481_);
  or _79653_ (_29484_, _29483_, _06019_);
  nand _79654_ (_29485_, _12021_, _06019_);
  and _79655_ (_29486_, _29485_, _10662_);
  and _79656_ (_29487_, _29486_, _29484_);
  and _79657_ (_29488_, _11875_, _10661_);
  or _79658_ (_29489_, _29488_, _12412_);
  or _79659_ (_29491_, _29489_, _29487_);
  nor _79660_ (_29492_, _12445_, \oc8051_golden_model_1.DPH [6]);
  nor _79661_ (_29493_, _29492_, _12446_);
  or _79662_ (_29494_, _29493_, _12413_);
  and _79663_ (_29495_, _29494_, _12415_);
  and _79664_ (_29496_, _29495_, _29491_);
  nor _79665_ (_29497_, _12415_, _15457_);
  or _79666_ (_29498_, _29497_, _29496_);
  and _79667_ (_29499_, _29498_, _12454_);
  or _79668_ (_29500_, _29356_, _11071_);
  or _79669_ (_29502_, _11875_, _12459_);
  and _79670_ (_29503_, _29502_, _12453_);
  and _79671_ (_29504_, _29503_, _29500_);
  or _79672_ (_29505_, _29504_, _12006_);
  or _79673_ (_29506_, _29505_, _29499_);
  nand _79674_ (_29507_, _29346_, _12006_);
  and _79675_ (_29508_, _29507_, _12466_);
  and _79676_ (_29509_, _29508_, _29506_);
  nor _79677_ (_29510_, _12466_, _15457_);
  or _79678_ (_29511_, _29510_, _06112_);
  or _79679_ (_29513_, _29511_, _29509_);
  nand _79680_ (_29514_, _12021_, _06112_);
  and _79681_ (_29515_, _29514_, _12473_);
  and _79682_ (_29516_, _29515_, _29513_);
  or _79683_ (_29517_, _29516_, _29351_);
  and _79684_ (_29518_, _29517_, _12477_);
  or _79685_ (_29519_, _29356_, _12459_);
  or _79686_ (_29520_, _11875_, _11071_);
  and _79687_ (_29521_, _29520_, _12476_);
  and _79688_ (_29522_, _29521_, _29519_);
  or _79689_ (_29523_, _29522_, _12481_);
  or _79690_ (_29524_, _29523_, _29518_);
  or _79691_ (_29525_, _29345_, _12002_);
  and _79692_ (_29526_, _29525_, _10742_);
  and _79693_ (_29527_, _29526_, _29524_);
  nor _79694_ (_29528_, _15457_, _10742_);
  or _79695_ (_29529_, _29528_, _06108_);
  or _79696_ (_29530_, _29529_, _29527_);
  nand _79697_ (_29531_, _12021_, _06108_);
  and _79698_ (_29532_, _29531_, _12494_);
  and _79699_ (_29535_, _29532_, _29530_);
  or _79700_ (_29536_, _29535_, _29350_);
  and _79701_ (_29537_, _29536_, _12498_);
  or _79702_ (_29538_, _29356_, \oc8051_golden_model_1.PSW [7]);
  or _79703_ (_29539_, _11875_, _10606_);
  and _79704_ (_29540_, _29539_, _12497_);
  and _79705_ (_29541_, _29540_, _29538_);
  or _79706_ (_29542_, _29541_, _12502_);
  or _79707_ (_29543_, _29542_, _29537_);
  or _79708_ (_29544_, _29345_, _11993_);
  and _79709_ (_29546_, _29544_, _11986_);
  and _79710_ (_29547_, _29546_, _29543_);
  nor _79711_ (_29548_, _15457_, _11986_);
  or _79712_ (_29549_, _29548_, _06130_);
  or _79713_ (_29550_, _29549_, _29547_);
  nand _79714_ (_29551_, _12021_, _06130_);
  and _79715_ (_29552_, _29551_, _12515_);
  and _79716_ (_29553_, _29552_, _29550_);
  or _79717_ (_29554_, _29553_, _29349_);
  and _79718_ (_29555_, _29554_, _12518_);
  or _79719_ (_29557_, _29356_, _10606_);
  or _79720_ (_29558_, _11875_, \oc8051_golden_model_1.PSW [7]);
  and _79721_ (_29559_, _29558_, _11982_);
  and _79722_ (_29560_, _29559_, _29557_);
  or _79723_ (_29561_, _29560_, _12525_);
  or _79724_ (_29562_, _29561_, _29555_);
  or _79725_ (_29563_, _29345_, _12523_);
  and _79726_ (_29564_, _29563_, _10825_);
  and _79727_ (_29565_, _29564_, _29562_);
  nor _79728_ (_29566_, _15457_, _10825_);
  or _79729_ (_29568_, _29566_, _10854_);
  or _79730_ (_29569_, _29568_, _29565_);
  nand _79731_ (_29570_, _29346_, _10854_);
  and _79732_ (_29571_, _29570_, _13619_);
  and _79733_ (_29572_, _29571_, _29569_);
  nor _79734_ (_29573_, _07883_, _13619_);
  or _79735_ (_29574_, _29573_, _05732_);
  or _79736_ (_29575_, _29574_, _29572_);
  nand _79737_ (_29576_, _15457_, _05732_);
  and _79738_ (_29577_, _29576_, _06306_);
  and _79739_ (_29579_, _29577_, _29575_);
  or _79740_ (_29580_, _12020_, _12722_);
  nand _79741_ (_29581_, _29409_, _12722_);
  and _79742_ (_29582_, _29581_, _06129_);
  and _79743_ (_29583_, _29582_, _29580_);
  or _79744_ (_29584_, _29583_, _12541_);
  or _79745_ (_29585_, _29584_, _29579_);
  or _79746_ (_29586_, _29345_, _11872_);
  and _79747_ (_29587_, _29586_, _10975_);
  and _79748_ (_29588_, _29587_, _29585_);
  nor _79749_ (_29590_, _15457_, _10975_);
  or _79750_ (_29591_, _29590_, _11015_);
  or _79751_ (_29592_, _29591_, _29588_);
  and _79752_ (_29593_, _29592_, _29348_);
  or _79753_ (_29594_, _29593_, _06049_);
  nand _79754_ (_29595_, _07883_, _06049_);
  and _79755_ (_29596_, _29595_, _05748_);
  and _79756_ (_29597_, _29596_, _29594_);
  and _79757_ (_29598_, _11875_, _05747_);
  or _79758_ (_29599_, _29598_, _06126_);
  or _79759_ (_29601_, _29599_, _29597_);
  and _79760_ (_29602_, _12021_, _12722_);
  nor _79761_ (_29603_, _29383_, _12722_);
  nor _79762_ (_29604_, _29603_, _29602_);
  or _79763_ (_29605_, _29604_, _06704_);
  and _79764_ (_29606_, _29605_, _29601_);
  nor _79765_ (_29607_, _29606_, _12750_);
  nor _79766_ (_29608_, _29345_, _12749_);
  nor _79767_ (_29609_, _29608_, _29607_);
  nor _79768_ (_29610_, _29609_, _06316_);
  nand _79769_ (_29612_, _15457_, _06316_);
  and _79770_ (_29613_, _29612_, _12756_);
  not _79771_ (_29614_, _29613_);
  nor _79772_ (_29615_, _29614_, _29610_);
  nor _79773_ (_29616_, _29346_, _12756_);
  nor _79774_ (_29617_, _29616_, _06127_);
  not _79775_ (_29618_, _29617_);
  nor _79776_ (_29619_, _29618_, _29615_);
  and _79777_ (_29620_, _06127_, _06084_);
  or _79778_ (_29621_, _29620_, _05752_);
  nor _79779_ (_29623_, _29621_, _29619_);
  and _79780_ (_29624_, _11875_, _05752_);
  or _79781_ (_29625_, _29624_, _05652_);
  nor _79782_ (_29626_, _29625_, _29623_);
  nor _79783_ (_29627_, _29604_, _05653_);
  nor _79784_ (_29628_, _29627_, _12772_);
  not _79785_ (_29629_, _29628_);
  nor _79786_ (_29630_, _29629_, _29626_);
  nor _79787_ (_29631_, _29346_, _12771_);
  nor _79788_ (_29632_, _29631_, _06047_);
  not _79789_ (_29634_, _29632_);
  nor _79790_ (_29635_, _29634_, _29630_);
  or _79791_ (_29636_, _29635_, _26405_);
  nor _79792_ (_29637_, _29636_, _29343_);
  nor _79793_ (_29638_, _29346_, _12779_);
  or _79794_ (_29639_, _29638_, _29637_);
  and _79795_ (_29640_, _29639_, _12782_);
  nor _79796_ (_29641_, _12782_, _06084_);
  or _79797_ (_29642_, _29641_, _29640_);
  and _79798_ (_29643_, _29642_, _12791_);
  and _79799_ (_29645_, _11875_, _05751_);
  or _79800_ (_29646_, _29645_, _29643_);
  and _79801_ (_29647_, _29646_, _12790_);
  and _79802_ (_29648_, _29345_, _12789_);
  or _79803_ (_29649_, _29648_, _29647_);
  or _79804_ (_29650_, _29649_, _01340_);
  or _79805_ (_29651_, _01336_, \oc8051_golden_model_1.PC [14]);
  and _79806_ (_29652_, _29651_, _42882_);
  and _79807_ (_43432_, _29652_, _29650_);
  nor _79808_ (_29653_, \oc8051_golden_model_1.P2 [0], rst);
  nor _79809_ (_29655_, _29653_, _00000_);
  and _79810_ (_29656_, _12800_, \oc8051_golden_model_1.P2 [0]);
  and _79811_ (_29657_, _07686_, _08672_);
  or _79812_ (_29658_, _29657_, _29656_);
  or _79813_ (_29659_, _29658_, _06020_);
  and _79814_ (_29660_, _09120_, _07686_);
  or _79815_ (_29661_, _29656_, _07012_);
  or _79816_ (_29662_, _29661_, _29660_);
  nor _79817_ (_29663_, _08127_, _12800_);
  or _79818_ (_29664_, _29663_, _29656_);
  or _79819_ (_29666_, _29664_, _06954_);
  and _79820_ (_29667_, _07686_, \oc8051_golden_model_1.ACC [0]);
  or _79821_ (_29668_, _29667_, _29656_);
  and _79822_ (_29669_, _29668_, _06938_);
  and _79823_ (_29670_, _06939_, \oc8051_golden_model_1.P2 [0]);
  or _79824_ (_29671_, _29670_, _06102_);
  or _79825_ (_29672_, _29671_, _29669_);
  and _79826_ (_29673_, _29672_, _06044_);
  and _79827_ (_29674_, _29673_, _29666_);
  and _79828_ (_29675_, _12819_, \oc8051_golden_model_1.P2 [0]);
  and _79829_ (_29677_, _14102_, _08349_);
  or _79830_ (_29678_, _29677_, _29675_);
  and _79831_ (_29679_, _29678_, _06043_);
  or _79832_ (_29680_, _29679_, _29674_);
  and _79833_ (_29681_, _29680_, _06848_);
  and _79834_ (_29682_, _07686_, _06931_);
  or _79835_ (_29683_, _29682_, _29656_);
  and _79836_ (_29684_, _29683_, _06239_);
  or _79837_ (_29685_, _29684_, _06219_);
  or _79838_ (_29686_, _29685_, _29681_);
  or _79839_ (_29688_, _29668_, _06220_);
  and _79840_ (_29689_, _29688_, _06040_);
  and _79841_ (_29690_, _29689_, _29686_);
  and _79842_ (_29691_, _29656_, _06039_);
  or _79843_ (_29692_, _29691_, _06032_);
  or _79844_ (_29693_, _29692_, _29690_);
  or _79845_ (_29694_, _29664_, _06033_);
  and _79846_ (_29695_, _29694_, _06027_);
  and _79847_ (_29696_, _29695_, _29693_);
  or _79848_ (_29697_, _29675_, _14131_);
  and _79849_ (_29699_, _29697_, _06026_);
  and _79850_ (_29700_, _29699_, _29678_);
  or _79851_ (_29701_, _29700_, _09818_);
  or _79852_ (_29702_, _29701_, _29696_);
  or _79853_ (_29703_, _29683_, _09827_);
  and _79854_ (_29704_, _29703_, _05669_);
  and _79855_ (_29705_, _29704_, _29702_);
  and _79856_ (_29706_, _29705_, _29662_);
  and _79857_ (_29707_, _14186_, _07686_);
  or _79858_ (_29708_, _29707_, _29656_);
  and _79859_ (_29710_, _29708_, _09833_);
  or _79860_ (_29711_, _29710_, _06019_);
  or _79861_ (_29712_, _29711_, _29706_);
  and _79862_ (_29713_, _29712_, _29659_);
  or _79863_ (_29714_, _29713_, _06112_);
  and _79864_ (_29715_, _14086_, _07686_);
  or _79865_ (_29716_, _29656_, _08751_);
  or _79866_ (_29717_, _29716_, _29715_);
  and _79867_ (_29718_, _29717_, _08756_);
  and _79868_ (_29719_, _29718_, _29714_);
  nor _79869_ (_29721_, _12302_, _12800_);
  or _79870_ (_29722_, _29721_, _29656_);
  nand _79871_ (_29723_, _10995_, _07686_);
  and _79872_ (_29724_, _29723_, _06284_);
  and _79873_ (_29725_, _29724_, _29722_);
  or _79874_ (_29726_, _29725_, _29719_);
  and _79875_ (_29727_, _29726_, _07032_);
  nand _79876_ (_29728_, _29658_, _06108_);
  nor _79877_ (_29729_, _29728_, _29663_);
  or _79878_ (_29730_, _29729_, _06277_);
  or _79879_ (_29732_, _29730_, _29727_);
  nor _79880_ (_29733_, _29656_, _06278_);
  nand _79881_ (_29734_, _29733_, _29723_);
  and _79882_ (_29735_, _29734_, _29732_);
  or _79883_ (_29736_, _29735_, _06130_);
  and _79884_ (_29737_, _14083_, _07686_);
  or _79885_ (_29738_, _29656_, _08777_);
  or _79886_ (_29739_, _29738_, _29737_);
  and _79887_ (_29740_, _29739_, _08782_);
  and _79888_ (_29741_, _29740_, _29736_);
  and _79889_ (_29743_, _29722_, _06292_);
  or _79890_ (_29744_, _29743_, _06316_);
  or _79891_ (_29745_, _29744_, _29741_);
  or _79892_ (_29746_, _29664_, _06718_);
  and _79893_ (_29747_, _29746_, _29745_);
  or _79894_ (_29748_, _29747_, _05652_);
  or _79895_ (_29749_, _29656_, _05653_);
  and _79896_ (_29750_, _29749_, _29748_);
  or _79897_ (_29751_, _29750_, _06047_);
  or _79898_ (_29752_, _29664_, _06048_);
  and _79899_ (_29754_, _29752_, _01336_);
  and _79900_ (_29755_, _29754_, _29751_);
  or _79901_ (_43434_, _29755_, _29655_);
  nor _79902_ (_29756_, \oc8051_golden_model_1.P2 [1], rst);
  nor _79903_ (_29757_, _29756_, _00000_);
  and _79904_ (_29758_, _12800_, \oc8051_golden_model_1.P2 [1]);
  nor _79905_ (_29759_, _10993_, _12800_);
  or _79906_ (_29760_, _29759_, _29758_);
  or _79907_ (_29761_, _29760_, _08782_);
  nor _79908_ (_29762_, _12800_, _07132_);
  or _79909_ (_29764_, _29762_, _29758_);
  or _79910_ (_29765_, _29764_, _06848_);
  or _79911_ (_29766_, _07686_, \oc8051_golden_model_1.P2 [1]);
  and _79912_ (_29767_, _14284_, _07686_);
  not _79913_ (_29768_, _29767_);
  and _79914_ (_29769_, _29768_, _29766_);
  or _79915_ (_29770_, _29769_, _06954_);
  and _79916_ (_29771_, _07686_, \oc8051_golden_model_1.ACC [1]);
  or _79917_ (_29772_, _29771_, _29758_);
  and _79918_ (_29773_, _29772_, _06938_);
  and _79919_ (_29775_, _06939_, \oc8051_golden_model_1.P2 [1]);
  or _79920_ (_29776_, _29775_, _06102_);
  or _79921_ (_29777_, _29776_, _29773_);
  and _79922_ (_29778_, _29777_, _06044_);
  and _79923_ (_29779_, _29778_, _29770_);
  and _79924_ (_29780_, _12819_, \oc8051_golden_model_1.P2 [1]);
  and _79925_ (_29781_, _14266_, _08349_);
  or _79926_ (_29782_, _29781_, _29780_);
  and _79927_ (_29783_, _29782_, _06043_);
  or _79928_ (_29784_, _29783_, _06239_);
  or _79929_ (_29786_, _29784_, _29779_);
  and _79930_ (_29787_, _29786_, _29765_);
  or _79931_ (_29788_, _29787_, _06219_);
  or _79932_ (_29789_, _29772_, _06220_);
  and _79933_ (_29790_, _29789_, _06040_);
  and _79934_ (_29791_, _29790_, _29788_);
  and _79935_ (_29792_, _14273_, _08349_);
  or _79936_ (_29793_, _29792_, _29780_);
  and _79937_ (_29794_, _29793_, _06039_);
  or _79938_ (_29795_, _29794_, _06032_);
  or _79939_ (_29796_, _29795_, _29791_);
  and _79940_ (_29797_, _29781_, _14302_);
  or _79941_ (_29798_, _29780_, _06033_);
  or _79942_ (_29799_, _29798_, _29797_);
  and _79943_ (_29800_, _29799_, _06027_);
  and _79944_ (_29801_, _29800_, _29796_);
  or _79945_ (_29802_, _29780_, _14267_);
  and _79946_ (_29803_, _29802_, _06026_);
  and _79947_ (_29804_, _29803_, _29782_);
  or _79948_ (_29805_, _29804_, _09818_);
  or _79949_ (_29808_, _29805_, _29801_);
  and _79950_ (_29809_, _09075_, _07686_);
  or _79951_ (_29810_, _29758_, _07012_);
  or _79952_ (_29811_, _29810_, _29809_);
  or _79953_ (_29812_, _29764_, _09827_);
  and _79954_ (_29813_, _29812_, _05669_);
  and _79955_ (_29814_, _29813_, _29811_);
  and _79956_ (_29815_, _29814_, _29808_);
  and _79957_ (_29816_, _14367_, _07686_);
  or _79958_ (_29817_, _29816_, _29758_);
  and _79959_ (_29819_, _29817_, _09833_);
  or _79960_ (_29820_, _29819_, _29815_);
  and _79961_ (_29821_, _29820_, _06020_);
  nand _79962_ (_29822_, _07686_, _06832_);
  and _79963_ (_29823_, _29766_, _06019_);
  and _79964_ (_29824_, _29823_, _29822_);
  or _79965_ (_29825_, _29824_, _29821_);
  and _79966_ (_29826_, _29825_, _08751_);
  or _79967_ (_29827_, _14263_, _12800_);
  and _79968_ (_29828_, _29766_, _06112_);
  and _79969_ (_29830_, _29828_, _29827_);
  or _79970_ (_29831_, _29830_, _06284_);
  or _79971_ (_29832_, _29831_, _29826_);
  nand _79972_ (_29833_, _10992_, _07686_);
  and _79973_ (_29834_, _29833_, _29760_);
  or _79974_ (_29835_, _29834_, _08756_);
  and _79975_ (_29836_, _29835_, _07032_);
  and _79976_ (_29837_, _29836_, _29832_);
  or _79977_ (_29838_, _14261_, _12800_);
  and _79978_ (_29839_, _29766_, _06108_);
  and _79979_ (_29841_, _29839_, _29838_);
  or _79980_ (_29842_, _29841_, _06277_);
  or _79981_ (_29843_, _29842_, _29837_);
  nor _79982_ (_29844_, _29758_, _06278_);
  nand _79983_ (_29845_, _29844_, _29833_);
  and _79984_ (_29846_, _29845_, _08777_);
  and _79985_ (_29847_, _29846_, _29843_);
  or _79986_ (_29848_, _29822_, _08078_);
  and _79987_ (_29849_, _29766_, _06130_);
  and _79988_ (_29850_, _29849_, _29848_);
  or _79989_ (_29852_, _29850_, _06292_);
  or _79990_ (_29853_, _29852_, _29847_);
  and _79991_ (_29854_, _29853_, _29761_);
  or _79992_ (_29855_, _29854_, _06316_);
  or _79993_ (_29856_, _29769_, _06718_);
  and _79994_ (_29857_, _29856_, _05653_);
  and _79995_ (_29858_, _29857_, _29855_);
  and _79996_ (_29859_, _29793_, _05652_);
  or _79997_ (_29860_, _29859_, _06047_);
  or _79998_ (_29861_, _29860_, _29858_);
  or _79999_ (_29863_, _29758_, _06048_);
  or _80000_ (_29864_, _29863_, _29767_);
  and _80001_ (_29865_, _29864_, _01336_);
  and _80002_ (_29866_, _29865_, _29861_);
  or _80003_ (_43435_, _29866_, _29757_);
  nor _80004_ (_29867_, \oc8051_golden_model_1.P2 [2], rst);
  nor _80005_ (_29868_, _29867_, _00000_);
  and _80006_ (_29869_, _12800_, \oc8051_golden_model_1.P2 [2]);
  or _80007_ (_29870_, _29869_, _08177_);
  and _80008_ (_29871_, _07686_, _08730_);
  or _80009_ (_29873_, _29871_, _29869_);
  and _80010_ (_29874_, _29873_, _06108_);
  and _80011_ (_29875_, _29874_, _29870_);
  or _80012_ (_29876_, _29873_, _06020_);
  nor _80013_ (_29877_, _12800_, _07530_);
  or _80014_ (_29878_, _29877_, _29869_);
  or _80015_ (_29879_, _29878_, _06848_);
  and _80016_ (_29880_, _14493_, _07686_);
  or _80017_ (_29881_, _29880_, _29869_);
  or _80018_ (_29882_, _29881_, _06954_);
  and _80019_ (_29884_, _07686_, \oc8051_golden_model_1.ACC [2]);
  or _80020_ (_29885_, _29884_, _29869_);
  and _80021_ (_29886_, _29885_, _06938_);
  and _80022_ (_29887_, _06939_, \oc8051_golden_model_1.P2 [2]);
  or _80023_ (_29888_, _29887_, _06102_);
  or _80024_ (_29889_, _29888_, _29886_);
  and _80025_ (_29890_, _29889_, _06044_);
  and _80026_ (_29891_, _29890_, _29882_);
  and _80027_ (_29892_, _12819_, \oc8051_golden_model_1.P2 [2]);
  and _80028_ (_29893_, _14497_, _08349_);
  or _80029_ (_29895_, _29893_, _29892_);
  and _80030_ (_29896_, _29895_, _06043_);
  or _80031_ (_29897_, _29896_, _06239_);
  or _80032_ (_29898_, _29897_, _29891_);
  and _80033_ (_29899_, _29898_, _29879_);
  or _80034_ (_29900_, _29899_, _06219_);
  or _80035_ (_29901_, _29885_, _06220_);
  and _80036_ (_29902_, _29901_, _06040_);
  and _80037_ (_29903_, _29902_, _29900_);
  and _80038_ (_29904_, _14479_, _08349_);
  or _80039_ (_29906_, _29904_, _29892_);
  and _80040_ (_29907_, _29906_, _06039_);
  or _80041_ (_29908_, _29907_, _06032_);
  or _80042_ (_29909_, _29908_, _29903_);
  and _80043_ (_29910_, _29893_, _14512_);
  or _80044_ (_29911_, _29892_, _06033_);
  or _80045_ (_29912_, _29911_, _29910_);
  and _80046_ (_29913_, _29912_, _06027_);
  and _80047_ (_29914_, _29913_, _29909_);
  or _80048_ (_29915_, _29892_, _14525_);
  and _80049_ (_29917_, _29915_, _06026_);
  and _80050_ (_29918_, _29917_, _29895_);
  or _80051_ (_29919_, _29918_, _09818_);
  or _80052_ (_29920_, _29919_, _29914_);
  and _80053_ (_29921_, _09182_, _07686_);
  or _80054_ (_29922_, _29869_, _07012_);
  or _80055_ (_29923_, _29922_, _29921_);
  or _80056_ (_29924_, _29878_, _09827_);
  and _80057_ (_29925_, _29924_, _05669_);
  and _80058_ (_29926_, _29925_, _29923_);
  and _80059_ (_29928_, _29926_, _29920_);
  and _80060_ (_29929_, _14580_, _07686_);
  or _80061_ (_29930_, _29929_, _29869_);
  and _80062_ (_29931_, _29930_, _09833_);
  or _80063_ (_29932_, _29931_, _06019_);
  or _80064_ (_29933_, _29932_, _29928_);
  and _80065_ (_29934_, _29933_, _29876_);
  or _80066_ (_29935_, _29934_, _06112_);
  and _80067_ (_29936_, _14596_, _07686_);
  or _80068_ (_29937_, _29936_, _29869_);
  or _80069_ (_29939_, _29937_, _08751_);
  and _80070_ (_29940_, _29939_, _08756_);
  and _80071_ (_29941_, _29940_, _29935_);
  and _80072_ (_29942_, _10991_, _07686_);
  or _80073_ (_29943_, _29942_, _29869_);
  and _80074_ (_29944_, _29943_, _06284_);
  or _80075_ (_29945_, _29944_, _29941_);
  and _80076_ (_29946_, _29945_, _07032_);
  or _80077_ (_29947_, _29946_, _29875_);
  and _80078_ (_29948_, _29947_, _06278_);
  and _80079_ (_29950_, _29885_, _06277_);
  and _80080_ (_29951_, _29950_, _29870_);
  or _80081_ (_29952_, _29951_, _06130_);
  or _80082_ (_29953_, _29952_, _29948_);
  and _80083_ (_29954_, _14593_, _07686_);
  or _80084_ (_29955_, _29869_, _08777_);
  or _80085_ (_29956_, _29955_, _29954_);
  and _80086_ (_29957_, _29956_, _08782_);
  and _80087_ (_29958_, _29957_, _29953_);
  nor _80088_ (_29959_, _10990_, _12800_);
  or _80089_ (_29961_, _29959_, _29869_);
  and _80090_ (_29962_, _29961_, _06292_);
  or _80091_ (_29963_, _29962_, _06316_);
  or _80092_ (_29964_, _29963_, _29958_);
  or _80093_ (_29965_, _29881_, _06718_);
  and _80094_ (_29966_, _29965_, _05653_);
  and _80095_ (_29967_, _29966_, _29964_);
  and _80096_ (_29968_, _29906_, _05652_);
  or _80097_ (_29969_, _29968_, _06047_);
  or _80098_ (_29970_, _29969_, _29967_);
  and _80099_ (_29972_, _14657_, _07686_);
  or _80100_ (_29973_, _29869_, _06048_);
  or _80101_ (_29974_, _29973_, _29972_);
  and _80102_ (_29975_, _29974_, _01336_);
  and _80103_ (_29976_, _29975_, _29970_);
  or _80104_ (_43436_, _29976_, _29868_);
  and _80105_ (_29977_, _12800_, \oc8051_golden_model_1.P2 [3]);
  and _80106_ (_29978_, _07686_, _08662_);
  or _80107_ (_29979_, _29978_, _29977_);
  or _80108_ (_29980_, _29979_, _06020_);
  and _80109_ (_29982_, _14672_, _07686_);
  or _80110_ (_29983_, _29982_, _29977_);
  or _80111_ (_29984_, _29983_, _06954_);
  and _80112_ (_29985_, _07686_, \oc8051_golden_model_1.ACC [3]);
  or _80113_ (_29986_, _29985_, _29977_);
  and _80114_ (_29987_, _29986_, _06938_);
  and _80115_ (_29988_, _06939_, \oc8051_golden_model_1.P2 [3]);
  or _80116_ (_29989_, _29988_, _06102_);
  or _80117_ (_29990_, _29989_, _29987_);
  and _80118_ (_29991_, _29990_, _06044_);
  and _80119_ (_29993_, _29991_, _29984_);
  and _80120_ (_29994_, _12819_, \oc8051_golden_model_1.P2 [3]);
  and _80121_ (_29995_, _14683_, _08349_);
  or _80122_ (_29996_, _29995_, _29994_);
  and _80123_ (_29997_, _29996_, _06043_);
  or _80124_ (_29998_, _29997_, _06239_);
  or _80125_ (_29999_, _29998_, _29993_);
  nor _80126_ (_30000_, _12800_, _07353_);
  or _80127_ (_30001_, _30000_, _29977_);
  or _80128_ (_30002_, _30001_, _06848_);
  and _80129_ (_30004_, _30002_, _29999_);
  or _80130_ (_30005_, _30004_, _06219_);
  or _80131_ (_30006_, _29986_, _06220_);
  and _80132_ (_30007_, _30006_, _06040_);
  and _80133_ (_30008_, _30007_, _30005_);
  and _80134_ (_30009_, _14681_, _08349_);
  or _80135_ (_30010_, _30009_, _29994_);
  and _80136_ (_30011_, _30010_, _06039_);
  or _80137_ (_30012_, _30011_, _06032_);
  or _80138_ (_30013_, _30012_, _30008_);
  or _80139_ (_30015_, _29994_, _14708_);
  and _80140_ (_30016_, _30015_, _29996_);
  or _80141_ (_30017_, _30016_, _06033_);
  and _80142_ (_30018_, _30017_, _06027_);
  and _80143_ (_30019_, _30018_, _30013_);
  and _80144_ (_30020_, _14724_, _08349_);
  or _80145_ (_30021_, _30020_, _29994_);
  and _80146_ (_30022_, _30021_, _06026_);
  or _80147_ (_30023_, _30022_, _09818_);
  or _80148_ (_30024_, _30023_, _30019_);
  and _80149_ (_30026_, _09181_, _07686_);
  or _80150_ (_30027_, _29977_, _07012_);
  or _80151_ (_30028_, _30027_, _30026_);
  or _80152_ (_30029_, _30001_, _09827_);
  and _80153_ (_30030_, _30029_, _05669_);
  and _80154_ (_30031_, _30030_, _30028_);
  and _80155_ (_30032_, _30031_, _30024_);
  and _80156_ (_30033_, _14778_, _07686_);
  or _80157_ (_30034_, _30033_, _29977_);
  and _80158_ (_30035_, _30034_, _09833_);
  or _80159_ (_30037_, _30035_, _06019_);
  or _80160_ (_30038_, _30037_, _30032_);
  and _80161_ (_30039_, _30038_, _29980_);
  or _80162_ (_30040_, _30039_, _06112_);
  and _80163_ (_30041_, _14793_, _07686_);
  or _80164_ (_30042_, _29977_, _08751_);
  or _80165_ (_30043_, _30042_, _30041_);
  and _80166_ (_30044_, _30043_, _08756_);
  and _80167_ (_30045_, _30044_, _30040_);
  and _80168_ (_30046_, _12299_, _07686_);
  or _80169_ (_30048_, _30046_, _29977_);
  and _80170_ (_30049_, _30048_, _06284_);
  or _80171_ (_30050_, _30049_, _30045_);
  and _80172_ (_30051_, _30050_, _07032_);
  or _80173_ (_30052_, _29977_, _08029_);
  and _80174_ (_30053_, _29979_, _06108_);
  and _80175_ (_30054_, _30053_, _30052_);
  or _80176_ (_30055_, _30054_, _30051_);
  and _80177_ (_30056_, _30055_, _06278_);
  and _80178_ (_30057_, _29986_, _06277_);
  and _80179_ (_30059_, _30057_, _30052_);
  or _80180_ (_30060_, _30059_, _06130_);
  or _80181_ (_30061_, _30060_, _30056_);
  and _80182_ (_30062_, _14792_, _07686_);
  or _80183_ (_30063_, _29977_, _08777_);
  or _80184_ (_30064_, _30063_, _30062_);
  and _80185_ (_30065_, _30064_, _08782_);
  and _80186_ (_30066_, _30065_, _30061_);
  nor _80187_ (_30067_, _10988_, _12800_);
  or _80188_ (_30068_, _30067_, _29977_);
  and _80189_ (_30070_, _30068_, _06292_);
  or _80190_ (_30071_, _30070_, _06316_);
  or _80191_ (_30072_, _30071_, _30066_);
  or _80192_ (_30073_, _29983_, _06718_);
  and _80193_ (_30074_, _30073_, _05653_);
  and _80194_ (_30075_, _30074_, _30072_);
  and _80195_ (_30076_, _30010_, _05652_);
  or _80196_ (_30077_, _30076_, _06047_);
  or _80197_ (_30078_, _30077_, _30075_);
  and _80198_ (_30079_, _14849_, _07686_);
  or _80199_ (_30081_, _29977_, _06048_);
  or _80200_ (_30082_, _30081_, _30079_);
  and _80201_ (_30083_, _30082_, _01336_);
  and _80202_ (_30084_, _30083_, _30078_);
  nor _80203_ (_30085_, \oc8051_golden_model_1.P2 [3], rst);
  nor _80204_ (_30086_, _30085_, _00000_);
  or _80205_ (_43437_, _30086_, _30084_);
  and _80206_ (_30087_, _12800_, \oc8051_golden_model_1.P2 [4]);
  and _80207_ (_30088_, _08665_, _07686_);
  or _80208_ (_30089_, _30088_, _30087_);
  or _80209_ (_30091_, _30089_, _06020_);
  and _80210_ (_30092_, _14887_, _07686_);
  or _80211_ (_30093_, _30092_, _30087_);
  or _80212_ (_30094_, _30093_, _06954_);
  and _80213_ (_30095_, _07686_, \oc8051_golden_model_1.ACC [4]);
  or _80214_ (_30096_, _30095_, _30087_);
  and _80215_ (_30097_, _30096_, _06938_);
  and _80216_ (_30098_, _06939_, \oc8051_golden_model_1.P2 [4]);
  or _80217_ (_30099_, _30098_, _06102_);
  or _80218_ (_30100_, _30099_, _30097_);
  and _80219_ (_30102_, _30100_, _06044_);
  and _80220_ (_30103_, _30102_, _30094_);
  and _80221_ (_30104_, _12819_, \oc8051_golden_model_1.P2 [4]);
  and _80222_ (_30105_, _14878_, _08349_);
  or _80223_ (_30106_, _30105_, _30104_);
  and _80224_ (_30107_, _30106_, _06043_);
  or _80225_ (_30108_, _30107_, _06239_);
  or _80226_ (_30109_, _30108_, _30103_);
  nor _80227_ (_30110_, _08270_, _12800_);
  or _80228_ (_30111_, _30110_, _30087_);
  or _80229_ (_30113_, _30111_, _06848_);
  and _80230_ (_30114_, _30113_, _30109_);
  or _80231_ (_30115_, _30114_, _06219_);
  or _80232_ (_30116_, _30096_, _06220_);
  and _80233_ (_30117_, _30116_, _06040_);
  and _80234_ (_30118_, _30117_, _30115_);
  and _80235_ (_30119_, _14882_, _08349_);
  or _80236_ (_30120_, _30119_, _30104_);
  and _80237_ (_30121_, _30120_, _06039_);
  or _80238_ (_30122_, _30121_, _06032_);
  or _80239_ (_30124_, _30122_, _30118_);
  or _80240_ (_30125_, _30104_, _14914_);
  and _80241_ (_30126_, _30125_, _30106_);
  or _80242_ (_30127_, _30126_, _06033_);
  and _80243_ (_30128_, _30127_, _06027_);
  and _80244_ (_30129_, _30128_, _30124_);
  or _80245_ (_30130_, _30104_, _14879_);
  and _80246_ (_30131_, _30130_, _06026_);
  and _80247_ (_30132_, _30131_, _30106_);
  or _80248_ (_30133_, _30132_, _09818_);
  or _80249_ (_30135_, _30133_, _30129_);
  and _80250_ (_30136_, _09180_, _07686_);
  or _80251_ (_30137_, _30087_, _07012_);
  or _80252_ (_30138_, _30137_, _30136_);
  or _80253_ (_30139_, _30111_, _09827_);
  and _80254_ (_30140_, _30139_, _05669_);
  and _80255_ (_30141_, _30140_, _30138_);
  and _80256_ (_30142_, _30141_, _30135_);
  and _80257_ (_30143_, _14983_, _07686_);
  or _80258_ (_30144_, _30143_, _30087_);
  and _80259_ (_30146_, _30144_, _09833_);
  or _80260_ (_30147_, _30146_, _06019_);
  or _80261_ (_30148_, _30147_, _30142_);
  and _80262_ (_30149_, _30148_, _30091_);
  or _80263_ (_30150_, _30149_, _06112_);
  and _80264_ (_30151_, _14876_, _07686_);
  or _80265_ (_30152_, _30087_, _08751_);
  or _80266_ (_30153_, _30152_, _30151_);
  and _80267_ (_30154_, _30153_, _08756_);
  and _80268_ (_30155_, _30154_, _30150_);
  and _80269_ (_30157_, _10986_, _07686_);
  or _80270_ (_30158_, _30157_, _30087_);
  and _80271_ (_30159_, _30158_, _06284_);
  or _80272_ (_30160_, _30159_, _30155_);
  and _80273_ (_30161_, _30160_, _07032_);
  or _80274_ (_30162_, _30087_, _08273_);
  and _80275_ (_30163_, _30089_, _06108_);
  and _80276_ (_30164_, _30163_, _30162_);
  or _80277_ (_30165_, _30164_, _30161_);
  and _80278_ (_30166_, _30165_, _06278_);
  and _80279_ (_30168_, _30096_, _06277_);
  and _80280_ (_30169_, _30168_, _30162_);
  or _80281_ (_30170_, _30169_, _06130_);
  or _80282_ (_30171_, _30170_, _30166_);
  and _80283_ (_30172_, _14873_, _07686_);
  or _80284_ (_30173_, _30087_, _08777_);
  or _80285_ (_30174_, _30173_, _30172_);
  and _80286_ (_30175_, _30174_, _08782_);
  and _80287_ (_30176_, _30175_, _30171_);
  nor _80288_ (_30177_, _10985_, _12800_);
  or _80289_ (_30179_, _30177_, _30087_);
  and _80290_ (_30180_, _30179_, _06292_);
  or _80291_ (_30181_, _30180_, _06316_);
  or _80292_ (_30182_, _30181_, _30176_);
  or _80293_ (_30183_, _30093_, _06718_);
  and _80294_ (_30184_, _30183_, _05653_);
  and _80295_ (_30185_, _30184_, _30182_);
  and _80296_ (_30186_, _30120_, _05652_);
  or _80297_ (_30187_, _30186_, _06047_);
  or _80298_ (_30188_, _30187_, _30185_);
  and _80299_ (_30190_, _15055_, _07686_);
  or _80300_ (_30191_, _30087_, _06048_);
  or _80301_ (_30192_, _30191_, _30190_);
  and _80302_ (_30193_, _30192_, _01336_);
  and _80303_ (_30194_, _30193_, _30188_);
  nor _80304_ (_30195_, \oc8051_golden_model_1.P2 [4], rst);
  nor _80305_ (_30196_, _30195_, _00000_);
  or _80306_ (_43438_, _30196_, _30194_);
  and _80307_ (_30197_, _12800_, \oc8051_golden_model_1.P2 [5]);
  and _80308_ (_30198_, _08652_, _07686_);
  or _80309_ (_30200_, _30198_, _30197_);
  or _80310_ (_30201_, _30200_, _06020_);
  and _80311_ (_30202_, _15093_, _07686_);
  or _80312_ (_30203_, _30202_, _30197_);
  or _80313_ (_30204_, _30203_, _06954_);
  and _80314_ (_30205_, _07686_, \oc8051_golden_model_1.ACC [5]);
  or _80315_ (_30206_, _30205_, _30197_);
  and _80316_ (_30207_, _30206_, _06938_);
  and _80317_ (_30208_, _06939_, \oc8051_golden_model_1.P2 [5]);
  or _80318_ (_30209_, _30208_, _06102_);
  or _80319_ (_30211_, _30209_, _30207_);
  and _80320_ (_30212_, _30211_, _06044_);
  and _80321_ (_30213_, _30212_, _30204_);
  and _80322_ (_30214_, _12819_, \oc8051_golden_model_1.P2 [5]);
  and _80323_ (_30215_, _15073_, _08349_);
  or _80324_ (_30216_, _30215_, _30214_);
  and _80325_ (_30217_, _30216_, _06043_);
  or _80326_ (_30218_, _30217_, _06239_);
  or _80327_ (_30219_, _30218_, _30213_);
  nor _80328_ (_30220_, _07977_, _12800_);
  or _80329_ (_30222_, _30220_, _30197_);
  or _80330_ (_30223_, _30222_, _06848_);
  and _80331_ (_30224_, _30223_, _30219_);
  or _80332_ (_30225_, _30224_, _06219_);
  or _80333_ (_30226_, _30206_, _06220_);
  and _80334_ (_30227_, _30226_, _06040_);
  and _80335_ (_30228_, _30227_, _30225_);
  and _80336_ (_30229_, _15077_, _08349_);
  or _80337_ (_30230_, _30229_, _30214_);
  and _80338_ (_30231_, _30230_, _06039_);
  or _80339_ (_30233_, _30231_, _06032_);
  or _80340_ (_30234_, _30233_, _30228_);
  or _80341_ (_30235_, _30214_, _15110_);
  and _80342_ (_30236_, _30235_, _30216_);
  or _80343_ (_30237_, _30236_, _06033_);
  and _80344_ (_30238_, _30237_, _06027_);
  and _80345_ (_30239_, _30238_, _30234_);
  or _80346_ (_30240_, _30214_, _15074_);
  and _80347_ (_30241_, _30240_, _06026_);
  and _80348_ (_30242_, _30241_, _30216_);
  or _80349_ (_30244_, _30242_, _09818_);
  or _80350_ (_30245_, _30244_, _30239_);
  and _80351_ (_30246_, _09179_, _07686_);
  or _80352_ (_30247_, _30197_, _07012_);
  or _80353_ (_30248_, _30247_, _30246_);
  or _80354_ (_30249_, _30222_, _09827_);
  and _80355_ (_30250_, _30249_, _05669_);
  and _80356_ (_30251_, _30250_, _30248_);
  and _80357_ (_30252_, _30251_, _30245_);
  and _80358_ (_30253_, _15179_, _07686_);
  or _80359_ (_30255_, _30253_, _30197_);
  and _80360_ (_30256_, _30255_, _09833_);
  or _80361_ (_30257_, _30256_, _06019_);
  or _80362_ (_30258_, _30257_, _30252_);
  and _80363_ (_30259_, _30258_, _30201_);
  or _80364_ (_30260_, _30259_, _06112_);
  and _80365_ (_30261_, _15195_, _07686_);
  or _80366_ (_30262_, _30197_, _08751_);
  or _80367_ (_30263_, _30262_, _30261_);
  and _80368_ (_30264_, _30263_, _08756_);
  and _80369_ (_30266_, _30264_, _30260_);
  and _80370_ (_30267_, _12306_, _07686_);
  or _80371_ (_30268_, _30267_, _30197_);
  and _80372_ (_30269_, _30268_, _06284_);
  or _80373_ (_30270_, _30269_, _30266_);
  and _80374_ (_30271_, _30270_, _07032_);
  or _80375_ (_30272_, _30197_, _07980_);
  and _80376_ (_30273_, _30200_, _06108_);
  and _80377_ (_30274_, _30273_, _30272_);
  or _80378_ (_30275_, _30274_, _30271_);
  and _80379_ (_30277_, _30275_, _06278_);
  and _80380_ (_30278_, _30206_, _06277_);
  and _80381_ (_30279_, _30278_, _30272_);
  or _80382_ (_30280_, _30279_, _06130_);
  or _80383_ (_30281_, _30280_, _30277_);
  and _80384_ (_30282_, _15194_, _07686_);
  or _80385_ (_30283_, _30197_, _08777_);
  or _80386_ (_30284_, _30283_, _30282_);
  and _80387_ (_30285_, _30284_, _08782_);
  and _80388_ (_30286_, _30285_, _30281_);
  nor _80389_ (_30288_, _10982_, _12800_);
  or _80390_ (_30289_, _30288_, _30197_);
  and _80391_ (_30290_, _30289_, _06292_);
  or _80392_ (_30291_, _30290_, _06316_);
  or _80393_ (_30292_, _30291_, _30286_);
  or _80394_ (_30293_, _30203_, _06718_);
  and _80395_ (_30294_, _30293_, _05653_);
  and _80396_ (_30295_, _30294_, _30292_);
  and _80397_ (_30296_, _30230_, _05652_);
  or _80398_ (_30297_, _30296_, _06047_);
  or _80399_ (_30299_, _30297_, _30295_);
  and _80400_ (_30300_, _15253_, _07686_);
  or _80401_ (_30301_, _30197_, _06048_);
  or _80402_ (_30302_, _30301_, _30300_);
  and _80403_ (_30303_, _30302_, _01336_);
  and _80404_ (_30304_, _30303_, _30299_);
  nor _80405_ (_30305_, \oc8051_golden_model_1.P2 [5], rst);
  nor _80406_ (_30306_, _30305_, _00000_);
  or _80407_ (_43440_, _30306_, _30304_);
  nor _80408_ (_30307_, \oc8051_golden_model_1.P2 [6], rst);
  nor _80409_ (_30309_, _30307_, _00000_);
  and _80410_ (_30310_, _12800_, \oc8051_golden_model_1.P2 [6]);
  and _80411_ (_30311_, _15389_, _07686_);
  or _80412_ (_30312_, _30311_, _30310_);
  or _80413_ (_30313_, _30312_, _06020_);
  and _80414_ (_30314_, _15293_, _07686_);
  or _80415_ (_30315_, _30314_, _30310_);
  or _80416_ (_30316_, _30315_, _06954_);
  and _80417_ (_30317_, _07686_, \oc8051_golden_model_1.ACC [6]);
  or _80418_ (_30318_, _30317_, _30310_);
  and _80419_ (_30320_, _30318_, _06938_);
  and _80420_ (_30321_, _06939_, \oc8051_golden_model_1.P2 [6]);
  or _80421_ (_30322_, _30321_, _06102_);
  or _80422_ (_30323_, _30322_, _30320_);
  and _80423_ (_30324_, _30323_, _06044_);
  and _80424_ (_30325_, _30324_, _30316_);
  and _80425_ (_30326_, _12819_, \oc8051_golden_model_1.P2 [6]);
  and _80426_ (_30327_, _15280_, _08349_);
  or _80427_ (_30328_, _30327_, _30326_);
  and _80428_ (_30329_, _30328_, _06043_);
  or _80429_ (_30331_, _30329_, _06239_);
  or _80430_ (_30332_, _30331_, _30325_);
  nor _80431_ (_30333_, _07883_, _12800_);
  or _80432_ (_30334_, _30333_, _30310_);
  or _80433_ (_30335_, _30334_, _06848_);
  and _80434_ (_30336_, _30335_, _30332_);
  or _80435_ (_30337_, _30336_, _06219_);
  or _80436_ (_30338_, _30318_, _06220_);
  and _80437_ (_30339_, _30338_, _06040_);
  and _80438_ (_30340_, _30339_, _30337_);
  and _80439_ (_30342_, _15278_, _08349_);
  or _80440_ (_30343_, _30342_, _30326_);
  and _80441_ (_30344_, _30343_, _06039_);
  or _80442_ (_30345_, _30344_, _06032_);
  or _80443_ (_30346_, _30345_, _30340_);
  or _80444_ (_30347_, _30326_, _15310_);
  and _80445_ (_30348_, _30347_, _30328_);
  or _80446_ (_30349_, _30348_, _06033_);
  and _80447_ (_30350_, _30349_, _06027_);
  and _80448_ (_30351_, _30350_, _30346_);
  or _80449_ (_30353_, _30326_, _15326_);
  and _80450_ (_30354_, _30353_, _06026_);
  and _80451_ (_30355_, _30354_, _30328_);
  or _80452_ (_30356_, _30355_, _09818_);
  or _80453_ (_30357_, _30356_, _30351_);
  and _80454_ (_30358_, _09178_, _07686_);
  or _80455_ (_30359_, _30310_, _07012_);
  or _80456_ (_30360_, _30359_, _30358_);
  or _80457_ (_30361_, _30334_, _09827_);
  and _80458_ (_30362_, _30361_, _05669_);
  and _80459_ (_30364_, _30362_, _30360_);
  and _80460_ (_30365_, _30364_, _30357_);
  and _80461_ (_30366_, _15382_, _07686_);
  or _80462_ (_30367_, _30366_, _30310_);
  and _80463_ (_30368_, _30367_, _09833_);
  or _80464_ (_30369_, _30368_, _06019_);
  or _80465_ (_30370_, _30369_, _30365_);
  and _80466_ (_30371_, _30370_, _30313_);
  or _80467_ (_30372_, _30371_, _06112_);
  and _80468_ (_30373_, _15399_, _07686_);
  or _80469_ (_30375_, _30373_, _30310_);
  or _80470_ (_30376_, _30375_, _08751_);
  and _80471_ (_30377_, _30376_, _08756_);
  and _80472_ (_30378_, _30377_, _30372_);
  and _80473_ (_30379_, _10980_, _07686_);
  or _80474_ (_30380_, _30379_, _30310_);
  and _80475_ (_30381_, _30380_, _06284_);
  or _80476_ (_30382_, _30381_, _30378_);
  and _80477_ (_30383_, _30382_, _07032_);
  or _80478_ (_30384_, _30310_, _07886_);
  and _80479_ (_30386_, _30312_, _06108_);
  and _80480_ (_30387_, _30386_, _30384_);
  or _80481_ (_30388_, _30387_, _30383_);
  and _80482_ (_30389_, _30388_, _06278_);
  and _80483_ (_30390_, _30318_, _06277_);
  and _80484_ (_30391_, _30390_, _30384_);
  or _80485_ (_30392_, _30391_, _06130_);
  or _80486_ (_30393_, _30392_, _30389_);
  and _80487_ (_30394_, _15396_, _07686_);
  or _80488_ (_30395_, _30310_, _08777_);
  or _80489_ (_30397_, _30395_, _30394_);
  and _80490_ (_30398_, _30397_, _08782_);
  and _80491_ (_30399_, _30398_, _30393_);
  nor _80492_ (_30400_, _10979_, _12800_);
  or _80493_ (_30401_, _30400_, _30310_);
  and _80494_ (_30402_, _30401_, _06292_);
  or _80495_ (_30403_, _30402_, _06316_);
  or _80496_ (_30404_, _30403_, _30399_);
  or _80497_ (_30405_, _30315_, _06718_);
  and _80498_ (_30406_, _30405_, _05653_);
  and _80499_ (_30408_, _30406_, _30404_);
  and _80500_ (_30409_, _30343_, _05652_);
  or _80501_ (_30410_, _30409_, _06047_);
  or _80502_ (_30411_, _30410_, _30408_);
  and _80503_ (_30412_, _15451_, _07686_);
  or _80504_ (_30413_, _30310_, _06048_);
  or _80505_ (_30414_, _30413_, _30412_);
  and _80506_ (_30415_, _30414_, _01336_);
  and _80507_ (_30416_, _30415_, _30411_);
  or _80508_ (_43441_, _30416_, _30309_);
  nand _80509_ (_30417_, _10995_, _07692_);
  and _80510_ (_30418_, _12902_, \oc8051_golden_model_1.P3 [0]);
  nor _80511_ (_30419_, _30418_, _06278_);
  nand _80512_ (_30420_, _30419_, _30417_);
  and _80513_ (_30421_, _07692_, _08672_);
  or _80514_ (_30422_, _30421_, _30418_);
  or _80515_ (_30423_, _30422_, _06020_);
  and _80516_ (_30424_, _09120_, _07692_);
  or _80517_ (_30425_, _30418_, _07012_);
  or _80518_ (_30426_, _30425_, _30424_);
  nor _80519_ (_30429_, _08127_, _12902_);
  or _80520_ (_30430_, _30429_, _30418_);
  or _80521_ (_30431_, _30430_, _06954_);
  and _80522_ (_30432_, _07692_, \oc8051_golden_model_1.ACC [0]);
  or _80523_ (_30433_, _30432_, _30418_);
  and _80524_ (_30434_, _30433_, _06938_);
  and _80525_ (_30435_, _06939_, \oc8051_golden_model_1.P3 [0]);
  or _80526_ (_30436_, _30435_, _06102_);
  or _80527_ (_30437_, _30436_, _30434_);
  and _80528_ (_30438_, _30437_, _06044_);
  and _80529_ (_30440_, _30438_, _30431_);
  and _80530_ (_30441_, _12921_, \oc8051_golden_model_1.P3 [0]);
  and _80531_ (_30442_, _14102_, _08353_);
  or _80532_ (_30443_, _30442_, _30441_);
  and _80533_ (_30444_, _30443_, _06043_);
  or _80534_ (_30445_, _30444_, _30440_);
  and _80535_ (_30446_, _30445_, _06848_);
  and _80536_ (_30447_, _07692_, _06931_);
  or _80537_ (_30448_, _30447_, _30418_);
  and _80538_ (_30449_, _30448_, _06239_);
  or _80539_ (_30451_, _30449_, _06219_);
  or _80540_ (_30452_, _30451_, _30446_);
  or _80541_ (_30453_, _30433_, _06220_);
  and _80542_ (_30454_, _30453_, _06040_);
  and _80543_ (_30455_, _30454_, _30452_);
  and _80544_ (_30456_, _30418_, _06039_);
  or _80545_ (_30457_, _30456_, _06032_);
  or _80546_ (_30458_, _30457_, _30455_);
  or _80547_ (_30459_, _30430_, _06033_);
  and _80548_ (_30460_, _30459_, _06027_);
  and _80549_ (_30462_, _30460_, _30458_);
  or _80550_ (_30463_, _30441_, _14131_);
  and _80551_ (_30464_, _30463_, _06026_);
  and _80552_ (_30465_, _30464_, _30443_);
  or _80553_ (_30466_, _30465_, _09818_);
  or _80554_ (_30467_, _30466_, _30462_);
  or _80555_ (_30468_, _30448_, _09827_);
  and _80556_ (_30469_, _30468_, _05669_);
  and _80557_ (_30470_, _30469_, _30467_);
  and _80558_ (_30471_, _30470_, _30426_);
  and _80559_ (_30473_, _14186_, _07692_);
  or _80560_ (_30474_, _30473_, _30418_);
  and _80561_ (_30475_, _30474_, _09833_);
  or _80562_ (_30476_, _30475_, _06019_);
  or _80563_ (_30477_, _30476_, _30471_);
  and _80564_ (_30478_, _30477_, _30423_);
  or _80565_ (_30479_, _30478_, _06112_);
  and _80566_ (_30480_, _14086_, _07692_);
  or _80567_ (_30481_, _30418_, _08751_);
  or _80568_ (_30482_, _30481_, _30480_);
  and _80569_ (_30484_, _30482_, _08756_);
  and _80570_ (_30485_, _30484_, _30479_);
  nor _80571_ (_30486_, _12302_, _12902_);
  or _80572_ (_30487_, _30486_, _30418_);
  and _80573_ (_30488_, _30417_, _06284_);
  and _80574_ (_30489_, _30488_, _30487_);
  or _80575_ (_30490_, _30489_, _30485_);
  and _80576_ (_30491_, _30490_, _07032_);
  nand _80577_ (_30492_, _30422_, _06108_);
  nor _80578_ (_30493_, _30492_, _30429_);
  or _80579_ (_30495_, _30493_, _06277_);
  or _80580_ (_30496_, _30495_, _30491_);
  and _80581_ (_30497_, _30496_, _30420_);
  or _80582_ (_30498_, _30497_, _06130_);
  and _80583_ (_30499_, _14083_, _07692_);
  or _80584_ (_30500_, _30418_, _08777_);
  or _80585_ (_30501_, _30500_, _30499_);
  and _80586_ (_30502_, _30501_, _08782_);
  and _80587_ (_30503_, _30502_, _30498_);
  and _80588_ (_30504_, _30487_, _06292_);
  or _80589_ (_30506_, _30504_, _06316_);
  or _80590_ (_30507_, _30506_, _30503_);
  or _80591_ (_30508_, _30430_, _06718_);
  and _80592_ (_30509_, _30508_, _30507_);
  or _80593_ (_30510_, _30509_, _05652_);
  or _80594_ (_30511_, _30418_, _05653_);
  and _80595_ (_30512_, _30511_, _30510_);
  or _80596_ (_30513_, _30512_, _06047_);
  or _80597_ (_30514_, _30430_, _06048_);
  and _80598_ (_30515_, _30514_, _01336_);
  and _80599_ (_30517_, _30515_, _30513_);
  nor _80600_ (_30518_, \oc8051_golden_model_1.P3 [0], rst);
  nor _80601_ (_30519_, _30518_, _00000_);
  or _80602_ (_43442_, _30519_, _30517_);
  and _80603_ (_30520_, _12902_, \oc8051_golden_model_1.P3 [1]);
  nor _80604_ (_30521_, _10993_, _12902_);
  or _80605_ (_30522_, _30521_, _30520_);
  or _80606_ (_30523_, _30522_, _08782_);
  nor _80607_ (_30524_, _12902_, _07132_);
  or _80608_ (_30525_, _30524_, _30520_);
  or _80609_ (_30527_, _30525_, _06848_);
  or _80610_ (_30528_, _07692_, \oc8051_golden_model_1.P3 [1]);
  and _80611_ (_30529_, _14284_, _07692_);
  not _80612_ (_30530_, _30529_);
  and _80613_ (_30531_, _30530_, _30528_);
  or _80614_ (_30532_, _30531_, _06954_);
  and _80615_ (_30533_, _07692_, \oc8051_golden_model_1.ACC [1]);
  or _80616_ (_30534_, _30533_, _30520_);
  and _80617_ (_30535_, _30534_, _06938_);
  and _80618_ (_30536_, _06939_, \oc8051_golden_model_1.P3 [1]);
  or _80619_ (_30538_, _30536_, _06102_);
  or _80620_ (_30539_, _30538_, _30535_);
  and _80621_ (_30540_, _30539_, _06044_);
  and _80622_ (_30541_, _30540_, _30532_);
  and _80623_ (_30542_, _12921_, \oc8051_golden_model_1.P3 [1]);
  and _80624_ (_30543_, _14266_, _08353_);
  or _80625_ (_30544_, _30543_, _30542_);
  and _80626_ (_30545_, _30544_, _06043_);
  or _80627_ (_30546_, _30545_, _06239_);
  or _80628_ (_30547_, _30546_, _30541_);
  and _80629_ (_30549_, _30547_, _30527_);
  or _80630_ (_30550_, _30549_, _06219_);
  or _80631_ (_30551_, _30534_, _06220_);
  and _80632_ (_30552_, _30551_, _06040_);
  and _80633_ (_30553_, _30552_, _30550_);
  and _80634_ (_30554_, _14273_, _08353_);
  or _80635_ (_30555_, _30554_, _30542_);
  and _80636_ (_30556_, _30555_, _06039_);
  or _80637_ (_30557_, _30556_, _06032_);
  or _80638_ (_30558_, _30557_, _30553_);
  and _80639_ (_30560_, _30543_, _14302_);
  or _80640_ (_30561_, _30542_, _06033_);
  or _80641_ (_30562_, _30561_, _30560_);
  and _80642_ (_30563_, _30562_, _06027_);
  and _80643_ (_30564_, _30563_, _30558_);
  or _80644_ (_30565_, _30542_, _14267_);
  and _80645_ (_30566_, _30565_, _06026_);
  and _80646_ (_30567_, _30566_, _30544_);
  or _80647_ (_30568_, _30567_, _09818_);
  or _80648_ (_30569_, _30568_, _30564_);
  and _80649_ (_30571_, _09075_, _07692_);
  or _80650_ (_30572_, _30520_, _07012_);
  or _80651_ (_30573_, _30572_, _30571_);
  or _80652_ (_30574_, _30525_, _09827_);
  and _80653_ (_30575_, _30574_, _05669_);
  and _80654_ (_30576_, _30575_, _30573_);
  and _80655_ (_30577_, _30576_, _30569_);
  and _80656_ (_30578_, _14367_, _07692_);
  or _80657_ (_30579_, _30578_, _30520_);
  and _80658_ (_30580_, _30579_, _09833_);
  or _80659_ (_30582_, _30580_, _30577_);
  and _80660_ (_30583_, _30582_, _06020_);
  nand _80661_ (_30584_, _07692_, _06832_);
  and _80662_ (_30585_, _30528_, _06019_);
  and _80663_ (_30586_, _30585_, _30584_);
  or _80664_ (_30587_, _30586_, _30583_);
  and _80665_ (_30588_, _30587_, _08751_);
  or _80666_ (_30589_, _14263_, _12902_);
  and _80667_ (_30590_, _30528_, _06112_);
  and _80668_ (_30591_, _30590_, _30589_);
  or _80669_ (_30593_, _30591_, _06284_);
  or _80670_ (_30594_, _30593_, _30588_);
  nand _80671_ (_30595_, _10992_, _07692_);
  and _80672_ (_30596_, _30595_, _30522_);
  or _80673_ (_30597_, _30596_, _08756_);
  and _80674_ (_30598_, _30597_, _07032_);
  and _80675_ (_30599_, _30598_, _30594_);
  or _80676_ (_30600_, _14261_, _12902_);
  and _80677_ (_30601_, _30528_, _06108_);
  and _80678_ (_30602_, _30601_, _30600_);
  or _80679_ (_30604_, _30602_, _06277_);
  or _80680_ (_30605_, _30604_, _30599_);
  nor _80681_ (_30606_, _30520_, _06278_);
  nand _80682_ (_30607_, _30606_, _30595_);
  and _80683_ (_30608_, _30607_, _08777_);
  and _80684_ (_30609_, _30608_, _30605_);
  or _80685_ (_30610_, _30584_, _08078_);
  and _80686_ (_30611_, _30528_, _06130_);
  and _80687_ (_30612_, _30611_, _30610_);
  or _80688_ (_30613_, _30612_, _06292_);
  or _80689_ (_30615_, _30613_, _30609_);
  and _80690_ (_30616_, _30615_, _30523_);
  or _80691_ (_30617_, _30616_, _06316_);
  or _80692_ (_30618_, _30531_, _06718_);
  and _80693_ (_30619_, _30618_, _05653_);
  and _80694_ (_30620_, _30619_, _30617_);
  and _80695_ (_30621_, _30555_, _05652_);
  or _80696_ (_30622_, _30621_, _06047_);
  or _80697_ (_30623_, _30622_, _30620_);
  or _80698_ (_30624_, _30520_, _06048_);
  or _80699_ (_30626_, _30624_, _30529_);
  and _80700_ (_30627_, _30626_, _01336_);
  and _80701_ (_30628_, _30627_, _30623_);
  nor _80702_ (_30629_, \oc8051_golden_model_1.P3 [1], rst);
  nor _80703_ (_30630_, _30629_, _00000_);
  or _80704_ (_43444_, _30630_, _30628_);
  nor _80705_ (_30631_, \oc8051_golden_model_1.P3 [2], rst);
  nor _80706_ (_30632_, _30631_, _00000_);
  and _80707_ (_30633_, _12902_, \oc8051_golden_model_1.P3 [2]);
  and _80708_ (_30634_, _07692_, _08730_);
  or _80709_ (_30636_, _30634_, _30633_);
  or _80710_ (_30637_, _30636_, _06020_);
  nor _80711_ (_30638_, _12902_, _07530_);
  or _80712_ (_30639_, _30638_, _30633_);
  and _80713_ (_30640_, _30639_, _06239_);
  and _80714_ (_30641_, _12921_, \oc8051_golden_model_1.P3 [2]);
  and _80715_ (_30642_, _14497_, _08353_);
  or _80716_ (_30643_, _30642_, _30641_);
  or _80717_ (_30644_, _30643_, _06044_);
  and _80718_ (_30645_, _14493_, _07692_);
  or _80719_ (_30647_, _30645_, _30633_);
  and _80720_ (_30648_, _30647_, _06102_);
  and _80721_ (_30649_, _06939_, \oc8051_golden_model_1.P3 [2]);
  and _80722_ (_30650_, _07692_, \oc8051_golden_model_1.ACC [2]);
  or _80723_ (_30651_, _30650_, _30633_);
  and _80724_ (_30652_, _30651_, _06938_);
  or _80725_ (_30653_, _30652_, _30649_);
  and _80726_ (_30654_, _30653_, _06954_);
  or _80727_ (_30655_, _30654_, _06043_);
  or _80728_ (_30656_, _30655_, _30648_);
  and _80729_ (_30658_, _30656_, _30644_);
  and _80730_ (_30659_, _30658_, _06848_);
  or _80731_ (_30660_, _30659_, _30640_);
  or _80732_ (_30661_, _30660_, _06219_);
  or _80733_ (_30662_, _30651_, _06220_);
  and _80734_ (_30663_, _30662_, _06040_);
  and _80735_ (_30664_, _30663_, _30661_);
  and _80736_ (_30665_, _14479_, _08353_);
  or _80737_ (_30666_, _30665_, _30641_);
  and _80738_ (_30667_, _30666_, _06039_);
  or _80739_ (_30669_, _30667_, _06032_);
  or _80740_ (_30670_, _30669_, _30664_);
  or _80741_ (_30671_, _30641_, _14512_);
  and _80742_ (_30672_, _30671_, _30643_);
  or _80743_ (_30673_, _30672_, _06033_);
  and _80744_ (_30674_, _30673_, _06027_);
  and _80745_ (_30675_, _30674_, _30670_);
  or _80746_ (_30676_, _30641_, _14525_);
  and _80747_ (_30677_, _30676_, _06026_);
  and _80748_ (_30678_, _30677_, _30643_);
  or _80749_ (_30680_, _30678_, _09818_);
  or _80750_ (_30681_, _30680_, _30675_);
  and _80751_ (_30682_, _09182_, _07692_);
  or _80752_ (_30683_, _30633_, _07012_);
  or _80753_ (_30684_, _30683_, _30682_);
  or _80754_ (_30685_, _30639_, _09827_);
  and _80755_ (_30686_, _30685_, _05669_);
  and _80756_ (_30687_, _30686_, _30684_);
  and _80757_ (_30688_, _30687_, _30681_);
  and _80758_ (_30689_, _14580_, _07692_);
  or _80759_ (_30691_, _30689_, _30633_);
  and _80760_ (_30692_, _30691_, _09833_);
  or _80761_ (_30693_, _30692_, _06019_);
  or _80762_ (_30694_, _30693_, _30688_);
  and _80763_ (_30695_, _30694_, _30637_);
  or _80764_ (_30696_, _30695_, _06112_);
  and _80765_ (_30697_, _14596_, _07692_);
  or _80766_ (_30698_, _30633_, _08751_);
  or _80767_ (_30699_, _30698_, _30697_);
  and _80768_ (_30700_, _30699_, _08756_);
  and _80769_ (_30702_, _30700_, _30696_);
  and _80770_ (_30703_, _10991_, _07692_);
  or _80771_ (_30704_, _30703_, _30633_);
  and _80772_ (_30705_, _30704_, _06284_);
  or _80773_ (_30706_, _30705_, _30702_);
  and _80774_ (_30707_, _30706_, _07032_);
  or _80775_ (_30708_, _30633_, _08177_);
  and _80776_ (_30709_, _30636_, _06108_);
  and _80777_ (_30710_, _30709_, _30708_);
  or _80778_ (_30711_, _30710_, _30707_);
  and _80779_ (_30713_, _30711_, _06278_);
  and _80780_ (_30714_, _30651_, _06277_);
  and _80781_ (_30715_, _30714_, _30708_);
  or _80782_ (_30716_, _30715_, _06130_);
  or _80783_ (_30717_, _30716_, _30713_);
  and _80784_ (_30718_, _14593_, _07692_);
  or _80785_ (_30719_, _30633_, _08777_);
  or _80786_ (_30720_, _30719_, _30718_);
  and _80787_ (_30721_, _30720_, _08782_);
  and _80788_ (_30722_, _30721_, _30717_);
  nor _80789_ (_30724_, _10990_, _12902_);
  or _80790_ (_30725_, _30724_, _30633_);
  and _80791_ (_30726_, _30725_, _06292_);
  or _80792_ (_30727_, _30726_, _06316_);
  or _80793_ (_30728_, _30727_, _30722_);
  or _80794_ (_30729_, _30647_, _06718_);
  and _80795_ (_30730_, _30729_, _05653_);
  and _80796_ (_30731_, _30730_, _30728_);
  and _80797_ (_30732_, _30666_, _05652_);
  or _80798_ (_30733_, _30732_, _06047_);
  or _80799_ (_30735_, _30733_, _30731_);
  and _80800_ (_30736_, _14657_, _07692_);
  or _80801_ (_30737_, _30633_, _06048_);
  or _80802_ (_30738_, _30737_, _30736_);
  and _80803_ (_30739_, _30738_, _01336_);
  and _80804_ (_30740_, _30739_, _30735_);
  or _80805_ (_43445_, _30740_, _30632_);
  nor _80806_ (_30741_, \oc8051_golden_model_1.P3 [3], rst);
  nor _80807_ (_30742_, _30741_, _00000_);
  and _80808_ (_30743_, _12902_, \oc8051_golden_model_1.P3 [3]);
  and _80809_ (_30745_, _07692_, _08662_);
  or _80810_ (_30746_, _30745_, _30743_);
  or _80811_ (_30747_, _30746_, _06020_);
  and _80812_ (_30748_, _14672_, _07692_);
  or _80813_ (_30749_, _30748_, _30743_);
  or _80814_ (_30750_, _30749_, _06954_);
  and _80815_ (_30751_, _07692_, \oc8051_golden_model_1.ACC [3]);
  or _80816_ (_30752_, _30751_, _30743_);
  and _80817_ (_30753_, _30752_, _06938_);
  and _80818_ (_30754_, _06939_, \oc8051_golden_model_1.P3 [3]);
  or _80819_ (_30756_, _30754_, _06102_);
  or _80820_ (_30757_, _30756_, _30753_);
  and _80821_ (_30758_, _30757_, _06044_);
  and _80822_ (_30759_, _30758_, _30750_);
  and _80823_ (_30760_, _12921_, \oc8051_golden_model_1.P3 [3]);
  and _80824_ (_30761_, _14683_, _08353_);
  or _80825_ (_30762_, _30761_, _30760_);
  and _80826_ (_30763_, _30762_, _06043_);
  or _80827_ (_30764_, _30763_, _06239_);
  or _80828_ (_30765_, _30764_, _30759_);
  nor _80829_ (_30767_, _12902_, _07353_);
  or _80830_ (_30768_, _30767_, _30743_);
  or _80831_ (_30769_, _30768_, _06848_);
  and _80832_ (_30770_, _30769_, _30765_);
  or _80833_ (_30771_, _30770_, _06219_);
  or _80834_ (_30772_, _30752_, _06220_);
  and _80835_ (_30773_, _30772_, _06040_);
  and _80836_ (_30774_, _30773_, _30771_);
  and _80837_ (_30775_, _14681_, _08353_);
  or _80838_ (_30776_, _30775_, _30760_);
  and _80839_ (_30778_, _30776_, _06039_);
  or _80840_ (_30779_, _30778_, _06032_);
  or _80841_ (_30780_, _30779_, _30774_);
  or _80842_ (_30781_, _30760_, _14708_);
  and _80843_ (_30782_, _30781_, _30762_);
  or _80844_ (_30783_, _30782_, _06033_);
  and _80845_ (_30784_, _30783_, _06027_);
  and _80846_ (_30785_, _30784_, _30780_);
  and _80847_ (_30786_, _14724_, _08353_);
  or _80848_ (_30787_, _30786_, _30760_);
  and _80849_ (_30789_, _30787_, _06026_);
  or _80850_ (_30790_, _30789_, _09818_);
  or _80851_ (_30791_, _30790_, _30785_);
  and _80852_ (_30792_, _09181_, _07692_);
  or _80853_ (_30793_, _30743_, _07012_);
  or _80854_ (_30794_, _30793_, _30792_);
  or _80855_ (_30795_, _30768_, _09827_);
  and _80856_ (_30796_, _30795_, _05669_);
  and _80857_ (_30797_, _30796_, _30794_);
  and _80858_ (_30798_, _30797_, _30791_);
  and _80859_ (_30800_, _14778_, _07692_);
  or _80860_ (_30801_, _30800_, _30743_);
  and _80861_ (_30802_, _30801_, _09833_);
  or _80862_ (_30803_, _30802_, _06019_);
  or _80863_ (_30804_, _30803_, _30798_);
  and _80864_ (_30805_, _30804_, _30747_);
  or _80865_ (_30806_, _30805_, _06112_);
  and _80866_ (_30807_, _14793_, _07692_);
  or _80867_ (_30808_, _30743_, _08751_);
  or _80868_ (_30809_, _30808_, _30807_);
  and _80869_ (_30811_, _30809_, _08756_);
  and _80870_ (_30812_, _30811_, _30806_);
  and _80871_ (_30813_, _12299_, _07692_);
  or _80872_ (_30814_, _30813_, _30743_);
  and _80873_ (_30815_, _30814_, _06284_);
  or _80874_ (_30816_, _30815_, _30812_);
  and _80875_ (_30817_, _30816_, _07032_);
  or _80876_ (_30818_, _30743_, _08029_);
  and _80877_ (_30819_, _30746_, _06108_);
  and _80878_ (_30820_, _30819_, _30818_);
  or _80879_ (_30822_, _30820_, _30817_);
  and _80880_ (_30823_, _30822_, _06278_);
  and _80881_ (_30824_, _30752_, _06277_);
  and _80882_ (_30825_, _30824_, _30818_);
  or _80883_ (_30826_, _30825_, _06130_);
  or _80884_ (_30827_, _30826_, _30823_);
  and _80885_ (_30828_, _14792_, _07692_);
  or _80886_ (_30829_, _30743_, _08777_);
  or _80887_ (_30830_, _30829_, _30828_);
  and _80888_ (_30831_, _30830_, _08782_);
  and _80889_ (_30833_, _30831_, _30827_);
  nor _80890_ (_30834_, _10988_, _12902_);
  or _80891_ (_30835_, _30834_, _30743_);
  and _80892_ (_30836_, _30835_, _06292_);
  or _80893_ (_30837_, _30836_, _06316_);
  or _80894_ (_30838_, _30837_, _30833_);
  or _80895_ (_30839_, _30749_, _06718_);
  and _80896_ (_30840_, _30839_, _05653_);
  and _80897_ (_30841_, _30840_, _30838_);
  and _80898_ (_30842_, _30776_, _05652_);
  or _80899_ (_30844_, _30842_, _06047_);
  or _80900_ (_30845_, _30844_, _30841_);
  and _80901_ (_30846_, _14849_, _07692_);
  or _80902_ (_30847_, _30743_, _06048_);
  or _80903_ (_30848_, _30847_, _30846_);
  and _80904_ (_30849_, _30848_, _01336_);
  and _80905_ (_30850_, _30849_, _30845_);
  or _80906_ (_43446_, _30850_, _30742_);
  and _80907_ (_30851_, _12902_, \oc8051_golden_model_1.P3 [4]);
  and _80908_ (_30852_, _08665_, _07692_);
  or _80909_ (_30854_, _30852_, _30851_);
  or _80910_ (_30855_, _30854_, _06020_);
  and _80911_ (_30856_, _14887_, _07692_);
  or _80912_ (_30857_, _30856_, _30851_);
  or _80913_ (_30858_, _30857_, _06954_);
  and _80914_ (_30859_, _07692_, \oc8051_golden_model_1.ACC [4]);
  or _80915_ (_30860_, _30859_, _30851_);
  and _80916_ (_30861_, _30860_, _06938_);
  and _80917_ (_30862_, _06939_, \oc8051_golden_model_1.P3 [4]);
  or _80918_ (_30863_, _30862_, _06102_);
  or _80919_ (_30865_, _30863_, _30861_);
  and _80920_ (_30866_, _30865_, _06044_);
  and _80921_ (_30867_, _30866_, _30858_);
  and _80922_ (_30868_, _12921_, \oc8051_golden_model_1.P3 [4]);
  and _80923_ (_30869_, _14878_, _08353_);
  or _80924_ (_30870_, _30869_, _30868_);
  and _80925_ (_30871_, _30870_, _06043_);
  or _80926_ (_30872_, _30871_, _06239_);
  or _80927_ (_30873_, _30872_, _30867_);
  nor _80928_ (_30874_, _08270_, _12902_);
  or _80929_ (_30876_, _30874_, _30851_);
  or _80930_ (_30877_, _30876_, _06848_);
  and _80931_ (_30878_, _30877_, _30873_);
  or _80932_ (_30879_, _30878_, _06219_);
  or _80933_ (_30880_, _30860_, _06220_);
  and _80934_ (_30881_, _30880_, _06040_);
  and _80935_ (_30882_, _30881_, _30879_);
  and _80936_ (_30883_, _14882_, _08353_);
  or _80937_ (_30884_, _30883_, _30868_);
  and _80938_ (_30885_, _30884_, _06039_);
  or _80939_ (_30887_, _30885_, _06032_);
  or _80940_ (_30888_, _30887_, _30882_);
  or _80941_ (_30889_, _30868_, _14914_);
  and _80942_ (_30890_, _30889_, _30870_);
  or _80943_ (_30891_, _30890_, _06033_);
  and _80944_ (_30892_, _30891_, _06027_);
  and _80945_ (_30893_, _30892_, _30888_);
  or _80946_ (_30894_, _30868_, _14879_);
  and _80947_ (_30895_, _30894_, _06026_);
  and _80948_ (_30896_, _30895_, _30870_);
  or _80949_ (_30898_, _30896_, _09818_);
  or _80950_ (_30899_, _30898_, _30893_);
  and _80951_ (_30900_, _09180_, _07692_);
  or _80952_ (_30901_, _30851_, _07012_);
  or _80953_ (_30902_, _30901_, _30900_);
  or _80954_ (_30903_, _30876_, _09827_);
  and _80955_ (_30904_, _30903_, _05669_);
  and _80956_ (_30905_, _30904_, _30902_);
  and _80957_ (_30906_, _30905_, _30899_);
  and _80958_ (_30907_, _14983_, _07692_);
  or _80959_ (_30909_, _30907_, _30851_);
  and _80960_ (_30910_, _30909_, _09833_);
  or _80961_ (_30911_, _30910_, _06019_);
  or _80962_ (_30912_, _30911_, _30906_);
  and _80963_ (_30913_, _30912_, _30855_);
  or _80964_ (_30914_, _30913_, _06112_);
  and _80965_ (_30915_, _14876_, _07692_);
  or _80966_ (_30916_, _30915_, _30851_);
  or _80967_ (_30917_, _30916_, _08751_);
  and _80968_ (_30918_, _30917_, _08756_);
  and _80969_ (_30920_, _30918_, _30914_);
  and _80970_ (_30921_, _10986_, _07692_);
  or _80971_ (_30922_, _30921_, _30851_);
  and _80972_ (_30923_, _30922_, _06284_);
  or _80973_ (_30924_, _30923_, _30920_);
  and _80974_ (_30925_, _30924_, _07032_);
  or _80975_ (_30926_, _30851_, _08273_);
  and _80976_ (_30927_, _30854_, _06108_);
  and _80977_ (_30928_, _30927_, _30926_);
  or _80978_ (_30929_, _30928_, _30925_);
  and _80979_ (_30931_, _30929_, _06278_);
  and _80980_ (_30932_, _30860_, _06277_);
  and _80981_ (_30933_, _30932_, _30926_);
  or _80982_ (_30934_, _30933_, _06130_);
  or _80983_ (_30935_, _30934_, _30931_);
  and _80984_ (_30936_, _14873_, _07692_);
  or _80985_ (_30937_, _30851_, _08777_);
  or _80986_ (_30938_, _30937_, _30936_);
  and _80987_ (_30939_, _30938_, _08782_);
  and _80988_ (_30940_, _30939_, _30935_);
  nor _80989_ (_30942_, _10985_, _12902_);
  or _80990_ (_30943_, _30942_, _30851_);
  and _80991_ (_30944_, _30943_, _06292_);
  or _80992_ (_30945_, _30944_, _06316_);
  or _80993_ (_30946_, _30945_, _30940_);
  or _80994_ (_30947_, _30857_, _06718_);
  and _80995_ (_30948_, _30947_, _05653_);
  and _80996_ (_30949_, _30948_, _30946_);
  and _80997_ (_30950_, _30884_, _05652_);
  or _80998_ (_30951_, _30950_, _06047_);
  or _80999_ (_30953_, _30951_, _30949_);
  and _81000_ (_30954_, _15055_, _07692_);
  or _81001_ (_30955_, _30851_, _06048_);
  or _81002_ (_30956_, _30955_, _30954_);
  and _81003_ (_30957_, _30956_, _01336_);
  and _81004_ (_30958_, _30957_, _30953_);
  nor _81005_ (_30959_, \oc8051_golden_model_1.P3 [4], rst);
  nor _81006_ (_30960_, _30959_, _00000_);
  or _81007_ (_43447_, _30960_, _30958_);
  nor _81008_ (_30961_, \oc8051_golden_model_1.P3 [5], rst);
  nor _81009_ (_30963_, _30961_, _00000_);
  and _81010_ (_30964_, _12902_, \oc8051_golden_model_1.P3 [5]);
  and _81011_ (_30965_, _08652_, _07692_);
  or _81012_ (_30966_, _30965_, _30964_);
  or _81013_ (_30967_, _30966_, _06020_);
  and _81014_ (_30968_, _15093_, _07692_);
  or _81015_ (_30969_, _30968_, _30964_);
  or _81016_ (_30970_, _30969_, _06954_);
  and _81017_ (_30971_, _07692_, \oc8051_golden_model_1.ACC [5]);
  or _81018_ (_30972_, _30971_, _30964_);
  and _81019_ (_30974_, _30972_, _06938_);
  and _81020_ (_30975_, _06939_, \oc8051_golden_model_1.P3 [5]);
  or _81021_ (_30976_, _30975_, _06102_);
  or _81022_ (_30977_, _30976_, _30974_);
  and _81023_ (_30978_, _30977_, _06044_);
  and _81024_ (_30979_, _30978_, _30970_);
  and _81025_ (_30980_, _12921_, \oc8051_golden_model_1.P3 [5]);
  and _81026_ (_30981_, _15073_, _08353_);
  or _81027_ (_30982_, _30981_, _30980_);
  and _81028_ (_30983_, _30982_, _06043_);
  or _81029_ (_30985_, _30983_, _06239_);
  or _81030_ (_30986_, _30985_, _30979_);
  nor _81031_ (_30987_, _07977_, _12902_);
  or _81032_ (_30988_, _30987_, _30964_);
  or _81033_ (_30989_, _30988_, _06848_);
  and _81034_ (_30990_, _30989_, _30986_);
  or _81035_ (_30991_, _30990_, _06219_);
  or _81036_ (_30992_, _30972_, _06220_);
  and _81037_ (_30993_, _30992_, _06040_);
  and _81038_ (_30994_, _30993_, _30991_);
  and _81039_ (_30996_, _15077_, _08353_);
  or _81040_ (_30997_, _30996_, _30980_);
  and _81041_ (_30998_, _30997_, _06039_);
  or _81042_ (_30999_, _30998_, _06032_);
  or _81043_ (_31000_, _30999_, _30994_);
  or _81044_ (_31001_, _30980_, _15110_);
  and _81045_ (_31002_, _31001_, _30982_);
  or _81046_ (_31003_, _31002_, _06033_);
  and _81047_ (_31004_, _31003_, _06027_);
  and _81048_ (_31005_, _31004_, _31000_);
  or _81049_ (_31007_, _30980_, _15074_);
  and _81050_ (_31008_, _31007_, _06026_);
  and _81051_ (_31009_, _31008_, _30982_);
  or _81052_ (_31010_, _31009_, _09818_);
  or _81053_ (_31011_, _31010_, _31005_);
  and _81054_ (_31012_, _09179_, _07692_);
  or _81055_ (_31013_, _30964_, _07012_);
  or _81056_ (_31014_, _31013_, _31012_);
  or _81057_ (_31015_, _30988_, _09827_);
  and _81058_ (_31016_, _31015_, _05669_);
  and _81059_ (_31018_, _31016_, _31014_);
  and _81060_ (_31019_, _31018_, _31011_);
  and _81061_ (_31020_, _15179_, _07692_);
  or _81062_ (_31021_, _31020_, _30964_);
  and _81063_ (_31022_, _31021_, _09833_);
  or _81064_ (_31023_, _31022_, _06019_);
  or _81065_ (_31024_, _31023_, _31019_);
  and _81066_ (_31025_, _31024_, _30967_);
  or _81067_ (_31026_, _31025_, _06112_);
  and _81068_ (_31027_, _15195_, _07692_);
  or _81069_ (_31029_, _30964_, _08751_);
  or _81070_ (_31030_, _31029_, _31027_);
  and _81071_ (_31031_, _31030_, _08756_);
  and _81072_ (_31032_, _31031_, _31026_);
  and _81073_ (_31033_, _12306_, _07692_);
  or _81074_ (_31034_, _31033_, _30964_);
  and _81075_ (_31035_, _31034_, _06284_);
  or _81076_ (_31036_, _31035_, _31032_);
  and _81077_ (_31037_, _31036_, _07032_);
  or _81078_ (_31038_, _30964_, _07980_);
  and _81079_ (_31040_, _30966_, _06108_);
  and _81080_ (_31041_, _31040_, _31038_);
  or _81081_ (_31042_, _31041_, _31037_);
  and _81082_ (_31043_, _31042_, _06278_);
  and _81083_ (_31044_, _30972_, _06277_);
  and _81084_ (_31045_, _31044_, _31038_);
  or _81085_ (_31046_, _31045_, _06130_);
  or _81086_ (_31047_, _31046_, _31043_);
  and _81087_ (_31048_, _15194_, _07692_);
  or _81088_ (_31049_, _30964_, _08777_);
  or _81089_ (_31051_, _31049_, _31048_);
  and _81090_ (_31052_, _31051_, _08782_);
  and _81091_ (_31053_, _31052_, _31047_);
  nor _81092_ (_31054_, _10982_, _12902_);
  or _81093_ (_31055_, _31054_, _30964_);
  and _81094_ (_31056_, _31055_, _06292_);
  or _81095_ (_31057_, _31056_, _06316_);
  or _81096_ (_31058_, _31057_, _31053_);
  or _81097_ (_31059_, _30969_, _06718_);
  and _81098_ (_31060_, _31059_, _05653_);
  and _81099_ (_31062_, _31060_, _31058_);
  and _81100_ (_31063_, _30997_, _05652_);
  or _81101_ (_31064_, _31063_, _06047_);
  or _81102_ (_31065_, _31064_, _31062_);
  and _81103_ (_31066_, _15253_, _07692_);
  or _81104_ (_31067_, _30964_, _06048_);
  or _81105_ (_31068_, _31067_, _31066_);
  and _81106_ (_31069_, _31068_, _01336_);
  and _81107_ (_31070_, _31069_, _31065_);
  or _81108_ (_43448_, _31070_, _30963_);
  and _81109_ (_31072_, _12902_, \oc8051_golden_model_1.P3 [6]);
  and _81110_ (_31073_, _15389_, _07692_);
  or _81111_ (_31074_, _31073_, _31072_);
  or _81112_ (_31075_, _31074_, _06020_);
  and _81113_ (_31076_, _15293_, _07692_);
  or _81114_ (_31077_, _31076_, _31072_);
  or _81115_ (_31078_, _31077_, _06954_);
  and _81116_ (_31079_, _07692_, \oc8051_golden_model_1.ACC [6]);
  or _81117_ (_31080_, _31079_, _31072_);
  and _81118_ (_31081_, _31080_, _06938_);
  and _81119_ (_31083_, _06939_, \oc8051_golden_model_1.P3 [6]);
  or _81120_ (_31084_, _31083_, _06102_);
  or _81121_ (_31085_, _31084_, _31081_);
  and _81122_ (_31086_, _31085_, _06044_);
  and _81123_ (_31087_, _31086_, _31078_);
  and _81124_ (_31088_, _12921_, \oc8051_golden_model_1.P3 [6]);
  and _81125_ (_31089_, _15280_, _08353_);
  or _81126_ (_31090_, _31089_, _31088_);
  and _81127_ (_31091_, _31090_, _06043_);
  or _81128_ (_31092_, _31091_, _06239_);
  or _81129_ (_31094_, _31092_, _31087_);
  nor _81130_ (_31095_, _07883_, _12902_);
  or _81131_ (_31096_, _31095_, _31072_);
  or _81132_ (_31097_, _31096_, _06848_);
  and _81133_ (_31098_, _31097_, _31094_);
  or _81134_ (_31099_, _31098_, _06219_);
  or _81135_ (_31100_, _31080_, _06220_);
  and _81136_ (_31101_, _31100_, _06040_);
  and _81137_ (_31102_, _31101_, _31099_);
  and _81138_ (_31103_, _15278_, _08353_);
  or _81139_ (_31105_, _31103_, _31088_);
  and _81140_ (_31106_, _31105_, _06039_);
  or _81141_ (_31107_, _31106_, _06032_);
  or _81142_ (_31108_, _31107_, _31102_);
  or _81143_ (_31109_, _31088_, _15310_);
  and _81144_ (_31110_, _31109_, _31090_);
  or _81145_ (_31111_, _31110_, _06033_);
  and _81146_ (_31112_, _31111_, _06027_);
  and _81147_ (_31113_, _31112_, _31108_);
  or _81148_ (_31114_, _31088_, _15326_);
  and _81149_ (_31116_, _31114_, _06026_);
  and _81150_ (_31117_, _31116_, _31090_);
  or _81151_ (_31118_, _31117_, _09818_);
  or _81152_ (_31119_, _31118_, _31113_);
  and _81153_ (_31120_, _09178_, _07692_);
  or _81154_ (_31121_, _31072_, _07012_);
  or _81155_ (_31122_, _31121_, _31120_);
  or _81156_ (_31123_, _31096_, _09827_);
  and _81157_ (_31124_, _31123_, _05669_);
  and _81158_ (_31125_, _31124_, _31122_);
  and _81159_ (_31127_, _31125_, _31119_);
  and _81160_ (_31128_, _15382_, _07692_);
  or _81161_ (_31129_, _31128_, _31072_);
  and _81162_ (_31130_, _31129_, _09833_);
  or _81163_ (_31131_, _31130_, _06019_);
  or _81164_ (_31132_, _31131_, _31127_);
  and _81165_ (_31133_, _31132_, _31075_);
  or _81166_ (_31134_, _31133_, _06112_);
  and _81167_ (_31135_, _15399_, _07692_);
  or _81168_ (_31136_, _31072_, _08751_);
  or _81169_ (_31139_, _31136_, _31135_);
  and _81170_ (_31140_, _31139_, _08756_);
  and _81171_ (_31141_, _31140_, _31134_);
  and _81172_ (_31142_, _10980_, _07692_);
  or _81173_ (_31143_, _31142_, _31072_);
  and _81174_ (_31144_, _31143_, _06284_);
  or _81175_ (_31145_, _31144_, _31141_);
  and _81176_ (_31146_, _31145_, _07032_);
  or _81177_ (_31147_, _31072_, _07886_);
  and _81178_ (_31148_, _31074_, _06108_);
  and _81179_ (_31150_, _31148_, _31147_);
  or _81180_ (_31151_, _31150_, _31146_);
  and _81181_ (_31152_, _31151_, _06278_);
  and _81182_ (_31153_, _31080_, _06277_);
  and _81183_ (_31154_, _31153_, _31147_);
  or _81184_ (_31155_, _31154_, _06130_);
  or _81185_ (_31156_, _31155_, _31152_);
  and _81186_ (_31157_, _15396_, _07692_);
  or _81187_ (_31158_, _31072_, _08777_);
  or _81188_ (_31159_, _31158_, _31157_);
  and _81189_ (_31162_, _31159_, _08782_);
  and _81190_ (_31163_, _31162_, _31156_);
  nor _81191_ (_31164_, _10979_, _12902_);
  or _81192_ (_31165_, _31164_, _31072_);
  and _81193_ (_31166_, _31165_, _06292_);
  or _81194_ (_31167_, _31166_, _06316_);
  or _81195_ (_31168_, _31167_, _31163_);
  or _81196_ (_31169_, _31077_, _06718_);
  and _81197_ (_31170_, _31169_, _05653_);
  and _81198_ (_31171_, _31170_, _31168_);
  and _81199_ (_31173_, _31105_, _05652_);
  or _81200_ (_31174_, _31173_, _06047_);
  or _81201_ (_31175_, _31174_, _31171_);
  and _81202_ (_31176_, _15451_, _07692_);
  or _81203_ (_31177_, _31072_, _06048_);
  or _81204_ (_31178_, _31177_, _31176_);
  and _81205_ (_31179_, _31178_, _01336_);
  and _81206_ (_31180_, _31179_, _31175_);
  nor _81207_ (_31181_, \oc8051_golden_model_1.P3 [6], rst);
  nor _81208_ (_31182_, _31181_, _00000_);
  or _81209_ (_43449_, _31182_, _31180_);
  nor _81210_ (_31185_, \oc8051_golden_model_1.P0 [0], rst);
  nor _81211_ (_31186_, _31185_, _00000_);
  nand _81212_ (_31187_, _10995_, _07730_);
  not _81213_ (_31188_, \oc8051_golden_model_1.P0 [0]);
  nor _81214_ (_31189_, _07730_, _31188_);
  nor _81215_ (_31190_, _31189_, _06278_);
  nand _81216_ (_31191_, _31190_, _31187_);
  and _81217_ (_31192_, _07730_, _08672_);
  or _81218_ (_31193_, _31192_, _31189_);
  or _81219_ (_31195_, _31193_, _06020_);
  and _81220_ (_31196_, _09120_, _07730_);
  or _81221_ (_31197_, _31189_, _07012_);
  or _81222_ (_31198_, _31197_, _31196_);
  nor _81223_ (_31199_, _08127_, _13006_);
  or _81224_ (_31200_, _31199_, _31189_);
  or _81225_ (_31201_, _31200_, _06954_);
  and _81226_ (_31202_, _07730_, \oc8051_golden_model_1.ACC [0]);
  or _81227_ (_31203_, _31202_, _31189_);
  and _81228_ (_31204_, _31203_, _06938_);
  nor _81229_ (_31207_, _06938_, _31188_);
  or _81230_ (_31208_, _31207_, _06102_);
  or _81231_ (_31209_, _31208_, _31204_);
  and _81232_ (_31210_, _31209_, _06044_);
  and _81233_ (_31211_, _31210_, _31201_);
  nor _81234_ (_31212_, _07638_, _31188_);
  and _81235_ (_31213_, _14102_, _07638_);
  or _81236_ (_31214_, _31213_, _31212_);
  and _81237_ (_31215_, _31214_, _06043_);
  or _81238_ (_31216_, _31215_, _31211_);
  and _81239_ (_31218_, _31216_, _06848_);
  and _81240_ (_31219_, _07730_, _06931_);
  or _81241_ (_31220_, _31219_, _31189_);
  and _81242_ (_31221_, _31220_, _06239_);
  or _81243_ (_31222_, _31221_, _06219_);
  or _81244_ (_31223_, _31222_, _31218_);
  or _81245_ (_31224_, _31203_, _06220_);
  and _81246_ (_31225_, _31224_, _06040_);
  and _81247_ (_31226_, _31225_, _31223_);
  and _81248_ (_31227_, _31189_, _06039_);
  or _81249_ (_31229_, _31227_, _06032_);
  or _81250_ (_31230_, _31229_, _31226_);
  or _81251_ (_31231_, _31200_, _06033_);
  and _81252_ (_31232_, _31231_, _06027_);
  and _81253_ (_31233_, _31232_, _31230_);
  or _81254_ (_31234_, _31212_, _14131_);
  and _81255_ (_31235_, _31234_, _06026_);
  and _81256_ (_31236_, _31235_, _31214_);
  or _81257_ (_31237_, _31236_, _09818_);
  or _81258_ (_31238_, _31237_, _31233_);
  or _81259_ (_31240_, _31220_, _09827_);
  and _81260_ (_31241_, _31240_, _05669_);
  and _81261_ (_31242_, _31241_, _31238_);
  and _81262_ (_31243_, _31242_, _31198_);
  and _81263_ (_31244_, _14186_, _07730_);
  or _81264_ (_31245_, _31244_, _31189_);
  and _81265_ (_31246_, _31245_, _09833_);
  or _81266_ (_31247_, _31246_, _06019_);
  or _81267_ (_31248_, _31247_, _31243_);
  and _81268_ (_31249_, _31248_, _31195_);
  or _81269_ (_31250_, _31249_, _06112_);
  and _81270_ (_31251_, _14086_, _07730_);
  or _81271_ (_31252_, _31251_, _31189_);
  or _81272_ (_31253_, _31252_, _08751_);
  and _81273_ (_31254_, _31253_, _08756_);
  and _81274_ (_31255_, _31254_, _31250_);
  nor _81275_ (_31256_, _12302_, _13006_);
  or _81276_ (_31257_, _31256_, _31189_);
  and _81277_ (_31258_, _31187_, _06284_);
  and _81278_ (_31259_, _31258_, _31257_);
  or _81279_ (_31262_, _31259_, _31255_);
  and _81280_ (_31263_, _31262_, _07032_);
  nand _81281_ (_31264_, _31193_, _06108_);
  nor _81282_ (_31265_, _31264_, _31199_);
  or _81283_ (_31266_, _31265_, _06277_);
  or _81284_ (_31267_, _31266_, _31263_);
  and _81285_ (_31268_, _31267_, _31191_);
  or _81286_ (_31269_, _31268_, _06130_);
  and _81287_ (_31270_, _14083_, _07730_);
  or _81288_ (_31271_, _31189_, _08777_);
  or _81289_ (_31272_, _31271_, _31270_);
  and _81290_ (_31273_, _31272_, _08782_);
  and _81291_ (_31274_, _31273_, _31269_);
  and _81292_ (_31275_, _31257_, _06292_);
  or _81293_ (_31276_, _31275_, _06316_);
  or _81294_ (_31277_, _31276_, _31274_);
  or _81295_ (_31278_, _31200_, _06718_);
  and _81296_ (_31279_, _31278_, _31277_);
  or _81297_ (_31280_, _31279_, _05652_);
  or _81298_ (_31281_, _31189_, _05653_);
  and _81299_ (_31284_, _31281_, _31280_);
  or _81300_ (_31285_, _31284_, _06047_);
  or _81301_ (_31286_, _31200_, _06048_);
  and _81302_ (_31287_, _31286_, _01336_);
  and _81303_ (_31288_, _31287_, _31285_);
  or _81304_ (_43451_, _31288_, _31186_);
  nor _81305_ (_31289_, \oc8051_golden_model_1.P0 [1], rst);
  nor _81306_ (_31290_, _31289_, _00000_);
  and _81307_ (_31291_, _13006_, \oc8051_golden_model_1.P0 [1]);
  nor _81308_ (_31292_, _10993_, _13006_);
  or _81309_ (_31293_, _31292_, _31291_);
  or _81310_ (_31294_, _31293_, _08782_);
  or _81311_ (_31295_, _14367_, _13006_);
  or _81312_ (_31296_, _07730_, \oc8051_golden_model_1.P0 [1]);
  and _81313_ (_31297_, _31296_, _09833_);
  and _81314_ (_31298_, _31297_, _31295_);
  nor _81315_ (_31299_, _13006_, _07132_);
  or _81316_ (_31300_, _31299_, _31291_);
  or _81317_ (_31301_, _31300_, _06848_);
  and _81318_ (_31302_, _14284_, _07730_);
  not _81319_ (_31305_, _31302_);
  and _81320_ (_31306_, _31305_, _31296_);
  or _81321_ (_31307_, _31306_, _06954_);
  and _81322_ (_31308_, _07730_, \oc8051_golden_model_1.ACC [1]);
  or _81323_ (_31309_, _31308_, _31291_);
  and _81324_ (_31310_, _31309_, _06938_);
  and _81325_ (_31311_, _06939_, \oc8051_golden_model_1.P0 [1]);
  or _81326_ (_31312_, _31311_, _06102_);
  or _81327_ (_31313_, _31312_, _31310_);
  and _81328_ (_31314_, _31313_, _06044_);
  and _81329_ (_31315_, _31314_, _31307_);
  and _81330_ (_31316_, _13025_, \oc8051_golden_model_1.P0 [1]);
  and _81331_ (_31317_, _14266_, _07638_);
  or _81332_ (_31318_, _31317_, _31316_);
  and _81333_ (_31319_, _31318_, _06043_);
  or _81334_ (_31320_, _31319_, _06239_);
  or _81335_ (_31321_, _31320_, _31315_);
  and _81336_ (_31322_, _31321_, _31301_);
  or _81337_ (_31323_, _31322_, _06219_);
  or _81338_ (_31324_, _31309_, _06220_);
  and _81339_ (_31327_, _31324_, _06040_);
  and _81340_ (_31328_, _31327_, _31323_);
  and _81341_ (_31329_, _14273_, _07638_);
  or _81342_ (_31330_, _31329_, _31316_);
  and _81343_ (_31331_, _31330_, _06039_);
  or _81344_ (_31332_, _31331_, _06032_);
  or _81345_ (_31333_, _31332_, _31328_);
  and _81346_ (_31334_, _31317_, _14302_);
  or _81347_ (_31335_, _31316_, _06033_);
  or _81348_ (_31336_, _31335_, _31334_);
  and _81349_ (_31337_, _31336_, _06027_);
  and _81350_ (_31338_, _31337_, _31333_);
  or _81351_ (_31339_, _31316_, _14267_);
  and _81352_ (_31340_, _31339_, _06026_);
  and _81353_ (_31341_, _31340_, _31318_);
  or _81354_ (_31342_, _31341_, _09818_);
  or _81355_ (_31343_, _31342_, _31338_);
  and _81356_ (_31344_, _09075_, _07730_);
  or _81357_ (_31345_, _31344_, _31291_);
  or _81358_ (_31346_, _31345_, _07012_);
  or _81359_ (_31349_, _31300_, _09827_);
  and _81360_ (_31350_, _31349_, _05669_);
  and _81361_ (_31351_, _31350_, _31346_);
  and _81362_ (_31352_, _31351_, _31343_);
  or _81363_ (_31353_, _31352_, _31298_);
  and _81364_ (_31354_, _31353_, _06020_);
  nand _81365_ (_31355_, _07730_, _06832_);
  and _81366_ (_31356_, _31296_, _06019_);
  and _81367_ (_31357_, _31356_, _31355_);
  or _81368_ (_31358_, _31357_, _31354_);
  and _81369_ (_31359_, _31358_, _08751_);
  or _81370_ (_31360_, _14263_, _13006_);
  and _81371_ (_31361_, _31296_, _06112_);
  and _81372_ (_31362_, _31361_, _31360_);
  or _81373_ (_31363_, _31362_, _06284_);
  or _81374_ (_31364_, _31363_, _31359_);
  and _81375_ (_31365_, _10994_, _07730_);
  or _81376_ (_31366_, _31365_, _31291_);
  or _81377_ (_31367_, _31366_, _08756_);
  and _81378_ (_31368_, _31367_, _07032_);
  and _81379_ (_31371_, _31368_, _31364_);
  or _81380_ (_31372_, _14261_, _13006_);
  and _81381_ (_31373_, _31296_, _06108_);
  and _81382_ (_31374_, _31373_, _31372_);
  or _81383_ (_31375_, _31374_, _06277_);
  or _81384_ (_31376_, _31375_, _31371_);
  and _81385_ (_31377_, _31308_, _08078_);
  or _81386_ (_31378_, _31291_, _06278_);
  or _81387_ (_31379_, _31378_, _31377_);
  and _81388_ (_31380_, _31379_, _08777_);
  and _81389_ (_31381_, _31380_, _31376_);
  or _81390_ (_31382_, _31355_, _08078_);
  and _81391_ (_31383_, _31296_, _06130_);
  and _81392_ (_31384_, _31383_, _31382_);
  or _81393_ (_31385_, _31384_, _06292_);
  or _81394_ (_31386_, _31385_, _31381_);
  and _81395_ (_31387_, _31386_, _31294_);
  or _81396_ (_31388_, _31387_, _06316_);
  or _81397_ (_31389_, _31306_, _06718_);
  and _81398_ (_31390_, _31389_, _05653_);
  and _81399_ (_31393_, _31390_, _31388_);
  and _81400_ (_31394_, _31330_, _05652_);
  or _81401_ (_31395_, _31394_, _06047_);
  or _81402_ (_31396_, _31395_, _31393_);
  or _81403_ (_31397_, _31291_, _06048_);
  or _81404_ (_31398_, _31397_, _31302_);
  and _81405_ (_31399_, _31398_, _01336_);
  and _81406_ (_31400_, _31399_, _31396_);
  or _81407_ (_43452_, _31400_, _31290_);
  nor _81408_ (_31401_, \oc8051_golden_model_1.P0 [2], rst);
  nor _81409_ (_31402_, _31401_, _00000_);
  and _81410_ (_31403_, _13006_, \oc8051_golden_model_1.P0 [2]);
  or _81411_ (_31404_, _31403_, _08177_);
  and _81412_ (_31405_, _07730_, _08730_);
  or _81413_ (_31406_, _31405_, _31403_);
  and _81414_ (_31407_, _31406_, _06108_);
  and _81415_ (_31408_, _31407_, _31404_);
  or _81416_ (_31409_, _31406_, _06020_);
  nor _81417_ (_31410_, _13006_, _07530_);
  or _81418_ (_31411_, _31410_, _31403_);
  or _81419_ (_31413_, _31411_, _06848_);
  and _81420_ (_31414_, _14493_, _07730_);
  or _81421_ (_31415_, _31414_, _31403_);
  or _81422_ (_31416_, _31415_, _06954_);
  and _81423_ (_31417_, _07730_, \oc8051_golden_model_1.ACC [2]);
  or _81424_ (_31418_, _31417_, _31403_);
  and _81425_ (_31419_, _31418_, _06938_);
  and _81426_ (_31420_, _06939_, \oc8051_golden_model_1.P0 [2]);
  or _81427_ (_31421_, _31420_, _06102_);
  or _81428_ (_31422_, _31421_, _31419_);
  and _81429_ (_31423_, _31422_, _06044_);
  and _81430_ (_31424_, _31423_, _31416_);
  and _81431_ (_31425_, _13025_, \oc8051_golden_model_1.P0 [2]);
  and _81432_ (_31426_, _14497_, _07638_);
  or _81433_ (_31427_, _31426_, _31425_);
  and _81434_ (_31428_, _31427_, _06043_);
  or _81435_ (_31429_, _31428_, _06239_);
  or _81436_ (_31430_, _31429_, _31424_);
  and _81437_ (_31431_, _31430_, _31413_);
  or _81438_ (_31432_, _31431_, _06219_);
  or _81439_ (_31435_, _31418_, _06220_);
  and _81440_ (_31436_, _31435_, _06040_);
  and _81441_ (_31437_, _31436_, _31432_);
  and _81442_ (_31438_, _14479_, _07638_);
  or _81443_ (_31439_, _31438_, _31425_);
  and _81444_ (_31440_, _31439_, _06039_);
  or _81445_ (_31441_, _31440_, _06032_);
  or _81446_ (_31442_, _31441_, _31437_);
  and _81447_ (_31443_, _31426_, _14512_);
  or _81448_ (_31444_, _31425_, _06033_);
  or _81449_ (_31445_, _31444_, _31443_);
  and _81450_ (_31446_, _31445_, _06027_);
  and _81451_ (_31447_, _31446_, _31442_);
  or _81452_ (_31448_, _31425_, _14525_);
  and _81453_ (_31449_, _31448_, _06026_);
  and _81454_ (_31450_, _31449_, _31427_);
  or _81455_ (_31451_, _31450_, _09818_);
  or _81456_ (_31452_, _31451_, _31447_);
  and _81457_ (_31453_, _09182_, _07730_);
  or _81458_ (_31454_, _31403_, _07012_);
  or _81459_ (_31457_, _31454_, _31453_);
  or _81460_ (_31458_, _31411_, _09827_);
  and _81461_ (_31459_, _31458_, _05669_);
  and _81462_ (_31460_, _31459_, _31457_);
  and _81463_ (_31461_, _31460_, _31452_);
  and _81464_ (_31462_, _14580_, _07730_);
  or _81465_ (_31463_, _31462_, _31403_);
  and _81466_ (_31464_, _31463_, _09833_);
  or _81467_ (_31465_, _31464_, _06019_);
  or _81468_ (_31466_, _31465_, _31461_);
  and _81469_ (_31467_, _31466_, _31409_);
  or _81470_ (_31468_, _31467_, _06112_);
  and _81471_ (_31469_, _14596_, _07730_);
  or _81472_ (_31470_, _31403_, _08751_);
  or _81473_ (_31471_, _31470_, _31469_);
  and _81474_ (_31472_, _31471_, _08756_);
  and _81475_ (_31473_, _31472_, _31468_);
  and _81476_ (_31474_, _10991_, _07730_);
  or _81477_ (_31475_, _31474_, _31403_);
  and _81478_ (_31476_, _31475_, _06284_);
  or _81479_ (_31479_, _31476_, _31473_);
  and _81480_ (_31480_, _31479_, _07032_);
  or _81481_ (_31481_, _31480_, _31408_);
  and _81482_ (_31482_, _31481_, _06278_);
  and _81483_ (_31483_, _31418_, _06277_);
  and _81484_ (_31484_, _31483_, _31404_);
  or _81485_ (_31485_, _31484_, _06130_);
  or _81486_ (_31486_, _31485_, _31482_);
  and _81487_ (_31487_, _14593_, _07730_);
  or _81488_ (_31488_, _31403_, _08777_);
  or _81489_ (_31489_, _31488_, _31487_);
  and _81490_ (_31490_, _31489_, _08782_);
  and _81491_ (_31491_, _31490_, _31486_);
  nor _81492_ (_31492_, _10990_, _13006_);
  or _81493_ (_31493_, _31492_, _31403_);
  and _81494_ (_31494_, _31493_, _06292_);
  or _81495_ (_31495_, _31494_, _06316_);
  or _81496_ (_31496_, _31495_, _31491_);
  or _81497_ (_31497_, _31415_, _06718_);
  and _81498_ (_31498_, _31497_, _05653_);
  and _81499_ (_31501_, _31498_, _31496_);
  and _81500_ (_31502_, _31439_, _05652_);
  or _81501_ (_31503_, _31502_, _06047_);
  or _81502_ (_31504_, _31503_, _31501_);
  and _81503_ (_31505_, _14657_, _07730_);
  or _81504_ (_31506_, _31403_, _06048_);
  or _81505_ (_31507_, _31506_, _31505_);
  and _81506_ (_31508_, _31507_, _01336_);
  and _81507_ (_31509_, _31508_, _31504_);
  or _81508_ (_43453_, _31509_, _31402_);
  and _81509_ (_31510_, _13006_, \oc8051_golden_model_1.P0 [3]);
  and _81510_ (_31511_, _07730_, _08662_);
  or _81511_ (_31512_, _31511_, _31510_);
  or _81512_ (_31513_, _31512_, _06020_);
  and _81513_ (_31514_, _14672_, _07730_);
  or _81514_ (_31515_, _31514_, _31510_);
  or _81515_ (_31516_, _31515_, _06954_);
  and _81516_ (_31517_, _07730_, \oc8051_golden_model_1.ACC [3]);
  or _81517_ (_31518_, _31517_, _31510_);
  and _81518_ (_31519_, _31518_, _06938_);
  and _81519_ (_31522_, _06939_, \oc8051_golden_model_1.P0 [3]);
  or _81520_ (_31523_, _31522_, _06102_);
  or _81521_ (_31524_, _31523_, _31519_);
  and _81522_ (_31525_, _31524_, _06044_);
  and _81523_ (_31526_, _31525_, _31516_);
  and _81524_ (_31527_, _13025_, \oc8051_golden_model_1.P0 [3]);
  and _81525_ (_31528_, _14683_, _07638_);
  or _81526_ (_31529_, _31528_, _31527_);
  and _81527_ (_31530_, _31529_, _06043_);
  or _81528_ (_31531_, _31530_, _06239_);
  or _81529_ (_31532_, _31531_, _31526_);
  nor _81530_ (_31533_, _13006_, _07353_);
  or _81531_ (_31534_, _31533_, _31510_);
  or _81532_ (_31535_, _31534_, _06848_);
  and _81533_ (_31536_, _31535_, _31532_);
  or _81534_ (_31537_, _31536_, _06219_);
  or _81535_ (_31538_, _31518_, _06220_);
  and _81536_ (_31539_, _31538_, _06040_);
  and _81537_ (_31540_, _31539_, _31537_);
  and _81538_ (_31541_, _14681_, _07638_);
  or _81539_ (_31544_, _31541_, _31527_);
  and _81540_ (_31545_, _31544_, _06039_);
  or _81541_ (_31546_, _31545_, _06032_);
  or _81542_ (_31547_, _31546_, _31540_);
  or _81543_ (_31548_, _31527_, _14708_);
  and _81544_ (_31549_, _31548_, _31529_);
  or _81545_ (_31550_, _31549_, _06033_);
  and _81546_ (_31551_, _31550_, _06027_);
  and _81547_ (_31552_, _31551_, _31547_);
  and _81548_ (_31553_, _14724_, _07638_);
  or _81549_ (_31554_, _31553_, _31527_);
  and _81550_ (_31555_, _31554_, _06026_);
  or _81551_ (_31556_, _31555_, _09818_);
  or _81552_ (_31557_, _31556_, _31552_);
  and _81553_ (_31558_, _09181_, _07730_);
  or _81554_ (_31559_, _31510_, _07012_);
  or _81555_ (_31560_, _31559_, _31558_);
  or _81556_ (_31561_, _31534_, _09827_);
  and _81557_ (_31562_, _31561_, _05669_);
  and _81558_ (_31563_, _31562_, _31560_);
  and _81559_ (_31566_, _31563_, _31557_);
  and _81560_ (_31567_, _14778_, _07730_);
  or _81561_ (_31568_, _31567_, _31510_);
  and _81562_ (_31569_, _31568_, _09833_);
  or _81563_ (_31570_, _31569_, _06019_);
  or _81564_ (_31571_, _31570_, _31566_);
  and _81565_ (_31572_, _31571_, _31513_);
  or _81566_ (_31573_, _31572_, _06112_);
  and _81567_ (_31574_, _14793_, _07730_);
  or _81568_ (_31575_, _31510_, _08751_);
  or _81569_ (_31576_, _31575_, _31574_);
  and _81570_ (_31577_, _31576_, _08756_);
  and _81571_ (_31578_, _31577_, _31573_);
  and _81572_ (_31579_, _12299_, _07730_);
  or _81573_ (_31580_, _31579_, _31510_);
  and _81574_ (_31581_, _31580_, _06284_);
  or _81575_ (_31582_, _31581_, _31578_);
  and _81576_ (_31583_, _31582_, _07032_);
  or _81577_ (_31584_, _31510_, _08029_);
  and _81578_ (_31585_, _31512_, _06108_);
  and _81579_ (_31588_, _31585_, _31584_);
  or _81580_ (_31589_, _31588_, _31583_);
  and _81581_ (_31590_, _31589_, _06278_);
  and _81582_ (_31591_, _31518_, _06277_);
  and _81583_ (_31592_, _31591_, _31584_);
  or _81584_ (_31593_, _31592_, _06130_);
  or _81585_ (_31594_, _31593_, _31590_);
  and _81586_ (_31595_, _14792_, _07730_);
  or _81587_ (_31596_, _31510_, _08777_);
  or _81588_ (_31597_, _31596_, _31595_);
  and _81589_ (_31598_, _31597_, _08782_);
  and _81590_ (_31599_, _31598_, _31594_);
  nor _81591_ (_31600_, _10988_, _13006_);
  or _81592_ (_31601_, _31600_, _31510_);
  and _81593_ (_31602_, _31601_, _06292_);
  or _81594_ (_31603_, _31602_, _06316_);
  or _81595_ (_31604_, _31603_, _31599_);
  or _81596_ (_31605_, _31515_, _06718_);
  and _81597_ (_31606_, _31605_, _05653_);
  and _81598_ (_31607_, _31606_, _31604_);
  and _81599_ (_31610_, _31544_, _05652_);
  or _81600_ (_31611_, _31610_, _06047_);
  or _81601_ (_31612_, _31611_, _31607_);
  and _81602_ (_31613_, _14849_, _07730_);
  or _81603_ (_31614_, _31510_, _06048_);
  or _81604_ (_31615_, _31614_, _31613_);
  and _81605_ (_31616_, _31615_, _01336_);
  and _81606_ (_31617_, _31616_, _31612_);
  nor _81607_ (_31618_, \oc8051_golden_model_1.P0 [3], rst);
  nor _81608_ (_31619_, _31618_, _00000_);
  or _81609_ (_43454_, _31619_, _31617_);
  nor _81610_ (_31620_, \oc8051_golden_model_1.P0 [4], rst);
  nor _81611_ (_31621_, _31620_, _00000_);
  and _81612_ (_31622_, _13006_, \oc8051_golden_model_1.P0 [4]);
  and _81613_ (_31623_, _08665_, _07730_);
  or _81614_ (_31624_, _31623_, _31622_);
  or _81615_ (_31625_, _31624_, _06020_);
  and _81616_ (_31626_, _14887_, _07730_);
  or _81617_ (_31627_, _31626_, _31622_);
  or _81618_ (_31628_, _31627_, _06954_);
  and _81619_ (_31631_, _07730_, \oc8051_golden_model_1.ACC [4]);
  or _81620_ (_31632_, _31631_, _31622_);
  and _81621_ (_31633_, _31632_, _06938_);
  and _81622_ (_31634_, _06939_, \oc8051_golden_model_1.P0 [4]);
  or _81623_ (_31635_, _31634_, _06102_);
  or _81624_ (_31636_, _31635_, _31633_);
  and _81625_ (_31637_, _31636_, _06044_);
  and _81626_ (_31638_, _31637_, _31628_);
  and _81627_ (_31639_, _13025_, \oc8051_golden_model_1.P0 [4]);
  and _81628_ (_31640_, _14878_, _07638_);
  or _81629_ (_31641_, _31640_, _31639_);
  and _81630_ (_31642_, _31641_, _06043_);
  or _81631_ (_31643_, _31642_, _06239_);
  or _81632_ (_31644_, _31643_, _31638_);
  nor _81633_ (_31645_, _08270_, _13006_);
  or _81634_ (_31646_, _31645_, _31622_);
  or _81635_ (_31647_, _31646_, _06848_);
  and _81636_ (_31648_, _31647_, _31644_);
  or _81637_ (_31649_, _31648_, _06219_);
  or _81638_ (_31650_, _31632_, _06220_);
  and _81639_ (_31653_, _31650_, _06040_);
  and _81640_ (_31654_, _31653_, _31649_);
  and _81641_ (_31655_, _14882_, _07638_);
  or _81642_ (_31656_, _31655_, _31639_);
  and _81643_ (_31657_, _31656_, _06039_);
  or _81644_ (_31658_, _31657_, _06032_);
  or _81645_ (_31659_, _31658_, _31654_);
  or _81646_ (_31660_, _31639_, _14914_);
  and _81647_ (_31661_, _31660_, _31641_);
  or _81648_ (_31662_, _31661_, _06033_);
  and _81649_ (_31663_, _31662_, _06027_);
  and _81650_ (_31664_, _31663_, _31659_);
  or _81651_ (_31665_, _31639_, _14879_);
  and _81652_ (_31666_, _31665_, _06026_);
  and _81653_ (_31667_, _31666_, _31641_);
  or _81654_ (_31668_, _31667_, _09818_);
  or _81655_ (_31669_, _31668_, _31664_);
  and _81656_ (_31670_, _09180_, _07730_);
  or _81657_ (_31671_, _31622_, _07012_);
  or _81658_ (_31672_, _31671_, _31670_);
  or _81659_ (_31675_, _31646_, _09827_);
  and _81660_ (_31676_, _31675_, _05669_);
  and _81661_ (_31677_, _31676_, _31672_);
  and _81662_ (_31678_, _31677_, _31669_);
  and _81663_ (_31679_, _14983_, _07730_);
  or _81664_ (_31680_, _31679_, _31622_);
  and _81665_ (_31681_, _31680_, _09833_);
  or _81666_ (_31682_, _31681_, _06019_);
  or _81667_ (_31683_, _31682_, _31678_);
  and _81668_ (_31684_, _31683_, _31625_);
  or _81669_ (_31685_, _31684_, _06112_);
  and _81670_ (_31686_, _14876_, _07730_);
  or _81671_ (_31687_, _31686_, _31622_);
  or _81672_ (_31688_, _31687_, _08751_);
  and _81673_ (_31689_, _31688_, _08756_);
  and _81674_ (_31690_, _31689_, _31685_);
  and _81675_ (_31691_, _10986_, _07730_);
  or _81676_ (_31692_, _31691_, _31622_);
  and _81677_ (_31693_, _31692_, _06284_);
  or _81678_ (_31694_, _31693_, _31690_);
  and _81679_ (_31697_, _31694_, _07032_);
  or _81680_ (_31698_, _31622_, _08273_);
  and _81681_ (_31699_, _31624_, _06108_);
  and _81682_ (_31700_, _31699_, _31698_);
  or _81683_ (_31701_, _31700_, _31697_);
  and _81684_ (_31702_, _31701_, _06278_);
  and _81685_ (_31703_, _31632_, _06277_);
  and _81686_ (_31704_, _31703_, _31698_);
  or _81687_ (_31705_, _31704_, _06130_);
  or _81688_ (_31706_, _31705_, _31702_);
  and _81689_ (_31707_, _14873_, _07730_);
  or _81690_ (_31708_, _31622_, _08777_);
  or _81691_ (_31709_, _31708_, _31707_);
  and _81692_ (_31710_, _31709_, _08782_);
  and _81693_ (_31711_, _31710_, _31706_);
  nor _81694_ (_31712_, _10985_, _13006_);
  or _81695_ (_31713_, _31712_, _31622_);
  and _81696_ (_31714_, _31713_, _06292_);
  or _81697_ (_31715_, _31714_, _06316_);
  or _81698_ (_31716_, _31715_, _31711_);
  or _81699_ (_31719_, _31627_, _06718_);
  and _81700_ (_31720_, _31719_, _05653_);
  and _81701_ (_31721_, _31720_, _31716_);
  and _81702_ (_31722_, _31656_, _05652_);
  or _81703_ (_31723_, _31722_, _06047_);
  or _81704_ (_31724_, _31723_, _31721_);
  and _81705_ (_31725_, _15055_, _07730_);
  or _81706_ (_31726_, _31622_, _06048_);
  or _81707_ (_31727_, _31726_, _31725_);
  and _81708_ (_31728_, _31727_, _01336_);
  and _81709_ (_31729_, _31728_, _31724_);
  or _81710_ (_43455_, _31729_, _31621_);
  and _81711_ (_31730_, _13006_, \oc8051_golden_model_1.P0 [5]);
  and _81712_ (_31731_, _08652_, _07730_);
  or _81713_ (_31732_, _31731_, _31730_);
  or _81714_ (_31733_, _31732_, _06020_);
  and _81715_ (_31734_, _15093_, _07730_);
  or _81716_ (_31735_, _31734_, _31730_);
  or _81717_ (_31736_, _31735_, _06954_);
  and _81718_ (_31737_, _07730_, \oc8051_golden_model_1.ACC [5]);
  or _81719_ (_31740_, _31737_, _31730_);
  and _81720_ (_31741_, _31740_, _06938_);
  and _81721_ (_31742_, _06939_, \oc8051_golden_model_1.P0 [5]);
  or _81722_ (_31743_, _31742_, _06102_);
  or _81723_ (_31744_, _31743_, _31741_);
  and _81724_ (_31745_, _31744_, _06044_);
  and _81725_ (_31746_, _31745_, _31736_);
  and _81726_ (_31747_, _13025_, \oc8051_golden_model_1.P0 [5]);
  and _81727_ (_31748_, _15073_, _07638_);
  or _81728_ (_31749_, _31748_, _31747_);
  and _81729_ (_31750_, _31749_, _06043_);
  or _81730_ (_31751_, _31750_, _06239_);
  or _81731_ (_31752_, _31751_, _31746_);
  nor _81732_ (_31753_, _07977_, _13006_);
  or _81733_ (_31754_, _31753_, _31730_);
  or _81734_ (_31755_, _31754_, _06848_);
  and _81735_ (_31756_, _31755_, _31752_);
  or _81736_ (_31757_, _31756_, _06219_);
  or _81737_ (_31758_, _31740_, _06220_);
  and _81738_ (_31759_, _31758_, _06040_);
  and _81739_ (_31762_, _31759_, _31757_);
  and _81740_ (_31763_, _15077_, _07638_);
  or _81741_ (_31764_, _31763_, _31747_);
  and _81742_ (_31765_, _31764_, _06039_);
  or _81743_ (_31766_, _31765_, _06032_);
  or _81744_ (_31767_, _31766_, _31762_);
  or _81745_ (_31768_, _31747_, _15110_);
  and _81746_ (_31769_, _31768_, _31749_);
  or _81747_ (_31770_, _31769_, _06033_);
  and _81748_ (_31771_, _31770_, _06027_);
  and _81749_ (_31772_, _31771_, _31767_);
  or _81750_ (_31773_, _31747_, _15074_);
  and _81751_ (_31774_, _31773_, _06026_);
  and _81752_ (_31775_, _31774_, _31749_);
  or _81753_ (_31776_, _31775_, _09818_);
  or _81754_ (_31777_, _31776_, _31772_);
  and _81755_ (_31778_, _09179_, _07730_);
  or _81756_ (_31779_, _31730_, _07012_);
  or _81757_ (_31780_, _31779_, _31778_);
  or _81758_ (_31781_, _31754_, _09827_);
  and _81759_ (_31784_, _31781_, _05669_);
  and _81760_ (_31785_, _31784_, _31780_);
  and _81761_ (_31786_, _31785_, _31777_);
  and _81762_ (_31787_, _15179_, _07730_);
  or _81763_ (_31788_, _31787_, _31730_);
  and _81764_ (_31789_, _31788_, _09833_);
  or _81765_ (_31790_, _31789_, _06019_);
  or _81766_ (_31791_, _31790_, _31786_);
  and _81767_ (_31792_, _31791_, _31733_);
  or _81768_ (_31793_, _31792_, _06112_);
  and _81769_ (_31794_, _15195_, _07730_);
  or _81770_ (_31795_, _31794_, _31730_);
  or _81771_ (_31796_, _31795_, _08751_);
  and _81772_ (_31797_, _31796_, _08756_);
  and _81773_ (_31798_, _31797_, _31793_);
  and _81774_ (_31799_, _12306_, _07730_);
  or _81775_ (_31800_, _31799_, _31730_);
  and _81776_ (_31801_, _31800_, _06284_);
  or _81777_ (_31802_, _31801_, _31798_);
  and _81778_ (_31803_, _31802_, _07032_);
  or _81779_ (_31806_, _31730_, _07980_);
  and _81780_ (_31807_, _31732_, _06108_);
  and _81781_ (_31808_, _31807_, _31806_);
  or _81782_ (_31809_, _31808_, _31803_);
  and _81783_ (_31810_, _31809_, _06278_);
  and _81784_ (_31811_, _31740_, _06277_);
  and _81785_ (_31812_, _31811_, _31806_);
  or _81786_ (_31813_, _31812_, _06130_);
  or _81787_ (_31814_, _31813_, _31810_);
  and _81788_ (_31815_, _15194_, _07730_);
  or _81789_ (_31816_, _31730_, _08777_);
  or _81790_ (_31817_, _31816_, _31815_);
  and _81791_ (_31818_, _31817_, _08782_);
  and _81792_ (_31819_, _31818_, _31814_);
  nor _81793_ (_31820_, _10982_, _13006_);
  or _81794_ (_31821_, _31820_, _31730_);
  and _81795_ (_31822_, _31821_, _06292_);
  or _81796_ (_31823_, _31822_, _06316_);
  or _81797_ (_31824_, _31823_, _31819_);
  or _81798_ (_31825_, _31735_, _06718_);
  and _81799_ (_31828_, _31825_, _05653_);
  and _81800_ (_31829_, _31828_, _31824_);
  and _81801_ (_31830_, _31764_, _05652_);
  or _81802_ (_31831_, _31830_, _06047_);
  or _81803_ (_31832_, _31831_, _31829_);
  and _81804_ (_31833_, _15253_, _07730_);
  or _81805_ (_31834_, _31730_, _06048_);
  or _81806_ (_31835_, _31834_, _31833_);
  and _81807_ (_31836_, _31835_, _01336_);
  and _81808_ (_31837_, _31836_, _31832_);
  nor _81809_ (_31838_, \oc8051_golden_model_1.P0 [5], rst);
  nor _81810_ (_31839_, _31838_, _00000_);
  or _81811_ (_43456_, _31839_, _31837_);
  nor _81812_ (_31840_, \oc8051_golden_model_1.P0 [6], rst);
  nor _81813_ (_31841_, _31840_, _00000_);
  and _81814_ (_31842_, _13006_, \oc8051_golden_model_1.P0 [6]);
  and _81815_ (_31843_, _15389_, _07730_);
  or _81816_ (_31844_, _31843_, _31842_);
  or _81817_ (_31845_, _31844_, _06020_);
  and _81818_ (_31846_, _15293_, _07730_);
  or _81819_ (_31849_, _31846_, _31842_);
  or _81820_ (_31850_, _31849_, _06954_);
  and _81821_ (_31851_, _07730_, \oc8051_golden_model_1.ACC [6]);
  or _81822_ (_31852_, _31851_, _31842_);
  and _81823_ (_31853_, _31852_, _06938_);
  and _81824_ (_31854_, _06939_, \oc8051_golden_model_1.P0 [6]);
  or _81825_ (_31855_, _31854_, _06102_);
  or _81826_ (_31856_, _31855_, _31853_);
  and _81827_ (_31857_, _31856_, _06044_);
  and _81828_ (_31858_, _31857_, _31850_);
  and _81829_ (_31860_, _13025_, \oc8051_golden_model_1.P0 [6]);
  and _81830_ (_31861_, _15280_, _07638_);
  or _81831_ (_31862_, _31861_, _31860_);
  and _81832_ (_31863_, _31862_, _06043_);
  or _81833_ (_31864_, _31863_, _06239_);
  or _81834_ (_31865_, _31864_, _31858_);
  nor _81835_ (_31866_, _07883_, _13006_);
  or _81836_ (_31867_, _31866_, _31842_);
  or _81837_ (_31868_, _31867_, _06848_);
  and _81838_ (_31869_, _31868_, _31865_);
  or _81839_ (_31871_, _31869_, _06219_);
  or _81840_ (_31872_, _31852_, _06220_);
  and _81841_ (_31873_, _31872_, _06040_);
  and _81842_ (_31874_, _31873_, _31871_);
  and _81843_ (_31875_, _15278_, _07638_);
  or _81844_ (_31876_, _31875_, _31860_);
  and _81845_ (_31877_, _31876_, _06039_);
  or _81846_ (_31878_, _31877_, _06032_);
  or _81847_ (_31879_, _31878_, _31874_);
  or _81848_ (_31880_, _31860_, _15310_);
  and _81849_ (_31882_, _31880_, _31862_);
  or _81850_ (_31883_, _31882_, _06033_);
  and _81851_ (_31884_, _31883_, _06027_);
  and _81852_ (_31885_, _31884_, _31879_);
  or _81853_ (_31886_, _31860_, _15326_);
  and _81854_ (_31887_, _31886_, _06026_);
  and _81855_ (_31888_, _31887_, _31862_);
  or _81856_ (_31889_, _31888_, _09818_);
  or _81857_ (_31890_, _31889_, _31885_);
  and _81858_ (_31891_, _09178_, _07730_);
  or _81859_ (_31893_, _31842_, _07012_);
  or _81860_ (_31894_, _31893_, _31891_);
  or _81861_ (_31895_, _31867_, _09827_);
  and _81862_ (_31896_, _31895_, _05669_);
  and _81863_ (_31897_, _31896_, _31894_);
  and _81864_ (_31898_, _31897_, _31890_);
  and _81865_ (_31899_, _15382_, _07730_);
  or _81866_ (_31900_, _31899_, _31842_);
  and _81867_ (_31901_, _31900_, _09833_);
  or _81868_ (_31902_, _31901_, _06019_);
  or _81869_ (_31904_, _31902_, _31898_);
  and _81870_ (_31905_, _31904_, _31845_);
  or _81871_ (_31906_, _31905_, _06112_);
  and _81872_ (_31907_, _15399_, _07730_);
  or _81873_ (_31908_, _31842_, _08751_);
  or _81874_ (_31909_, _31908_, _31907_);
  and _81875_ (_31910_, _31909_, _08756_);
  and _81876_ (_31911_, _31910_, _31906_);
  and _81877_ (_31912_, _10980_, _07730_);
  or _81878_ (_31913_, _31912_, _31842_);
  and _81879_ (_31915_, _31913_, _06284_);
  or _81880_ (_31916_, _31915_, _31911_);
  and _81881_ (_31917_, _31916_, _07032_);
  or _81882_ (_31918_, _31842_, _07886_);
  and _81883_ (_31919_, _31844_, _06108_);
  and _81884_ (_31920_, _31919_, _31918_);
  or _81885_ (_31921_, _31920_, _31917_);
  and _81886_ (_31922_, _31921_, _06278_);
  and _81887_ (_31923_, _31852_, _06277_);
  and _81888_ (_31924_, _31923_, _31918_);
  or _81889_ (_31925_, _31924_, _06130_);
  or _81890_ (_31926_, _31925_, _31922_);
  and _81891_ (_31927_, _15396_, _07730_);
  or _81892_ (_31928_, _31842_, _08777_);
  or _81893_ (_31929_, _31928_, _31927_);
  and _81894_ (_31930_, _31929_, _08782_);
  and _81895_ (_31931_, _31930_, _31926_);
  nor _81896_ (_31932_, _10979_, _13006_);
  or _81897_ (_31933_, _31932_, _31842_);
  and _81898_ (_31934_, _31933_, _06292_);
  or _81899_ (_31936_, _31934_, _06316_);
  or _81900_ (_31937_, _31936_, _31931_);
  or _81901_ (_31938_, _31849_, _06718_);
  and _81902_ (_31939_, _31938_, _05653_);
  and _81903_ (_31940_, _31939_, _31937_);
  and _81904_ (_31941_, _31876_, _05652_);
  or _81905_ (_31942_, _31941_, _06047_);
  or _81906_ (_31943_, _31942_, _31940_);
  and _81907_ (_31944_, _15451_, _07730_);
  or _81908_ (_31945_, _31842_, _06048_);
  or _81909_ (_31947_, _31945_, _31944_);
  and _81910_ (_31948_, _31947_, _01336_);
  and _81911_ (_31949_, _31948_, _31943_);
  or _81912_ (_43457_, _31949_, _31841_);
  nor _81913_ (_31950_, \oc8051_golden_model_1.P1 [0], rst);
  nor _81914_ (_31951_, _31950_, _00000_);
  and _81915_ (_31952_, _07677_, \oc8051_golden_model_1.ACC [0]);
  and _81916_ (_31953_, _31952_, _08127_);
  and _81917_ (_31954_, _13108_, \oc8051_golden_model_1.P1 [0]);
  or _81918_ (_31955_, _31954_, _06278_);
  or _81919_ (_31957_, _31955_, _31953_);
  and _81920_ (_31958_, _07677_, _08672_);
  or _81921_ (_31959_, _31958_, _31954_);
  or _81922_ (_31960_, _31959_, _06020_);
  and _81923_ (_31961_, _09120_, _07677_);
  or _81924_ (_31962_, _31954_, _07012_);
  or _81925_ (_31963_, _31962_, _31961_);
  nor _81926_ (_31964_, _08127_, _13108_);
  or _81927_ (_31965_, _31964_, _31954_);
  and _81928_ (_31966_, _31965_, _06102_);
  and _81929_ (_31968_, _06939_, \oc8051_golden_model_1.P1 [0]);
  or _81930_ (_31969_, _31952_, _31954_);
  and _81931_ (_31970_, _31969_, _06938_);
  or _81932_ (_31971_, _31970_, _31968_);
  and _81933_ (_31972_, _31971_, _06954_);
  or _81934_ (_31973_, _31972_, _06043_);
  or _81935_ (_31974_, _31973_, _31966_);
  and _81936_ (_31975_, _14102_, _08345_);
  and _81937_ (_31976_, _13127_, \oc8051_golden_model_1.P1 [0]);
  or _81938_ (_31977_, _31976_, _06044_);
  or _81939_ (_31979_, _31977_, _31975_);
  and _81940_ (_31980_, _31979_, _06848_);
  and _81941_ (_31981_, _31980_, _31974_);
  and _81942_ (_31982_, _07677_, _06931_);
  or _81943_ (_31983_, _31982_, _31954_);
  and _81944_ (_31984_, _31983_, _06239_);
  or _81945_ (_31985_, _31984_, _06219_);
  or _81946_ (_31986_, _31985_, _31981_);
  or _81947_ (_31987_, _31969_, _06220_);
  and _81948_ (_31988_, _31987_, _06040_);
  and _81949_ (_31990_, _31988_, _31986_);
  and _81950_ (_31991_, _31954_, _06039_);
  or _81951_ (_31992_, _31991_, _06032_);
  or _81952_ (_31993_, _31992_, _31990_);
  or _81953_ (_31994_, _31965_, _06033_);
  and _81954_ (_31995_, _31994_, _06027_);
  and _81955_ (_31996_, _31995_, _31993_);
  and _81956_ (_31997_, _14132_, _08345_);
  or _81957_ (_31998_, _31997_, _31976_);
  and _81958_ (_31999_, _31998_, _06026_);
  or _81959_ (_32001_, _31999_, _09818_);
  or _81960_ (_32002_, _32001_, _31996_);
  or _81961_ (_32003_, _31983_, _09827_);
  and _81962_ (_32004_, _32003_, _05669_);
  and _81963_ (_32005_, _32004_, _32002_);
  and _81964_ (_32006_, _32005_, _31963_);
  and _81965_ (_32007_, _14186_, _07677_);
  or _81966_ (_32008_, _32007_, _31954_);
  and _81967_ (_32009_, _32008_, _09833_);
  or _81968_ (_32010_, _32009_, _06019_);
  or _81969_ (_32012_, _32010_, _32006_);
  and _81970_ (_32013_, _32012_, _31960_);
  or _81971_ (_32014_, _32013_, _06112_);
  and _81972_ (_32015_, _14086_, _07677_);
  or _81973_ (_32016_, _32015_, _31954_);
  or _81974_ (_32017_, _32016_, _08751_);
  and _81975_ (_32018_, _32017_, _08756_);
  and _81976_ (_32019_, _32018_, _32014_);
  nor _81977_ (_32020_, _12302_, _13108_);
  or _81978_ (_32021_, _32020_, _31954_);
  nor _81979_ (_32023_, _31953_, _08756_);
  and _81980_ (_32024_, _32023_, _32021_);
  or _81981_ (_32025_, _32024_, _32019_);
  and _81982_ (_32026_, _32025_, _07032_);
  nand _81983_ (_32027_, _31959_, _06108_);
  nor _81984_ (_32028_, _32027_, _31964_);
  or _81985_ (_32029_, _32028_, _06277_);
  or _81986_ (_32030_, _32029_, _32026_);
  and _81987_ (_32031_, _32030_, _31957_);
  or _81988_ (_32032_, _32031_, _06130_);
  and _81989_ (_32034_, _14083_, _07677_);
  or _81990_ (_32035_, _31954_, _08777_);
  or _81991_ (_32036_, _32035_, _32034_);
  and _81992_ (_32037_, _32036_, _08782_);
  and _81993_ (_32038_, _32037_, _32032_);
  and _81994_ (_32039_, _32021_, _06292_);
  or _81995_ (_32040_, _32039_, _06316_);
  or _81996_ (_32041_, _32040_, _32038_);
  or _81997_ (_32042_, _31965_, _06718_);
  and _81998_ (_32043_, _32042_, _32041_);
  or _81999_ (_32045_, _32043_, _05652_);
  or _82000_ (_32046_, _31954_, _05653_);
  and _82001_ (_32047_, _32046_, _32045_);
  or _82002_ (_32048_, _32047_, _06047_);
  or _82003_ (_32049_, _31965_, _06048_);
  and _82004_ (_32050_, _32049_, _01336_);
  and _82005_ (_32051_, _32050_, _32048_);
  or _82006_ (_43459_, _32051_, _31951_);
  and _82007_ (_32052_, _13108_, \oc8051_golden_model_1.P1 [1]);
  nor _82008_ (_32053_, _10993_, _13108_);
  or _82009_ (_32055_, _32053_, _32052_);
  or _82010_ (_32056_, _32055_, _08782_);
  or _82011_ (_32057_, _14367_, _13108_);
  or _82012_ (_32058_, _07677_, \oc8051_golden_model_1.P1 [1]);
  and _82013_ (_32059_, _32058_, _09833_);
  and _82014_ (_32060_, _32059_, _32057_);
  nor _82015_ (_32061_, _13108_, _07132_);
  or _82016_ (_32062_, _32061_, _32052_);
  and _82017_ (_32063_, _32062_, _06239_);
  and _82018_ (_32064_, _13127_, \oc8051_golden_model_1.P1 [1]);
  and _82019_ (_32066_, _14266_, _08345_);
  or _82020_ (_32067_, _32066_, _32064_);
  or _82021_ (_32068_, _32067_, _06044_);
  and _82022_ (_32069_, _14284_, _07677_);
  not _82023_ (_32070_, _32069_);
  and _82024_ (_32071_, _32070_, _32058_);
  and _82025_ (_32072_, _32071_, _06102_);
  and _82026_ (_32073_, _06939_, \oc8051_golden_model_1.P1 [1]);
  and _82027_ (_32074_, _07677_, \oc8051_golden_model_1.ACC [1]);
  or _82028_ (_32075_, _32074_, _32052_);
  and _82029_ (_32077_, _32075_, _06938_);
  or _82030_ (_32078_, _32077_, _32073_);
  and _82031_ (_32079_, _32078_, _06954_);
  or _82032_ (_32080_, _32079_, _06043_);
  or _82033_ (_32081_, _32080_, _32072_);
  and _82034_ (_32082_, _32081_, _32068_);
  and _82035_ (_32083_, _32082_, _06848_);
  or _82036_ (_32084_, _32083_, _32063_);
  or _82037_ (_32085_, _32084_, _06219_);
  or _82038_ (_32086_, _32075_, _06220_);
  and _82039_ (_32088_, _32086_, _06040_);
  and _82040_ (_32089_, _32088_, _32085_);
  and _82041_ (_32090_, _14273_, _08345_);
  or _82042_ (_32091_, _32090_, _32064_);
  and _82043_ (_32092_, _32091_, _06039_);
  or _82044_ (_32093_, _32092_, _06032_);
  or _82045_ (_32094_, _32093_, _32089_);
  or _82046_ (_32095_, _32064_, _14302_);
  and _82047_ (_32096_, _32095_, _32067_);
  or _82048_ (_32097_, _32096_, _06033_);
  and _82049_ (_32099_, _32097_, _06027_);
  and _82050_ (_32100_, _32099_, _32094_);
  or _82051_ (_32101_, _32064_, _14267_);
  and _82052_ (_32102_, _32101_, _06026_);
  and _82053_ (_32103_, _32102_, _32067_);
  or _82054_ (_32104_, _32103_, _09815_);
  or _82055_ (_32105_, _32104_, _32100_);
  or _82056_ (_32106_, _32062_, _09827_);
  and _82057_ (_32107_, _32106_, _32105_);
  or _82058_ (_32108_, _32107_, _07011_);
  and _82059_ (_32110_, _09075_, _07677_);
  or _82060_ (_32111_, _32052_, _07012_);
  or _82061_ (_32112_, _32111_, _32110_);
  and _82062_ (_32113_, _32112_, _05669_);
  and _82063_ (_32114_, _32113_, _32108_);
  or _82064_ (_32115_, _32114_, _32060_);
  and _82065_ (_32116_, _32115_, _06020_);
  nand _82066_ (_32117_, _07677_, _06832_);
  and _82067_ (_32118_, _32058_, _06019_);
  and _82068_ (_32119_, _32118_, _32117_);
  or _82069_ (_32121_, _32119_, _32116_);
  and _82070_ (_32122_, _32121_, _08751_);
  or _82071_ (_32123_, _14263_, _13108_);
  and _82072_ (_32124_, _32058_, _06112_);
  and _82073_ (_32125_, _32124_, _32123_);
  or _82074_ (_32126_, _32125_, _06284_);
  or _82075_ (_32127_, _32126_, _32122_);
  nand _82076_ (_32128_, _10992_, _07677_);
  and _82077_ (_32129_, _32128_, _32055_);
  or _82078_ (_32130_, _32129_, _08756_);
  and _82079_ (_32132_, _32130_, _07032_);
  and _82080_ (_32133_, _32132_, _32127_);
  or _82081_ (_32134_, _14261_, _13108_);
  and _82082_ (_32135_, _32058_, _06108_);
  and _82083_ (_32136_, _32135_, _32134_);
  or _82084_ (_32137_, _32136_, _06277_);
  or _82085_ (_32138_, _32137_, _32133_);
  nor _82086_ (_32139_, _32052_, _06278_);
  nand _82087_ (_32140_, _32139_, _32128_);
  and _82088_ (_32141_, _32140_, _08777_);
  and _82089_ (_32143_, _32141_, _32138_);
  or _82090_ (_32144_, _32117_, _08078_);
  and _82091_ (_32145_, _32058_, _06130_);
  and _82092_ (_32146_, _32145_, _32144_);
  or _82093_ (_32147_, _32146_, _06292_);
  or _82094_ (_32148_, _32147_, _32143_);
  and _82095_ (_32149_, _32148_, _32056_);
  or _82096_ (_32150_, _32149_, _06316_);
  or _82097_ (_32151_, _32071_, _06718_);
  and _82098_ (_32152_, _32151_, _05653_);
  and _82099_ (_32154_, _32152_, _32150_);
  and _82100_ (_32155_, _32091_, _05652_);
  or _82101_ (_32156_, _32155_, _06047_);
  or _82102_ (_32157_, _32156_, _32154_);
  or _82103_ (_32158_, _32052_, _06048_);
  or _82104_ (_32159_, _32158_, _32069_);
  and _82105_ (_32160_, _32159_, _01336_);
  and _82106_ (_32161_, _32160_, _32157_);
  nor _82107_ (_32162_, \oc8051_golden_model_1.P1 [1], rst);
  nor _82108_ (_32163_, _32162_, _00000_);
  or _82109_ (_43460_, _32163_, _32161_);
  nor _82110_ (_32165_, \oc8051_golden_model_1.P1 [2], rst);
  nor _82111_ (_32166_, _32165_, _00000_);
  and _82112_ (_32167_, _13108_, \oc8051_golden_model_1.P1 [2]);
  and _82113_ (_32168_, _07677_, _08730_);
  or _82114_ (_32169_, _32168_, _32167_);
  or _82115_ (_32170_, _32169_, _06020_);
  nor _82116_ (_32171_, _13108_, _07530_);
  or _82117_ (_32172_, _32171_, _32167_);
  and _82118_ (_32173_, _32172_, _06239_);
  and _82119_ (_32175_, _13127_, \oc8051_golden_model_1.P1 [2]);
  and _82120_ (_32176_, _14497_, _08345_);
  or _82121_ (_32177_, _32176_, _32175_);
  or _82122_ (_32178_, _32177_, _06044_);
  and _82123_ (_32179_, _14493_, _07677_);
  or _82124_ (_32180_, _32179_, _32167_);
  and _82125_ (_32181_, _32180_, _06102_);
  and _82126_ (_32182_, _06939_, \oc8051_golden_model_1.P1 [2]);
  and _82127_ (_32183_, _07677_, \oc8051_golden_model_1.ACC [2]);
  or _82128_ (_32184_, _32183_, _32167_);
  and _82129_ (_32186_, _32184_, _06938_);
  or _82130_ (_32187_, _32186_, _32182_);
  and _82131_ (_32188_, _32187_, _06954_);
  or _82132_ (_32189_, _32188_, _06043_);
  or _82133_ (_32190_, _32189_, _32181_);
  and _82134_ (_32191_, _32190_, _32178_);
  and _82135_ (_32192_, _32191_, _06848_);
  or _82136_ (_32193_, _32192_, _32173_);
  or _82137_ (_32194_, _32193_, _06219_);
  or _82138_ (_32195_, _32184_, _06220_);
  and _82139_ (_32197_, _32195_, _06040_);
  and _82140_ (_32198_, _32197_, _32194_);
  and _82141_ (_32199_, _14479_, _08345_);
  or _82142_ (_32200_, _32199_, _32175_);
  and _82143_ (_32201_, _32200_, _06039_);
  or _82144_ (_32202_, _32201_, _06032_);
  or _82145_ (_32203_, _32202_, _32198_);
  or _82146_ (_32204_, _32175_, _14512_);
  and _82147_ (_32205_, _32204_, _32177_);
  or _82148_ (_32206_, _32205_, _06033_);
  and _82149_ (_32208_, _32206_, _06027_);
  and _82150_ (_32209_, _32208_, _32203_);
  or _82151_ (_32210_, _32175_, _14525_);
  and _82152_ (_32211_, _32210_, _06026_);
  and _82153_ (_32212_, _32211_, _32177_);
  or _82154_ (_32213_, _32212_, _09818_);
  or _82155_ (_32214_, _32213_, _32209_);
  and _82156_ (_32215_, _09182_, _07677_);
  or _82157_ (_32216_, _32167_, _07012_);
  or _82158_ (_32217_, _32216_, _32215_);
  or _82159_ (_32219_, _32172_, _09827_);
  and _82160_ (_32220_, _32219_, _05669_);
  and _82161_ (_32221_, _32220_, _32217_);
  and _82162_ (_32222_, _32221_, _32214_);
  and _82163_ (_32223_, _14580_, _07677_);
  or _82164_ (_32224_, _32223_, _32167_);
  and _82165_ (_32225_, _32224_, _09833_);
  or _82166_ (_32226_, _32225_, _06019_);
  or _82167_ (_32227_, _32226_, _32222_);
  and _82168_ (_32228_, _32227_, _32170_);
  or _82169_ (_32230_, _32228_, _06112_);
  and _82170_ (_32231_, _14596_, _07677_);
  or _82171_ (_32232_, _32167_, _08751_);
  or _82172_ (_32233_, _32232_, _32231_);
  and _82173_ (_32234_, _32233_, _08756_);
  and _82174_ (_32235_, _32234_, _32230_);
  and _82175_ (_32236_, _10991_, _07677_);
  or _82176_ (_32237_, _32236_, _32167_);
  and _82177_ (_32238_, _32237_, _06284_);
  or _82178_ (_32239_, _32238_, _32235_);
  and _82179_ (_32241_, _32239_, _07032_);
  or _82180_ (_32242_, _32167_, _08177_);
  and _82181_ (_32243_, _32169_, _06108_);
  and _82182_ (_32244_, _32243_, _32242_);
  or _82183_ (_32245_, _32244_, _32241_);
  and _82184_ (_32246_, _32245_, _06278_);
  and _82185_ (_32247_, _32184_, _06277_);
  and _82186_ (_32248_, _32247_, _32242_);
  or _82187_ (_32249_, _32248_, _06130_);
  or _82188_ (_32250_, _32249_, _32246_);
  and _82189_ (_32252_, _14593_, _07677_);
  or _82190_ (_32253_, _32167_, _08777_);
  or _82191_ (_32254_, _32253_, _32252_);
  and _82192_ (_32255_, _32254_, _08782_);
  and _82193_ (_32256_, _32255_, _32250_);
  nor _82194_ (_32257_, _10990_, _13108_);
  or _82195_ (_32258_, _32257_, _32167_);
  and _82196_ (_32259_, _32258_, _06292_);
  or _82197_ (_32260_, _32259_, _06316_);
  or _82198_ (_32261_, _32260_, _32256_);
  or _82199_ (_32263_, _32180_, _06718_);
  and _82200_ (_32264_, _32263_, _05653_);
  and _82201_ (_32265_, _32264_, _32261_);
  and _82202_ (_32266_, _32200_, _05652_);
  or _82203_ (_32267_, _32266_, _06047_);
  or _82204_ (_32268_, _32267_, _32265_);
  and _82205_ (_32269_, _14657_, _07677_);
  or _82206_ (_32270_, _32167_, _06048_);
  or _82207_ (_32271_, _32270_, _32269_);
  and _82208_ (_32272_, _32271_, _01336_);
  and _82209_ (_32274_, _32272_, _32268_);
  or _82210_ (_43461_, _32274_, _32166_);
  and _82211_ (_32275_, _13108_, \oc8051_golden_model_1.P1 [3]);
  and _82212_ (_32276_, _07677_, _08662_);
  or _82213_ (_32277_, _32276_, _32275_);
  or _82214_ (_32278_, _32277_, _06020_);
  and _82215_ (_32279_, _14672_, _07677_);
  or _82216_ (_32280_, _32279_, _32275_);
  or _82217_ (_32281_, _32280_, _06954_);
  and _82218_ (_32282_, _07677_, \oc8051_golden_model_1.ACC [3]);
  or _82219_ (_32284_, _32282_, _32275_);
  and _82220_ (_32285_, _32284_, _06938_);
  and _82221_ (_32286_, _06939_, \oc8051_golden_model_1.P1 [3]);
  or _82222_ (_32287_, _32286_, _06102_);
  or _82223_ (_32288_, _32287_, _32285_);
  and _82224_ (_32289_, _32288_, _06044_);
  and _82225_ (_32290_, _32289_, _32281_);
  and _82226_ (_32291_, _13127_, \oc8051_golden_model_1.P1 [3]);
  and _82227_ (_32292_, _14683_, _08345_);
  or _82228_ (_32293_, _32292_, _32291_);
  and _82229_ (_32295_, _32293_, _06043_);
  or _82230_ (_32296_, _32295_, _06239_);
  or _82231_ (_32297_, _32296_, _32290_);
  nor _82232_ (_32298_, _13108_, _07353_);
  or _82233_ (_32299_, _32298_, _32275_);
  or _82234_ (_32300_, _32299_, _06848_);
  and _82235_ (_32301_, _32300_, _32297_);
  or _82236_ (_32302_, _32301_, _06219_);
  or _82237_ (_32303_, _32284_, _06220_);
  and _82238_ (_32304_, _32303_, _06040_);
  and _82239_ (_32306_, _32304_, _32302_);
  and _82240_ (_32307_, _14681_, _08345_);
  or _82241_ (_32308_, _32307_, _32291_);
  and _82242_ (_32309_, _32308_, _06039_);
  or _82243_ (_32310_, _32309_, _06032_);
  or _82244_ (_32311_, _32310_, _32306_);
  or _82245_ (_32312_, _32291_, _14708_);
  and _82246_ (_32313_, _32312_, _32293_);
  or _82247_ (_32314_, _32313_, _06033_);
  and _82248_ (_32315_, _32314_, _06027_);
  and _82249_ (_32317_, _32315_, _32311_);
  and _82250_ (_32318_, _14724_, _08345_);
  or _82251_ (_32319_, _32318_, _32291_);
  and _82252_ (_32320_, _32319_, _06026_);
  or _82253_ (_32321_, _32320_, _09818_);
  or _82254_ (_32322_, _32321_, _32317_);
  and _82255_ (_32323_, _09181_, _07677_);
  or _82256_ (_32324_, _32275_, _07012_);
  or _82257_ (_32325_, _32324_, _32323_);
  or _82258_ (_32326_, _32299_, _09827_);
  and _82259_ (_32328_, _32326_, _05669_);
  and _82260_ (_32329_, _32328_, _32325_);
  and _82261_ (_32330_, _32329_, _32322_);
  and _82262_ (_32331_, _14778_, _07677_);
  or _82263_ (_32332_, _32331_, _32275_);
  and _82264_ (_32333_, _32332_, _09833_);
  or _82265_ (_32334_, _32333_, _06019_);
  or _82266_ (_32335_, _32334_, _32330_);
  and _82267_ (_32336_, _32335_, _32278_);
  or _82268_ (_32337_, _32336_, _06112_);
  and _82269_ (_32339_, _14793_, _07677_);
  or _82270_ (_32340_, _32275_, _08751_);
  or _82271_ (_32341_, _32340_, _32339_);
  and _82272_ (_32342_, _32341_, _08756_);
  and _82273_ (_32343_, _32342_, _32337_);
  and _82274_ (_32344_, _12299_, _07677_);
  or _82275_ (_32345_, _32344_, _32275_);
  and _82276_ (_32346_, _32345_, _06284_);
  or _82277_ (_32347_, _32346_, _32343_);
  and _82278_ (_32348_, _32347_, _07032_);
  or _82279_ (_32350_, _32275_, _08029_);
  and _82280_ (_32351_, _32277_, _06108_);
  and _82281_ (_32352_, _32351_, _32350_);
  or _82282_ (_32353_, _32352_, _32348_);
  and _82283_ (_32354_, _32353_, _06278_);
  and _82284_ (_32355_, _32284_, _06277_);
  and _82285_ (_32356_, _32355_, _32350_);
  or _82286_ (_32357_, _32356_, _06130_);
  or _82287_ (_32358_, _32357_, _32354_);
  and _82288_ (_32359_, _14792_, _07677_);
  or _82289_ (_32361_, _32275_, _08777_);
  or _82290_ (_32362_, _32361_, _32359_);
  and _82291_ (_32363_, _32362_, _08782_);
  and _82292_ (_32364_, _32363_, _32358_);
  nor _82293_ (_32365_, _10988_, _13108_);
  or _82294_ (_32366_, _32365_, _32275_);
  and _82295_ (_32367_, _32366_, _06292_);
  or _82296_ (_32368_, _32367_, _06316_);
  or _82297_ (_32369_, _32368_, _32364_);
  or _82298_ (_32370_, _32280_, _06718_);
  and _82299_ (_32372_, _32370_, _05653_);
  and _82300_ (_32373_, _32372_, _32369_);
  and _82301_ (_32374_, _32308_, _05652_);
  or _82302_ (_32375_, _32374_, _06047_);
  or _82303_ (_32376_, _32375_, _32373_);
  and _82304_ (_32377_, _14849_, _07677_);
  or _82305_ (_32378_, _32275_, _06048_);
  or _82306_ (_32379_, _32378_, _32377_);
  and _82307_ (_32380_, _32379_, _01336_);
  and _82308_ (_32381_, _32380_, _32376_);
  nor _82309_ (_32383_, \oc8051_golden_model_1.P1 [3], rst);
  nor _82310_ (_32384_, _32383_, _00000_);
  or _82311_ (_43463_, _32384_, _32381_);
  and _82312_ (_32385_, _13108_, \oc8051_golden_model_1.P1 [4]);
  and _82313_ (_32386_, _08665_, _07677_);
  or _82314_ (_32387_, _32386_, _32385_);
  or _82315_ (_32388_, _32387_, _06020_);
  and _82316_ (_32389_, _14887_, _07677_);
  or _82317_ (_32390_, _32389_, _32385_);
  or _82318_ (_32391_, _32390_, _06954_);
  and _82319_ (_32393_, _07677_, \oc8051_golden_model_1.ACC [4]);
  or _82320_ (_32394_, _32393_, _32385_);
  and _82321_ (_32395_, _32394_, _06938_);
  and _82322_ (_32396_, _06939_, \oc8051_golden_model_1.P1 [4]);
  or _82323_ (_32397_, _32396_, _06102_);
  or _82324_ (_32398_, _32397_, _32395_);
  and _82325_ (_32399_, _32398_, _06044_);
  and _82326_ (_32400_, _32399_, _32391_);
  and _82327_ (_32401_, _13127_, \oc8051_golden_model_1.P1 [4]);
  and _82328_ (_32402_, _14878_, _08345_);
  or _82329_ (_32404_, _32402_, _32401_);
  and _82330_ (_32405_, _32404_, _06043_);
  or _82331_ (_32406_, _32405_, _06239_);
  or _82332_ (_32407_, _32406_, _32400_);
  nor _82333_ (_32408_, _08270_, _13108_);
  or _82334_ (_32409_, _32408_, _32385_);
  or _82335_ (_32410_, _32409_, _06848_);
  and _82336_ (_32411_, _32410_, _32407_);
  or _82337_ (_32412_, _32411_, _06219_);
  or _82338_ (_32413_, _32394_, _06220_);
  and _82339_ (_32415_, _32413_, _06040_);
  and _82340_ (_32416_, _32415_, _32412_);
  and _82341_ (_32417_, _14882_, _08345_);
  or _82342_ (_32418_, _32417_, _32401_);
  and _82343_ (_32419_, _32418_, _06039_);
  or _82344_ (_32420_, _32419_, _06032_);
  or _82345_ (_32421_, _32420_, _32416_);
  or _82346_ (_32422_, _32401_, _14914_);
  and _82347_ (_32423_, _32422_, _32404_);
  or _82348_ (_32424_, _32423_, _06033_);
  and _82349_ (_32426_, _32424_, _06027_);
  and _82350_ (_32427_, _32426_, _32421_);
  or _82351_ (_32428_, _32401_, _14879_);
  and _82352_ (_32429_, _32428_, _06026_);
  and _82353_ (_32430_, _32429_, _32404_);
  or _82354_ (_32431_, _32430_, _09818_);
  or _82355_ (_32432_, _32431_, _32427_);
  and _82356_ (_32433_, _09180_, _07677_);
  or _82357_ (_32434_, _32385_, _07012_);
  or _82358_ (_32435_, _32434_, _32433_);
  or _82359_ (_32437_, _32409_, _09827_);
  and _82360_ (_32438_, _32437_, _05669_);
  and _82361_ (_32439_, _32438_, _32435_);
  and _82362_ (_32440_, _32439_, _32432_);
  and _82363_ (_32441_, _14983_, _07677_);
  or _82364_ (_32442_, _32441_, _32385_);
  and _82365_ (_32443_, _32442_, _09833_);
  or _82366_ (_32444_, _32443_, _06019_);
  or _82367_ (_32445_, _32444_, _32440_);
  and _82368_ (_32446_, _32445_, _32388_);
  or _82369_ (_32448_, _32446_, _06112_);
  and _82370_ (_32449_, _14876_, _07677_);
  or _82371_ (_32450_, _32449_, _32385_);
  or _82372_ (_32451_, _32450_, _08751_);
  and _82373_ (_32452_, _32451_, _08756_);
  and _82374_ (_32453_, _32452_, _32448_);
  and _82375_ (_32454_, _10986_, _07677_);
  or _82376_ (_32455_, _32454_, _32385_);
  and _82377_ (_32456_, _32455_, _06284_);
  or _82378_ (_32457_, _32456_, _32453_);
  and _82379_ (_32459_, _32457_, _07032_);
  or _82380_ (_32460_, _32385_, _08273_);
  and _82381_ (_32461_, _32387_, _06108_);
  and _82382_ (_32462_, _32461_, _32460_);
  or _82383_ (_32463_, _32462_, _32459_);
  and _82384_ (_32464_, _32463_, _06278_);
  and _82385_ (_32465_, _32394_, _06277_);
  and _82386_ (_32466_, _32465_, _32460_);
  or _82387_ (_32467_, _32466_, _06130_);
  or _82388_ (_32468_, _32467_, _32464_);
  and _82389_ (_32470_, _14873_, _07677_);
  or _82390_ (_32471_, _32385_, _08777_);
  or _82391_ (_32472_, _32471_, _32470_);
  and _82392_ (_32473_, _32472_, _08782_);
  and _82393_ (_32474_, _32473_, _32468_);
  nor _82394_ (_32475_, _10985_, _13108_);
  or _82395_ (_32476_, _32475_, _32385_);
  and _82396_ (_32477_, _32476_, _06292_);
  or _82397_ (_32478_, _32477_, _06316_);
  or _82398_ (_32479_, _32478_, _32474_);
  or _82399_ (_32481_, _32390_, _06718_);
  and _82400_ (_32482_, _32481_, _05653_);
  and _82401_ (_32483_, _32482_, _32479_);
  and _82402_ (_32484_, _32418_, _05652_);
  or _82403_ (_32485_, _32484_, _06047_);
  or _82404_ (_32486_, _32485_, _32483_);
  and _82405_ (_32487_, _15055_, _07677_);
  or _82406_ (_32488_, _32385_, _06048_);
  or _82407_ (_32489_, _32488_, _32487_);
  and _82408_ (_32490_, _32489_, _01336_);
  and _82409_ (_32492_, _32490_, _32486_);
  nor _82410_ (_32493_, \oc8051_golden_model_1.P1 [4], rst);
  nor _82411_ (_32494_, _32493_, _00000_);
  or _82412_ (_43464_, _32494_, _32492_);
  and _82413_ (_32495_, _13108_, \oc8051_golden_model_1.P1 [5]);
  and _82414_ (_32496_, _08652_, _07677_);
  or _82415_ (_32497_, _32496_, _32495_);
  or _82416_ (_32498_, _32497_, _06020_);
  and _82417_ (_32499_, _15093_, _07677_);
  or _82418_ (_32500_, _32499_, _32495_);
  or _82419_ (_32502_, _32500_, _06954_);
  and _82420_ (_32503_, _07677_, \oc8051_golden_model_1.ACC [5]);
  or _82421_ (_32504_, _32503_, _32495_);
  and _82422_ (_32505_, _32504_, _06938_);
  and _82423_ (_32506_, _06939_, \oc8051_golden_model_1.P1 [5]);
  or _82424_ (_32507_, _32506_, _06102_);
  or _82425_ (_32508_, _32507_, _32505_);
  and _82426_ (_32509_, _32508_, _06044_);
  and _82427_ (_32510_, _32509_, _32502_);
  and _82428_ (_32511_, _13127_, \oc8051_golden_model_1.P1 [5]);
  and _82429_ (_32513_, _15073_, _08345_);
  or _82430_ (_32514_, _32513_, _32511_);
  and _82431_ (_32515_, _32514_, _06043_);
  or _82432_ (_32516_, _32515_, _06239_);
  or _82433_ (_32517_, _32516_, _32510_);
  nor _82434_ (_32518_, _07977_, _13108_);
  or _82435_ (_32519_, _32518_, _32495_);
  or _82436_ (_32520_, _32519_, _06848_);
  and _82437_ (_32521_, _32520_, _32517_);
  or _82438_ (_32522_, _32521_, _06219_);
  or _82439_ (_32524_, _32504_, _06220_);
  and _82440_ (_32525_, _32524_, _06040_);
  and _82441_ (_32526_, _32525_, _32522_);
  and _82442_ (_32527_, _15077_, _08345_);
  or _82443_ (_32528_, _32527_, _32511_);
  and _82444_ (_32529_, _32528_, _06039_);
  or _82445_ (_32530_, _32529_, _06032_);
  or _82446_ (_32531_, _32530_, _32526_);
  or _82447_ (_32532_, _32511_, _15110_);
  and _82448_ (_32533_, _32532_, _32514_);
  or _82449_ (_32535_, _32533_, _06033_);
  and _82450_ (_32536_, _32535_, _06027_);
  and _82451_ (_32537_, _32536_, _32531_);
  or _82452_ (_32538_, _32511_, _15074_);
  and _82453_ (_32539_, _32538_, _06026_);
  and _82454_ (_32540_, _32539_, _32514_);
  or _82455_ (_32541_, _32540_, _09818_);
  or _82456_ (_32542_, _32541_, _32537_);
  and _82457_ (_32543_, _09179_, _07677_);
  or _82458_ (_32544_, _32495_, _07012_);
  or _82459_ (_32546_, _32544_, _32543_);
  or _82460_ (_32547_, _32519_, _09827_);
  and _82461_ (_32548_, _32547_, _05669_);
  and _82462_ (_32549_, _32548_, _32546_);
  and _82463_ (_32550_, _32549_, _32542_);
  and _82464_ (_32551_, _15179_, _07677_);
  or _82465_ (_32552_, _32551_, _32495_);
  and _82466_ (_32553_, _32552_, _09833_);
  or _82467_ (_32554_, _32553_, _06019_);
  or _82468_ (_32555_, _32554_, _32550_);
  and _82469_ (_32557_, _32555_, _32498_);
  or _82470_ (_32558_, _32557_, _06112_);
  and _82471_ (_32559_, _15195_, _07677_);
  or _82472_ (_32560_, _32495_, _08751_);
  or _82473_ (_32561_, _32560_, _32559_);
  and _82474_ (_32562_, _32561_, _08756_);
  and _82475_ (_32563_, _32562_, _32558_);
  and _82476_ (_32564_, _12306_, _07677_);
  or _82477_ (_32565_, _32564_, _32495_);
  and _82478_ (_32566_, _32565_, _06284_);
  or _82479_ (_32568_, _32566_, _32563_);
  and _82480_ (_32569_, _32568_, _07032_);
  or _82481_ (_32570_, _32495_, _07980_);
  and _82482_ (_32571_, _32497_, _06108_);
  and _82483_ (_32572_, _32571_, _32570_);
  or _82484_ (_32573_, _32572_, _32569_);
  and _82485_ (_32574_, _32573_, _06278_);
  and _82486_ (_32575_, _32504_, _06277_);
  and _82487_ (_32576_, _32575_, _32570_);
  or _82488_ (_32577_, _32576_, _06130_);
  or _82489_ (_32579_, _32577_, _32574_);
  and _82490_ (_32580_, _15194_, _07677_);
  or _82491_ (_32581_, _32495_, _08777_);
  or _82492_ (_32582_, _32581_, _32580_);
  and _82493_ (_32583_, _32582_, _08782_);
  and _82494_ (_32584_, _32583_, _32579_);
  nor _82495_ (_32585_, _10982_, _13108_);
  or _82496_ (_32586_, _32585_, _32495_);
  and _82497_ (_32587_, _32586_, _06292_);
  or _82498_ (_32588_, _32587_, _06316_);
  or _82499_ (_32590_, _32588_, _32584_);
  or _82500_ (_32591_, _32500_, _06718_);
  and _82501_ (_32592_, _32591_, _05653_);
  and _82502_ (_32593_, _32592_, _32590_);
  and _82503_ (_32594_, _32528_, _05652_);
  or _82504_ (_32595_, _32594_, _06047_);
  or _82505_ (_32596_, _32595_, _32593_);
  and _82506_ (_32597_, _15253_, _07677_);
  or _82507_ (_32598_, _32495_, _06048_);
  or _82508_ (_32599_, _32598_, _32597_);
  and _82509_ (_32601_, _32599_, _01336_);
  and _82510_ (_32602_, _32601_, _32596_);
  nor _82511_ (_32603_, \oc8051_golden_model_1.P1 [5], rst);
  nor _82512_ (_32604_, _32603_, _00000_);
  or _82513_ (_43465_, _32604_, _32602_);
  and _82514_ (_32605_, _13108_, \oc8051_golden_model_1.P1 [6]);
  and _82515_ (_32606_, _15389_, _07677_);
  or _82516_ (_32607_, _32606_, _32605_);
  or _82517_ (_32608_, _32607_, _06020_);
  and _82518_ (_32609_, _15293_, _07677_);
  or _82519_ (_32611_, _32609_, _32605_);
  or _82520_ (_32612_, _32611_, _06954_);
  and _82521_ (_32613_, _07677_, \oc8051_golden_model_1.ACC [6]);
  or _82522_ (_32614_, _32613_, _32605_);
  and _82523_ (_32615_, _32614_, _06938_);
  and _82524_ (_32616_, _06939_, \oc8051_golden_model_1.P1 [6]);
  or _82525_ (_32617_, _32616_, _06102_);
  or _82526_ (_32618_, _32617_, _32615_);
  and _82527_ (_32619_, _32618_, _06044_);
  and _82528_ (_32620_, _32619_, _32612_);
  and _82529_ (_32622_, _13127_, \oc8051_golden_model_1.P1 [6]);
  and _82530_ (_32623_, _15280_, _08345_);
  or _82531_ (_32624_, _32623_, _32622_);
  and _82532_ (_32625_, _32624_, _06043_);
  or _82533_ (_32626_, _32625_, _06239_);
  or _82534_ (_32627_, _32626_, _32620_);
  nor _82535_ (_32628_, _07883_, _13108_);
  or _82536_ (_32629_, _32628_, _32605_);
  or _82537_ (_32630_, _32629_, _06848_);
  and _82538_ (_32631_, _32630_, _32627_);
  or _82539_ (_32633_, _32631_, _06219_);
  or _82540_ (_32634_, _32614_, _06220_);
  and _82541_ (_32635_, _32634_, _06040_);
  and _82542_ (_32636_, _32635_, _32633_);
  and _82543_ (_32637_, _15278_, _08345_);
  or _82544_ (_32638_, _32637_, _32622_);
  and _82545_ (_32639_, _32638_, _06039_);
  or _82546_ (_32640_, _32639_, _06032_);
  or _82547_ (_32641_, _32640_, _32636_);
  or _82548_ (_32642_, _32622_, _15310_);
  and _82549_ (_32644_, _32642_, _32624_);
  or _82550_ (_32645_, _32644_, _06033_);
  and _82551_ (_32646_, _32645_, _06027_);
  and _82552_ (_32647_, _32646_, _32641_);
  or _82553_ (_32648_, _32622_, _15326_);
  and _82554_ (_32649_, _32648_, _06026_);
  and _82555_ (_32650_, _32649_, _32624_);
  or _82556_ (_32651_, _32650_, _09818_);
  or _82557_ (_32652_, _32651_, _32647_);
  and _82558_ (_32653_, _09178_, _07677_);
  or _82559_ (_32654_, _32605_, _07012_);
  or _82560_ (_32655_, _32654_, _32653_);
  or _82561_ (_32656_, _32629_, _09827_);
  and _82562_ (_32657_, _32656_, _05669_);
  and _82563_ (_32658_, _32657_, _32655_);
  and _82564_ (_32659_, _32658_, _32652_);
  and _82565_ (_32660_, _15382_, _07677_);
  or _82566_ (_32661_, _32660_, _32605_);
  and _82567_ (_32662_, _32661_, _09833_);
  or _82568_ (_32663_, _32662_, _06019_);
  or _82569_ (_32665_, _32663_, _32659_);
  and _82570_ (_32666_, _32665_, _32608_);
  or _82571_ (_32667_, _32666_, _06112_);
  and _82572_ (_32668_, _15399_, _07677_);
  or _82573_ (_32669_, _32605_, _08751_);
  or _82574_ (_32670_, _32669_, _32668_);
  and _82575_ (_32671_, _32670_, _08756_);
  and _82576_ (_32672_, _32671_, _32667_);
  and _82577_ (_32673_, _10980_, _07677_);
  or _82578_ (_32674_, _32673_, _32605_);
  and _82579_ (_32676_, _32674_, _06284_);
  or _82580_ (_32677_, _32676_, _32672_);
  and _82581_ (_32678_, _32677_, _07032_);
  or _82582_ (_32679_, _32605_, _07886_);
  and _82583_ (_32680_, _32607_, _06108_);
  and _82584_ (_32681_, _32680_, _32679_);
  or _82585_ (_32682_, _32681_, _32678_);
  and _82586_ (_32683_, _32682_, _06278_);
  and _82587_ (_32684_, _32614_, _06277_);
  and _82588_ (_32685_, _32684_, _32679_);
  or _82589_ (_32687_, _32685_, _06130_);
  or _82590_ (_32688_, _32687_, _32683_);
  and _82591_ (_32689_, _15396_, _07677_);
  or _82592_ (_32690_, _32605_, _08777_);
  or _82593_ (_32691_, _32690_, _32689_);
  and _82594_ (_32692_, _32691_, _08782_);
  and _82595_ (_32693_, _32692_, _32688_);
  nor _82596_ (_32694_, _10979_, _13108_);
  or _82597_ (_32695_, _32694_, _32605_);
  and _82598_ (_32696_, _32695_, _06292_);
  or _82599_ (_32698_, _32696_, _06316_);
  or _82600_ (_32699_, _32698_, _32693_);
  or _82601_ (_32700_, _32611_, _06718_);
  and _82602_ (_32701_, _32700_, _05653_);
  and _82603_ (_32702_, _32701_, _32699_);
  and _82604_ (_32703_, _32638_, _05652_);
  or _82605_ (_32704_, _32703_, _06047_);
  or _82606_ (_32705_, _32704_, _32702_);
  and _82607_ (_32706_, _15451_, _07677_);
  or _82608_ (_32707_, _32605_, _06048_);
  or _82609_ (_32709_, _32707_, _32706_);
  and _82610_ (_32710_, _32709_, _01336_);
  and _82611_ (_32711_, _32710_, _32705_);
  nor _82612_ (_32712_, \oc8051_golden_model_1.P1 [6], rst);
  nor _82613_ (_32713_, _32712_, _00000_);
  or _82614_ (_43466_, _32713_, _32711_);
  not _82615_ (_32714_, \oc8051_golden_model_1.IP [0]);
  nor _82616_ (_32715_, _01336_, _32714_);
  nand _82617_ (_32716_, _10995_, _07694_);
  nor _82618_ (_32717_, _07694_, _32714_);
  nor _82619_ (_32719_, _32717_, _06278_);
  nand _82620_ (_32720_, _32719_, _32716_);
  and _82621_ (_32721_, _07694_, _08672_);
  or _82622_ (_32722_, _32721_, _32717_);
  or _82623_ (_32723_, _32722_, _06020_);
  and _82624_ (_32724_, _09120_, _07694_);
  or _82625_ (_32725_, _32717_, _07012_);
  or _82626_ (_32726_, _32725_, _32724_);
  nor _82627_ (_32727_, _08127_, _13209_);
  or _82628_ (_32728_, _32727_, _32717_);
  or _82629_ (_32730_, _32728_, _06954_);
  and _82630_ (_32731_, _07694_, \oc8051_golden_model_1.ACC [0]);
  or _82631_ (_32732_, _32731_, _32717_);
  and _82632_ (_32733_, _32732_, _06938_);
  nor _82633_ (_32734_, _06938_, _32714_);
  or _82634_ (_32735_, _32734_, _06102_);
  or _82635_ (_32736_, _32735_, _32733_);
  and _82636_ (_32737_, _32736_, _06044_);
  and _82637_ (_32738_, _32737_, _32730_);
  nor _82638_ (_32739_, _08357_, _32714_);
  and _82639_ (_32741_, _14102_, _08357_);
  or _82640_ (_32742_, _32741_, _32739_);
  and _82641_ (_32743_, _32742_, _06043_);
  or _82642_ (_32744_, _32743_, _32738_);
  and _82643_ (_32745_, _32744_, _06848_);
  and _82644_ (_32746_, _07694_, _06931_);
  or _82645_ (_32747_, _32746_, _32717_);
  and _82646_ (_32748_, _32747_, _06239_);
  or _82647_ (_32749_, _32748_, _06219_);
  or _82648_ (_32750_, _32749_, _32745_);
  or _82649_ (_32752_, _32732_, _06220_);
  and _82650_ (_32753_, _32752_, _06040_);
  and _82651_ (_32754_, _32753_, _32750_);
  and _82652_ (_32755_, _32717_, _06039_);
  or _82653_ (_32756_, _32755_, _06032_);
  or _82654_ (_32757_, _32756_, _32754_);
  or _82655_ (_32758_, _32728_, _06033_);
  and _82656_ (_32759_, _32758_, _06027_);
  and _82657_ (_32760_, _32759_, _32757_);
  or _82658_ (_32761_, _32739_, _14131_);
  and _82659_ (_32763_, _32761_, _06026_);
  and _82660_ (_32764_, _32763_, _32742_);
  or _82661_ (_32765_, _32764_, _09818_);
  or _82662_ (_32766_, _32765_, _32760_);
  or _82663_ (_32767_, _32747_, _09827_);
  and _82664_ (_32768_, _32767_, _05669_);
  and _82665_ (_32769_, _32768_, _32766_);
  and _82666_ (_32770_, _32769_, _32726_);
  and _82667_ (_32771_, _14186_, _07694_);
  or _82668_ (_32772_, _32771_, _32717_);
  and _82669_ (_32774_, _32772_, _09833_);
  or _82670_ (_32775_, _32774_, _06019_);
  or _82671_ (_32776_, _32775_, _32770_);
  and _82672_ (_32777_, _32776_, _32723_);
  or _82673_ (_32778_, _32777_, _06112_);
  and _82674_ (_32779_, _14086_, _07694_);
  or _82675_ (_32780_, _32717_, _08751_);
  or _82676_ (_32781_, _32780_, _32779_);
  and _82677_ (_32782_, _32781_, _08756_);
  and _82678_ (_32783_, _32782_, _32778_);
  nor _82679_ (_32785_, _12302_, _13209_);
  or _82680_ (_32786_, _32785_, _32717_);
  and _82681_ (_32787_, _32716_, _06284_);
  and _82682_ (_32788_, _32787_, _32786_);
  or _82683_ (_32789_, _32788_, _32783_);
  and _82684_ (_32790_, _32789_, _07032_);
  nand _82685_ (_32791_, _32722_, _06108_);
  nor _82686_ (_32792_, _32791_, _32727_);
  or _82687_ (_32793_, _32792_, _06277_);
  or _82688_ (_32794_, _32793_, _32790_);
  and _82689_ (_32796_, _32794_, _32720_);
  or _82690_ (_32797_, _32796_, _06130_);
  and _82691_ (_32798_, _14083_, _07694_);
  or _82692_ (_32799_, _32717_, _08777_);
  or _82693_ (_32800_, _32799_, _32798_);
  and _82694_ (_32801_, _32800_, _08782_);
  and _82695_ (_32802_, _32801_, _32797_);
  and _82696_ (_32803_, _32786_, _06292_);
  or _82697_ (_32804_, _32803_, _06316_);
  or _82698_ (_32805_, _32804_, _32802_);
  or _82699_ (_32807_, _32728_, _06718_);
  and _82700_ (_32808_, _32807_, _32805_);
  or _82701_ (_32809_, _32808_, _05652_);
  or _82702_ (_32810_, _32717_, _05653_);
  and _82703_ (_32811_, _32810_, _32809_);
  or _82704_ (_32812_, _32811_, _06047_);
  or _82705_ (_32813_, _32728_, _06048_);
  and _82706_ (_32814_, _32813_, _01336_);
  and _82707_ (_32815_, _32814_, _32812_);
  or _82708_ (_32816_, _32815_, _32715_);
  and _82709_ (_43468_, _32816_, _42882_);
  not _82710_ (_32818_, \oc8051_golden_model_1.IP [1]);
  nor _82711_ (_32819_, _01336_, _32818_);
  nor _82712_ (_32820_, _07694_, _32818_);
  nor _82713_ (_32821_, _10993_, _13209_);
  or _82714_ (_32822_, _32821_, _32820_);
  or _82715_ (_32823_, _32822_, _08782_);
  or _82716_ (_32824_, _14367_, _13209_);
  or _82717_ (_32825_, _07694_, \oc8051_golden_model_1.IP [1]);
  and _82718_ (_32826_, _32825_, _09833_);
  and _82719_ (_32828_, _32826_, _32824_);
  nor _82720_ (_32829_, _13209_, _07132_);
  or _82721_ (_32830_, _32829_, _32820_);
  and _82722_ (_32831_, _32830_, _06239_);
  nor _82723_ (_32832_, _08357_, _32818_);
  and _82724_ (_32833_, _14266_, _08357_);
  or _82725_ (_32834_, _32833_, _32832_);
  or _82726_ (_32835_, _32834_, _06044_);
  and _82727_ (_32836_, _14284_, _07694_);
  not _82728_ (_32837_, _32836_);
  and _82729_ (_32839_, _32837_, _32825_);
  and _82730_ (_32840_, _32839_, _06102_);
  nor _82731_ (_32841_, _06938_, _32818_);
  and _82732_ (_32842_, _07694_, \oc8051_golden_model_1.ACC [1]);
  or _82733_ (_32843_, _32842_, _32820_);
  and _82734_ (_32844_, _32843_, _06938_);
  or _82735_ (_32845_, _32844_, _32841_);
  and _82736_ (_32846_, _32845_, _06954_);
  or _82737_ (_32847_, _32846_, _06043_);
  or _82738_ (_32848_, _32847_, _32840_);
  and _82739_ (_32850_, _32848_, _32835_);
  and _82740_ (_32851_, _32850_, _06848_);
  or _82741_ (_32852_, _32851_, _32831_);
  or _82742_ (_32853_, _32852_, _06219_);
  or _82743_ (_32854_, _32843_, _06220_);
  and _82744_ (_32855_, _32854_, _06040_);
  and _82745_ (_32856_, _32855_, _32853_);
  and _82746_ (_32857_, _14273_, _08357_);
  or _82747_ (_32858_, _32857_, _32832_);
  and _82748_ (_32859_, _32858_, _06039_);
  or _82749_ (_32861_, _32859_, _06032_);
  or _82750_ (_32862_, _32861_, _32856_);
  or _82751_ (_32863_, _32832_, _14302_);
  and _82752_ (_32864_, _32863_, _32834_);
  or _82753_ (_32865_, _32864_, _06033_);
  and _82754_ (_32866_, _32865_, _06027_);
  and _82755_ (_32867_, _32866_, _32862_);
  or _82756_ (_32868_, _32832_, _14267_);
  and _82757_ (_32869_, _32868_, _06026_);
  and _82758_ (_32870_, _32869_, _32834_);
  or _82759_ (_32872_, _32870_, _09815_);
  or _82760_ (_32873_, _32872_, _32867_);
  or _82761_ (_32874_, _32830_, _09827_);
  and _82762_ (_32875_, _32874_, _32873_);
  or _82763_ (_32876_, _32875_, _07011_);
  and _82764_ (_32877_, _09075_, _07694_);
  or _82765_ (_32878_, _32820_, _07012_);
  or _82766_ (_32879_, _32878_, _32877_);
  and _82767_ (_32880_, _32879_, _05669_);
  and _82768_ (_32881_, _32880_, _32876_);
  or _82769_ (_32883_, _32881_, _32828_);
  and _82770_ (_32884_, _32883_, _06020_);
  nand _82771_ (_32885_, _07694_, _06832_);
  and _82772_ (_32886_, _32825_, _06019_);
  and _82773_ (_32887_, _32886_, _32885_);
  or _82774_ (_32888_, _32887_, _32884_);
  and _82775_ (_32889_, _32888_, _08751_);
  or _82776_ (_32890_, _14263_, _13209_);
  and _82777_ (_32891_, _32825_, _06112_);
  and _82778_ (_32892_, _32891_, _32890_);
  or _82779_ (_32894_, _32892_, _06284_);
  or _82780_ (_32895_, _32894_, _32889_);
  nand _82781_ (_32896_, _10992_, _07694_);
  and _82782_ (_32897_, _32896_, _32822_);
  or _82783_ (_32898_, _32897_, _08756_);
  and _82784_ (_32899_, _32898_, _07032_);
  and _82785_ (_32900_, _32899_, _32895_);
  or _82786_ (_32901_, _14261_, _13209_);
  and _82787_ (_32902_, _32825_, _06108_);
  and _82788_ (_32903_, _32902_, _32901_);
  or _82789_ (_32905_, _32903_, _06277_);
  or _82790_ (_32906_, _32905_, _32900_);
  nor _82791_ (_32907_, _32820_, _06278_);
  nand _82792_ (_32908_, _32907_, _32896_);
  and _82793_ (_32909_, _32908_, _08777_);
  and _82794_ (_32910_, _32909_, _32906_);
  or _82795_ (_32911_, _32885_, _08078_);
  and _82796_ (_32912_, _32825_, _06130_);
  and _82797_ (_32913_, _32912_, _32911_);
  or _82798_ (_32914_, _32913_, _06292_);
  or _82799_ (_32916_, _32914_, _32910_);
  and _82800_ (_32917_, _32916_, _32823_);
  or _82801_ (_32918_, _32917_, _06316_);
  or _82802_ (_32919_, _32839_, _06718_);
  and _82803_ (_32920_, _32919_, _05653_);
  and _82804_ (_32921_, _32920_, _32918_);
  and _82805_ (_32922_, _32858_, _05652_);
  or _82806_ (_32923_, _32922_, _06047_);
  or _82807_ (_32924_, _32923_, _32921_);
  or _82808_ (_32925_, _32820_, _06048_);
  or _82809_ (_32927_, _32925_, _32836_);
  and _82810_ (_32928_, _32927_, _01336_);
  and _82811_ (_32929_, _32928_, _32924_);
  or _82812_ (_32930_, _32929_, _32819_);
  and _82813_ (_43469_, _32930_, _42882_);
  and _82814_ (_32931_, _01340_, \oc8051_golden_model_1.IP [2]);
  and _82815_ (_32932_, _13209_, \oc8051_golden_model_1.IP [2]);
  or _82816_ (_32933_, _32932_, _08177_);
  and _82817_ (_32934_, _07694_, _08730_);
  or _82818_ (_32935_, _32934_, _32932_);
  and _82819_ (_32937_, _32935_, _06108_);
  and _82820_ (_32938_, _32937_, _32933_);
  or _82821_ (_32939_, _32935_, _06020_);
  nor _82822_ (_32940_, _13209_, _07530_);
  or _82823_ (_32941_, _32940_, _32932_);
  or _82824_ (_32942_, _32941_, _06848_);
  and _82825_ (_32943_, _14493_, _07694_);
  or _82826_ (_32944_, _32943_, _32932_);
  or _82827_ (_32945_, _32944_, _06954_);
  and _82828_ (_32946_, _07694_, \oc8051_golden_model_1.ACC [2]);
  or _82829_ (_32948_, _32946_, _32932_);
  and _82830_ (_32949_, _32948_, _06938_);
  and _82831_ (_32950_, _06939_, \oc8051_golden_model_1.IP [2]);
  or _82832_ (_32951_, _32950_, _06102_);
  or _82833_ (_32952_, _32951_, _32949_);
  and _82834_ (_32953_, _32952_, _06044_);
  and _82835_ (_32954_, _32953_, _32945_);
  and _82836_ (_32955_, _13228_, \oc8051_golden_model_1.IP [2]);
  and _82837_ (_32956_, _14497_, _08357_);
  or _82838_ (_32957_, _32956_, _32955_);
  and _82839_ (_32959_, _32957_, _06043_);
  or _82840_ (_32960_, _32959_, _06239_);
  or _82841_ (_32961_, _32960_, _32954_);
  and _82842_ (_32962_, _32961_, _32942_);
  or _82843_ (_32963_, _32962_, _06219_);
  or _82844_ (_32964_, _32948_, _06220_);
  and _82845_ (_32965_, _32964_, _06040_);
  and _82846_ (_32966_, _32965_, _32963_);
  and _82847_ (_32967_, _14479_, _08357_);
  or _82848_ (_32968_, _32967_, _32955_);
  and _82849_ (_32970_, _32968_, _06039_);
  or _82850_ (_32971_, _32970_, _06032_);
  or _82851_ (_32972_, _32971_, _32966_);
  and _82852_ (_32973_, _32956_, _14512_);
  or _82853_ (_32974_, _32955_, _06033_);
  or _82854_ (_32975_, _32974_, _32973_);
  and _82855_ (_32976_, _32975_, _06027_);
  and _82856_ (_32977_, _32976_, _32972_);
  or _82857_ (_32978_, _32955_, _14525_);
  and _82858_ (_32979_, _32978_, _06026_);
  and _82859_ (_32981_, _32979_, _32957_);
  or _82860_ (_32982_, _32981_, _09818_);
  or _82861_ (_32983_, _32982_, _32977_);
  and _82862_ (_32984_, _09182_, _07694_);
  or _82863_ (_32985_, _32932_, _07012_);
  or _82864_ (_32986_, _32985_, _32984_);
  or _82865_ (_32987_, _32941_, _09827_);
  and _82866_ (_32988_, _32987_, _05669_);
  and _82867_ (_32989_, _32988_, _32986_);
  and _82868_ (_32990_, _32989_, _32983_);
  and _82869_ (_32992_, _14580_, _07694_);
  or _82870_ (_32993_, _32992_, _32932_);
  and _82871_ (_32994_, _32993_, _09833_);
  or _82872_ (_32995_, _32994_, _06019_);
  or _82873_ (_32996_, _32995_, _32990_);
  and _82874_ (_32997_, _32996_, _32939_);
  or _82875_ (_32998_, _32997_, _06112_);
  and _82876_ (_32999_, _14596_, _07694_);
  or _82877_ (_33000_, _32932_, _08751_);
  or _82878_ (_33001_, _33000_, _32999_);
  and _82879_ (_33003_, _33001_, _08756_);
  and _82880_ (_33004_, _33003_, _32998_);
  and _82881_ (_33005_, _10991_, _07694_);
  or _82882_ (_33006_, _33005_, _32932_);
  and _82883_ (_33007_, _33006_, _06284_);
  or _82884_ (_33008_, _33007_, _33004_);
  and _82885_ (_33009_, _33008_, _07032_);
  or _82886_ (_33010_, _33009_, _32938_);
  and _82887_ (_33011_, _33010_, _06278_);
  and _82888_ (_33012_, _32948_, _06277_);
  and _82889_ (_33014_, _33012_, _32933_);
  or _82890_ (_33015_, _33014_, _06130_);
  or _82891_ (_33016_, _33015_, _33011_);
  and _82892_ (_33017_, _14593_, _07694_);
  or _82893_ (_33018_, _32932_, _08777_);
  or _82894_ (_33019_, _33018_, _33017_);
  and _82895_ (_33020_, _33019_, _08782_);
  and _82896_ (_33021_, _33020_, _33016_);
  nor _82897_ (_33022_, _10990_, _13209_);
  or _82898_ (_33023_, _33022_, _32932_);
  and _82899_ (_33025_, _33023_, _06292_);
  or _82900_ (_33026_, _33025_, _06316_);
  or _82901_ (_33027_, _33026_, _33021_);
  or _82902_ (_33028_, _32944_, _06718_);
  and _82903_ (_33029_, _33028_, _05653_);
  and _82904_ (_33030_, _33029_, _33027_);
  and _82905_ (_33031_, _32968_, _05652_);
  or _82906_ (_33032_, _33031_, _06047_);
  or _82907_ (_33033_, _33032_, _33030_);
  and _82908_ (_33034_, _14657_, _07694_);
  or _82909_ (_33036_, _32932_, _06048_);
  or _82910_ (_33037_, _33036_, _33034_);
  and _82911_ (_33038_, _33037_, _01336_);
  and _82912_ (_33039_, _33038_, _33033_);
  or _82913_ (_33040_, _33039_, _32931_);
  and _82914_ (_43470_, _33040_, _42882_);
  and _82915_ (_33041_, _01340_, \oc8051_golden_model_1.IP [3]);
  and _82916_ (_33042_, _13209_, \oc8051_golden_model_1.IP [3]);
  and _82917_ (_33043_, _07694_, _08662_);
  or _82918_ (_33044_, _33043_, _33042_);
  or _82919_ (_33046_, _33044_, _06020_);
  and _82920_ (_33047_, _14672_, _07694_);
  or _82921_ (_33048_, _33047_, _33042_);
  or _82922_ (_33049_, _33048_, _06954_);
  and _82923_ (_33050_, _07694_, \oc8051_golden_model_1.ACC [3]);
  or _82924_ (_33051_, _33050_, _33042_);
  and _82925_ (_33052_, _33051_, _06938_);
  and _82926_ (_33053_, _06939_, \oc8051_golden_model_1.IP [3]);
  or _82927_ (_33054_, _33053_, _06102_);
  or _82928_ (_33055_, _33054_, _33052_);
  and _82929_ (_33057_, _33055_, _06044_);
  and _82930_ (_33058_, _33057_, _33049_);
  and _82931_ (_33059_, _13228_, \oc8051_golden_model_1.IP [3]);
  and _82932_ (_33060_, _14683_, _08357_);
  or _82933_ (_33061_, _33060_, _33059_);
  and _82934_ (_33062_, _33061_, _06043_);
  or _82935_ (_33063_, _33062_, _06239_);
  or _82936_ (_33064_, _33063_, _33058_);
  nor _82937_ (_33065_, _13209_, _07353_);
  or _82938_ (_33066_, _33065_, _33042_);
  or _82939_ (_33068_, _33066_, _06848_);
  and _82940_ (_33069_, _33068_, _33064_);
  or _82941_ (_33070_, _33069_, _06219_);
  or _82942_ (_33071_, _33051_, _06220_);
  and _82943_ (_33072_, _33071_, _06040_);
  and _82944_ (_33073_, _33072_, _33070_);
  and _82945_ (_33074_, _14681_, _08357_);
  or _82946_ (_33075_, _33074_, _33059_);
  and _82947_ (_33076_, _33075_, _06039_);
  or _82948_ (_33077_, _33076_, _06032_);
  or _82949_ (_33079_, _33077_, _33073_);
  or _82950_ (_33080_, _33059_, _14708_);
  and _82951_ (_33081_, _33080_, _33061_);
  or _82952_ (_33082_, _33081_, _06033_);
  and _82953_ (_33083_, _33082_, _06027_);
  and _82954_ (_33084_, _33083_, _33079_);
  and _82955_ (_33085_, _14724_, _08357_);
  or _82956_ (_33086_, _33085_, _33059_);
  and _82957_ (_33087_, _33086_, _06026_);
  or _82958_ (_33088_, _33087_, _09818_);
  or _82959_ (_33090_, _33088_, _33084_);
  and _82960_ (_33091_, _09181_, _07694_);
  or _82961_ (_33092_, _33042_, _07012_);
  or _82962_ (_33093_, _33092_, _33091_);
  or _82963_ (_33094_, _33066_, _09827_);
  and _82964_ (_33095_, _33094_, _05669_);
  and _82965_ (_33096_, _33095_, _33093_);
  and _82966_ (_33097_, _33096_, _33090_);
  and _82967_ (_33098_, _14778_, _07694_);
  or _82968_ (_33099_, _33098_, _33042_);
  and _82969_ (_33101_, _33099_, _09833_);
  or _82970_ (_33102_, _33101_, _06019_);
  or _82971_ (_33103_, _33102_, _33097_);
  and _82972_ (_33104_, _33103_, _33046_);
  or _82973_ (_33105_, _33104_, _06112_);
  and _82974_ (_33106_, _14793_, _07694_);
  or _82975_ (_33107_, _33042_, _08751_);
  or _82976_ (_33108_, _33107_, _33106_);
  and _82977_ (_33109_, _33108_, _08756_);
  and _82978_ (_33110_, _33109_, _33105_);
  and _82979_ (_33112_, _12299_, _07694_);
  or _82980_ (_33113_, _33112_, _33042_);
  and _82981_ (_33114_, _33113_, _06284_);
  or _82982_ (_33115_, _33114_, _33110_);
  and _82983_ (_33116_, _33115_, _07032_);
  or _82984_ (_33117_, _33042_, _08029_);
  and _82985_ (_33118_, _33044_, _06108_);
  and _82986_ (_33119_, _33118_, _33117_);
  or _82987_ (_33120_, _33119_, _33116_);
  and _82988_ (_33121_, _33120_, _06278_);
  and _82989_ (_33123_, _33051_, _06277_);
  and _82990_ (_33124_, _33123_, _33117_);
  or _82991_ (_33125_, _33124_, _06130_);
  or _82992_ (_33126_, _33125_, _33121_);
  and _82993_ (_33127_, _14792_, _07694_);
  or _82994_ (_33128_, _33042_, _08777_);
  or _82995_ (_33129_, _33128_, _33127_);
  and _82996_ (_33130_, _33129_, _08782_);
  and _82997_ (_33131_, _33130_, _33126_);
  nor _82998_ (_33132_, _10988_, _13209_);
  or _82999_ (_33134_, _33132_, _33042_);
  and _83000_ (_33135_, _33134_, _06292_);
  or _83001_ (_33136_, _33135_, _06316_);
  or _83002_ (_33137_, _33136_, _33131_);
  or _83003_ (_33138_, _33048_, _06718_);
  and _83004_ (_33139_, _33138_, _05653_);
  and _83005_ (_33140_, _33139_, _33137_);
  and _83006_ (_33141_, _33075_, _05652_);
  or _83007_ (_33142_, _33141_, _06047_);
  or _83008_ (_33143_, _33142_, _33140_);
  and _83009_ (_33145_, _14849_, _07694_);
  or _83010_ (_33146_, _33042_, _06048_);
  or _83011_ (_33147_, _33146_, _33145_);
  and _83012_ (_33148_, _33147_, _01336_);
  and _83013_ (_33149_, _33148_, _33143_);
  or _83014_ (_33150_, _33149_, _33041_);
  and _83015_ (_43471_, _33150_, _42882_);
  and _83016_ (_33151_, _01340_, \oc8051_golden_model_1.IP [4]);
  and _83017_ (_33152_, _13209_, \oc8051_golden_model_1.IP [4]);
  and _83018_ (_33153_, _08665_, _07694_);
  or _83019_ (_33155_, _33153_, _33152_);
  or _83020_ (_33156_, _33155_, _06020_);
  and _83021_ (_33157_, _14887_, _07694_);
  or _83022_ (_33158_, _33157_, _33152_);
  or _83023_ (_33159_, _33158_, _06954_);
  and _83024_ (_33160_, _07694_, \oc8051_golden_model_1.ACC [4]);
  or _83025_ (_33161_, _33160_, _33152_);
  and _83026_ (_33162_, _33161_, _06938_);
  and _83027_ (_33163_, _06939_, \oc8051_golden_model_1.IP [4]);
  or _83028_ (_33164_, _33163_, _06102_);
  or _83029_ (_33166_, _33164_, _33162_);
  and _83030_ (_33167_, _33166_, _06044_);
  and _83031_ (_33168_, _33167_, _33159_);
  and _83032_ (_33169_, _13228_, \oc8051_golden_model_1.IP [4]);
  and _83033_ (_33170_, _14878_, _08357_);
  or _83034_ (_33171_, _33170_, _33169_);
  and _83035_ (_33172_, _33171_, _06043_);
  or _83036_ (_33173_, _33172_, _06239_);
  or _83037_ (_33174_, _33173_, _33168_);
  nor _83038_ (_33175_, _08270_, _13209_);
  or _83039_ (_33177_, _33175_, _33152_);
  or _83040_ (_33178_, _33177_, _06848_);
  and _83041_ (_33179_, _33178_, _33174_);
  or _83042_ (_33180_, _33179_, _06219_);
  or _83043_ (_33181_, _33161_, _06220_);
  and _83044_ (_33182_, _33181_, _06040_);
  and _83045_ (_33183_, _33182_, _33180_);
  and _83046_ (_33184_, _14882_, _08357_);
  or _83047_ (_33185_, _33184_, _33169_);
  and _83048_ (_33186_, _33185_, _06039_);
  or _83049_ (_33188_, _33186_, _06032_);
  or _83050_ (_33189_, _33188_, _33183_);
  or _83051_ (_33190_, _33169_, _14914_);
  and _83052_ (_33191_, _33190_, _33171_);
  or _83053_ (_33192_, _33191_, _06033_);
  and _83054_ (_33193_, _33192_, _06027_);
  and _83055_ (_33194_, _33193_, _33189_);
  or _83056_ (_33195_, _33169_, _14879_);
  and _83057_ (_33196_, _33195_, _06026_);
  and _83058_ (_33197_, _33196_, _33171_);
  or _83059_ (_33199_, _33197_, _09818_);
  or _83060_ (_33200_, _33199_, _33194_);
  and _83061_ (_33201_, _09180_, _07694_);
  or _83062_ (_33202_, _33152_, _07012_);
  or _83063_ (_33203_, _33202_, _33201_);
  or _83064_ (_33204_, _33177_, _09827_);
  and _83065_ (_33205_, _33204_, _05669_);
  and _83066_ (_33206_, _33205_, _33203_);
  and _83067_ (_33207_, _33206_, _33200_);
  and _83068_ (_33208_, _14983_, _07694_);
  or _83069_ (_33210_, _33208_, _33152_);
  and _83070_ (_33211_, _33210_, _09833_);
  or _83071_ (_33212_, _33211_, _06019_);
  or _83072_ (_33213_, _33212_, _33207_);
  and _83073_ (_33214_, _33213_, _33156_);
  or _83074_ (_33215_, _33214_, _06112_);
  and _83075_ (_33216_, _14876_, _07694_);
  or _83076_ (_33217_, _33216_, _33152_);
  or _83077_ (_33218_, _33217_, _08751_);
  and _83078_ (_33219_, _33218_, _08756_);
  and _83079_ (_33221_, _33219_, _33215_);
  and _83080_ (_33222_, _10986_, _07694_);
  or _83081_ (_33223_, _33222_, _33152_);
  and _83082_ (_33224_, _33223_, _06284_);
  or _83083_ (_33225_, _33224_, _33221_);
  and _83084_ (_33226_, _33225_, _07032_);
  or _83085_ (_33227_, _33152_, _08273_);
  and _83086_ (_33228_, _33155_, _06108_);
  and _83087_ (_33229_, _33228_, _33227_);
  or _83088_ (_33230_, _33229_, _33226_);
  and _83089_ (_33232_, _33230_, _06278_);
  and _83090_ (_33233_, _33161_, _06277_);
  and _83091_ (_33234_, _33233_, _33227_);
  or _83092_ (_33235_, _33234_, _06130_);
  or _83093_ (_33236_, _33235_, _33232_);
  and _83094_ (_33237_, _14873_, _07694_);
  or _83095_ (_33238_, _33152_, _08777_);
  or _83096_ (_33239_, _33238_, _33237_);
  and _83097_ (_33240_, _33239_, _08782_);
  and _83098_ (_33241_, _33240_, _33236_);
  nor _83099_ (_33243_, _10985_, _13209_);
  or _83100_ (_33244_, _33243_, _33152_);
  and _83101_ (_33245_, _33244_, _06292_);
  or _83102_ (_33246_, _33245_, _06316_);
  or _83103_ (_33247_, _33246_, _33241_);
  or _83104_ (_33248_, _33158_, _06718_);
  and _83105_ (_33249_, _33248_, _05653_);
  and _83106_ (_33250_, _33249_, _33247_);
  and _83107_ (_33251_, _33185_, _05652_);
  or _83108_ (_33252_, _33251_, _06047_);
  or _83109_ (_33254_, _33252_, _33250_);
  and _83110_ (_33255_, _15055_, _07694_);
  or _83111_ (_33256_, _33152_, _06048_);
  or _83112_ (_33257_, _33256_, _33255_);
  and _83113_ (_33258_, _33257_, _01336_);
  and _83114_ (_33259_, _33258_, _33254_);
  or _83115_ (_33260_, _33259_, _33151_);
  and _83116_ (_43472_, _33260_, _42882_);
  and _83117_ (_33261_, _01340_, \oc8051_golden_model_1.IP [5]);
  and _83118_ (_33262_, _13209_, \oc8051_golden_model_1.IP [5]);
  and _83119_ (_33264_, _08652_, _07694_);
  or _83120_ (_33265_, _33264_, _33262_);
  or _83121_ (_33266_, _33265_, _06020_);
  and _83122_ (_33267_, _15093_, _07694_);
  or _83123_ (_33268_, _33267_, _33262_);
  or _83124_ (_33269_, _33268_, _06954_);
  and _83125_ (_33270_, _07694_, \oc8051_golden_model_1.ACC [5]);
  or _83126_ (_33271_, _33270_, _33262_);
  and _83127_ (_33272_, _33271_, _06938_);
  and _83128_ (_33273_, _06939_, \oc8051_golden_model_1.IP [5]);
  or _83129_ (_33275_, _33273_, _06102_);
  or _83130_ (_33276_, _33275_, _33272_);
  and _83131_ (_33277_, _33276_, _06044_);
  and _83132_ (_33278_, _33277_, _33269_);
  and _83133_ (_33279_, _13228_, \oc8051_golden_model_1.IP [5]);
  and _83134_ (_33280_, _15073_, _08357_);
  or _83135_ (_33281_, _33280_, _33279_);
  and _83136_ (_33282_, _33281_, _06043_);
  or _83137_ (_33283_, _33282_, _06239_);
  or _83138_ (_33284_, _33283_, _33278_);
  nor _83139_ (_33286_, _07977_, _13209_);
  or _83140_ (_33287_, _33286_, _33262_);
  or _83141_ (_33288_, _33287_, _06848_);
  and _83142_ (_33289_, _33288_, _33284_);
  or _83143_ (_33290_, _33289_, _06219_);
  or _83144_ (_33291_, _33271_, _06220_);
  and _83145_ (_33292_, _33291_, _06040_);
  and _83146_ (_33293_, _33292_, _33290_);
  and _83147_ (_33294_, _15077_, _08357_);
  or _83148_ (_33295_, _33294_, _33279_);
  and _83149_ (_33297_, _33295_, _06039_);
  or _83150_ (_33298_, _33297_, _06032_);
  or _83151_ (_33299_, _33298_, _33293_);
  or _83152_ (_33300_, _33279_, _15110_);
  and _83153_ (_33301_, _33300_, _33281_);
  or _83154_ (_33302_, _33301_, _06033_);
  and _83155_ (_33303_, _33302_, _06027_);
  and _83156_ (_33304_, _33303_, _33299_);
  or _83157_ (_33305_, _33279_, _15074_);
  and _83158_ (_33306_, _33305_, _06026_);
  and _83159_ (_33308_, _33306_, _33281_);
  or _83160_ (_33309_, _33308_, _09818_);
  or _83161_ (_33310_, _33309_, _33304_);
  and _83162_ (_33311_, _09179_, _07694_);
  or _83163_ (_33312_, _33262_, _07012_);
  or _83164_ (_33313_, _33312_, _33311_);
  or _83165_ (_33314_, _33287_, _09827_);
  and _83166_ (_33315_, _33314_, _05669_);
  and _83167_ (_33316_, _33315_, _33313_);
  and _83168_ (_33317_, _33316_, _33310_);
  and _83169_ (_33319_, _15179_, _07694_);
  or _83170_ (_33320_, _33319_, _33262_);
  and _83171_ (_33321_, _33320_, _09833_);
  or _83172_ (_33322_, _33321_, _06019_);
  or _83173_ (_33323_, _33322_, _33317_);
  and _83174_ (_33324_, _33323_, _33266_);
  or _83175_ (_33325_, _33324_, _06112_);
  and _83176_ (_33326_, _15195_, _07694_);
  or _83177_ (_33327_, _33262_, _08751_);
  or _83178_ (_33328_, _33327_, _33326_);
  and _83179_ (_33330_, _33328_, _08756_);
  and _83180_ (_33331_, _33330_, _33325_);
  and _83181_ (_33332_, _12306_, _07694_);
  or _83182_ (_33333_, _33332_, _33262_);
  and _83183_ (_33334_, _33333_, _06284_);
  or _83184_ (_33335_, _33334_, _33331_);
  and _83185_ (_33336_, _33335_, _07032_);
  or _83186_ (_33337_, _33262_, _07980_);
  and _83187_ (_33338_, _33265_, _06108_);
  and _83188_ (_33339_, _33338_, _33337_);
  or _83189_ (_33341_, _33339_, _33336_);
  and _83190_ (_33342_, _33341_, _06278_);
  and _83191_ (_33343_, _33271_, _06277_);
  and _83192_ (_33344_, _33343_, _33337_);
  or _83193_ (_33345_, _33344_, _06130_);
  or _83194_ (_33346_, _33345_, _33342_);
  and _83195_ (_33347_, _15194_, _07694_);
  or _83196_ (_33348_, _33262_, _08777_);
  or _83197_ (_33349_, _33348_, _33347_);
  and _83198_ (_33350_, _33349_, _08782_);
  and _83199_ (_33352_, _33350_, _33346_);
  nor _83200_ (_33353_, _10982_, _13209_);
  or _83201_ (_33354_, _33353_, _33262_);
  and _83202_ (_33355_, _33354_, _06292_);
  or _83203_ (_33356_, _33355_, _06316_);
  or _83204_ (_33357_, _33356_, _33352_);
  or _83205_ (_33358_, _33268_, _06718_);
  and _83206_ (_33359_, _33358_, _05653_);
  and _83207_ (_33360_, _33359_, _33357_);
  and _83208_ (_33361_, _33295_, _05652_);
  or _83209_ (_33363_, _33361_, _06047_);
  or _83210_ (_33364_, _33363_, _33360_);
  and _83211_ (_33365_, _15253_, _07694_);
  or _83212_ (_33366_, _33262_, _06048_);
  or _83213_ (_33367_, _33366_, _33365_);
  and _83214_ (_33368_, _33367_, _01336_);
  and _83215_ (_33369_, _33368_, _33364_);
  or _83216_ (_33370_, _33369_, _33261_);
  and _83217_ (_43473_, _33370_, _42882_);
  and _83218_ (_33371_, _01340_, \oc8051_golden_model_1.IP [6]);
  and _83219_ (_33373_, _13209_, \oc8051_golden_model_1.IP [6]);
  and _83220_ (_33374_, _15389_, _07694_);
  or _83221_ (_33375_, _33374_, _33373_);
  or _83222_ (_33376_, _33375_, _06020_);
  and _83223_ (_33377_, _15293_, _07694_);
  or _83224_ (_33378_, _33377_, _33373_);
  or _83225_ (_33379_, _33378_, _06954_);
  and _83226_ (_33380_, _07694_, \oc8051_golden_model_1.ACC [6]);
  or _83227_ (_33381_, _33380_, _33373_);
  and _83228_ (_33382_, _33381_, _06938_);
  and _83229_ (_33384_, _06939_, \oc8051_golden_model_1.IP [6]);
  or _83230_ (_33385_, _33384_, _06102_);
  or _83231_ (_33386_, _33385_, _33382_);
  and _83232_ (_33387_, _33386_, _06044_);
  and _83233_ (_33388_, _33387_, _33379_);
  and _83234_ (_33389_, _13228_, \oc8051_golden_model_1.IP [6]);
  and _83235_ (_33390_, _15280_, _08357_);
  or _83236_ (_33391_, _33390_, _33389_);
  and _83237_ (_33392_, _33391_, _06043_);
  or _83238_ (_33393_, _33392_, _06239_);
  or _83239_ (_33395_, _33393_, _33388_);
  nor _83240_ (_33396_, _07883_, _13209_);
  or _83241_ (_33397_, _33396_, _33373_);
  or _83242_ (_33398_, _33397_, _06848_);
  and _83243_ (_33399_, _33398_, _33395_);
  or _83244_ (_33400_, _33399_, _06219_);
  or _83245_ (_33401_, _33381_, _06220_);
  and _83246_ (_33402_, _33401_, _06040_);
  and _83247_ (_33403_, _33402_, _33400_);
  and _83248_ (_33404_, _15278_, _08357_);
  or _83249_ (_33406_, _33404_, _33389_);
  and _83250_ (_33407_, _33406_, _06039_);
  or _83251_ (_33408_, _33407_, _06032_);
  or _83252_ (_33409_, _33408_, _33403_);
  or _83253_ (_33410_, _33389_, _15310_);
  and _83254_ (_33411_, _33410_, _33391_);
  or _83255_ (_33412_, _33411_, _06033_);
  and _83256_ (_33413_, _33412_, _06027_);
  and _83257_ (_33414_, _33413_, _33409_);
  or _83258_ (_33415_, _33389_, _15326_);
  and _83259_ (_33416_, _33415_, _06026_);
  and _83260_ (_33417_, _33416_, _33391_);
  or _83261_ (_33418_, _33417_, _09818_);
  or _83262_ (_33419_, _33418_, _33414_);
  and _83263_ (_33420_, _09178_, _07694_);
  or _83264_ (_33421_, _33373_, _07012_);
  or _83265_ (_33422_, _33421_, _33420_);
  or _83266_ (_33423_, _33397_, _09827_);
  and _83267_ (_33424_, _33423_, _05669_);
  and _83268_ (_33425_, _33424_, _33422_);
  and _83269_ (_33427_, _33425_, _33419_);
  and _83270_ (_33428_, _15382_, _07694_);
  or _83271_ (_33429_, _33428_, _33373_);
  and _83272_ (_33430_, _33429_, _09833_);
  or _83273_ (_33431_, _33430_, _06019_);
  or _83274_ (_33432_, _33431_, _33427_);
  and _83275_ (_33433_, _33432_, _33376_);
  or _83276_ (_33434_, _33433_, _06112_);
  and _83277_ (_33435_, _15399_, _07694_);
  or _83278_ (_33436_, _33435_, _33373_);
  or _83279_ (_33438_, _33436_, _08751_);
  and _83280_ (_33439_, _33438_, _08756_);
  and _83281_ (_33440_, _33439_, _33434_);
  and _83282_ (_33441_, _10980_, _07694_);
  or _83283_ (_33442_, _33441_, _33373_);
  and _83284_ (_33443_, _33442_, _06284_);
  or _83285_ (_33444_, _33443_, _33440_);
  and _83286_ (_33445_, _33444_, _07032_);
  or _83287_ (_33446_, _33373_, _07886_);
  and _83288_ (_33447_, _33375_, _06108_);
  and _83289_ (_33449_, _33447_, _33446_);
  or _83290_ (_33450_, _33449_, _33445_);
  and _83291_ (_33451_, _33450_, _06278_);
  and _83292_ (_33452_, _33381_, _06277_);
  and _83293_ (_33453_, _33452_, _33446_);
  or _83294_ (_33454_, _33453_, _06130_);
  or _83295_ (_33455_, _33454_, _33451_);
  and _83296_ (_33456_, _15396_, _07694_);
  or _83297_ (_33457_, _33373_, _08777_);
  or _83298_ (_33458_, _33457_, _33456_);
  and _83299_ (_33460_, _33458_, _08782_);
  and _83300_ (_33461_, _33460_, _33455_);
  nor _83301_ (_33462_, _10979_, _13209_);
  or _83302_ (_33463_, _33462_, _33373_);
  and _83303_ (_33464_, _33463_, _06292_);
  or _83304_ (_33465_, _33464_, _06316_);
  or _83305_ (_33466_, _33465_, _33461_);
  or _83306_ (_33467_, _33378_, _06718_);
  and _83307_ (_33468_, _33467_, _05653_);
  and _83308_ (_33469_, _33468_, _33466_);
  and _83309_ (_33471_, _33406_, _05652_);
  or _83310_ (_33472_, _33471_, _06047_);
  or _83311_ (_33473_, _33472_, _33469_);
  and _83312_ (_33474_, _15451_, _07694_);
  or _83313_ (_33475_, _33373_, _06048_);
  or _83314_ (_33476_, _33475_, _33474_);
  and _83315_ (_33477_, _33476_, _01336_);
  and _83316_ (_33478_, _33477_, _33473_);
  or _83317_ (_33479_, _33478_, _33371_);
  and _83318_ (_43474_, _33479_, _42882_);
  not _83319_ (_33481_, \oc8051_golden_model_1.IE [0]);
  nor _83320_ (_33482_, _01336_, _33481_);
  nor _83321_ (_33483_, _07688_, _33481_);
  and _83322_ (_33484_, _07688_, _08672_);
  or _83323_ (_33485_, _33484_, _33483_);
  or _83324_ (_33486_, _33485_, _06020_);
  and _83325_ (_33487_, _09120_, _07688_);
  or _83326_ (_33488_, _33483_, _07012_);
  or _83327_ (_33489_, _33488_, _33487_);
  nor _83328_ (_33490_, _08127_, _13311_);
  or _83329_ (_33492_, _33490_, _33483_);
  or _83330_ (_33493_, _33492_, _06954_);
  and _83331_ (_33494_, _07688_, \oc8051_golden_model_1.ACC [0]);
  or _83332_ (_33495_, _33494_, _33483_);
  and _83333_ (_33496_, _33495_, _06938_);
  nor _83334_ (_33497_, _06938_, _33481_);
  or _83335_ (_33498_, _33497_, _06102_);
  or _83336_ (_33499_, _33498_, _33496_);
  and _83337_ (_33500_, _33499_, _06044_);
  and _83338_ (_33501_, _33500_, _33493_);
  nor _83339_ (_33503_, _08351_, _33481_);
  and _83340_ (_33504_, _14102_, _08351_);
  or _83341_ (_33505_, _33504_, _33503_);
  and _83342_ (_33506_, _33505_, _06043_);
  or _83343_ (_33507_, _33506_, _33501_);
  and _83344_ (_33508_, _33507_, _06848_);
  and _83345_ (_33509_, _07688_, _06931_);
  or _83346_ (_33510_, _33509_, _33483_);
  and _83347_ (_33511_, _33510_, _06239_);
  or _83348_ (_33512_, _33511_, _06219_);
  or _83349_ (_33514_, _33512_, _33508_);
  or _83350_ (_33515_, _33495_, _06220_);
  and _83351_ (_33516_, _33515_, _06040_);
  and _83352_ (_33517_, _33516_, _33514_);
  and _83353_ (_33518_, _33483_, _06039_);
  or _83354_ (_33519_, _33518_, _06032_);
  or _83355_ (_33520_, _33519_, _33517_);
  or _83356_ (_33521_, _33492_, _06033_);
  and _83357_ (_33522_, _33521_, _06027_);
  and _83358_ (_33523_, _33522_, _33520_);
  or _83359_ (_33525_, _33503_, _14131_);
  and _83360_ (_33526_, _33525_, _06026_);
  and _83361_ (_33527_, _33526_, _33505_);
  or _83362_ (_33528_, _33527_, _09818_);
  or _83363_ (_33529_, _33528_, _33523_);
  or _83364_ (_33530_, _33510_, _09827_);
  and _83365_ (_33531_, _33530_, _05669_);
  and _83366_ (_33532_, _33531_, _33529_);
  and _83367_ (_33533_, _33532_, _33489_);
  and _83368_ (_33534_, _14186_, _07688_);
  or _83369_ (_33536_, _33534_, _33483_);
  and _83370_ (_33537_, _33536_, _09833_);
  or _83371_ (_33538_, _33537_, _06019_);
  or _83372_ (_33539_, _33538_, _33533_);
  and _83373_ (_33540_, _33539_, _33486_);
  or _83374_ (_33541_, _33540_, _06112_);
  and _83375_ (_33542_, _14086_, _07688_);
  or _83376_ (_33543_, _33483_, _08751_);
  or _83377_ (_33544_, _33543_, _33542_);
  and _83378_ (_33545_, _33544_, _08756_);
  and _83379_ (_33547_, _33545_, _33541_);
  nor _83380_ (_33548_, _12302_, _13311_);
  or _83381_ (_33549_, _33548_, _33483_);
  nand _83382_ (_33550_, _10995_, _07688_);
  and _83383_ (_33551_, _33550_, _06284_);
  and _83384_ (_33552_, _33551_, _33549_);
  or _83385_ (_33553_, _33552_, _33547_);
  and _83386_ (_33554_, _33553_, _07032_);
  nand _83387_ (_33555_, _33485_, _06108_);
  nor _83388_ (_33556_, _33555_, _33490_);
  or _83389_ (_33558_, _33556_, _06277_);
  or _83390_ (_33559_, _33558_, _33554_);
  nor _83391_ (_33560_, _33483_, _06278_);
  nand _83392_ (_33561_, _33560_, _33550_);
  and _83393_ (_33562_, _33561_, _33559_);
  or _83394_ (_33563_, _33562_, _06130_);
  and _83395_ (_33564_, _14083_, _07688_);
  or _83396_ (_33565_, _33483_, _08777_);
  or _83397_ (_33566_, _33565_, _33564_);
  and _83398_ (_33567_, _33566_, _08782_);
  and _83399_ (_33569_, _33567_, _33563_);
  and _83400_ (_33570_, _33549_, _06292_);
  or _83401_ (_33571_, _33570_, _06316_);
  or _83402_ (_33572_, _33571_, _33569_);
  or _83403_ (_33573_, _33492_, _06718_);
  and _83404_ (_33574_, _33573_, _33572_);
  or _83405_ (_33575_, _33574_, _05652_);
  or _83406_ (_33576_, _33483_, _05653_);
  and _83407_ (_33577_, _33576_, _33575_);
  or _83408_ (_33578_, _33577_, _06047_);
  or _83409_ (_33580_, _33492_, _06048_);
  and _83410_ (_33581_, _33580_, _01336_);
  and _83411_ (_33582_, _33581_, _33578_);
  or _83412_ (_33583_, _33582_, _33482_);
  and _83413_ (_43476_, _33583_, _42882_);
  not _83414_ (_33584_, \oc8051_golden_model_1.IE [1]);
  nor _83415_ (_33585_, _01336_, _33584_);
  nor _83416_ (_33586_, _07688_, _33584_);
  nor _83417_ (_33587_, _10993_, _13311_);
  or _83418_ (_33588_, _33587_, _33586_);
  or _83419_ (_33590_, _33588_, _08782_);
  or _83420_ (_33591_, _14367_, _13311_);
  or _83421_ (_33592_, _07688_, \oc8051_golden_model_1.IE [1]);
  and _83422_ (_33593_, _33592_, _09833_);
  and _83423_ (_33594_, _33593_, _33591_);
  nor _83424_ (_33595_, _13311_, _07132_);
  or _83425_ (_33596_, _33595_, _33586_);
  or _83426_ (_33597_, _33596_, _06848_);
  and _83427_ (_33598_, _14284_, _07688_);
  not _83428_ (_33599_, _33598_);
  and _83429_ (_33601_, _33599_, _33592_);
  or _83430_ (_33602_, _33601_, _06954_);
  and _83431_ (_33603_, _07688_, \oc8051_golden_model_1.ACC [1]);
  or _83432_ (_33604_, _33603_, _33586_);
  and _83433_ (_33605_, _33604_, _06938_);
  nor _83434_ (_33606_, _06938_, _33584_);
  or _83435_ (_33607_, _33606_, _06102_);
  or _83436_ (_33608_, _33607_, _33605_);
  and _83437_ (_33609_, _33608_, _06044_);
  and _83438_ (_33610_, _33609_, _33602_);
  nor _83439_ (_33612_, _08351_, _33584_);
  and _83440_ (_33613_, _14266_, _08351_);
  or _83441_ (_33614_, _33613_, _33612_);
  and _83442_ (_33615_, _33614_, _06043_);
  or _83443_ (_33616_, _33615_, _06239_);
  or _83444_ (_33617_, _33616_, _33610_);
  and _83445_ (_33618_, _33617_, _33597_);
  or _83446_ (_33619_, _33618_, _06219_);
  or _83447_ (_33620_, _33604_, _06220_);
  and _83448_ (_33621_, _33620_, _06040_);
  and _83449_ (_33623_, _33621_, _33619_);
  and _83450_ (_33624_, _14273_, _08351_);
  or _83451_ (_33625_, _33624_, _33612_);
  and _83452_ (_33626_, _33625_, _06039_);
  or _83453_ (_33627_, _33626_, _06032_);
  or _83454_ (_33628_, _33627_, _33623_);
  and _83455_ (_33629_, _33613_, _14302_);
  or _83456_ (_33630_, _33612_, _06033_);
  or _83457_ (_33631_, _33630_, _33629_);
  and _83458_ (_33632_, _33631_, _06027_);
  and _83459_ (_33634_, _33632_, _33628_);
  or _83460_ (_33635_, _33612_, _14267_);
  and _83461_ (_33636_, _33635_, _06026_);
  and _83462_ (_33637_, _33636_, _33614_);
  or _83463_ (_33638_, _33637_, _09818_);
  or _83464_ (_33639_, _33638_, _33634_);
  and _83465_ (_33640_, _09075_, _07688_);
  or _83466_ (_33641_, _33586_, _07012_);
  or _83467_ (_33642_, _33641_, _33640_);
  or _83468_ (_33643_, _33596_, _09827_);
  and _83469_ (_33645_, _33643_, _05669_);
  and _83470_ (_33646_, _33645_, _33642_);
  and _83471_ (_33647_, _33646_, _33639_);
  or _83472_ (_33648_, _33647_, _33594_);
  and _83473_ (_33649_, _33648_, _06020_);
  nand _83474_ (_33650_, _07688_, _06832_);
  and _83475_ (_33651_, _33592_, _06019_);
  and _83476_ (_33652_, _33651_, _33650_);
  or _83477_ (_33653_, _33652_, _33649_);
  and _83478_ (_33654_, _33653_, _08751_);
  or _83479_ (_33656_, _14263_, _13311_);
  and _83480_ (_33657_, _33592_, _06112_);
  and _83481_ (_33658_, _33657_, _33656_);
  or _83482_ (_33659_, _33658_, _06284_);
  or _83483_ (_33660_, _33659_, _33654_);
  nand _83484_ (_33661_, _10992_, _07688_);
  and _83485_ (_33662_, _33661_, _33588_);
  or _83486_ (_33663_, _33662_, _08756_);
  and _83487_ (_33664_, _33663_, _07032_);
  and _83488_ (_33665_, _33664_, _33660_);
  or _83489_ (_33667_, _14261_, _13311_);
  and _83490_ (_33668_, _33592_, _06108_);
  and _83491_ (_33669_, _33668_, _33667_);
  or _83492_ (_33670_, _33669_, _06277_);
  or _83493_ (_33671_, _33670_, _33665_);
  nor _83494_ (_33672_, _33586_, _06278_);
  nand _83495_ (_33673_, _33672_, _33661_);
  and _83496_ (_33674_, _33673_, _08777_);
  and _83497_ (_33675_, _33674_, _33671_);
  or _83498_ (_33676_, _33650_, _08078_);
  and _83499_ (_33678_, _33592_, _06130_);
  and _83500_ (_33679_, _33678_, _33676_);
  or _83501_ (_33680_, _33679_, _06292_);
  or _83502_ (_33681_, _33680_, _33675_);
  and _83503_ (_33682_, _33681_, _33590_);
  or _83504_ (_33683_, _33682_, _06316_);
  or _83505_ (_33684_, _33601_, _06718_);
  and _83506_ (_33685_, _33684_, _05653_);
  and _83507_ (_33686_, _33685_, _33683_);
  and _83508_ (_33687_, _33625_, _05652_);
  or _83509_ (_33689_, _33687_, _06047_);
  or _83510_ (_33690_, _33689_, _33686_);
  or _83511_ (_33691_, _33586_, _06048_);
  or _83512_ (_33692_, _33691_, _33598_);
  and _83513_ (_33693_, _33692_, _01336_);
  and _83514_ (_33694_, _33693_, _33690_);
  or _83515_ (_33695_, _33694_, _33585_);
  and _83516_ (_43477_, _33695_, _42882_);
  and _83517_ (_33696_, _01340_, \oc8051_golden_model_1.IE [2]);
  and _83518_ (_33697_, _13311_, \oc8051_golden_model_1.IE [2]);
  and _83519_ (_33699_, _07688_, _08730_);
  or _83520_ (_33700_, _33699_, _33697_);
  or _83521_ (_33701_, _33700_, _06020_);
  nor _83522_ (_33702_, _13311_, _07530_);
  or _83523_ (_33703_, _33702_, _33697_);
  and _83524_ (_33704_, _33703_, _06239_);
  and _83525_ (_33705_, _13330_, \oc8051_golden_model_1.IE [2]);
  and _83526_ (_33706_, _14497_, _08351_);
  or _83527_ (_33707_, _33706_, _33705_);
  or _83528_ (_33708_, _33707_, _06044_);
  and _83529_ (_33710_, _14493_, _07688_);
  or _83530_ (_33711_, _33710_, _33697_);
  and _83531_ (_33712_, _33711_, _06102_);
  and _83532_ (_33713_, _06939_, \oc8051_golden_model_1.IE [2]);
  and _83533_ (_33714_, _07688_, \oc8051_golden_model_1.ACC [2]);
  or _83534_ (_33715_, _33714_, _33697_);
  and _83535_ (_33716_, _33715_, _06938_);
  or _83536_ (_33717_, _33716_, _33713_);
  and _83537_ (_33718_, _33717_, _06954_);
  or _83538_ (_33719_, _33718_, _06043_);
  or _83539_ (_33721_, _33719_, _33712_);
  and _83540_ (_33722_, _33721_, _33708_);
  and _83541_ (_33723_, _33722_, _06848_);
  or _83542_ (_33724_, _33723_, _33704_);
  or _83543_ (_33725_, _33724_, _06219_);
  or _83544_ (_33726_, _33715_, _06220_);
  and _83545_ (_33727_, _33726_, _06040_);
  and _83546_ (_33728_, _33727_, _33725_);
  and _83547_ (_33729_, _14479_, _08351_);
  or _83548_ (_33730_, _33729_, _33705_);
  and _83549_ (_33732_, _33730_, _06039_);
  or _83550_ (_33733_, _33732_, _06032_);
  or _83551_ (_33734_, _33733_, _33728_);
  or _83552_ (_33735_, _33705_, _14512_);
  and _83553_ (_33736_, _33735_, _33707_);
  or _83554_ (_33737_, _33736_, _06033_);
  and _83555_ (_33738_, _33737_, _06027_);
  and _83556_ (_33739_, _33738_, _33734_);
  or _83557_ (_33740_, _33705_, _14525_);
  and _83558_ (_33741_, _33740_, _06026_);
  and _83559_ (_33743_, _33741_, _33707_);
  or _83560_ (_33744_, _33743_, _09818_);
  or _83561_ (_33745_, _33744_, _33739_);
  and _83562_ (_33746_, _09182_, _07688_);
  or _83563_ (_33747_, _33697_, _07012_);
  or _83564_ (_33748_, _33747_, _33746_);
  or _83565_ (_33749_, _33703_, _09827_);
  and _83566_ (_33750_, _33749_, _05669_);
  and _83567_ (_33751_, _33750_, _33748_);
  and _83568_ (_33752_, _33751_, _33745_);
  and _83569_ (_33754_, _14580_, _07688_);
  or _83570_ (_33755_, _33754_, _33697_);
  and _83571_ (_33756_, _33755_, _09833_);
  or _83572_ (_33757_, _33756_, _06019_);
  or _83573_ (_33758_, _33757_, _33752_);
  and _83574_ (_33759_, _33758_, _33701_);
  or _83575_ (_33760_, _33759_, _06112_);
  and _83576_ (_33761_, _14596_, _07688_);
  or _83577_ (_33762_, _33697_, _08751_);
  or _83578_ (_33763_, _33762_, _33761_);
  and _83579_ (_33765_, _33763_, _08756_);
  and _83580_ (_33766_, _33765_, _33760_);
  and _83581_ (_33767_, _10991_, _07688_);
  or _83582_ (_33768_, _33767_, _33697_);
  and _83583_ (_33769_, _33768_, _06284_);
  or _83584_ (_33770_, _33769_, _33766_);
  and _83585_ (_33771_, _33770_, _07032_);
  or _83586_ (_33772_, _33697_, _08177_);
  and _83587_ (_33773_, _33700_, _06108_);
  and _83588_ (_33774_, _33773_, _33772_);
  or _83589_ (_33776_, _33774_, _33771_);
  and _83590_ (_33777_, _33776_, _06278_);
  and _83591_ (_33778_, _33715_, _06277_);
  and _83592_ (_33779_, _33778_, _33772_);
  or _83593_ (_33780_, _33779_, _06130_);
  or _83594_ (_33781_, _33780_, _33777_);
  and _83595_ (_33782_, _14593_, _07688_);
  or _83596_ (_33783_, _33697_, _08777_);
  or _83597_ (_33784_, _33783_, _33782_);
  and _83598_ (_33785_, _33784_, _08782_);
  and _83599_ (_33787_, _33785_, _33781_);
  nor _83600_ (_33788_, _10990_, _13311_);
  or _83601_ (_33789_, _33788_, _33697_);
  and _83602_ (_33790_, _33789_, _06292_);
  or _83603_ (_33791_, _33790_, _06316_);
  or _83604_ (_33792_, _33791_, _33787_);
  or _83605_ (_33793_, _33711_, _06718_);
  and _83606_ (_33794_, _33793_, _05653_);
  and _83607_ (_33795_, _33794_, _33792_);
  and _83608_ (_33796_, _33730_, _05652_);
  or _83609_ (_33798_, _33796_, _06047_);
  or _83610_ (_33799_, _33798_, _33795_);
  and _83611_ (_33800_, _14657_, _07688_);
  or _83612_ (_33801_, _33697_, _06048_);
  or _83613_ (_33802_, _33801_, _33800_);
  and _83614_ (_33803_, _33802_, _01336_);
  and _83615_ (_33804_, _33803_, _33799_);
  or _83616_ (_33805_, _33804_, _33696_);
  and _83617_ (_43478_, _33805_, _42882_);
  and _83618_ (_33806_, _01340_, \oc8051_golden_model_1.IE [3]);
  and _83619_ (_33808_, _13311_, \oc8051_golden_model_1.IE [3]);
  and _83620_ (_33809_, _07688_, _08662_);
  or _83621_ (_33810_, _33809_, _33808_);
  or _83622_ (_33811_, _33810_, _06020_);
  and _83623_ (_33812_, _14672_, _07688_);
  or _83624_ (_33813_, _33812_, _33808_);
  or _83625_ (_33814_, _33813_, _06954_);
  and _83626_ (_33815_, _07688_, \oc8051_golden_model_1.ACC [3]);
  or _83627_ (_33816_, _33815_, _33808_);
  and _83628_ (_33817_, _33816_, _06938_);
  and _83629_ (_33819_, _06939_, \oc8051_golden_model_1.IE [3]);
  or _83630_ (_33820_, _33819_, _06102_);
  or _83631_ (_33821_, _33820_, _33817_);
  and _83632_ (_33822_, _33821_, _06044_);
  and _83633_ (_33823_, _33822_, _33814_);
  and _83634_ (_33824_, _13330_, \oc8051_golden_model_1.IE [3]);
  and _83635_ (_33825_, _14683_, _08351_);
  or _83636_ (_33826_, _33825_, _33824_);
  and _83637_ (_33827_, _33826_, _06043_);
  or _83638_ (_33828_, _33827_, _06239_);
  or _83639_ (_33830_, _33828_, _33823_);
  nor _83640_ (_33831_, _13311_, _07353_);
  or _83641_ (_33832_, _33831_, _33808_);
  or _83642_ (_33833_, _33832_, _06848_);
  and _83643_ (_33834_, _33833_, _33830_);
  or _83644_ (_33835_, _33834_, _06219_);
  or _83645_ (_33836_, _33816_, _06220_);
  and _83646_ (_33837_, _33836_, _06040_);
  and _83647_ (_33838_, _33837_, _33835_);
  and _83648_ (_33839_, _14681_, _08351_);
  or _83649_ (_33841_, _33839_, _33824_);
  and _83650_ (_33842_, _33841_, _06039_);
  or _83651_ (_33843_, _33842_, _06032_);
  or _83652_ (_33844_, _33843_, _33838_);
  or _83653_ (_33845_, _33824_, _14708_);
  and _83654_ (_33846_, _33845_, _33826_);
  or _83655_ (_33847_, _33846_, _06033_);
  and _83656_ (_33848_, _33847_, _06027_);
  and _83657_ (_33849_, _33848_, _33844_);
  and _83658_ (_33850_, _14724_, _08351_);
  or _83659_ (_33852_, _33850_, _33824_);
  and _83660_ (_33853_, _33852_, _06026_);
  or _83661_ (_33854_, _33853_, _09818_);
  or _83662_ (_33855_, _33854_, _33849_);
  and _83663_ (_33856_, _09181_, _07688_);
  or _83664_ (_33857_, _33808_, _07012_);
  or _83665_ (_33858_, _33857_, _33856_);
  or _83666_ (_33859_, _33832_, _09827_);
  and _83667_ (_33860_, _33859_, _05669_);
  and _83668_ (_33861_, _33860_, _33858_);
  and _83669_ (_33863_, _33861_, _33855_);
  and _83670_ (_33864_, _14778_, _07688_);
  or _83671_ (_33865_, _33864_, _33808_);
  and _83672_ (_33866_, _33865_, _09833_);
  or _83673_ (_33867_, _33866_, _06019_);
  or _83674_ (_33868_, _33867_, _33863_);
  and _83675_ (_33869_, _33868_, _33811_);
  or _83676_ (_33870_, _33869_, _06112_);
  and _83677_ (_33871_, _14793_, _07688_);
  or _83678_ (_33872_, _33808_, _08751_);
  or _83679_ (_33874_, _33872_, _33871_);
  and _83680_ (_33875_, _33874_, _08756_);
  and _83681_ (_33876_, _33875_, _33870_);
  and _83682_ (_33877_, _12299_, _07688_);
  or _83683_ (_33878_, _33877_, _33808_);
  and _83684_ (_33879_, _33878_, _06284_);
  or _83685_ (_33880_, _33879_, _33876_);
  and _83686_ (_33881_, _33880_, _07032_);
  or _83687_ (_33882_, _33808_, _08029_);
  and _83688_ (_33883_, _33810_, _06108_);
  and _83689_ (_33885_, _33883_, _33882_);
  or _83690_ (_33886_, _33885_, _33881_);
  and _83691_ (_33887_, _33886_, _06278_);
  and _83692_ (_33888_, _33816_, _06277_);
  and _83693_ (_33889_, _33888_, _33882_);
  or _83694_ (_33890_, _33889_, _06130_);
  or _83695_ (_33891_, _33890_, _33887_);
  and _83696_ (_33892_, _14792_, _07688_);
  or _83697_ (_33893_, _33808_, _08777_);
  or _83698_ (_33894_, _33893_, _33892_);
  and _83699_ (_33896_, _33894_, _08782_);
  and _83700_ (_33897_, _33896_, _33891_);
  nor _83701_ (_33898_, _10988_, _13311_);
  or _83702_ (_33899_, _33898_, _33808_);
  and _83703_ (_33900_, _33899_, _06292_);
  or _83704_ (_33901_, _33900_, _06316_);
  or _83705_ (_33902_, _33901_, _33897_);
  or _83706_ (_33903_, _33813_, _06718_);
  and _83707_ (_33904_, _33903_, _05653_);
  and _83708_ (_33905_, _33904_, _33902_);
  and _83709_ (_33907_, _33841_, _05652_);
  or _83710_ (_33908_, _33907_, _06047_);
  or _83711_ (_33909_, _33908_, _33905_);
  and _83712_ (_33910_, _14849_, _07688_);
  or _83713_ (_33911_, _33808_, _06048_);
  or _83714_ (_33912_, _33911_, _33910_);
  and _83715_ (_33913_, _33912_, _01336_);
  and _83716_ (_33914_, _33913_, _33909_);
  or _83717_ (_33915_, _33914_, _33806_);
  and _83718_ (_43479_, _33915_, _42882_);
  and _83719_ (_33917_, _01340_, \oc8051_golden_model_1.IE [4]);
  and _83720_ (_33918_, _13311_, \oc8051_golden_model_1.IE [4]);
  and _83721_ (_33919_, _08665_, _07688_);
  or _83722_ (_33920_, _33919_, _33918_);
  or _83723_ (_33921_, _33920_, _06020_);
  and _83724_ (_33922_, _14887_, _07688_);
  or _83725_ (_33923_, _33922_, _33918_);
  or _83726_ (_33924_, _33923_, _06954_);
  and _83727_ (_33925_, _07688_, \oc8051_golden_model_1.ACC [4]);
  or _83728_ (_33926_, _33925_, _33918_);
  and _83729_ (_33928_, _33926_, _06938_);
  and _83730_ (_33929_, _06939_, \oc8051_golden_model_1.IE [4]);
  or _83731_ (_33930_, _33929_, _06102_);
  or _83732_ (_33931_, _33930_, _33928_);
  and _83733_ (_33932_, _33931_, _06044_);
  and _83734_ (_33933_, _33932_, _33924_);
  and _83735_ (_33934_, _13330_, \oc8051_golden_model_1.IE [4]);
  and _83736_ (_33935_, _14878_, _08351_);
  or _83737_ (_33936_, _33935_, _33934_);
  and _83738_ (_33937_, _33936_, _06043_);
  or _83739_ (_33939_, _33937_, _06239_);
  or _83740_ (_33940_, _33939_, _33933_);
  nor _83741_ (_33941_, _08270_, _13311_);
  or _83742_ (_33942_, _33941_, _33918_);
  or _83743_ (_33943_, _33942_, _06848_);
  and _83744_ (_33944_, _33943_, _33940_);
  or _83745_ (_33945_, _33944_, _06219_);
  or _83746_ (_33946_, _33926_, _06220_);
  and _83747_ (_33947_, _33946_, _06040_);
  and _83748_ (_33948_, _33947_, _33945_);
  and _83749_ (_33950_, _14882_, _08351_);
  or _83750_ (_33951_, _33950_, _33934_);
  and _83751_ (_33952_, _33951_, _06039_);
  or _83752_ (_33953_, _33952_, _06032_);
  or _83753_ (_33954_, _33953_, _33948_);
  or _83754_ (_33955_, _33934_, _14914_);
  and _83755_ (_33956_, _33955_, _33936_);
  or _83756_ (_33957_, _33956_, _06033_);
  and _83757_ (_33958_, _33957_, _06027_);
  and _83758_ (_33959_, _33958_, _33954_);
  or _83759_ (_33961_, _33934_, _14879_);
  and _83760_ (_33962_, _33961_, _06026_);
  and _83761_ (_33963_, _33962_, _33936_);
  or _83762_ (_33964_, _33963_, _09818_);
  or _83763_ (_33965_, _33964_, _33959_);
  and _83764_ (_33966_, _09180_, _07688_);
  or _83765_ (_33967_, _33918_, _07012_);
  or _83766_ (_33968_, _33967_, _33966_);
  or _83767_ (_33969_, _33942_, _09827_);
  and _83768_ (_33970_, _33969_, _05669_);
  and _83769_ (_33972_, _33970_, _33968_);
  and _83770_ (_33973_, _33972_, _33965_);
  and _83771_ (_33974_, _14983_, _07688_);
  or _83772_ (_33975_, _33974_, _33918_);
  and _83773_ (_33976_, _33975_, _09833_);
  or _83774_ (_33977_, _33976_, _06019_);
  or _83775_ (_33978_, _33977_, _33973_);
  and _83776_ (_33979_, _33978_, _33921_);
  or _83777_ (_33980_, _33979_, _06112_);
  and _83778_ (_33981_, _14876_, _07688_);
  or _83779_ (_33983_, _33918_, _08751_);
  or _83780_ (_33984_, _33983_, _33981_);
  and _83781_ (_33985_, _33984_, _08756_);
  and _83782_ (_33986_, _33985_, _33980_);
  and _83783_ (_33987_, _10986_, _07688_);
  or _83784_ (_33988_, _33987_, _33918_);
  and _83785_ (_33989_, _33988_, _06284_);
  or _83786_ (_33990_, _33989_, _33986_);
  and _83787_ (_33991_, _33990_, _07032_);
  or _83788_ (_33992_, _33918_, _08273_);
  and _83789_ (_33994_, _33920_, _06108_);
  and _83790_ (_33995_, _33994_, _33992_);
  or _83791_ (_33996_, _33995_, _33991_);
  and _83792_ (_33997_, _33996_, _06278_);
  and _83793_ (_33998_, _33926_, _06277_);
  and _83794_ (_33999_, _33998_, _33992_);
  or _83795_ (_34000_, _33999_, _06130_);
  or _83796_ (_34001_, _34000_, _33997_);
  and _83797_ (_34002_, _14873_, _07688_);
  or _83798_ (_34003_, _33918_, _08777_);
  or _83799_ (_34005_, _34003_, _34002_);
  and _83800_ (_34006_, _34005_, _08782_);
  and _83801_ (_34007_, _34006_, _34001_);
  nor _83802_ (_34008_, _10985_, _13311_);
  or _83803_ (_34009_, _34008_, _33918_);
  and _83804_ (_34010_, _34009_, _06292_);
  or _83805_ (_34011_, _34010_, _06316_);
  or _83806_ (_34012_, _34011_, _34007_);
  or _83807_ (_34013_, _33923_, _06718_);
  and _83808_ (_34014_, _34013_, _05653_);
  and _83809_ (_34016_, _34014_, _34012_);
  and _83810_ (_34017_, _33951_, _05652_);
  or _83811_ (_34018_, _34017_, _06047_);
  or _83812_ (_34019_, _34018_, _34016_);
  and _83813_ (_34020_, _15055_, _07688_);
  or _83814_ (_34021_, _33918_, _06048_);
  or _83815_ (_34022_, _34021_, _34020_);
  and _83816_ (_34023_, _34022_, _01336_);
  and _83817_ (_34024_, _34023_, _34019_);
  or _83818_ (_34025_, _34024_, _33917_);
  and _83819_ (_43480_, _34025_, _42882_);
  and _83820_ (_34027_, _01340_, \oc8051_golden_model_1.IE [5]);
  and _83821_ (_34028_, _13311_, \oc8051_golden_model_1.IE [5]);
  and _83822_ (_34029_, _08652_, _07688_);
  or _83823_ (_34030_, _34029_, _34028_);
  or _83824_ (_34031_, _34030_, _06020_);
  and _83825_ (_34032_, _15093_, _07688_);
  or _83826_ (_34033_, _34032_, _34028_);
  or _83827_ (_34034_, _34033_, _06954_);
  and _83828_ (_34035_, _07688_, \oc8051_golden_model_1.ACC [5]);
  or _83829_ (_34037_, _34035_, _34028_);
  and _83830_ (_34038_, _34037_, _06938_);
  and _83831_ (_34039_, _06939_, \oc8051_golden_model_1.IE [5]);
  or _83832_ (_34040_, _34039_, _06102_);
  or _83833_ (_34041_, _34040_, _34038_);
  and _83834_ (_34042_, _34041_, _06044_);
  and _83835_ (_34043_, _34042_, _34034_);
  and _83836_ (_34044_, _13330_, \oc8051_golden_model_1.IE [5]);
  and _83837_ (_34045_, _15073_, _08351_);
  or _83838_ (_34046_, _34045_, _34044_);
  and _83839_ (_34048_, _34046_, _06043_);
  or _83840_ (_34049_, _34048_, _06239_);
  or _83841_ (_34050_, _34049_, _34043_);
  nor _83842_ (_34051_, _07977_, _13311_);
  or _83843_ (_34052_, _34051_, _34028_);
  or _83844_ (_34053_, _34052_, _06848_);
  and _83845_ (_34054_, _34053_, _34050_);
  or _83846_ (_34055_, _34054_, _06219_);
  or _83847_ (_34056_, _34037_, _06220_);
  and _83848_ (_34057_, _34056_, _06040_);
  and _83849_ (_34059_, _34057_, _34055_);
  and _83850_ (_34060_, _15077_, _08351_);
  or _83851_ (_34061_, _34060_, _34044_);
  and _83852_ (_34062_, _34061_, _06039_);
  or _83853_ (_34063_, _34062_, _06032_);
  or _83854_ (_34064_, _34063_, _34059_);
  or _83855_ (_34065_, _34044_, _15110_);
  and _83856_ (_34066_, _34065_, _34046_);
  or _83857_ (_34067_, _34066_, _06033_);
  and _83858_ (_34068_, _34067_, _06027_);
  and _83859_ (_34070_, _34068_, _34064_);
  or _83860_ (_34071_, _34044_, _15074_);
  and _83861_ (_34072_, _34071_, _06026_);
  and _83862_ (_34073_, _34072_, _34046_);
  or _83863_ (_34074_, _34073_, _09818_);
  or _83864_ (_34075_, _34074_, _34070_);
  and _83865_ (_34076_, _09179_, _07688_);
  or _83866_ (_34077_, _34028_, _07012_);
  or _83867_ (_34078_, _34077_, _34076_);
  or _83868_ (_34079_, _34052_, _09827_);
  and _83869_ (_34081_, _34079_, _05669_);
  and _83870_ (_34082_, _34081_, _34078_);
  and _83871_ (_34083_, _34082_, _34075_);
  and _83872_ (_34084_, _15179_, _07688_);
  or _83873_ (_34085_, _34084_, _34028_);
  and _83874_ (_34086_, _34085_, _09833_);
  or _83875_ (_34087_, _34086_, _06019_);
  or _83876_ (_34088_, _34087_, _34083_);
  and _83877_ (_34089_, _34088_, _34031_);
  or _83878_ (_34090_, _34089_, _06112_);
  and _83879_ (_34092_, _15195_, _07688_);
  or _83880_ (_34093_, _34092_, _34028_);
  or _83881_ (_34094_, _34093_, _08751_);
  and _83882_ (_34095_, _34094_, _08756_);
  and _83883_ (_34096_, _34095_, _34090_);
  and _83884_ (_34097_, _12306_, _07688_);
  or _83885_ (_34098_, _34097_, _34028_);
  and _83886_ (_34099_, _34098_, _06284_);
  or _83887_ (_34100_, _34099_, _34096_);
  and _83888_ (_34101_, _34100_, _07032_);
  or _83889_ (_34103_, _34028_, _07980_);
  and _83890_ (_34104_, _34030_, _06108_);
  and _83891_ (_34105_, _34104_, _34103_);
  or _83892_ (_34106_, _34105_, _34101_);
  and _83893_ (_34107_, _34106_, _06278_);
  and _83894_ (_34108_, _34037_, _06277_);
  and _83895_ (_34109_, _34108_, _34103_);
  or _83896_ (_34110_, _34109_, _06130_);
  or _83897_ (_34111_, _34110_, _34107_);
  and _83898_ (_34112_, _15194_, _07688_);
  or _83899_ (_34113_, _34028_, _08777_);
  or _83900_ (_34114_, _34113_, _34112_);
  and _83901_ (_34115_, _34114_, _08782_);
  and _83902_ (_34116_, _34115_, _34111_);
  nor _83903_ (_34117_, _10982_, _13311_);
  or _83904_ (_34118_, _34117_, _34028_);
  and _83905_ (_34119_, _34118_, _06292_);
  or _83906_ (_34120_, _34119_, _06316_);
  or _83907_ (_34121_, _34120_, _34116_);
  or _83908_ (_34122_, _34033_, _06718_);
  and _83909_ (_34124_, _34122_, _05653_);
  and _83910_ (_34125_, _34124_, _34121_);
  and _83911_ (_34126_, _34061_, _05652_);
  or _83912_ (_34127_, _34126_, _06047_);
  or _83913_ (_34128_, _34127_, _34125_);
  and _83914_ (_34129_, _15253_, _07688_);
  or _83915_ (_34130_, _34028_, _06048_);
  or _83916_ (_34131_, _34130_, _34129_);
  and _83917_ (_34132_, _34131_, _01336_);
  and _83918_ (_34133_, _34132_, _34128_);
  or _83919_ (_34135_, _34133_, _34027_);
  and _83920_ (_43482_, _34135_, _42882_);
  and _83921_ (_34136_, _01340_, \oc8051_golden_model_1.IE [6]);
  and _83922_ (_34137_, _13311_, \oc8051_golden_model_1.IE [6]);
  and _83923_ (_34138_, _15389_, _07688_);
  or _83924_ (_34139_, _34138_, _34137_);
  or _83925_ (_34140_, _34139_, _06020_);
  and _83926_ (_34141_, _15293_, _07688_);
  or _83927_ (_34142_, _34141_, _34137_);
  or _83928_ (_34143_, _34142_, _06954_);
  and _83929_ (_34145_, _07688_, \oc8051_golden_model_1.ACC [6]);
  or _83930_ (_34146_, _34145_, _34137_);
  and _83931_ (_34147_, _34146_, _06938_);
  and _83932_ (_34148_, _06939_, \oc8051_golden_model_1.IE [6]);
  or _83933_ (_34149_, _34148_, _06102_);
  or _83934_ (_34150_, _34149_, _34147_);
  and _83935_ (_34151_, _34150_, _06044_);
  and _83936_ (_34152_, _34151_, _34143_);
  and _83937_ (_34153_, _13330_, \oc8051_golden_model_1.IE [6]);
  and _83938_ (_34154_, _15280_, _08351_);
  or _83939_ (_34156_, _34154_, _34153_);
  and _83940_ (_34157_, _34156_, _06043_);
  or _83941_ (_34158_, _34157_, _06239_);
  or _83942_ (_34159_, _34158_, _34152_);
  nor _83943_ (_34160_, _07883_, _13311_);
  or _83944_ (_34161_, _34160_, _34137_);
  or _83945_ (_34162_, _34161_, _06848_);
  and _83946_ (_34163_, _34162_, _34159_);
  or _83947_ (_34164_, _34163_, _06219_);
  or _83948_ (_34165_, _34146_, _06220_);
  and _83949_ (_34167_, _34165_, _06040_);
  and _83950_ (_34168_, _34167_, _34164_);
  and _83951_ (_34169_, _15278_, _08351_);
  or _83952_ (_34170_, _34169_, _34153_);
  and _83953_ (_34171_, _34170_, _06039_);
  or _83954_ (_34172_, _34171_, _06032_);
  or _83955_ (_34173_, _34172_, _34168_);
  or _83956_ (_34174_, _34153_, _15310_);
  and _83957_ (_34175_, _34174_, _34156_);
  or _83958_ (_34176_, _34175_, _06033_);
  and _83959_ (_34178_, _34176_, _06027_);
  and _83960_ (_34179_, _34178_, _34173_);
  or _83961_ (_34180_, _34153_, _15326_);
  and _83962_ (_34181_, _34180_, _06026_);
  and _83963_ (_34182_, _34181_, _34156_);
  or _83964_ (_34183_, _34182_, _09818_);
  or _83965_ (_34184_, _34183_, _34179_);
  and _83966_ (_34185_, _09178_, _07688_);
  or _83967_ (_34186_, _34137_, _07012_);
  or _83968_ (_34187_, _34186_, _34185_);
  or _83969_ (_34189_, _34161_, _09827_);
  and _83970_ (_34190_, _34189_, _05669_);
  and _83971_ (_34191_, _34190_, _34187_);
  and _83972_ (_34192_, _34191_, _34184_);
  and _83973_ (_34193_, _15382_, _07688_);
  or _83974_ (_34194_, _34193_, _34137_);
  and _83975_ (_34195_, _34194_, _09833_);
  or _83976_ (_34196_, _34195_, _06019_);
  or _83977_ (_34197_, _34196_, _34192_);
  and _83978_ (_34198_, _34197_, _34140_);
  or _83979_ (_34200_, _34198_, _06112_);
  and _83980_ (_34201_, _15399_, _07688_);
  or _83981_ (_34202_, _34201_, _34137_);
  or _83982_ (_34203_, _34202_, _08751_);
  and _83983_ (_34204_, _34203_, _08756_);
  and _83984_ (_34205_, _34204_, _34200_);
  and _83985_ (_34206_, _10980_, _07688_);
  or _83986_ (_34207_, _34206_, _34137_);
  and _83987_ (_34208_, _34207_, _06284_);
  or _83988_ (_34209_, _34208_, _34205_);
  and _83989_ (_34211_, _34209_, _07032_);
  or _83990_ (_34212_, _34137_, _07886_);
  and _83991_ (_34213_, _34139_, _06108_);
  and _83992_ (_34214_, _34213_, _34212_);
  or _83993_ (_34215_, _34214_, _34211_);
  and _83994_ (_34216_, _34215_, _06278_);
  and _83995_ (_34217_, _34146_, _06277_);
  and _83996_ (_34218_, _34217_, _34212_);
  or _83997_ (_34219_, _34218_, _06130_);
  or _83998_ (_34220_, _34219_, _34216_);
  and _83999_ (_34222_, _15396_, _07688_);
  or _84000_ (_34223_, _34137_, _08777_);
  or _84001_ (_34224_, _34223_, _34222_);
  and _84002_ (_34225_, _34224_, _08782_);
  and _84003_ (_34226_, _34225_, _34220_);
  nor _84004_ (_34227_, _10979_, _13311_);
  or _84005_ (_34228_, _34227_, _34137_);
  and _84006_ (_34229_, _34228_, _06292_);
  or _84007_ (_34230_, _34229_, _06316_);
  or _84008_ (_34231_, _34230_, _34226_);
  or _84009_ (_34233_, _34142_, _06718_);
  and _84010_ (_34234_, _34233_, _05653_);
  and _84011_ (_34235_, _34234_, _34231_);
  and _84012_ (_34236_, _34170_, _05652_);
  or _84013_ (_34237_, _34236_, _06047_);
  or _84014_ (_34238_, _34237_, _34235_);
  and _84015_ (_34239_, _15451_, _07688_);
  or _84016_ (_34240_, _34137_, _06048_);
  or _84017_ (_34241_, _34240_, _34239_);
  and _84018_ (_34242_, _34241_, _01336_);
  and _84019_ (_34244_, _34242_, _34238_);
  or _84020_ (_34245_, _34244_, _34136_);
  and _84021_ (_43483_, _34245_, _42882_);
  and _84022_ (_34246_, _01340_, \oc8051_golden_model_1.SCON [0]);
  and _84023_ (_34247_, _07679_, \oc8051_golden_model_1.ACC [0]);
  and _84024_ (_34248_, _34247_, _08127_);
  and _84025_ (_34249_, _13413_, \oc8051_golden_model_1.SCON [0]);
  or _84026_ (_34250_, _34249_, _06278_);
  or _84027_ (_34251_, _34250_, _34248_);
  and _84028_ (_34252_, _07679_, _08672_);
  or _84029_ (_34254_, _34252_, _34249_);
  or _84030_ (_34255_, _34254_, _06020_);
  and _84031_ (_34256_, _09120_, _07679_);
  or _84032_ (_34257_, _34249_, _07012_);
  or _84033_ (_34258_, _34257_, _34256_);
  nor _84034_ (_34259_, _08127_, _13413_);
  or _84035_ (_34260_, _34259_, _34249_);
  or _84036_ (_34261_, _34260_, _06954_);
  or _84037_ (_34262_, _34247_, _34249_);
  and _84038_ (_34263_, _34262_, _06938_);
  and _84039_ (_34265_, _06939_, \oc8051_golden_model_1.SCON [0]);
  or _84040_ (_34266_, _34265_, _06102_);
  or _84041_ (_34267_, _34266_, _34263_);
  and _84042_ (_34268_, _34267_, _06044_);
  and _84043_ (_34269_, _34268_, _34261_);
  and _84044_ (_34270_, _13432_, \oc8051_golden_model_1.SCON [0]);
  and _84045_ (_34271_, _14102_, _08347_);
  or _84046_ (_34272_, _34271_, _34270_);
  and _84047_ (_34274_, _34272_, _06043_);
  or _84048_ (_34276_, _34274_, _34269_);
  and _84049_ (_34279_, _34276_, _06848_);
  and _84050_ (_34281_, _07679_, _06931_);
  or _84051_ (_34283_, _34281_, _34249_);
  and _84052_ (_34285_, _34283_, _06239_);
  or _84053_ (_34287_, _34285_, _06219_);
  or _84054_ (_34289_, _34287_, _34279_);
  or _84055_ (_34291_, _34262_, _06220_);
  and _84056_ (_34293_, _34291_, _06040_);
  and _84057_ (_34294_, _34293_, _34289_);
  and _84058_ (_34295_, _34249_, _06039_);
  or _84059_ (_34297_, _34295_, _06032_);
  or _84060_ (_34298_, _34297_, _34294_);
  or _84061_ (_34299_, _34260_, _06033_);
  and _84062_ (_34300_, _34299_, _06027_);
  and _84063_ (_34301_, _34300_, _34298_);
  or _84064_ (_34302_, _34270_, _14131_);
  and _84065_ (_34303_, _34302_, _06026_);
  and _84066_ (_34304_, _34303_, _34272_);
  or _84067_ (_34305_, _34304_, _09818_);
  or _84068_ (_34306_, _34305_, _34301_);
  or _84069_ (_34308_, _34283_, _09827_);
  and _84070_ (_34309_, _34308_, _05669_);
  and _84071_ (_34310_, _34309_, _34306_);
  and _84072_ (_34311_, _34310_, _34258_);
  and _84073_ (_34312_, _14186_, _07679_);
  or _84074_ (_34313_, _34312_, _34249_);
  and _84075_ (_34314_, _34313_, _09833_);
  or _84076_ (_34315_, _34314_, _06019_);
  or _84077_ (_34316_, _34315_, _34311_);
  and _84078_ (_34317_, _34316_, _34255_);
  or _84079_ (_34319_, _34317_, _06112_);
  and _84080_ (_34320_, _14086_, _07679_);
  or _84081_ (_34321_, _34249_, _08751_);
  or _84082_ (_34322_, _34321_, _34320_);
  and _84083_ (_34323_, _34322_, _08756_);
  and _84084_ (_34324_, _34323_, _34319_);
  nor _84085_ (_34325_, _12302_, _13413_);
  or _84086_ (_34326_, _34325_, _34249_);
  nor _84087_ (_34327_, _34248_, _08756_);
  and _84088_ (_34328_, _34327_, _34326_);
  or _84089_ (_34330_, _34328_, _34324_);
  and _84090_ (_34331_, _34330_, _07032_);
  nand _84091_ (_34332_, _34254_, _06108_);
  nor _84092_ (_34333_, _34332_, _34259_);
  or _84093_ (_34334_, _34333_, _06277_);
  or _84094_ (_34335_, _34334_, _34331_);
  and _84095_ (_34336_, _34335_, _34251_);
  or _84096_ (_34337_, _34336_, _06130_);
  and _84097_ (_34338_, _14083_, _07679_);
  or _84098_ (_34339_, _34249_, _08777_);
  or _84099_ (_34341_, _34339_, _34338_);
  and _84100_ (_34342_, _34341_, _08782_);
  and _84101_ (_34343_, _34342_, _34337_);
  and _84102_ (_34344_, _34326_, _06292_);
  or _84103_ (_34345_, _34344_, _06316_);
  or _84104_ (_34346_, _34345_, _34343_);
  or _84105_ (_34347_, _34260_, _06718_);
  and _84106_ (_34348_, _34347_, _34346_);
  or _84107_ (_34349_, _34348_, _05652_);
  or _84108_ (_34350_, _34249_, _05653_);
  and _84109_ (_34352_, _34350_, _34349_);
  or _84110_ (_34353_, _34352_, _06047_);
  or _84111_ (_34354_, _34260_, _06048_);
  and _84112_ (_34355_, _34354_, _01336_);
  and _84113_ (_34356_, _34355_, _34353_);
  or _84114_ (_34357_, _34356_, _34246_);
  and _84115_ (_43484_, _34357_, _42882_);
  not _84116_ (_34358_, \oc8051_golden_model_1.SCON [1]);
  nor _84117_ (_34359_, _01336_, _34358_);
  nor _84118_ (_34360_, _07679_, _34358_);
  nor _84119_ (_34362_, _10993_, _13413_);
  or _84120_ (_34363_, _34362_, _34360_);
  or _84121_ (_34364_, _34363_, _08782_);
  nor _84122_ (_34365_, _13413_, _07132_);
  or _84123_ (_34366_, _34365_, _34360_);
  or _84124_ (_34367_, _34366_, _06848_);
  or _84125_ (_34368_, _07679_, \oc8051_golden_model_1.SCON [1]);
  and _84126_ (_34369_, _14284_, _07679_);
  not _84127_ (_34370_, _34369_);
  and _84128_ (_34371_, _34370_, _34368_);
  or _84129_ (_34373_, _34371_, _06954_);
  and _84130_ (_34374_, _07679_, \oc8051_golden_model_1.ACC [1]);
  or _84131_ (_34375_, _34374_, _34360_);
  and _84132_ (_34376_, _34375_, _06938_);
  nor _84133_ (_34377_, _06938_, _34358_);
  or _84134_ (_34378_, _34377_, _06102_);
  or _84135_ (_34379_, _34378_, _34376_);
  and _84136_ (_34380_, _34379_, _06044_);
  and _84137_ (_34381_, _34380_, _34373_);
  nor _84138_ (_34382_, _08347_, _34358_);
  and _84139_ (_34384_, _14266_, _08347_);
  or _84140_ (_34385_, _34384_, _34382_);
  and _84141_ (_34386_, _34385_, _06043_);
  or _84142_ (_34387_, _34386_, _06239_);
  or _84143_ (_34388_, _34387_, _34381_);
  and _84144_ (_34389_, _34388_, _34367_);
  or _84145_ (_34390_, _34389_, _06219_);
  or _84146_ (_34391_, _34375_, _06220_);
  and _84147_ (_34392_, _34391_, _06040_);
  and _84148_ (_34393_, _34392_, _34390_);
  and _84149_ (_34395_, _14273_, _08347_);
  or _84150_ (_34396_, _34395_, _34382_);
  and _84151_ (_34397_, _34396_, _06039_);
  or _84152_ (_34398_, _34397_, _06032_);
  or _84153_ (_34399_, _34398_, _34393_);
  and _84154_ (_34400_, _34384_, _14302_);
  or _84155_ (_34401_, _34382_, _06033_);
  or _84156_ (_34402_, _34401_, _34400_);
  and _84157_ (_34403_, _34402_, _06027_);
  and _84158_ (_34404_, _34403_, _34399_);
  or _84159_ (_34406_, _34382_, _14267_);
  and _84160_ (_34407_, _34406_, _06026_);
  and _84161_ (_34408_, _34407_, _34385_);
  or _84162_ (_34409_, _34408_, _09818_);
  or _84163_ (_34410_, _34409_, _34404_);
  and _84164_ (_34411_, _09075_, _07679_);
  or _84165_ (_34412_, _34360_, _07012_);
  or _84166_ (_34413_, _34412_, _34411_);
  or _84167_ (_34414_, _34366_, _09827_);
  and _84168_ (_34415_, _34414_, _05669_);
  and _84169_ (_34417_, _34415_, _34413_);
  and _84170_ (_34418_, _34417_, _34410_);
  and _84171_ (_34419_, _14367_, _07679_);
  or _84172_ (_34420_, _34419_, _34360_);
  and _84173_ (_34421_, _34420_, _09833_);
  or _84174_ (_34422_, _34421_, _34418_);
  and _84175_ (_34423_, _34422_, _06020_);
  nand _84176_ (_34424_, _07679_, _06832_);
  and _84177_ (_34425_, _34368_, _06019_);
  and _84178_ (_34426_, _34425_, _34424_);
  or _84179_ (_34428_, _34426_, _34423_);
  and _84180_ (_34429_, _34428_, _08751_);
  or _84181_ (_34430_, _14263_, _13413_);
  and _84182_ (_34431_, _34368_, _06112_);
  and _84183_ (_34432_, _34431_, _34430_);
  or _84184_ (_34433_, _34432_, _06284_);
  or _84185_ (_34434_, _34433_, _34429_);
  nand _84186_ (_34435_, _10992_, _07679_);
  and _84187_ (_34436_, _34435_, _34363_);
  or _84188_ (_34437_, _34436_, _08756_);
  and _84189_ (_34439_, _34437_, _07032_);
  and _84190_ (_34440_, _34439_, _34434_);
  or _84191_ (_34441_, _14261_, _13413_);
  and _84192_ (_34442_, _34368_, _06108_);
  and _84193_ (_34443_, _34442_, _34441_);
  or _84194_ (_34444_, _34443_, _06277_);
  or _84195_ (_34445_, _34444_, _34440_);
  nor _84196_ (_34446_, _34360_, _06278_);
  nand _84197_ (_34447_, _34446_, _34435_);
  and _84198_ (_34448_, _34447_, _08777_);
  and _84199_ (_34450_, _34448_, _34445_);
  or _84200_ (_34451_, _34424_, _08078_);
  and _84201_ (_34452_, _34368_, _06130_);
  and _84202_ (_34453_, _34452_, _34451_);
  or _84203_ (_34454_, _34453_, _06292_);
  or _84204_ (_34455_, _34454_, _34450_);
  and _84205_ (_34456_, _34455_, _34364_);
  or _84206_ (_34457_, _34456_, _06316_);
  or _84207_ (_34458_, _34371_, _06718_);
  and _84208_ (_34459_, _34458_, _05653_);
  and _84209_ (_34461_, _34459_, _34457_);
  and _84210_ (_34462_, _34396_, _05652_);
  or _84211_ (_34463_, _34462_, _06047_);
  or _84212_ (_34464_, _34463_, _34461_);
  or _84213_ (_34465_, _34360_, _06048_);
  or _84214_ (_34466_, _34465_, _34369_);
  and _84215_ (_34467_, _34466_, _01336_);
  and _84216_ (_34468_, _34467_, _34464_);
  or _84217_ (_34469_, _34468_, _34359_);
  and _84218_ (_43486_, _34469_, _42882_);
  and _84219_ (_34471_, _01340_, \oc8051_golden_model_1.SCON [2]);
  and _84220_ (_34472_, _13413_, \oc8051_golden_model_1.SCON [2]);
  and _84221_ (_34473_, _07679_, _08730_);
  or _84222_ (_34474_, _34473_, _34472_);
  or _84223_ (_34475_, _34474_, _06020_);
  nor _84224_ (_34476_, _13413_, _07530_);
  or _84225_ (_34477_, _34476_, _34472_);
  and _84226_ (_34478_, _34477_, _06239_);
  and _84227_ (_34479_, _13432_, \oc8051_golden_model_1.SCON [2]);
  and _84228_ (_34480_, _14497_, _08347_);
  or _84229_ (_34482_, _34480_, _34479_);
  or _84230_ (_34483_, _34482_, _06044_);
  and _84231_ (_34484_, _14493_, _07679_);
  or _84232_ (_34485_, _34484_, _34472_);
  and _84233_ (_34486_, _34485_, _06102_);
  and _84234_ (_34487_, _06939_, \oc8051_golden_model_1.SCON [2]);
  and _84235_ (_34488_, _07679_, \oc8051_golden_model_1.ACC [2]);
  or _84236_ (_34489_, _34488_, _34472_);
  and _84237_ (_34490_, _34489_, _06938_);
  or _84238_ (_34491_, _34490_, _34487_);
  and _84239_ (_34493_, _34491_, _06954_);
  or _84240_ (_34494_, _34493_, _06043_);
  or _84241_ (_34495_, _34494_, _34486_);
  and _84242_ (_34496_, _34495_, _34483_);
  and _84243_ (_34497_, _34496_, _06848_);
  or _84244_ (_34498_, _34497_, _34478_);
  or _84245_ (_34499_, _34498_, _06219_);
  or _84246_ (_34500_, _34489_, _06220_);
  and _84247_ (_34501_, _34500_, _06040_);
  and _84248_ (_34502_, _34501_, _34499_);
  and _84249_ (_34504_, _14479_, _08347_);
  or _84250_ (_34505_, _34504_, _34479_);
  and _84251_ (_34506_, _34505_, _06039_);
  or _84252_ (_34507_, _34506_, _06032_);
  or _84253_ (_34508_, _34507_, _34502_);
  or _84254_ (_34509_, _34479_, _14512_);
  and _84255_ (_34510_, _34509_, _34482_);
  or _84256_ (_34511_, _34510_, _06033_);
  and _84257_ (_34512_, _34511_, _06027_);
  and _84258_ (_34513_, _34512_, _34508_);
  or _84259_ (_34515_, _34479_, _14525_);
  and _84260_ (_34516_, _34515_, _06026_);
  and _84261_ (_34517_, _34516_, _34482_);
  or _84262_ (_34518_, _34517_, _09818_);
  or _84263_ (_34519_, _34518_, _34513_);
  and _84264_ (_34520_, _09182_, _07679_);
  or _84265_ (_34521_, _34472_, _07012_);
  or _84266_ (_34522_, _34521_, _34520_);
  or _84267_ (_34523_, _34477_, _09827_);
  and _84268_ (_34524_, _34523_, _05669_);
  and _84269_ (_34526_, _34524_, _34522_);
  and _84270_ (_34527_, _34526_, _34519_);
  and _84271_ (_34528_, _14580_, _07679_);
  or _84272_ (_34529_, _34528_, _34472_);
  and _84273_ (_34530_, _34529_, _09833_);
  or _84274_ (_34531_, _34530_, _06019_);
  or _84275_ (_34532_, _34531_, _34527_);
  and _84276_ (_34533_, _34532_, _34475_);
  or _84277_ (_34534_, _34533_, _06112_);
  and _84278_ (_34535_, _14596_, _07679_);
  or _84279_ (_34537_, _34535_, _34472_);
  or _84280_ (_34538_, _34537_, _08751_);
  and _84281_ (_34539_, _34538_, _08756_);
  and _84282_ (_34540_, _34539_, _34534_);
  and _84283_ (_34541_, _10991_, _07679_);
  or _84284_ (_34542_, _34541_, _34472_);
  and _84285_ (_34543_, _34542_, _06284_);
  or _84286_ (_34544_, _34543_, _34540_);
  and _84287_ (_34545_, _34544_, _07032_);
  or _84288_ (_34546_, _34472_, _08177_);
  and _84289_ (_34548_, _34474_, _06108_);
  and _84290_ (_34549_, _34548_, _34546_);
  or _84291_ (_34550_, _34549_, _34545_);
  and _84292_ (_34551_, _34550_, _06278_);
  and _84293_ (_34552_, _34489_, _06277_);
  and _84294_ (_34553_, _34552_, _34546_);
  or _84295_ (_34554_, _34553_, _06130_);
  or _84296_ (_34555_, _34554_, _34551_);
  and _84297_ (_34556_, _14593_, _07679_);
  or _84298_ (_34557_, _34472_, _08777_);
  or _84299_ (_34559_, _34557_, _34556_);
  and _84300_ (_34560_, _34559_, _08782_);
  and _84301_ (_34561_, _34560_, _34555_);
  nor _84302_ (_34562_, _10990_, _13413_);
  or _84303_ (_34563_, _34562_, _34472_);
  and _84304_ (_34564_, _34563_, _06292_);
  or _84305_ (_34565_, _34564_, _06316_);
  or _84306_ (_34566_, _34565_, _34561_);
  or _84307_ (_34567_, _34485_, _06718_);
  and _84308_ (_34568_, _34567_, _05653_);
  and _84309_ (_34570_, _34568_, _34566_);
  and _84310_ (_34571_, _34505_, _05652_);
  or _84311_ (_34572_, _34571_, _06047_);
  or _84312_ (_34573_, _34572_, _34570_);
  and _84313_ (_34574_, _14657_, _07679_);
  or _84314_ (_34575_, _34472_, _06048_);
  or _84315_ (_34576_, _34575_, _34574_);
  and _84316_ (_34577_, _34576_, _01336_);
  and _84317_ (_34578_, _34577_, _34573_);
  or _84318_ (_34579_, _34578_, _34471_);
  and _84319_ (_43487_, _34579_, _42882_);
  and _84320_ (_34581_, _01340_, \oc8051_golden_model_1.SCON [3]);
  and _84321_ (_34582_, _13413_, \oc8051_golden_model_1.SCON [3]);
  and _84322_ (_34583_, _07679_, _08662_);
  or _84323_ (_34584_, _34583_, _34582_);
  or _84324_ (_34585_, _34584_, _06020_);
  and _84325_ (_34586_, _14672_, _07679_);
  or _84326_ (_34587_, _34586_, _34582_);
  or _84327_ (_34588_, _34587_, _06954_);
  and _84328_ (_34589_, _07679_, \oc8051_golden_model_1.ACC [3]);
  or _84329_ (_34591_, _34589_, _34582_);
  and _84330_ (_34592_, _34591_, _06938_);
  and _84331_ (_34593_, _06939_, \oc8051_golden_model_1.SCON [3]);
  or _84332_ (_34594_, _34593_, _06102_);
  or _84333_ (_34595_, _34594_, _34592_);
  and _84334_ (_34596_, _34595_, _06044_);
  and _84335_ (_34597_, _34596_, _34588_);
  and _84336_ (_34598_, _13432_, \oc8051_golden_model_1.SCON [3]);
  and _84337_ (_34599_, _14683_, _08347_);
  or _84338_ (_34600_, _34599_, _34598_);
  and _84339_ (_34602_, _34600_, _06043_);
  or _84340_ (_34603_, _34602_, _06239_);
  or _84341_ (_34604_, _34603_, _34597_);
  nor _84342_ (_34605_, _13413_, _07353_);
  or _84343_ (_34606_, _34605_, _34582_);
  or _84344_ (_34607_, _34606_, _06848_);
  and _84345_ (_34608_, _34607_, _34604_);
  or _84346_ (_34609_, _34608_, _06219_);
  or _84347_ (_34610_, _34591_, _06220_);
  and _84348_ (_34611_, _34610_, _06040_);
  and _84349_ (_34613_, _34611_, _34609_);
  and _84350_ (_34614_, _14681_, _08347_);
  or _84351_ (_34615_, _34614_, _34598_);
  and _84352_ (_34616_, _34615_, _06039_);
  or _84353_ (_34617_, _34616_, _06032_);
  or _84354_ (_34618_, _34617_, _34613_);
  or _84355_ (_34619_, _34598_, _14708_);
  and _84356_ (_34620_, _34619_, _34600_);
  or _84357_ (_34621_, _34620_, _06033_);
  and _84358_ (_34622_, _34621_, _06027_);
  and _84359_ (_34624_, _34622_, _34618_);
  and _84360_ (_34625_, _14724_, _08347_);
  or _84361_ (_34626_, _34625_, _34598_);
  and _84362_ (_34627_, _34626_, _06026_);
  or _84363_ (_34628_, _34627_, _09818_);
  or _84364_ (_34629_, _34628_, _34624_);
  and _84365_ (_34630_, _09181_, _07679_);
  or _84366_ (_34631_, _34582_, _07012_);
  or _84367_ (_34632_, _34631_, _34630_);
  or _84368_ (_34633_, _34606_, _09827_);
  and _84369_ (_34635_, _34633_, _05669_);
  and _84370_ (_34636_, _34635_, _34632_);
  and _84371_ (_34637_, _34636_, _34629_);
  and _84372_ (_34638_, _14778_, _07679_);
  or _84373_ (_34639_, _34638_, _34582_);
  and _84374_ (_34640_, _34639_, _09833_);
  or _84375_ (_34641_, _34640_, _06019_);
  or _84376_ (_34642_, _34641_, _34637_);
  and _84377_ (_34643_, _34642_, _34585_);
  or _84378_ (_34644_, _34643_, _06112_);
  and _84379_ (_34646_, _14793_, _07679_);
  or _84380_ (_34647_, _34582_, _08751_);
  or _84381_ (_34648_, _34647_, _34646_);
  and _84382_ (_34649_, _34648_, _08756_);
  and _84383_ (_34650_, _34649_, _34644_);
  and _84384_ (_34651_, _12299_, _07679_);
  or _84385_ (_34652_, _34651_, _34582_);
  and _84386_ (_34653_, _34652_, _06284_);
  or _84387_ (_34654_, _34653_, _34650_);
  and _84388_ (_34655_, _34654_, _07032_);
  or _84389_ (_34657_, _34582_, _08029_);
  and _84390_ (_34658_, _34584_, _06108_);
  and _84391_ (_34659_, _34658_, _34657_);
  or _84392_ (_34660_, _34659_, _34655_);
  and _84393_ (_34661_, _34660_, _06278_);
  and _84394_ (_34662_, _34591_, _06277_);
  and _84395_ (_34663_, _34662_, _34657_);
  or _84396_ (_34664_, _34663_, _06130_);
  or _84397_ (_34665_, _34664_, _34661_);
  and _84398_ (_34666_, _14792_, _07679_);
  or _84399_ (_34668_, _34582_, _08777_);
  or _84400_ (_34669_, _34668_, _34666_);
  and _84401_ (_34670_, _34669_, _08782_);
  and _84402_ (_34671_, _34670_, _34665_);
  nor _84403_ (_34672_, _10988_, _13413_);
  or _84404_ (_34673_, _34672_, _34582_);
  and _84405_ (_34674_, _34673_, _06292_);
  or _84406_ (_34675_, _34674_, _06316_);
  or _84407_ (_34676_, _34675_, _34671_);
  or _84408_ (_34677_, _34587_, _06718_);
  and _84409_ (_34679_, _34677_, _05653_);
  and _84410_ (_34680_, _34679_, _34676_);
  and _84411_ (_34681_, _34615_, _05652_);
  or _84412_ (_34682_, _34681_, _06047_);
  or _84413_ (_34683_, _34682_, _34680_);
  and _84414_ (_34684_, _14849_, _07679_);
  or _84415_ (_34685_, _34582_, _06048_);
  or _84416_ (_34686_, _34685_, _34684_);
  and _84417_ (_34687_, _34686_, _01336_);
  and _84418_ (_34688_, _34687_, _34683_);
  or _84419_ (_34690_, _34688_, _34581_);
  and _84420_ (_43488_, _34690_, _42882_);
  and _84421_ (_34691_, _01340_, \oc8051_golden_model_1.SCON [4]);
  and _84422_ (_34692_, _13413_, \oc8051_golden_model_1.SCON [4]);
  and _84423_ (_34693_, _08665_, _07679_);
  or _84424_ (_34694_, _34693_, _34692_);
  or _84425_ (_34695_, _34694_, _06020_);
  and _84426_ (_34696_, _14887_, _07679_);
  or _84427_ (_34697_, _34696_, _34692_);
  or _84428_ (_34698_, _34697_, _06954_);
  and _84429_ (_34700_, _07679_, \oc8051_golden_model_1.ACC [4]);
  or _84430_ (_34701_, _34700_, _34692_);
  and _84431_ (_34702_, _34701_, _06938_);
  and _84432_ (_34703_, _06939_, \oc8051_golden_model_1.SCON [4]);
  or _84433_ (_34704_, _34703_, _06102_);
  or _84434_ (_34705_, _34704_, _34702_);
  and _84435_ (_34706_, _34705_, _06044_);
  and _84436_ (_34707_, _34706_, _34698_);
  and _84437_ (_34708_, _13432_, \oc8051_golden_model_1.SCON [4]);
  and _84438_ (_34709_, _14878_, _08347_);
  or _84439_ (_34711_, _34709_, _34708_);
  and _84440_ (_34712_, _34711_, _06043_);
  or _84441_ (_34713_, _34712_, _06239_);
  or _84442_ (_34714_, _34713_, _34707_);
  nor _84443_ (_34715_, _08270_, _13413_);
  or _84444_ (_34716_, _34715_, _34692_);
  or _84445_ (_34717_, _34716_, _06848_);
  and _84446_ (_34718_, _34717_, _34714_);
  or _84447_ (_34719_, _34718_, _06219_);
  or _84448_ (_34720_, _34701_, _06220_);
  and _84449_ (_34722_, _34720_, _06040_);
  and _84450_ (_34723_, _34722_, _34719_);
  and _84451_ (_34724_, _14882_, _08347_);
  or _84452_ (_34725_, _34724_, _34708_);
  and _84453_ (_34726_, _34725_, _06039_);
  or _84454_ (_34727_, _34726_, _06032_);
  or _84455_ (_34728_, _34727_, _34723_);
  or _84456_ (_34729_, _34708_, _14914_);
  and _84457_ (_34730_, _34729_, _34711_);
  or _84458_ (_34731_, _34730_, _06033_);
  and _84459_ (_34733_, _34731_, _06027_);
  and _84460_ (_34734_, _34733_, _34728_);
  or _84461_ (_34735_, _34708_, _14879_);
  and _84462_ (_34736_, _34735_, _06026_);
  and _84463_ (_34737_, _34736_, _34711_);
  or _84464_ (_34738_, _34737_, _09818_);
  or _84465_ (_34739_, _34738_, _34734_);
  and _84466_ (_34740_, _09180_, _07679_);
  or _84467_ (_34741_, _34692_, _07012_);
  or _84468_ (_34742_, _34741_, _34740_);
  or _84469_ (_34744_, _34716_, _09827_);
  and _84470_ (_34745_, _34744_, _05669_);
  and _84471_ (_34746_, _34745_, _34742_);
  and _84472_ (_34747_, _34746_, _34739_);
  and _84473_ (_34748_, _14983_, _07679_);
  or _84474_ (_34749_, _34748_, _34692_);
  and _84475_ (_34750_, _34749_, _09833_);
  or _84476_ (_34751_, _34750_, _06019_);
  or _84477_ (_34752_, _34751_, _34747_);
  and _84478_ (_34753_, _34752_, _34695_);
  or _84479_ (_34755_, _34753_, _06112_);
  and _84480_ (_34756_, _14876_, _07679_);
  or _84481_ (_34757_, _34756_, _34692_);
  or _84482_ (_34758_, _34757_, _08751_);
  and _84483_ (_34759_, _34758_, _08756_);
  and _84484_ (_34760_, _34759_, _34755_);
  and _84485_ (_34761_, _10986_, _07679_);
  or _84486_ (_34762_, _34761_, _34692_);
  and _84487_ (_34763_, _34762_, _06284_);
  or _84488_ (_34764_, _34763_, _34760_);
  and _84489_ (_34766_, _34764_, _07032_);
  or _84490_ (_34767_, _34692_, _08273_);
  and _84491_ (_34768_, _34694_, _06108_);
  and _84492_ (_34769_, _34768_, _34767_);
  or _84493_ (_34770_, _34769_, _34766_);
  and _84494_ (_34771_, _34770_, _06278_);
  and _84495_ (_34772_, _34701_, _06277_);
  and _84496_ (_34773_, _34772_, _34767_);
  or _84497_ (_34774_, _34773_, _06130_);
  or _84498_ (_34775_, _34774_, _34771_);
  and _84499_ (_34777_, _14873_, _07679_);
  or _84500_ (_34778_, _34692_, _08777_);
  or _84501_ (_34779_, _34778_, _34777_);
  and _84502_ (_34780_, _34779_, _08782_);
  and _84503_ (_34781_, _34780_, _34775_);
  nor _84504_ (_34782_, _10985_, _13413_);
  or _84505_ (_34783_, _34782_, _34692_);
  and _84506_ (_34784_, _34783_, _06292_);
  or _84507_ (_34785_, _34784_, _06316_);
  or _84508_ (_34786_, _34785_, _34781_);
  or _84509_ (_34788_, _34697_, _06718_);
  and _84510_ (_34789_, _34788_, _05653_);
  and _84511_ (_34790_, _34789_, _34786_);
  and _84512_ (_34791_, _34725_, _05652_);
  or _84513_ (_34792_, _34791_, _06047_);
  or _84514_ (_34793_, _34792_, _34790_);
  and _84515_ (_34794_, _15055_, _07679_);
  or _84516_ (_34795_, _34692_, _06048_);
  or _84517_ (_34796_, _34795_, _34794_);
  and _84518_ (_34797_, _34796_, _01336_);
  and _84519_ (_34799_, _34797_, _34793_);
  or _84520_ (_34800_, _34799_, _34691_);
  and _84521_ (_43489_, _34800_, _42882_);
  and _84522_ (_34801_, _01340_, \oc8051_golden_model_1.SCON [5]);
  and _84523_ (_34802_, _13413_, \oc8051_golden_model_1.SCON [5]);
  and _84524_ (_34803_, _08652_, _07679_);
  or _84525_ (_34804_, _34803_, _34802_);
  or _84526_ (_34805_, _34804_, _06020_);
  and _84527_ (_34806_, _15093_, _07679_);
  or _84528_ (_34807_, _34806_, _34802_);
  or _84529_ (_34809_, _34807_, _06954_);
  and _84530_ (_34810_, _07679_, \oc8051_golden_model_1.ACC [5]);
  or _84531_ (_34811_, _34810_, _34802_);
  and _84532_ (_34812_, _34811_, _06938_);
  and _84533_ (_34813_, _06939_, \oc8051_golden_model_1.SCON [5]);
  or _84534_ (_34814_, _34813_, _06102_);
  or _84535_ (_34815_, _34814_, _34812_);
  and _84536_ (_34816_, _34815_, _06044_);
  and _84537_ (_34817_, _34816_, _34809_);
  and _84538_ (_34818_, _13432_, \oc8051_golden_model_1.SCON [5]);
  and _84539_ (_34820_, _15073_, _08347_);
  or _84540_ (_34821_, _34820_, _34818_);
  and _84541_ (_34822_, _34821_, _06043_);
  or _84542_ (_34823_, _34822_, _06239_);
  or _84543_ (_34824_, _34823_, _34817_);
  nor _84544_ (_34825_, _07977_, _13413_);
  or _84545_ (_34826_, _34825_, _34802_);
  or _84546_ (_34827_, _34826_, _06848_);
  and _84547_ (_34828_, _34827_, _34824_);
  or _84548_ (_34829_, _34828_, _06219_);
  or _84549_ (_34831_, _34811_, _06220_);
  and _84550_ (_34832_, _34831_, _06040_);
  and _84551_ (_34833_, _34832_, _34829_);
  and _84552_ (_34834_, _15077_, _08347_);
  or _84553_ (_34835_, _34834_, _34818_);
  and _84554_ (_34836_, _34835_, _06039_);
  or _84555_ (_34837_, _34836_, _06032_);
  or _84556_ (_34838_, _34837_, _34833_);
  or _84557_ (_34839_, _34818_, _15110_);
  and _84558_ (_34840_, _34839_, _34821_);
  or _84559_ (_34842_, _34840_, _06033_);
  and _84560_ (_34843_, _34842_, _06027_);
  and _84561_ (_34844_, _34843_, _34838_);
  or _84562_ (_34845_, _34818_, _15074_);
  and _84563_ (_34846_, _34845_, _06026_);
  and _84564_ (_34847_, _34846_, _34821_);
  or _84565_ (_34848_, _34847_, _09818_);
  or _84566_ (_34849_, _34848_, _34844_);
  and _84567_ (_34850_, _09179_, _07679_);
  or _84568_ (_34851_, _34802_, _07012_);
  or _84569_ (_34853_, _34851_, _34850_);
  or _84570_ (_34854_, _34826_, _09827_);
  and _84571_ (_34855_, _34854_, _05669_);
  and _84572_ (_34856_, _34855_, _34853_);
  and _84573_ (_34857_, _34856_, _34849_);
  and _84574_ (_34858_, _15179_, _07679_);
  or _84575_ (_34859_, _34858_, _34802_);
  and _84576_ (_34860_, _34859_, _09833_);
  or _84577_ (_34861_, _34860_, _06019_);
  or _84578_ (_34862_, _34861_, _34857_);
  and _84579_ (_34864_, _34862_, _34805_);
  or _84580_ (_34865_, _34864_, _06112_);
  and _84581_ (_34866_, _15195_, _07679_);
  or _84582_ (_34867_, _34802_, _08751_);
  or _84583_ (_34868_, _34867_, _34866_);
  and _84584_ (_34869_, _34868_, _08756_);
  and _84585_ (_34870_, _34869_, _34865_);
  and _84586_ (_34871_, _12306_, _07679_);
  or _84587_ (_34872_, _34871_, _34802_);
  and _84588_ (_34873_, _34872_, _06284_);
  or _84589_ (_34875_, _34873_, _34870_);
  and _84590_ (_34876_, _34875_, _07032_);
  or _84591_ (_34877_, _34802_, _07980_);
  and _84592_ (_34878_, _34804_, _06108_);
  and _84593_ (_34879_, _34878_, _34877_);
  or _84594_ (_34880_, _34879_, _34876_);
  and _84595_ (_34881_, _34880_, _06278_);
  and _84596_ (_34882_, _34811_, _06277_);
  and _84597_ (_34883_, _34882_, _34877_);
  or _84598_ (_34884_, _34883_, _06130_);
  or _84599_ (_34886_, _34884_, _34881_);
  and _84600_ (_34887_, _15194_, _07679_);
  or _84601_ (_34888_, _34802_, _08777_);
  or _84602_ (_34889_, _34888_, _34887_);
  and _84603_ (_34890_, _34889_, _08782_);
  and _84604_ (_34891_, _34890_, _34886_);
  nor _84605_ (_34892_, _10982_, _13413_);
  or _84606_ (_34893_, _34892_, _34802_);
  and _84607_ (_34894_, _34893_, _06292_);
  or _84608_ (_34895_, _34894_, _06316_);
  or _84609_ (_34897_, _34895_, _34891_);
  or _84610_ (_34898_, _34807_, _06718_);
  and _84611_ (_34899_, _34898_, _05653_);
  and _84612_ (_34900_, _34899_, _34897_);
  and _84613_ (_34901_, _34835_, _05652_);
  or _84614_ (_34902_, _34901_, _06047_);
  or _84615_ (_34903_, _34902_, _34900_);
  and _84616_ (_34904_, _15253_, _07679_);
  or _84617_ (_34905_, _34802_, _06048_);
  or _84618_ (_34906_, _34905_, _34904_);
  and _84619_ (_34907_, _34906_, _01336_);
  and _84620_ (_34908_, _34907_, _34903_);
  or _84621_ (_34909_, _34908_, _34801_);
  and _84622_ (_43490_, _34909_, _42882_);
  and _84623_ (_34910_, _01340_, \oc8051_golden_model_1.SCON [6]);
  and _84624_ (_34911_, _13413_, \oc8051_golden_model_1.SCON [6]);
  and _84625_ (_34912_, _15389_, _07679_);
  or _84626_ (_34913_, _34912_, _34911_);
  or _84627_ (_34914_, _34913_, _06020_);
  and _84628_ (_34915_, _15293_, _07679_);
  or _84629_ (_34917_, _34915_, _34911_);
  or _84630_ (_34918_, _34917_, _06954_);
  and _84631_ (_34919_, _07679_, \oc8051_golden_model_1.ACC [6]);
  or _84632_ (_34920_, _34919_, _34911_);
  and _84633_ (_34921_, _34920_, _06938_);
  and _84634_ (_34922_, _06939_, \oc8051_golden_model_1.SCON [6]);
  or _84635_ (_34923_, _34922_, _06102_);
  or _84636_ (_34924_, _34923_, _34921_);
  and _84637_ (_34925_, _34924_, _06044_);
  and _84638_ (_34926_, _34925_, _34918_);
  and _84639_ (_34928_, _13432_, \oc8051_golden_model_1.SCON [6]);
  and _84640_ (_34929_, _15280_, _08347_);
  or _84641_ (_34930_, _34929_, _34928_);
  and _84642_ (_34931_, _34930_, _06043_);
  or _84643_ (_34932_, _34931_, _06239_);
  or _84644_ (_34933_, _34932_, _34926_);
  nor _84645_ (_34934_, _07883_, _13413_);
  or _84646_ (_34935_, _34934_, _34911_);
  or _84647_ (_34936_, _34935_, _06848_);
  and _84648_ (_34937_, _34936_, _34933_);
  or _84649_ (_34939_, _34937_, _06219_);
  or _84650_ (_34940_, _34920_, _06220_);
  and _84651_ (_34941_, _34940_, _06040_);
  and _84652_ (_34942_, _34941_, _34939_);
  and _84653_ (_34943_, _15278_, _08347_);
  or _84654_ (_34944_, _34943_, _34928_);
  and _84655_ (_34945_, _34944_, _06039_);
  or _84656_ (_34946_, _34945_, _06032_);
  or _84657_ (_34947_, _34946_, _34942_);
  or _84658_ (_34948_, _34928_, _15310_);
  and _84659_ (_34950_, _34948_, _34930_);
  or _84660_ (_34951_, _34950_, _06033_);
  and _84661_ (_34952_, _34951_, _06027_);
  and _84662_ (_34953_, _34952_, _34947_);
  or _84663_ (_34954_, _34928_, _15326_);
  and _84664_ (_34955_, _34954_, _06026_);
  and _84665_ (_34956_, _34955_, _34930_);
  or _84666_ (_34957_, _34956_, _09818_);
  or _84667_ (_34958_, _34957_, _34953_);
  and _84668_ (_34959_, _09178_, _07679_);
  or _84669_ (_34961_, _34911_, _07012_);
  or _84670_ (_34962_, _34961_, _34959_);
  or _84671_ (_34963_, _34935_, _09827_);
  and _84672_ (_34964_, _34963_, _05669_);
  and _84673_ (_34965_, _34964_, _34962_);
  and _84674_ (_34966_, _34965_, _34958_);
  and _84675_ (_34967_, _15382_, _07679_);
  or _84676_ (_34968_, _34967_, _34911_);
  and _84677_ (_34969_, _34968_, _09833_);
  or _84678_ (_34970_, _34969_, _06019_);
  or _84679_ (_34972_, _34970_, _34966_);
  and _84680_ (_34973_, _34972_, _34914_);
  or _84681_ (_34974_, _34973_, _06112_);
  and _84682_ (_34975_, _15399_, _07679_);
  or _84683_ (_34976_, _34975_, _34911_);
  or _84684_ (_34977_, _34976_, _08751_);
  and _84685_ (_34978_, _34977_, _08756_);
  and _84686_ (_34979_, _34978_, _34974_);
  and _84687_ (_34980_, _10980_, _07679_);
  or _84688_ (_34981_, _34980_, _34911_);
  and _84689_ (_34983_, _34981_, _06284_);
  or _84690_ (_34984_, _34983_, _34979_);
  and _84691_ (_34985_, _34984_, _07032_);
  or _84692_ (_34986_, _34911_, _07886_);
  and _84693_ (_34987_, _34913_, _06108_);
  and _84694_ (_34988_, _34987_, _34986_);
  or _84695_ (_34989_, _34988_, _34985_);
  and _84696_ (_34990_, _34989_, _06278_);
  and _84697_ (_34991_, _34920_, _06277_);
  and _84698_ (_34992_, _34991_, _34986_);
  or _84699_ (_34994_, _34992_, _06130_);
  or _84700_ (_34995_, _34994_, _34990_);
  and _84701_ (_34996_, _15396_, _07679_);
  or _84702_ (_34997_, _34911_, _08777_);
  or _84703_ (_34998_, _34997_, _34996_);
  and _84704_ (_34999_, _34998_, _08782_);
  and _84705_ (_35000_, _34999_, _34995_);
  nor _84706_ (_35001_, _10979_, _13413_);
  or _84707_ (_35002_, _35001_, _34911_);
  and _84708_ (_35003_, _35002_, _06292_);
  or _84709_ (_35005_, _35003_, _06316_);
  or _84710_ (_35006_, _35005_, _35000_);
  or _84711_ (_35007_, _34917_, _06718_);
  and _84712_ (_35008_, _35007_, _05653_);
  and _84713_ (_35009_, _35008_, _35006_);
  and _84714_ (_35010_, _34944_, _05652_);
  or _84715_ (_35011_, _35010_, _06047_);
  or _84716_ (_35012_, _35011_, _35009_);
  and _84717_ (_35013_, _15451_, _07679_);
  or _84718_ (_35014_, _34911_, _06048_);
  or _84719_ (_35016_, _35014_, _35013_);
  and _84720_ (_35017_, _35016_, _01336_);
  and _84721_ (_35018_, _35017_, _35012_);
  or _84722_ (_35019_, _35018_, _34910_);
  and _84723_ (_43491_, _35019_, _42882_);
  nor _84724_ (_35020_, _01336_, _06029_);
  nor _84725_ (_35021_, _07727_, _06029_);
  and _84726_ (_35022_, _07833_, \oc8051_golden_model_1.ACC [0]);
  and _84727_ (_35023_, _35022_, _08127_);
  or _84728_ (_35024_, _35023_, _35021_);
  or _84729_ (_35026_, _35024_, _06278_);
  or _84730_ (_35027_, _35021_, _07012_);
  and _84731_ (_35028_, _09120_, _07833_);
  or _84732_ (_35029_, _35028_, _35027_);
  and _84733_ (_35030_, _07727_, _06931_);
  or _84734_ (_35031_, _35021_, _09827_);
  or _84735_ (_35032_, _35031_, _35030_);
  nor _84736_ (_35033_, _08127_, _13575_);
  or _84737_ (_35034_, _35033_, _35021_);
  or _84738_ (_35035_, _35034_, _06954_);
  nor _84739_ (_35037_, _35022_, _35021_);
  nor _84740_ (_35038_, _35037_, _06939_);
  nor _84741_ (_35039_, _06938_, _06029_);
  or _84742_ (_35040_, _35039_, _06102_);
  or _84743_ (_35041_, _35040_, _35038_);
  and _84744_ (_35042_, _35041_, _06848_);
  nand _84745_ (_35043_, _35042_, _35035_);
  and _84746_ (_35044_, _35043_, _06544_);
  and _84747_ (_35045_, _35037_, _06219_);
  or _84748_ (_35046_, _35045_, _06038_);
  or _84749_ (_35048_, _35046_, _35044_);
  and _84750_ (_35049_, _07012_, _06982_);
  and _84751_ (_35050_, _35049_, _09827_);
  nand _84752_ (_35051_, _35050_, _35048_);
  and _84753_ (_35052_, _35051_, _35032_);
  and _84754_ (_35053_, _35052_, _35029_);
  or _84755_ (_35054_, _35053_, _09833_);
  and _84756_ (_35055_, _14186_, _07727_);
  or _84757_ (_35056_, _35021_, _05669_);
  or _84758_ (_35057_, _35056_, _35055_);
  and _84759_ (_35059_, _35057_, _06020_);
  and _84760_ (_35060_, _35059_, _35054_);
  and _84761_ (_35061_, _07833_, _08672_);
  or _84762_ (_35062_, _35061_, _35021_);
  and _84763_ (_35063_, _35062_, _06019_);
  or _84764_ (_35064_, _35063_, _06112_);
  or _84765_ (_35065_, _35064_, _35060_);
  and _84766_ (_35066_, _14086_, _07833_);
  or _84767_ (_35067_, _35066_, _35021_);
  or _84768_ (_35068_, _35067_, _08751_);
  and _84769_ (_35070_, _35068_, _08756_);
  and _84770_ (_35071_, _35070_, _35065_);
  nor _84771_ (_35072_, _12302_, _13575_);
  or _84772_ (_35073_, _35072_, _35021_);
  nor _84773_ (_35074_, _35023_, _08756_);
  and _84774_ (_35075_, _35074_, _35073_);
  or _84775_ (_35076_, _35075_, _35071_);
  and _84776_ (_35077_, _35076_, _07032_);
  nand _84777_ (_35078_, _35062_, _06108_);
  nor _84778_ (_35079_, _35078_, _35033_);
  or _84779_ (_35081_, _35079_, _06277_);
  or _84780_ (_35082_, _35081_, _35077_);
  and _84781_ (_35083_, _35082_, _35026_);
  or _84782_ (_35084_, _35083_, _06130_);
  and _84783_ (_35085_, _14083_, _07727_);
  or _84784_ (_35086_, _35021_, _08777_);
  or _84785_ (_35087_, _35086_, _35085_);
  and _84786_ (_35088_, _35087_, _08782_);
  and _84787_ (_35089_, _35088_, _35084_);
  and _84788_ (_35090_, _35073_, _06292_);
  or _84789_ (_35092_, _35090_, _19256_);
  or _84790_ (_35093_, _35092_, _35089_);
  or _84791_ (_35094_, _35034_, _06408_);
  and _84792_ (_35095_, _35094_, _01336_);
  and _84793_ (_35096_, _35095_, _35093_);
  or _84794_ (_35097_, _35096_, _35020_);
  and _84795_ (_43493_, _35097_, _42882_);
  nand _84796_ (_35098_, _06298_, \oc8051_golden_model_1.SP [1]);
  nand _84797_ (_35099_, _07727_, _06832_);
  or _84798_ (_35100_, _35099_, _08078_);
  or _84799_ (_35102_, _07727_, \oc8051_golden_model_1.SP [1]);
  and _84800_ (_35103_, _35102_, _06130_);
  and _84801_ (_35104_, _35103_, _35100_);
  and _84802_ (_35105_, _35102_, _09833_);
  or _84803_ (_35106_, _14367_, _13575_);
  and _84804_ (_35107_, _35106_, _35105_);
  and _84805_ (_35108_, _14284_, _07727_);
  not _84806_ (_35109_, _35108_);
  and _84807_ (_35110_, _35109_, _35102_);
  or _84808_ (_35111_, _35110_, _06954_);
  nand _84809_ (_35113_, _06943_, \oc8051_golden_model_1.SP [1]);
  nor _84810_ (_35114_, _07727_, _06847_);
  and _84811_ (_35115_, _07833_, \oc8051_golden_model_1.ACC [1]);
  or _84812_ (_35116_, _35115_, _35114_);
  and _84813_ (_35117_, _35116_, _06938_);
  nor _84814_ (_35118_, _06938_, _06847_);
  or _84815_ (_35119_, _35118_, _06943_);
  or _84816_ (_35120_, _35119_, _35117_);
  and _84817_ (_35121_, _35120_, _35113_);
  or _84818_ (_35122_, _35121_, _06102_);
  and _84819_ (_35124_, _35122_, _05690_);
  and _84820_ (_35125_, _35124_, _35111_);
  nor _84821_ (_35126_, _05690_, \oc8051_golden_model_1.SP [1]);
  or _84822_ (_35127_, _35126_, _06239_);
  or _84823_ (_35128_, _35127_, _35125_);
  nand _84824_ (_35129_, _07083_, _06239_);
  and _84825_ (_35130_, _35129_, _35128_);
  or _84826_ (_35131_, _35130_, _06219_);
  or _84827_ (_35132_, _35116_, _06220_);
  and _84828_ (_35133_, _35132_, _07364_);
  and _84829_ (_35135_, _35133_, _35131_);
  or _84830_ (_35136_, _13568_, _07169_);
  or _84831_ (_35137_, _35136_, _35135_);
  or _84832_ (_35138_, _07271_, _06847_);
  and _84833_ (_35139_, _35138_, _09827_);
  and _84834_ (_35140_, _35139_, _35137_);
  nand _84835_ (_35141_, _07727_, _07132_);
  and _84836_ (_35142_, _35102_, _09815_);
  and _84837_ (_35143_, _35142_, _35141_);
  or _84838_ (_35144_, _35143_, _07011_);
  or _84839_ (_35146_, _35144_, _35140_);
  or _84840_ (_35147_, _35114_, _07012_);
  and _84841_ (_35148_, _09075_, _07833_);
  or _84842_ (_35149_, _35148_, _35147_);
  and _84843_ (_35150_, _35149_, _05669_);
  and _84844_ (_35151_, _35150_, _35146_);
  or _84845_ (_35152_, _35151_, _35107_);
  and _84846_ (_35153_, _35152_, _06020_);
  and _84847_ (_35154_, _35102_, _06019_);
  and _84848_ (_35155_, _35154_, _35099_);
  or _84849_ (_35157_, _35155_, _05724_);
  or _84850_ (_35158_, _35157_, _35153_);
  and _84851_ (_35159_, _05724_, \oc8051_golden_model_1.SP [1]);
  nor _84852_ (_35160_, _35159_, _06112_);
  and _84853_ (_35161_, _35160_, _35158_);
  or _84854_ (_35162_, _14263_, _13575_);
  and _84855_ (_35163_, _35102_, _06112_);
  and _84856_ (_35164_, _35163_, _35162_);
  or _84857_ (_35165_, _35164_, _06284_);
  or _84858_ (_35166_, _35165_, _35161_);
  and _84859_ (_35168_, _10994_, _07833_);
  or _84860_ (_35169_, _35168_, _35114_);
  or _84861_ (_35170_, _35169_, _08756_);
  and _84862_ (_35171_, _35170_, _07032_);
  and _84863_ (_35172_, _35171_, _35166_);
  or _84864_ (_35173_, _14261_, _13575_);
  and _84865_ (_35174_, _35102_, _06108_);
  and _84866_ (_35175_, _35174_, _35173_);
  or _84867_ (_35176_, _35175_, _06277_);
  or _84868_ (_35177_, _35176_, _35172_);
  and _84869_ (_35179_, _35115_, _08078_);
  or _84870_ (_35180_, _35179_, _35114_);
  or _84871_ (_35181_, _35180_, _06278_);
  and _84872_ (_35182_, _35181_, _35177_);
  or _84873_ (_35183_, _35182_, _05736_);
  and _84874_ (_35184_, _05736_, \oc8051_golden_model_1.SP [1]);
  nor _84875_ (_35185_, _35184_, _06130_);
  and _84876_ (_35186_, _35185_, _35183_);
  or _84877_ (_35187_, _35186_, _35104_);
  and _84878_ (_35188_, _35187_, _08782_);
  nor _84879_ (_35190_, _10993_, _13575_);
  or _84880_ (_35191_, _35190_, _35114_);
  and _84881_ (_35192_, _35191_, _06292_);
  or _84882_ (_35193_, _35192_, _06298_);
  or _84883_ (_35194_, _35193_, _35188_);
  nand _84884_ (_35195_, _35194_, _35098_);
  nor _84885_ (_35196_, _06049_, _05732_);
  nand _84886_ (_35197_, _35196_, _35195_);
  or _84887_ (_35198_, _35196_, _06847_);
  and _84888_ (_35199_, _35198_, _06718_);
  and _84889_ (_35201_, _35199_, _35197_);
  and _84890_ (_35202_, _35110_, _06316_);
  or _84891_ (_35203_, _35202_, _07458_);
  or _84892_ (_35204_, _35203_, _35201_);
  or _84893_ (_35205_, _07059_, _06847_);
  and _84894_ (_35206_, _35205_, _06048_);
  and _84895_ (_35207_, _35206_, _35204_);
  or _84896_ (_35208_, _35108_, _35114_);
  and _84897_ (_35209_, _35208_, _06047_);
  or _84898_ (_35210_, _35209_, _01340_);
  or _84899_ (_35212_, _35210_, _35207_);
  or _84900_ (_35213_, _01336_, \oc8051_golden_model_1.SP [1]);
  and _84901_ (_35214_, _35213_, _42882_);
  and _84902_ (_43494_, _35214_, _35212_);
  nor _84903_ (_35215_, _01336_, _06447_);
  nand _84904_ (_35216_, _14449_, _05724_);
  nor _84905_ (_35217_, _13575_, _07530_);
  nor _84906_ (_35218_, _07727_, _06447_);
  or _84907_ (_35219_, _35218_, _09827_);
  or _84908_ (_35220_, _35219_, _35217_);
  and _84909_ (_35222_, _14493_, _07727_);
  or _84910_ (_35223_, _35222_, _35218_);
  or _84911_ (_35224_, _35223_, _06954_);
  and _84912_ (_35225_, _07833_, \oc8051_golden_model_1.ACC [2]);
  or _84913_ (_35226_, _35225_, _35218_);
  or _84914_ (_35227_, _35226_, _06939_);
  or _84915_ (_35228_, _06938_, \oc8051_golden_model_1.SP [2]);
  and _84916_ (_35229_, _35228_, _07233_);
  and _84917_ (_35230_, _35229_, _35227_);
  and _84918_ (_35231_, _07622_, _06943_);
  or _84919_ (_35233_, _35231_, _06102_);
  or _84920_ (_35234_, _35233_, _35230_);
  and _84921_ (_35235_, _35234_, _05690_);
  and _84922_ (_35236_, _35235_, _35224_);
  nor _84923_ (_35237_, _14449_, _05690_);
  or _84924_ (_35238_, _35237_, _06239_);
  or _84925_ (_35239_, _35238_, _35236_);
  nand _84926_ (_35240_, _08415_, _06239_);
  and _84927_ (_35241_, _35240_, _35239_);
  or _84928_ (_35242_, _35241_, _06219_);
  or _84929_ (_35244_, _35226_, _06220_);
  and _84930_ (_35245_, _35244_, _07364_);
  and _84931_ (_35246_, _35245_, _35242_);
  or _84932_ (_35247_, _07561_, _07355_);
  or _84933_ (_35248_, _35247_, _35246_);
  or _84934_ (_35249_, _07622_, _05686_);
  and _84935_ (_35250_, _35249_, _05673_);
  and _84936_ (_35251_, _35250_, _35248_);
  nor _84937_ (_35252_, _14449_, _05673_);
  or _84938_ (_35253_, _35252_, _09815_);
  or _84939_ (_35255_, _35253_, _35251_);
  and _84940_ (_35256_, _35255_, _35220_);
  or _84941_ (_35257_, _35256_, _07011_);
  or _84942_ (_35258_, _35218_, _07012_);
  and _84943_ (_35259_, _09182_, _07833_);
  or _84944_ (_35260_, _35259_, _35258_);
  and _84945_ (_35261_, _35260_, _05669_);
  and _84946_ (_35262_, _35261_, _35257_);
  and _84947_ (_35263_, _14580_, _07833_);
  or _84948_ (_35264_, _35263_, _35218_);
  and _84949_ (_35266_, _35264_, _09833_);
  or _84950_ (_35267_, _35266_, _06019_);
  or _84951_ (_35268_, _35267_, _35262_);
  and _84952_ (_35269_, _07833_, _08730_);
  or _84953_ (_35270_, _35269_, _35218_);
  or _84954_ (_35271_, _35270_, _06020_);
  and _84955_ (_35272_, _35271_, _35268_);
  or _84956_ (_35273_, _35272_, _05724_);
  and _84957_ (_35274_, _35273_, _35216_);
  or _84958_ (_35275_, _35274_, _06112_);
  and _84959_ (_35277_, _14596_, _07833_);
  or _84960_ (_35278_, _35277_, _35218_);
  or _84961_ (_35279_, _35278_, _08751_);
  and _84962_ (_35280_, _35279_, _08756_);
  and _84963_ (_35281_, _35280_, _35275_);
  and _84964_ (_35282_, _10991_, _07833_);
  or _84965_ (_35283_, _35282_, _35218_);
  and _84966_ (_35284_, _35283_, _06284_);
  or _84967_ (_35285_, _35284_, _35281_);
  and _84968_ (_35286_, _35285_, _07032_);
  or _84969_ (_35288_, _35218_, _08177_);
  and _84970_ (_35289_, _35270_, _06108_);
  and _84971_ (_35290_, _35289_, _35288_);
  or _84972_ (_35291_, _35290_, _35286_);
  and _84973_ (_35292_, _35291_, _12494_);
  and _84974_ (_35293_, _35226_, _06277_);
  and _84975_ (_35294_, _35293_, _35288_);
  and _84976_ (_35295_, _07622_, _05736_);
  or _84977_ (_35296_, _35295_, _06130_);
  or _84978_ (_35297_, _35296_, _35294_);
  or _84979_ (_35299_, _35297_, _35292_);
  and _84980_ (_35300_, _14593_, _07727_);
  or _84981_ (_35301_, _35218_, _08777_);
  or _84982_ (_35302_, _35301_, _35300_);
  and _84983_ (_35303_, _35302_, _35299_);
  or _84984_ (_35304_, _35303_, _06292_);
  nor _84985_ (_35305_, _10990_, _13575_);
  or _84986_ (_35306_, _35305_, _35218_);
  or _84987_ (_35307_, _35306_, _08782_);
  and _84988_ (_35308_, _35307_, _13619_);
  and _84989_ (_35310_, _35308_, _35304_);
  and _84990_ (_35311_, _14449_, _06298_);
  or _84991_ (_35312_, _35311_, _05732_);
  or _84992_ (_35313_, _35312_, _35310_);
  nand _84993_ (_35314_, _14449_, _05732_);
  and _84994_ (_35315_, _35314_, _06050_);
  and _84995_ (_35316_, _35315_, _35313_);
  and _84996_ (_35317_, _14449_, _06049_);
  or _84997_ (_35318_, _35317_, _06316_);
  or _84998_ (_35319_, _35318_, _35316_);
  or _84999_ (_35321_, _35223_, _06718_);
  and _85000_ (_35322_, _35321_, _07059_);
  and _85001_ (_35323_, _35322_, _35319_);
  nor _85002_ (_35324_, _14449_, _07059_);
  or _85003_ (_35325_, _35324_, _06047_);
  or _85004_ (_35326_, _35325_, _35323_);
  and _85005_ (_35327_, _14657_, _07727_);
  or _85006_ (_35328_, _35218_, _06048_);
  or _85007_ (_35329_, _35328_, _35327_);
  and _85008_ (_35330_, _35329_, _01336_);
  and _85009_ (_35332_, _35330_, _35326_);
  or _85010_ (_35333_, _35332_, _35215_);
  and _85011_ (_43495_, _35333_, _42882_);
  nor _85012_ (_35334_, _01336_, _06238_);
  or _85013_ (_35335_, _07625_, _07059_);
  nand _85014_ (_35336_, _14453_, _05724_);
  nor _85015_ (_35337_, _13575_, _07353_);
  nor _85016_ (_35338_, _07727_, _06238_);
  or _85017_ (_35339_, _35338_, _07011_);
  or _85018_ (_35340_, _35339_, _35337_);
  and _85019_ (_35342_, _35340_, _09818_);
  and _85020_ (_35343_, _14672_, _07727_);
  or _85021_ (_35344_, _35343_, _35338_);
  or _85022_ (_35345_, _35344_, _06954_);
  and _85023_ (_35346_, _07833_, \oc8051_golden_model_1.ACC [3]);
  or _85024_ (_35347_, _35346_, _35338_);
  or _85025_ (_35348_, _35347_, _06939_);
  or _85026_ (_35349_, _06938_, \oc8051_golden_model_1.SP [3]);
  and _85027_ (_35350_, _35349_, _07233_);
  and _85028_ (_35351_, _35350_, _35348_);
  and _85029_ (_35353_, _07625_, _06943_);
  or _85030_ (_35354_, _35353_, _06102_);
  or _85031_ (_35355_, _35354_, _35351_);
  and _85032_ (_35356_, _35355_, _05690_);
  and _85033_ (_35357_, _35356_, _35345_);
  nor _85034_ (_35358_, _14453_, _05690_);
  or _85035_ (_35359_, _35358_, _06239_);
  or _85036_ (_35360_, _35359_, _35357_);
  nand _85037_ (_35361_, _08405_, _06239_);
  and _85038_ (_35362_, _35361_, _35360_);
  or _85039_ (_35364_, _35362_, _06219_);
  or _85040_ (_35365_, _35347_, _06220_);
  and _85041_ (_35366_, _35365_, _07364_);
  and _85042_ (_35367_, _35366_, _35364_);
  or _85043_ (_35368_, _07404_, _13568_);
  or _85044_ (_35369_, _35368_, _35367_);
  or _85045_ (_35370_, _07625_, _07271_);
  and _85046_ (_35371_, _35370_, _09827_);
  and _85047_ (_35372_, _35371_, _35369_);
  or _85048_ (_35373_, _35372_, _35342_);
  or _85049_ (_35375_, _35338_, _07012_);
  and _85050_ (_35376_, _09181_, _07833_);
  or _85051_ (_35377_, _35376_, _35375_);
  and _85052_ (_35378_, _35377_, _05669_);
  and _85053_ (_35379_, _35378_, _35373_);
  and _85054_ (_35380_, _14778_, _07833_);
  or _85055_ (_35381_, _35380_, _35338_);
  and _85056_ (_35382_, _35381_, _09833_);
  or _85057_ (_35383_, _35382_, _06019_);
  or _85058_ (_35384_, _35383_, _35379_);
  and _85059_ (_35386_, _07833_, _08662_);
  or _85060_ (_35387_, _35386_, _35338_);
  or _85061_ (_35388_, _35387_, _06020_);
  and _85062_ (_35389_, _35388_, _35384_);
  or _85063_ (_35390_, _35389_, _05724_);
  and _85064_ (_35391_, _35390_, _35336_);
  or _85065_ (_35392_, _35391_, _06112_);
  and _85066_ (_35393_, _14793_, _07833_);
  or _85067_ (_35394_, _35393_, _35338_);
  or _85068_ (_35395_, _35394_, _08751_);
  and _85069_ (_35397_, _35395_, _08756_);
  and _85070_ (_35398_, _35397_, _35392_);
  and _85071_ (_35399_, _12299_, _07833_);
  or _85072_ (_35400_, _35399_, _35338_);
  and _85073_ (_35401_, _35400_, _06284_);
  or _85074_ (_35402_, _35401_, _35398_);
  and _85075_ (_35403_, _35402_, _07032_);
  or _85076_ (_35404_, _35338_, _08029_);
  and _85077_ (_35405_, _35387_, _06108_);
  and _85078_ (_35406_, _35405_, _35404_);
  or _85079_ (_35408_, _35406_, _35403_);
  and _85080_ (_35409_, _35408_, _12494_);
  and _85081_ (_35410_, _35347_, _06277_);
  and _85082_ (_35411_, _35410_, _35404_);
  and _85083_ (_35412_, _07625_, _05736_);
  or _85084_ (_35413_, _35412_, _06130_);
  or _85085_ (_35414_, _35413_, _35411_);
  or _85086_ (_35415_, _35414_, _35409_);
  and _85087_ (_35416_, _14792_, _07727_);
  or _85088_ (_35417_, _35338_, _08777_);
  or _85089_ (_35419_, _35417_, _35416_);
  and _85090_ (_35420_, _35419_, _35415_);
  or _85091_ (_35421_, _35420_, _06292_);
  nor _85092_ (_35422_, _10988_, _13575_);
  or _85093_ (_35423_, _35422_, _35338_);
  or _85094_ (_35424_, _35423_, _08782_);
  and _85095_ (_35425_, _35424_, _13619_);
  and _85096_ (_35426_, _35425_, _35421_);
  nor _85097_ (_35427_, _08402_, _06238_);
  or _85098_ (_35428_, _35427_, _08403_);
  and _85099_ (_35430_, _35428_, _06298_);
  or _85100_ (_35431_, _35430_, _05732_);
  or _85101_ (_35432_, _35431_, _35426_);
  nand _85102_ (_35433_, _14453_, _05732_);
  and _85103_ (_35434_, _35433_, _35432_);
  or _85104_ (_35435_, _35434_, _06049_);
  or _85105_ (_35436_, _35428_, _06050_);
  and _85106_ (_35437_, _35436_, _06718_);
  and _85107_ (_35438_, _35437_, _35435_);
  and _85108_ (_35439_, _35344_, _06316_);
  or _85109_ (_35441_, _35439_, _07458_);
  or _85110_ (_35442_, _35441_, _35438_);
  and _85111_ (_35443_, _35442_, _35335_);
  or _85112_ (_35444_, _35443_, _06047_);
  and _85113_ (_35445_, _14849_, _07727_);
  or _85114_ (_35446_, _35338_, _06048_);
  or _85115_ (_35447_, _35446_, _35445_);
  and _85116_ (_35448_, _35447_, _01336_);
  and _85117_ (_35449_, _35448_, _35444_);
  or _85118_ (_35450_, _35449_, _35334_);
  and _85119_ (_43496_, _35450_, _42882_);
  nor _85120_ (_35452_, _01336_, _13552_);
  nor _85121_ (_35453_, _07360_, \oc8051_golden_model_1.SP [4]);
  nor _85122_ (_35454_, _35453_, _13516_);
  or _85123_ (_35455_, _35454_, _07059_);
  or _85124_ (_35456_, _35454_, _05734_);
  or _85125_ (_35457_, _35454_, _07271_);
  nor _85126_ (_35458_, _07727_, _13552_);
  and _85127_ (_35459_, _14887_, _07727_);
  or _85128_ (_35460_, _35459_, _35458_);
  or _85129_ (_35462_, _35460_, _06954_);
  and _85130_ (_35463_, _07833_, \oc8051_golden_model_1.ACC [4]);
  or _85131_ (_35464_, _35463_, _35458_);
  or _85132_ (_35465_, _35464_, _06939_);
  or _85133_ (_35466_, _06938_, \oc8051_golden_model_1.SP [4]);
  and _85134_ (_35467_, _35466_, _07233_);
  and _85135_ (_35468_, _35467_, _35465_);
  and _85136_ (_35469_, _35454_, _06943_);
  or _85137_ (_35470_, _35469_, _06102_);
  or _85138_ (_35471_, _35470_, _35468_);
  and _85139_ (_35473_, _35471_, _05690_);
  and _85140_ (_35474_, _35473_, _35462_);
  and _85141_ (_35475_, _35454_, _07272_);
  or _85142_ (_35476_, _35475_, _06239_);
  or _85143_ (_35477_, _35476_, _35474_);
  and _85144_ (_35478_, _13553_, _06029_);
  nor _85145_ (_35479_, _08404_, _13552_);
  nor _85146_ (_35480_, _35479_, _35478_);
  nand _85147_ (_35481_, _35480_, _06239_);
  and _85148_ (_35482_, _35481_, _35477_);
  or _85149_ (_35484_, _35482_, _06219_);
  or _85150_ (_35485_, _35464_, _06220_);
  and _85151_ (_35486_, _35485_, _07364_);
  and _85152_ (_35487_, _35486_, _35484_);
  and _85153_ (_35488_, _07361_, \oc8051_golden_model_1.SP [4]);
  nor _85154_ (_35489_, _07361_, \oc8051_golden_model_1.SP [4]);
  nor _85155_ (_35490_, _35489_, _35488_);
  nand _85156_ (_35491_, _35490_, _06038_);
  nand _85157_ (_35492_, _35491_, _07271_);
  or _85158_ (_35493_, _35492_, _35487_);
  and _85159_ (_35495_, _35493_, _35457_);
  nor _85160_ (_35496_, _11995_, _05660_);
  and _85161_ (_35497_, _06227_, _05659_);
  and _85162_ (_35498_, _06133_, _05659_);
  nor _85163_ (_35499_, _35498_, _35497_);
  not _85164_ (_35500_, _35499_);
  or _85165_ (_35501_, _35500_, _35496_);
  or _85166_ (_35502_, _35501_, _35495_);
  and _85167_ (_35503_, _06096_, _05659_);
  not _85168_ (_35504_, _35501_);
  nor _85169_ (_35506_, _08270_, _13575_);
  or _85170_ (_35507_, _35506_, _35458_);
  nor _85171_ (_35508_, _35507_, _35504_);
  nor _85172_ (_35509_, _35508_, _35503_);
  and _85173_ (_35510_, _35509_, _35502_);
  and _85174_ (_35511_, _35507_, _35503_);
  or _85175_ (_35512_, _35511_, _07011_);
  or _85176_ (_35513_, _35512_, _35510_);
  or _85177_ (_35514_, _35458_, _07012_);
  and _85178_ (_35515_, _09180_, _07833_);
  or _85179_ (_35517_, _35515_, _35514_);
  and _85180_ (_35518_, _35517_, _35513_);
  or _85181_ (_35519_, _35518_, _09833_);
  and _85182_ (_35520_, _14983_, _07833_);
  or _85183_ (_35521_, _35520_, _35458_);
  or _85184_ (_35522_, _35521_, _05669_);
  and _85185_ (_35523_, _35522_, _06020_);
  and _85186_ (_35524_, _35523_, _35519_);
  and _85187_ (_35525_, _08665_, _07833_);
  or _85188_ (_35526_, _35525_, _35458_);
  and _85189_ (_35528_, _35526_, _06019_);
  or _85190_ (_35529_, _35528_, _05724_);
  or _85191_ (_35530_, _35529_, _35524_);
  or _85192_ (_35531_, _35454_, _13587_);
  and _85193_ (_35532_, _35531_, _35530_);
  or _85194_ (_35533_, _35532_, _06112_);
  and _85195_ (_35534_, _14876_, _07727_);
  or _85196_ (_35535_, _35458_, _08751_);
  or _85197_ (_35536_, _35535_, _35534_);
  and _85198_ (_35537_, _35536_, _08756_);
  and _85199_ (_35539_, _35537_, _35533_);
  and _85200_ (_35540_, _10986_, _07833_);
  or _85201_ (_35541_, _35540_, _35458_);
  and _85202_ (_35542_, _35541_, _06284_);
  or _85203_ (_35543_, _35542_, _35539_);
  and _85204_ (_35544_, _35543_, _07032_);
  or _85205_ (_35545_, _35458_, _08273_);
  and _85206_ (_35546_, _35526_, _06108_);
  and _85207_ (_35547_, _35546_, _35545_);
  or _85208_ (_35548_, _35547_, _35544_);
  and _85209_ (_35550_, _35548_, _12494_);
  and _85210_ (_35551_, _35464_, _06277_);
  and _85211_ (_35552_, _35551_, _35545_);
  and _85212_ (_35553_, _35454_, _05736_);
  or _85213_ (_35554_, _35553_, _06130_);
  or _85214_ (_35555_, _35554_, _35552_);
  or _85215_ (_35556_, _35555_, _35550_);
  and _85216_ (_35557_, _14873_, _07727_);
  or _85217_ (_35558_, _35458_, _08777_);
  or _85218_ (_35559_, _35558_, _35557_);
  and _85219_ (_35561_, _35559_, _35556_);
  or _85220_ (_35562_, _35561_, _06292_);
  nor _85221_ (_35563_, _10985_, _13575_);
  or _85222_ (_35564_, _35563_, _35458_);
  or _85223_ (_35565_, _35564_, _08782_);
  and _85224_ (_35566_, _35565_, _13619_);
  and _85225_ (_35567_, _35566_, _35562_);
  nor _85226_ (_35568_, _08403_, _13552_);
  or _85227_ (_35569_, _35568_, _13553_);
  and _85228_ (_35570_, _35569_, _06298_);
  or _85229_ (_35572_, _35570_, _05732_);
  or _85230_ (_35573_, _35572_, _35567_);
  and _85231_ (_35574_, _35573_, _35456_);
  or _85232_ (_35575_, _35574_, _06049_);
  or _85233_ (_35576_, _35569_, _06050_);
  and _85234_ (_35577_, _35576_, _06718_);
  and _85235_ (_35578_, _35577_, _35575_);
  and _85236_ (_35579_, _35460_, _06316_);
  or _85237_ (_35580_, _35579_, _07458_);
  or _85238_ (_35581_, _35580_, _35578_);
  and _85239_ (_35583_, _35581_, _35455_);
  or _85240_ (_35584_, _35583_, _06047_);
  and _85241_ (_35585_, _15055_, _07727_);
  or _85242_ (_35586_, _35458_, _06048_);
  or _85243_ (_35587_, _35586_, _35585_);
  and _85244_ (_35588_, _35587_, _01336_);
  and _85245_ (_35589_, _35588_, _35584_);
  or _85246_ (_35590_, _35589_, _35452_);
  and _85247_ (_43497_, _35590_, _42882_);
  nor _85248_ (_35591_, _01336_, _13551_);
  nor _85249_ (_35593_, _13516_, \oc8051_golden_model_1.SP [5]);
  nor _85250_ (_35594_, _35593_, _13517_);
  or _85251_ (_35595_, _35594_, _07059_);
  or _85252_ (_35596_, _35594_, _05734_);
  nor _85253_ (_35597_, _07977_, _13575_);
  nor _85254_ (_35598_, _07727_, _13551_);
  or _85255_ (_35599_, _35598_, _07011_);
  or _85256_ (_35600_, _35599_, _35597_);
  and _85257_ (_35601_, _35600_, _09818_);
  and _85258_ (_35602_, _15093_, _07727_);
  or _85259_ (_35604_, _35602_, _35598_);
  or _85260_ (_35605_, _35604_, _06954_);
  and _85261_ (_35606_, _07833_, \oc8051_golden_model_1.ACC [5]);
  or _85262_ (_35607_, _35606_, _35598_);
  or _85263_ (_35608_, _35607_, _06939_);
  or _85264_ (_35609_, _06938_, \oc8051_golden_model_1.SP [5]);
  and _85265_ (_35610_, _35609_, _07233_);
  and _85266_ (_35611_, _35610_, _35608_);
  and _85267_ (_35612_, _35594_, _06943_);
  or _85268_ (_35613_, _35612_, _06102_);
  or _85269_ (_35615_, _35613_, _35611_);
  and _85270_ (_35616_, _35615_, _05690_);
  and _85271_ (_35617_, _35616_, _35605_);
  and _85272_ (_35618_, _35594_, _07272_);
  or _85273_ (_35619_, _35618_, _06239_);
  or _85274_ (_35620_, _35619_, _35617_);
  and _85275_ (_35621_, _13554_, _06029_);
  nor _85276_ (_35622_, _35478_, _13551_);
  nor _85277_ (_35623_, _35622_, _35621_);
  nand _85278_ (_35624_, _35623_, _06239_);
  and _85279_ (_35626_, _35624_, _35620_);
  or _85280_ (_35627_, _35626_, _06219_);
  or _85281_ (_35628_, _35607_, _06220_);
  and _85282_ (_35629_, _35628_, _07364_);
  and _85283_ (_35630_, _35629_, _35627_);
  nor _85284_ (_35631_, _35488_, \oc8051_golden_model_1.SP [5]);
  nor _85285_ (_35632_, _35631_, _13527_);
  nand _85286_ (_35633_, _35632_, _06038_);
  nand _85287_ (_35634_, _35633_, _07271_);
  or _85288_ (_35635_, _35634_, _35630_);
  or _85289_ (_35636_, _35594_, _07271_);
  and _85290_ (_35637_, _35636_, _09827_);
  and _85291_ (_35638_, _35637_, _35635_);
  or _85292_ (_35639_, _35638_, _35601_);
  or _85293_ (_35640_, _35598_, _07012_);
  and _85294_ (_35641_, _09179_, _07833_);
  or _85295_ (_35642_, _35641_, _35640_);
  and _85296_ (_35643_, _35642_, _05669_);
  and _85297_ (_35644_, _35643_, _35639_);
  and _85298_ (_35645_, _15179_, _07833_);
  or _85299_ (_35647_, _35645_, _35598_);
  and _85300_ (_35648_, _35647_, _09833_);
  or _85301_ (_35649_, _35648_, _06019_);
  or _85302_ (_35650_, _35649_, _35644_);
  and _85303_ (_35651_, _08652_, _07833_);
  or _85304_ (_35652_, _35651_, _35598_);
  or _85305_ (_35653_, _35652_, _06020_);
  and _85306_ (_35654_, _35653_, _35650_);
  or _85307_ (_35655_, _35654_, _05724_);
  or _85308_ (_35656_, _35594_, _13587_);
  and _85309_ (_35658_, _35656_, _35655_);
  or _85310_ (_35659_, _35658_, _06112_);
  and _85311_ (_35660_, _15195_, _07727_);
  or _85312_ (_35661_, _35598_, _08751_);
  or _85313_ (_35662_, _35661_, _35660_);
  and _85314_ (_35663_, _35662_, _08756_);
  and _85315_ (_35664_, _35663_, _35659_);
  and _85316_ (_35665_, _12306_, _07833_);
  or _85317_ (_35666_, _35665_, _35598_);
  and _85318_ (_35667_, _35666_, _06284_);
  or _85319_ (_35669_, _35667_, _35664_);
  and _85320_ (_35670_, _35669_, _07032_);
  or _85321_ (_35671_, _35598_, _07980_);
  and _85322_ (_35672_, _35652_, _06108_);
  and _85323_ (_35673_, _35672_, _35671_);
  or _85324_ (_35674_, _35673_, _35670_);
  and _85325_ (_35675_, _35674_, _12494_);
  and _85326_ (_35676_, _35607_, _06277_);
  and _85327_ (_35677_, _35676_, _35671_);
  and _85328_ (_35678_, _35594_, _05736_);
  or _85329_ (_35680_, _35678_, _06130_);
  or _85330_ (_35681_, _35680_, _35677_);
  or _85331_ (_35682_, _35681_, _35675_);
  and _85332_ (_35683_, _15194_, _07727_);
  or _85333_ (_35684_, _35598_, _08777_);
  or _85334_ (_35685_, _35684_, _35683_);
  and _85335_ (_35686_, _35685_, _35682_);
  or _85336_ (_35687_, _35686_, _06292_);
  nor _85337_ (_35688_, _10982_, _13575_);
  or _85338_ (_35689_, _35688_, _35598_);
  or _85339_ (_35691_, _35689_, _08782_);
  and _85340_ (_35692_, _35691_, _13619_);
  and _85341_ (_35693_, _35692_, _35687_);
  nor _85342_ (_35694_, _13553_, _13551_);
  or _85343_ (_35695_, _35694_, _13554_);
  and _85344_ (_35696_, _35695_, _06298_);
  or _85345_ (_35697_, _35696_, _05732_);
  or _85346_ (_35698_, _35697_, _35693_);
  and _85347_ (_35699_, _35698_, _35596_);
  or _85348_ (_35700_, _35699_, _06049_);
  or _85349_ (_35702_, _35695_, _06050_);
  and _85350_ (_35703_, _35702_, _06718_);
  and _85351_ (_35704_, _35703_, _35700_);
  and _85352_ (_35705_, _35604_, _06316_);
  or _85353_ (_35706_, _35705_, _07458_);
  or _85354_ (_35707_, _35706_, _35704_);
  and _85355_ (_35708_, _35707_, _35595_);
  or _85356_ (_35709_, _35708_, _06047_);
  and _85357_ (_35710_, _15253_, _07727_);
  or _85358_ (_35711_, _35598_, _06048_);
  or _85359_ (_35713_, _35711_, _35710_);
  and _85360_ (_35714_, _35713_, _01336_);
  and _85361_ (_35715_, _35714_, _35709_);
  or _85362_ (_35716_, _35715_, _35591_);
  and _85363_ (_43498_, _35716_, _42882_);
  nor _85364_ (_35717_, _01336_, _13550_);
  nor _85365_ (_35718_, _07883_, _13575_);
  nor _85366_ (_35719_, _07727_, _13550_);
  or _85367_ (_35720_, _35719_, _09827_);
  or _85368_ (_35721_, _35720_, _35718_);
  and _85369_ (_35723_, _15293_, _07727_);
  or _85370_ (_35724_, _35723_, _35719_);
  or _85371_ (_35725_, _35724_, _06954_);
  and _85372_ (_35726_, _07833_, \oc8051_golden_model_1.ACC [6]);
  or _85373_ (_35727_, _35726_, _35719_);
  or _85374_ (_35728_, _35727_, _06939_);
  or _85375_ (_35729_, _06938_, \oc8051_golden_model_1.SP [6]);
  and _85376_ (_35730_, _35729_, _07233_);
  and _85377_ (_35731_, _35730_, _35728_);
  nor _85378_ (_35732_, _13517_, \oc8051_golden_model_1.SP [6]);
  nor _85379_ (_35734_, _35732_, _13518_);
  and _85380_ (_35735_, _35734_, _06943_);
  or _85381_ (_35736_, _35735_, _06102_);
  or _85382_ (_35737_, _35736_, _35731_);
  and _85383_ (_35738_, _35737_, _05690_);
  and _85384_ (_35739_, _35738_, _35725_);
  and _85385_ (_35740_, _35734_, _07272_);
  or _85386_ (_35741_, _35740_, _06239_);
  or _85387_ (_35742_, _35741_, _35739_);
  nor _85388_ (_35743_, _35621_, _13550_);
  nor _85389_ (_35745_, _35743_, _13556_);
  nand _85390_ (_35746_, _35745_, _06239_);
  and _85391_ (_35747_, _35746_, _35742_);
  or _85392_ (_35748_, _35747_, _06219_);
  or _85393_ (_35749_, _35727_, _06220_);
  and _85394_ (_35750_, _35749_, _07364_);
  and _85395_ (_35751_, _35750_, _35748_);
  nor _85396_ (_35752_, _13527_, \oc8051_golden_model_1.SP [6]);
  nor _85397_ (_35753_, _35752_, _13528_);
  and _85398_ (_35754_, _35753_, _06038_);
  or _85399_ (_35756_, _35754_, _35751_);
  and _85400_ (_35757_, _35756_, _07271_);
  and _85401_ (_35758_, _35734_, _13568_);
  or _85402_ (_35759_, _35758_, _09815_);
  or _85403_ (_35760_, _35759_, _35757_);
  and _85404_ (_35761_, _35760_, _35721_);
  or _85405_ (_35762_, _35761_, _07011_);
  or _85406_ (_35763_, _35719_, _07012_);
  and _85407_ (_35764_, _09178_, _07833_);
  or _85408_ (_35765_, _35764_, _35763_);
  and _85409_ (_35767_, _35765_, _05669_);
  and _85410_ (_35768_, _35767_, _35762_);
  and _85411_ (_35769_, _15382_, _07833_);
  or _85412_ (_35770_, _35769_, _35719_);
  and _85413_ (_35771_, _35770_, _09833_);
  or _85414_ (_35772_, _35771_, _06019_);
  or _85415_ (_35773_, _35772_, _35768_);
  and _85416_ (_35774_, _15389_, _07833_);
  or _85417_ (_35775_, _35774_, _35719_);
  or _85418_ (_35776_, _35775_, _06020_);
  and _85419_ (_35778_, _35776_, _35773_);
  or _85420_ (_35779_, _35778_, _05724_);
  or _85421_ (_35780_, _35734_, _13587_);
  and _85422_ (_35781_, _35780_, _35779_);
  or _85423_ (_35782_, _35781_, _06112_);
  and _85424_ (_35783_, _15399_, _07727_);
  or _85425_ (_35784_, _35719_, _08751_);
  or _85426_ (_35785_, _35784_, _35783_);
  and _85427_ (_35786_, _35785_, _08756_);
  and _85428_ (_35787_, _35786_, _35782_);
  and _85429_ (_35789_, _10980_, _07833_);
  or _85430_ (_35790_, _35789_, _35719_);
  and _85431_ (_35791_, _35790_, _06284_);
  or _85432_ (_35792_, _35791_, _35787_);
  and _85433_ (_35793_, _35792_, _07032_);
  or _85434_ (_35794_, _35719_, _07886_);
  and _85435_ (_35795_, _35775_, _06108_);
  and _85436_ (_35796_, _35795_, _35794_);
  or _85437_ (_35797_, _35796_, _35793_);
  and _85438_ (_35798_, _35797_, _12494_);
  and _85439_ (_35800_, _35727_, _06277_);
  and _85440_ (_35801_, _35800_, _35794_);
  and _85441_ (_35802_, _35734_, _05736_);
  or _85442_ (_35803_, _35802_, _06130_);
  or _85443_ (_35804_, _35803_, _35801_);
  or _85444_ (_35805_, _35804_, _35798_);
  and _85445_ (_35806_, _15396_, _07727_);
  or _85446_ (_35807_, _35719_, _08777_);
  or _85447_ (_35808_, _35807_, _35806_);
  and _85448_ (_35809_, _35808_, _35805_);
  or _85449_ (_35811_, _35809_, _06292_);
  nor _85450_ (_35812_, _10979_, _13575_);
  or _85451_ (_35813_, _35812_, _35719_);
  or _85452_ (_35814_, _35813_, _08782_);
  and _85453_ (_35815_, _35814_, _13619_);
  and _85454_ (_35816_, _35815_, _35811_);
  nor _85455_ (_35817_, _13554_, _13550_);
  or _85456_ (_35818_, _35817_, _13555_);
  and _85457_ (_35819_, _35818_, _06298_);
  or _85458_ (_35820_, _35819_, _05732_);
  or _85459_ (_35822_, _35820_, _35816_);
  or _85460_ (_35823_, _35734_, _05734_);
  and _85461_ (_35824_, _35823_, _35822_);
  or _85462_ (_35825_, _35824_, _06049_);
  or _85463_ (_35826_, _35818_, _06050_);
  and _85464_ (_35827_, _35826_, _35825_);
  or _85465_ (_35828_, _35827_, _06316_);
  or _85466_ (_35829_, _35724_, _06718_);
  and _85467_ (_35830_, _35829_, _07059_);
  and _85468_ (_35831_, _35830_, _35828_);
  and _85469_ (_35833_, _35734_, _07458_);
  or _85470_ (_35834_, _35833_, _06047_);
  or _85471_ (_35835_, _35834_, _35831_);
  and _85472_ (_35836_, _15451_, _07727_);
  or _85473_ (_35837_, _35719_, _06048_);
  or _85474_ (_35838_, _35837_, _35836_);
  and _85475_ (_35839_, _35838_, _01336_);
  and _85476_ (_35840_, _35839_, _35835_);
  or _85477_ (_35841_, _35840_, _35717_);
  and _85478_ (_43499_, _35841_, _42882_);
  not _85479_ (_35843_, \oc8051_golden_model_1.SBUF [0]);
  nor _85480_ (_35844_, _01336_, _35843_);
  nand _85481_ (_35845_, _10995_, _07681_);
  nor _85482_ (_35846_, _07681_, _35843_);
  nor _85483_ (_35847_, _35846_, _06278_);
  nand _85484_ (_35848_, _35847_, _35845_);
  and _85485_ (_35849_, _09120_, _07681_);
  or _85486_ (_35850_, _35846_, _07012_);
  or _85487_ (_35851_, _35850_, _35849_);
  and _85488_ (_35852_, _07681_, _06931_);
  nor _85489_ (_35854_, _35852_, _35846_);
  nand _85490_ (_35855_, _35854_, _09815_);
  nor _85491_ (_35856_, _08127_, _13650_);
  or _85492_ (_35857_, _35856_, _35846_);
  or _85493_ (_35858_, _35857_, _06954_);
  and _85494_ (_35859_, _07681_, \oc8051_golden_model_1.ACC [0]);
  nor _85495_ (_35860_, _35859_, _35846_);
  nor _85496_ (_35861_, _35860_, _06939_);
  nor _85497_ (_35862_, _06938_, _35843_);
  or _85498_ (_35863_, _35862_, _06102_);
  or _85499_ (_35865_, _35863_, _35861_);
  and _85500_ (_35866_, _35865_, _06848_);
  and _85501_ (_35867_, _35866_, _35858_);
  nor _85502_ (_35868_, _35854_, _06848_);
  or _85503_ (_35869_, _35868_, _35867_);
  nand _85504_ (_35870_, _35869_, _06220_);
  or _85505_ (_35871_, _35860_, _06220_);
  and _85506_ (_35872_, _35871_, _09817_);
  nand _85507_ (_35873_, _35872_, _35870_);
  and _85508_ (_35874_, _35873_, _35855_);
  and _85509_ (_35876_, _35874_, _35851_);
  or _85510_ (_35877_, _35876_, _09833_);
  and _85511_ (_35878_, _14186_, _07681_);
  or _85512_ (_35879_, _35878_, _35846_);
  or _85513_ (_35880_, _35879_, _05669_);
  and _85514_ (_35881_, _35880_, _06020_);
  and _85515_ (_35882_, _35881_, _35877_);
  and _85516_ (_35883_, _07681_, _08672_);
  or _85517_ (_35884_, _35883_, _35846_);
  and _85518_ (_35885_, _35884_, _06019_);
  or _85519_ (_35887_, _35885_, _06112_);
  or _85520_ (_35888_, _35887_, _35882_);
  and _85521_ (_35889_, _14086_, _07681_);
  or _85522_ (_35890_, _35846_, _08751_);
  or _85523_ (_35891_, _35890_, _35889_);
  and _85524_ (_35892_, _35891_, _08756_);
  and _85525_ (_35893_, _35892_, _35888_);
  nor _85526_ (_35894_, _12302_, _13650_);
  or _85527_ (_35895_, _35894_, _35846_);
  and _85528_ (_35896_, _35845_, _06284_);
  and _85529_ (_35898_, _35896_, _35895_);
  or _85530_ (_35899_, _35898_, _35893_);
  and _85531_ (_35900_, _35899_, _07032_);
  nand _85532_ (_35901_, _35884_, _06108_);
  nor _85533_ (_35902_, _35901_, _35856_);
  or _85534_ (_35903_, _35902_, _06277_);
  or _85535_ (_35904_, _35903_, _35900_);
  and _85536_ (_35905_, _35904_, _35848_);
  or _85537_ (_35906_, _35905_, _06130_);
  and _85538_ (_35907_, _14083_, _07681_);
  or _85539_ (_35909_, _35846_, _08777_);
  or _85540_ (_35910_, _35909_, _35907_);
  and _85541_ (_35911_, _35910_, _08782_);
  and _85542_ (_35912_, _35911_, _35906_);
  and _85543_ (_35913_, _35895_, _06292_);
  or _85544_ (_35914_, _35913_, _19256_);
  or _85545_ (_35915_, _35914_, _35912_);
  or _85546_ (_35916_, _35857_, _06408_);
  and _85547_ (_35917_, _35916_, _01336_);
  and _85548_ (_35918_, _35917_, _35915_);
  or _85549_ (_35920_, _35918_, _35844_);
  and _85550_ (_43501_, _35920_, _42882_);
  not _85551_ (_35921_, \oc8051_golden_model_1.SBUF [1]);
  nor _85552_ (_35922_, _01336_, _35921_);
  or _85553_ (_35923_, _14367_, _13650_);
  or _85554_ (_35924_, _07681_, \oc8051_golden_model_1.SBUF [1]);
  and _85555_ (_35925_, _35924_, _09833_);
  and _85556_ (_35926_, _35925_, _35923_);
  and _85557_ (_35927_, _09075_, _07681_);
  nor _85558_ (_35928_, _07681_, _35921_);
  or _85559_ (_35930_, _35928_, _07012_);
  or _85560_ (_35931_, _35930_, _35927_);
  and _85561_ (_35932_, _14284_, _07681_);
  not _85562_ (_35933_, _35932_);
  and _85563_ (_35934_, _35933_, _35924_);
  or _85564_ (_35935_, _35934_, _06954_);
  and _85565_ (_35936_, _07681_, \oc8051_golden_model_1.ACC [1]);
  or _85566_ (_35937_, _35936_, _35928_);
  and _85567_ (_35938_, _35937_, _06938_);
  nor _85568_ (_35939_, _06938_, _35921_);
  or _85569_ (_35941_, _35939_, _06102_);
  or _85570_ (_35942_, _35941_, _35938_);
  and _85571_ (_35943_, _35942_, _06848_);
  and _85572_ (_35944_, _35943_, _35935_);
  nor _85573_ (_35945_, _13650_, _07132_);
  or _85574_ (_35946_, _35945_, _35928_);
  and _85575_ (_35947_, _35946_, _06239_);
  or _85576_ (_35948_, _35947_, _35944_);
  and _85577_ (_35949_, _35948_, _06220_);
  and _85578_ (_35950_, _35937_, _06219_);
  or _85579_ (_35952_, _35950_, _09818_);
  or _85580_ (_35953_, _35952_, _35949_);
  or _85581_ (_35954_, _35946_, _09827_);
  and _85582_ (_35955_, _35954_, _05669_);
  and _85583_ (_35956_, _35955_, _35953_);
  and _85584_ (_35957_, _35956_, _35931_);
  or _85585_ (_35958_, _35957_, _35926_);
  and _85586_ (_35959_, _35958_, _06020_);
  nand _85587_ (_35960_, _07681_, _06832_);
  and _85588_ (_35961_, _35924_, _06019_);
  and _85589_ (_35963_, _35961_, _35960_);
  or _85590_ (_35964_, _35963_, _35959_);
  and _85591_ (_35965_, _35964_, _08751_);
  or _85592_ (_35966_, _14263_, _13650_);
  and _85593_ (_35967_, _35924_, _06112_);
  and _85594_ (_35968_, _35967_, _35966_);
  or _85595_ (_35969_, _35968_, _06284_);
  or _85596_ (_35970_, _35969_, _35965_);
  nor _85597_ (_35971_, _10993_, _13650_);
  or _85598_ (_35972_, _35971_, _35928_);
  nand _85599_ (_35974_, _10992_, _07681_);
  and _85600_ (_35975_, _35974_, _35972_);
  or _85601_ (_35976_, _35975_, _08756_);
  and _85602_ (_35977_, _35976_, _07032_);
  and _85603_ (_35978_, _35977_, _35970_);
  or _85604_ (_35979_, _14261_, _13650_);
  and _85605_ (_35980_, _35924_, _06108_);
  and _85606_ (_35981_, _35980_, _35979_);
  or _85607_ (_35982_, _35981_, _06277_);
  or _85608_ (_35983_, _35982_, _35978_);
  nor _85609_ (_35985_, _35928_, _06278_);
  nand _85610_ (_35986_, _35985_, _35974_);
  and _85611_ (_35987_, _35986_, _08777_);
  and _85612_ (_35988_, _35987_, _35983_);
  or _85613_ (_35989_, _35960_, _08078_);
  and _85614_ (_35990_, _35924_, _06130_);
  and _85615_ (_35991_, _35990_, _35989_);
  or _85616_ (_35992_, _35991_, _06292_);
  or _85617_ (_35993_, _35992_, _35988_);
  or _85618_ (_35994_, _35972_, _08782_);
  and _85619_ (_35996_, _35994_, _06718_);
  and _85620_ (_35997_, _35996_, _35993_);
  and _85621_ (_35998_, _35934_, _06316_);
  or _85622_ (_35999_, _35998_, _06047_);
  or _85623_ (_36000_, _35999_, _35997_);
  or _85624_ (_36001_, _35928_, _06048_);
  or _85625_ (_36002_, _36001_, _35932_);
  and _85626_ (_36003_, _36002_, _01336_);
  and _85627_ (_36004_, _36003_, _36000_);
  or _85628_ (_36005_, _36004_, _35922_);
  and _85629_ (_43502_, _36005_, _42882_);
  not _85630_ (_36007_, \oc8051_golden_model_1.SBUF [2]);
  nor _85631_ (_36008_, _01336_, _36007_);
  nor _85632_ (_36009_, _07681_, _36007_);
  or _85633_ (_36010_, _36009_, _08177_);
  and _85634_ (_36011_, _07681_, _08730_);
  or _85635_ (_36012_, _36011_, _36009_);
  and _85636_ (_36013_, _36012_, _06108_);
  and _85637_ (_36014_, _36013_, _36010_);
  and _85638_ (_36015_, _09182_, _07681_);
  or _85639_ (_36017_, _36009_, _07012_);
  or _85640_ (_36018_, _36017_, _36015_);
  nor _85641_ (_36019_, _13650_, _07530_);
  nor _85642_ (_36020_, _36019_, _36009_);
  nand _85643_ (_36021_, _36020_, _09815_);
  and _85644_ (_36022_, _14493_, _07681_);
  or _85645_ (_36023_, _36022_, _36009_);
  or _85646_ (_36024_, _36023_, _06954_);
  and _85647_ (_36025_, _07681_, \oc8051_golden_model_1.ACC [2]);
  nor _85648_ (_36026_, _36025_, _36009_);
  nor _85649_ (_36028_, _36026_, _06939_);
  nor _85650_ (_36029_, _06938_, _36007_);
  or _85651_ (_36030_, _36029_, _06102_);
  or _85652_ (_36031_, _36030_, _36028_);
  and _85653_ (_36032_, _36031_, _06848_);
  and _85654_ (_36033_, _36032_, _36024_);
  nor _85655_ (_36034_, _36020_, _06848_);
  or _85656_ (_36035_, _36034_, _36033_);
  nand _85657_ (_36036_, _36035_, _06220_);
  or _85658_ (_36037_, _36026_, _06220_);
  and _85659_ (_36039_, _36037_, _09817_);
  nand _85660_ (_36040_, _36039_, _36036_);
  and _85661_ (_36041_, _36040_, _36021_);
  and _85662_ (_36042_, _36041_, _36018_);
  or _85663_ (_36043_, _36042_, _09833_);
  and _85664_ (_36044_, _14580_, _07681_);
  or _85665_ (_36045_, _36044_, _36009_);
  or _85666_ (_36046_, _36045_, _05669_);
  and _85667_ (_36047_, _36046_, _06020_);
  and _85668_ (_36048_, _36047_, _36043_);
  and _85669_ (_36050_, _36012_, _06019_);
  or _85670_ (_36051_, _36050_, _06112_);
  or _85671_ (_36052_, _36051_, _36048_);
  and _85672_ (_36053_, _14596_, _07681_);
  or _85673_ (_36054_, _36009_, _08751_);
  or _85674_ (_36055_, _36054_, _36053_);
  and _85675_ (_36056_, _36055_, _08756_);
  and _85676_ (_36057_, _36056_, _36052_);
  and _85677_ (_36058_, _10991_, _07681_);
  or _85678_ (_36059_, _36058_, _36009_);
  and _85679_ (_36061_, _36059_, _06284_);
  or _85680_ (_36062_, _36061_, _36057_);
  and _85681_ (_36063_, _36062_, _07032_);
  or _85682_ (_36064_, _36063_, _36014_);
  and _85683_ (_36065_, _36064_, _06278_);
  nor _85684_ (_36066_, _36026_, _06278_);
  and _85685_ (_36067_, _36066_, _36010_);
  or _85686_ (_36068_, _36067_, _06130_);
  or _85687_ (_36069_, _36068_, _36065_);
  and _85688_ (_36070_, _14593_, _07681_);
  or _85689_ (_36072_, _36009_, _08777_);
  or _85690_ (_36073_, _36072_, _36070_);
  and _85691_ (_36074_, _36073_, _08782_);
  and _85692_ (_36075_, _36074_, _36069_);
  nor _85693_ (_36076_, _10990_, _13650_);
  or _85694_ (_36077_, _36076_, _36009_);
  and _85695_ (_36078_, _36077_, _06292_);
  or _85696_ (_36079_, _36078_, _36075_);
  and _85697_ (_36080_, _36079_, _06718_);
  and _85698_ (_36081_, _36023_, _06316_);
  or _85699_ (_36083_, _36081_, _06047_);
  or _85700_ (_36084_, _36083_, _36080_);
  and _85701_ (_36085_, _14657_, _07681_);
  or _85702_ (_36086_, _36009_, _06048_);
  or _85703_ (_36087_, _36086_, _36085_);
  and _85704_ (_36088_, _36087_, _01336_);
  and _85705_ (_36089_, _36088_, _36084_);
  or _85706_ (_36090_, _36089_, _36008_);
  and _85707_ (_43503_, _36090_, _42882_);
  and _85708_ (_36091_, _01340_, \oc8051_golden_model_1.SBUF [3]);
  and _85709_ (_36093_, _13650_, \oc8051_golden_model_1.SBUF [3]);
  and _85710_ (_36094_, _07681_, _08662_);
  or _85711_ (_36095_, _36094_, _36093_);
  or _85712_ (_36096_, _36095_, _06020_);
  and _85713_ (_36097_, _09181_, _07681_);
  or _85714_ (_36098_, _36093_, _07012_);
  or _85715_ (_36099_, _36098_, _36097_);
  and _85716_ (_36100_, _14672_, _07681_);
  or _85717_ (_36101_, _36100_, _36093_);
  or _85718_ (_36102_, _36101_, _06954_);
  and _85719_ (_36104_, _07681_, \oc8051_golden_model_1.ACC [3]);
  or _85720_ (_36105_, _36104_, _36093_);
  and _85721_ (_36106_, _36105_, _06938_);
  and _85722_ (_36107_, _06939_, \oc8051_golden_model_1.SBUF [3]);
  or _85723_ (_36108_, _36107_, _06102_);
  or _85724_ (_36109_, _36108_, _36106_);
  and _85725_ (_36110_, _36109_, _06848_);
  and _85726_ (_36111_, _36110_, _36102_);
  nor _85727_ (_36112_, _13650_, _07353_);
  or _85728_ (_36113_, _36112_, _36093_);
  and _85729_ (_36115_, _36113_, _06239_);
  or _85730_ (_36116_, _36115_, _36111_);
  and _85731_ (_36117_, _36116_, _06220_);
  and _85732_ (_36118_, _36105_, _06219_);
  or _85733_ (_36119_, _36118_, _09818_);
  or _85734_ (_36120_, _36119_, _36117_);
  or _85735_ (_36121_, _36113_, _09827_);
  and _85736_ (_36122_, _36121_, _05669_);
  and _85737_ (_36123_, _36122_, _36120_);
  and _85738_ (_36124_, _36123_, _36099_);
  and _85739_ (_36126_, _14778_, _07681_);
  or _85740_ (_36127_, _36126_, _36093_);
  and _85741_ (_36128_, _36127_, _09833_);
  or _85742_ (_36129_, _36128_, _06019_);
  or _85743_ (_36130_, _36129_, _36124_);
  and _85744_ (_36131_, _36130_, _36096_);
  or _85745_ (_36132_, _36131_, _06112_);
  and _85746_ (_36133_, _14793_, _07681_);
  or _85747_ (_36134_, _36133_, _36093_);
  or _85748_ (_36135_, _36134_, _08751_);
  and _85749_ (_36137_, _36135_, _08756_);
  and _85750_ (_36138_, _36137_, _36132_);
  and _85751_ (_36139_, _12299_, _07681_);
  or _85752_ (_36140_, _36139_, _36093_);
  and _85753_ (_36141_, _36140_, _06284_);
  or _85754_ (_36142_, _36141_, _36138_);
  and _85755_ (_36143_, _36142_, _07032_);
  or _85756_ (_36144_, _36093_, _08029_);
  and _85757_ (_36145_, _36095_, _06108_);
  and _85758_ (_36146_, _36145_, _36144_);
  or _85759_ (_36148_, _36146_, _36143_);
  and _85760_ (_36149_, _36148_, _06278_);
  and _85761_ (_36150_, _36105_, _06277_);
  and _85762_ (_36151_, _36150_, _36144_);
  or _85763_ (_36152_, _36151_, _06130_);
  or _85764_ (_36153_, _36152_, _36149_);
  and _85765_ (_36154_, _14792_, _07681_);
  or _85766_ (_36155_, _36093_, _08777_);
  or _85767_ (_36156_, _36155_, _36154_);
  and _85768_ (_36157_, _36156_, _08782_);
  and _85769_ (_36159_, _36157_, _36153_);
  nor _85770_ (_36160_, _10988_, _13650_);
  or _85771_ (_36161_, _36160_, _36093_);
  and _85772_ (_36162_, _36161_, _06292_);
  or _85773_ (_36163_, _36162_, _36159_);
  and _85774_ (_36164_, _36163_, _06718_);
  and _85775_ (_36165_, _36101_, _06316_);
  or _85776_ (_36166_, _36165_, _06047_);
  or _85777_ (_36167_, _36166_, _36164_);
  and _85778_ (_36168_, _14849_, _07681_);
  or _85779_ (_36170_, _36093_, _06048_);
  or _85780_ (_36171_, _36170_, _36168_);
  and _85781_ (_36172_, _36171_, _01336_);
  and _85782_ (_36173_, _36172_, _36167_);
  or _85783_ (_36174_, _36173_, _36091_);
  and _85784_ (_43505_, _36174_, _42882_);
  and _85785_ (_36175_, _01340_, \oc8051_golden_model_1.SBUF [4]);
  and _85786_ (_36176_, _13650_, \oc8051_golden_model_1.SBUF [4]);
  or _85787_ (_36177_, _36176_, _08273_);
  and _85788_ (_36178_, _08665_, _07681_);
  or _85789_ (_36180_, _36178_, _36176_);
  and _85790_ (_36181_, _36180_, _06108_);
  and _85791_ (_36182_, _36181_, _36177_);
  and _85792_ (_36183_, _14887_, _07681_);
  or _85793_ (_36184_, _36183_, _36176_);
  or _85794_ (_36185_, _36184_, _06954_);
  and _85795_ (_36186_, _07681_, \oc8051_golden_model_1.ACC [4]);
  or _85796_ (_36187_, _36186_, _36176_);
  and _85797_ (_36188_, _36187_, _06938_);
  and _85798_ (_36189_, _06939_, \oc8051_golden_model_1.SBUF [4]);
  or _85799_ (_36191_, _36189_, _06102_);
  or _85800_ (_36192_, _36191_, _36188_);
  and _85801_ (_36193_, _36192_, _06848_);
  and _85802_ (_36194_, _36193_, _36185_);
  nor _85803_ (_36195_, _08270_, _13650_);
  or _85804_ (_36196_, _36195_, _36176_);
  and _85805_ (_36197_, _36196_, _06239_);
  or _85806_ (_36198_, _36197_, _36194_);
  and _85807_ (_36199_, _36198_, _06220_);
  and _85808_ (_36200_, _36187_, _06219_);
  or _85809_ (_36202_, _36200_, _09815_);
  or _85810_ (_36203_, _36202_, _36199_);
  or _85811_ (_36204_, _36196_, _09827_);
  and _85812_ (_36205_, _36204_, _07012_);
  and _85813_ (_36206_, _36205_, _36203_);
  and _85814_ (_36207_, _09180_, _07681_);
  or _85815_ (_36208_, _36207_, _36176_);
  and _85816_ (_36209_, _36208_, _07011_);
  or _85817_ (_36210_, _36209_, _09833_);
  or _85818_ (_36211_, _36210_, _36206_);
  and _85819_ (_36213_, _14983_, _07681_);
  or _85820_ (_36214_, _36176_, _05669_);
  or _85821_ (_36215_, _36214_, _36213_);
  and _85822_ (_36216_, _36215_, _06020_);
  and _85823_ (_36217_, _36216_, _36211_);
  and _85824_ (_36218_, _36180_, _06019_);
  or _85825_ (_36219_, _36218_, _06112_);
  or _85826_ (_36220_, _36219_, _36217_);
  and _85827_ (_36221_, _14876_, _07681_);
  or _85828_ (_36222_, _36176_, _08751_);
  or _85829_ (_36224_, _36222_, _36221_);
  and _85830_ (_36225_, _36224_, _08756_);
  and _85831_ (_36226_, _36225_, _36220_);
  and _85832_ (_36227_, _10986_, _07681_);
  or _85833_ (_36228_, _36227_, _36176_);
  and _85834_ (_36229_, _36228_, _06284_);
  or _85835_ (_36230_, _36229_, _36226_);
  and _85836_ (_36231_, _36230_, _07032_);
  or _85837_ (_36232_, _36231_, _36182_);
  and _85838_ (_36233_, _36232_, _06278_);
  and _85839_ (_36235_, _36187_, _06277_);
  and _85840_ (_36236_, _36235_, _36177_);
  or _85841_ (_36237_, _36236_, _06130_);
  or _85842_ (_36238_, _36237_, _36233_);
  and _85843_ (_36239_, _14873_, _07681_);
  or _85844_ (_36240_, _36176_, _08777_);
  or _85845_ (_36241_, _36240_, _36239_);
  and _85846_ (_36242_, _36241_, _08782_);
  and _85847_ (_36243_, _36242_, _36238_);
  nor _85848_ (_36244_, _10985_, _13650_);
  or _85849_ (_36246_, _36244_, _36176_);
  and _85850_ (_36247_, _36246_, _06292_);
  or _85851_ (_36248_, _36247_, _36243_);
  and _85852_ (_36249_, _36248_, _06718_);
  and _85853_ (_36250_, _36184_, _06316_);
  or _85854_ (_36251_, _36250_, _06047_);
  or _85855_ (_36252_, _36251_, _36249_);
  and _85856_ (_36253_, _15055_, _07681_);
  or _85857_ (_36254_, _36176_, _06048_);
  or _85858_ (_36255_, _36254_, _36253_);
  and _85859_ (_36257_, _36255_, _01336_);
  and _85860_ (_36258_, _36257_, _36252_);
  or _85861_ (_36259_, _36258_, _36175_);
  and _85862_ (_43506_, _36259_, _42882_);
  and _85863_ (_36260_, _01340_, \oc8051_golden_model_1.SBUF [5]);
  and _85864_ (_36261_, _13650_, \oc8051_golden_model_1.SBUF [5]);
  or _85865_ (_36262_, _36261_, _07980_);
  and _85866_ (_36263_, _08652_, _07681_);
  or _85867_ (_36264_, _36263_, _36261_);
  and _85868_ (_36265_, _36264_, _06108_);
  and _85869_ (_36267_, _36265_, _36262_);
  or _85870_ (_36268_, _36264_, _06020_);
  and _85871_ (_36269_, _15093_, _07681_);
  or _85872_ (_36270_, _36269_, _36261_);
  or _85873_ (_36271_, _36270_, _06954_);
  and _85874_ (_36272_, _07681_, \oc8051_golden_model_1.ACC [5]);
  or _85875_ (_36273_, _36272_, _36261_);
  and _85876_ (_36274_, _36273_, _06938_);
  and _85877_ (_36275_, _06939_, \oc8051_golden_model_1.SBUF [5]);
  or _85878_ (_36276_, _36275_, _06102_);
  or _85879_ (_36278_, _36276_, _36274_);
  and _85880_ (_36279_, _36278_, _06848_);
  and _85881_ (_36280_, _36279_, _36271_);
  nor _85882_ (_36281_, _07977_, _13650_);
  or _85883_ (_36282_, _36281_, _36261_);
  and _85884_ (_36283_, _36282_, _06239_);
  or _85885_ (_36284_, _36283_, _36280_);
  and _85886_ (_36285_, _36284_, _06220_);
  and _85887_ (_36286_, _36273_, _06219_);
  or _85888_ (_36287_, _36286_, _09818_);
  or _85889_ (_36289_, _36287_, _36285_);
  and _85890_ (_36290_, _09179_, _07681_);
  or _85891_ (_36291_, _36261_, _07012_);
  or _85892_ (_36292_, _36291_, _36290_);
  or _85893_ (_36293_, _36282_, _09827_);
  and _85894_ (_36294_, _36293_, _05669_);
  and _85895_ (_36295_, _36294_, _36292_);
  and _85896_ (_36296_, _36295_, _36289_);
  and _85897_ (_36297_, _15179_, _07681_);
  or _85898_ (_36298_, _36297_, _36261_);
  and _85899_ (_36300_, _36298_, _09833_);
  or _85900_ (_36301_, _36300_, _06019_);
  or _85901_ (_36302_, _36301_, _36296_);
  and _85902_ (_36303_, _36302_, _36268_);
  or _85903_ (_36304_, _36303_, _06112_);
  and _85904_ (_36305_, _15195_, _07681_);
  or _85905_ (_36306_, _36305_, _36261_);
  or _85906_ (_36307_, _36306_, _08751_);
  and _85907_ (_36308_, _36307_, _08756_);
  and _85908_ (_36309_, _36308_, _36304_);
  and _85909_ (_36311_, _12306_, _07681_);
  or _85910_ (_36312_, _36311_, _36261_);
  and _85911_ (_36313_, _36312_, _06284_);
  or _85912_ (_36314_, _36313_, _36309_);
  and _85913_ (_36315_, _36314_, _07032_);
  or _85914_ (_36316_, _36315_, _36267_);
  and _85915_ (_36317_, _36316_, _06278_);
  and _85916_ (_36318_, _36273_, _06277_);
  and _85917_ (_36319_, _36318_, _36262_);
  or _85918_ (_36320_, _36319_, _06130_);
  or _85919_ (_36322_, _36320_, _36317_);
  and _85920_ (_36323_, _15194_, _07681_);
  or _85921_ (_36324_, _36261_, _08777_);
  or _85922_ (_36325_, _36324_, _36323_);
  and _85923_ (_36326_, _36325_, _08782_);
  and _85924_ (_36327_, _36326_, _36322_);
  nor _85925_ (_36328_, _10982_, _13650_);
  or _85926_ (_36329_, _36328_, _36261_);
  and _85927_ (_36330_, _36329_, _06292_);
  or _85928_ (_36331_, _36330_, _36327_);
  and _85929_ (_36333_, _36331_, _06718_);
  and _85930_ (_36334_, _36270_, _06316_);
  or _85931_ (_36335_, _36334_, _06047_);
  or _85932_ (_36336_, _36335_, _36333_);
  and _85933_ (_36337_, _15253_, _07681_);
  or _85934_ (_36338_, _36261_, _06048_);
  or _85935_ (_36339_, _36338_, _36337_);
  and _85936_ (_36340_, _36339_, _01336_);
  and _85937_ (_36341_, _36340_, _36336_);
  or _85938_ (_36342_, _36341_, _36260_);
  and _85939_ (_43507_, _36342_, _42882_);
  and _85940_ (_36344_, _01340_, \oc8051_golden_model_1.SBUF [6]);
  and _85941_ (_36345_, _13650_, \oc8051_golden_model_1.SBUF [6]);
  and _85942_ (_36346_, _15389_, _07681_);
  or _85943_ (_36347_, _36346_, _36345_);
  or _85944_ (_36348_, _36347_, _06020_);
  and _85945_ (_36349_, _15293_, _07681_);
  or _85946_ (_36350_, _36349_, _36345_);
  or _85947_ (_36351_, _36350_, _06954_);
  and _85948_ (_36352_, _07681_, \oc8051_golden_model_1.ACC [6]);
  or _85949_ (_36354_, _36352_, _36345_);
  and _85950_ (_36355_, _36354_, _06938_);
  and _85951_ (_36356_, _06939_, \oc8051_golden_model_1.SBUF [6]);
  or _85952_ (_36357_, _36356_, _06102_);
  or _85953_ (_36358_, _36357_, _36355_);
  and _85954_ (_36359_, _36358_, _06848_);
  and _85955_ (_36360_, _36359_, _36351_);
  nor _85956_ (_36361_, _07883_, _13650_);
  or _85957_ (_36362_, _36361_, _36345_);
  and _85958_ (_36363_, _36362_, _06239_);
  or _85959_ (_36364_, _36363_, _36360_);
  and _85960_ (_36365_, _36364_, _06220_);
  and _85961_ (_36366_, _36354_, _06219_);
  or _85962_ (_36367_, _36366_, _09818_);
  or _85963_ (_36368_, _36367_, _36365_);
  and _85964_ (_36369_, _09178_, _07681_);
  or _85965_ (_36370_, _36345_, _07012_);
  or _85966_ (_36371_, _36370_, _36369_);
  or _85967_ (_36372_, _36362_, _09827_);
  and _85968_ (_36373_, _36372_, _05669_);
  and _85969_ (_36375_, _36373_, _36371_);
  and _85970_ (_36376_, _36375_, _36368_);
  and _85971_ (_36377_, _15382_, _07681_);
  or _85972_ (_36378_, _36377_, _36345_);
  and _85973_ (_36379_, _36378_, _09833_);
  or _85974_ (_36380_, _36379_, _06019_);
  or _85975_ (_36381_, _36380_, _36376_);
  and _85976_ (_36382_, _36381_, _36348_);
  or _85977_ (_36383_, _36382_, _06112_);
  and _85978_ (_36384_, _15399_, _07681_);
  or _85979_ (_36386_, _36384_, _36345_);
  or _85980_ (_36387_, _36386_, _08751_);
  and _85981_ (_36388_, _36387_, _08756_);
  and _85982_ (_36389_, _36388_, _36383_);
  and _85983_ (_36390_, _10980_, _07681_);
  or _85984_ (_36391_, _36390_, _36345_);
  and _85985_ (_36392_, _36391_, _06284_);
  or _85986_ (_36393_, _36392_, _36389_);
  and _85987_ (_36394_, _36393_, _07032_);
  or _85988_ (_36395_, _36345_, _07886_);
  and _85989_ (_36397_, _36347_, _06108_);
  and _85990_ (_36398_, _36397_, _36395_);
  or _85991_ (_36399_, _36398_, _36394_);
  and _85992_ (_36400_, _36399_, _06278_);
  and _85993_ (_36401_, _36354_, _06277_);
  and _85994_ (_36402_, _36401_, _36395_);
  or _85995_ (_36403_, _36402_, _06130_);
  or _85996_ (_36404_, _36403_, _36400_);
  and _85997_ (_36405_, _15396_, _07681_);
  or _85998_ (_36406_, _36345_, _08777_);
  or _85999_ (_36408_, _36406_, _36405_);
  and _86000_ (_36409_, _36408_, _08782_);
  and _86001_ (_36410_, _36409_, _36404_);
  nor _86002_ (_36411_, _10979_, _13650_);
  or _86003_ (_36412_, _36411_, _36345_);
  and _86004_ (_36413_, _36412_, _06292_);
  or _86005_ (_36414_, _36413_, _36410_);
  and _86006_ (_36415_, _36414_, _06718_);
  and _86007_ (_36416_, _36350_, _06316_);
  or _86008_ (_36417_, _36416_, _06047_);
  or _86009_ (_36419_, _36417_, _36415_);
  and _86010_ (_36420_, _15451_, _07681_);
  or _86011_ (_36421_, _36345_, _06048_);
  or _86012_ (_36422_, _36421_, _36420_);
  and _86013_ (_36423_, _36422_, _01336_);
  and _86014_ (_36424_, _36423_, _36419_);
  or _86015_ (_36425_, _36424_, _36344_);
  and _86016_ (_43508_, _36425_, _42882_);
  not _86017_ (_36426_, \oc8051_golden_model_1.PSW [0]);
  nor _86018_ (_36427_, _01336_, _36426_);
  nand _86019_ (_36429_, _10995_, _07705_);
  nor _86020_ (_36430_, _07705_, _36426_);
  nor _86021_ (_36431_, _36430_, _06278_);
  nand _86022_ (_36432_, _36431_, _36429_);
  and _86023_ (_36433_, _07705_, _08672_);
  or _86024_ (_36434_, _36433_, _36430_);
  or _86025_ (_36435_, _36434_, _06020_);
  and _86026_ (_36436_, _09120_, _07705_);
  or _86027_ (_36437_, _36430_, _07012_);
  or _86028_ (_36438_, _36437_, _36436_);
  nor _86029_ (_36440_, _08127_, _13745_);
  or _86030_ (_36441_, _36440_, _36430_);
  or _86031_ (_36442_, _36441_, _06954_);
  and _86032_ (_36443_, _07705_, \oc8051_golden_model_1.ACC [0]);
  or _86033_ (_36444_, _36443_, _36430_);
  and _86034_ (_36445_, _36444_, _06938_);
  nor _86035_ (_36446_, _06938_, _36426_);
  or _86036_ (_36447_, _36446_, _06102_);
  or _86037_ (_36448_, _36447_, _36445_);
  and _86038_ (_36449_, _36448_, _06044_);
  and _86039_ (_36451_, _36449_, _36442_);
  nor _86040_ (_36452_, _08355_, _36426_);
  and _86041_ (_36453_, _14102_, _08355_);
  or _86042_ (_36454_, _36453_, _36452_);
  and _86043_ (_36455_, _36454_, _06043_);
  or _86044_ (_36456_, _36455_, _36451_);
  and _86045_ (_36457_, _36456_, _06848_);
  and _86046_ (_36458_, _07705_, _06931_);
  or _86047_ (_36459_, _36458_, _36430_);
  and _86048_ (_36460_, _36459_, _06239_);
  or _86049_ (_36462_, _36460_, _06219_);
  or _86050_ (_36463_, _36462_, _36457_);
  or _86051_ (_36464_, _36444_, _06220_);
  and _86052_ (_36465_, _36464_, _06040_);
  and _86053_ (_36466_, _36465_, _36463_);
  and _86054_ (_36467_, _36430_, _06039_);
  or _86055_ (_36468_, _36467_, _06032_);
  or _86056_ (_36469_, _36468_, _36466_);
  or _86057_ (_36470_, _36441_, _06033_);
  and _86058_ (_36471_, _36470_, _06027_);
  and _86059_ (_36473_, _36471_, _36469_);
  or _86060_ (_36474_, _36452_, _14131_);
  and _86061_ (_36475_, _36474_, _06026_);
  and _86062_ (_36476_, _36475_, _36454_);
  or _86063_ (_36477_, _36476_, _09818_);
  or _86064_ (_36478_, _36477_, _36473_);
  or _86065_ (_36479_, _36459_, _09827_);
  and _86066_ (_36480_, _36479_, _05669_);
  and _86067_ (_36481_, _36480_, _36478_);
  and _86068_ (_36482_, _36481_, _36438_);
  and _86069_ (_36484_, _14186_, _07705_);
  or _86070_ (_36485_, _36484_, _36430_);
  and _86071_ (_36486_, _36485_, _09833_);
  or _86072_ (_36487_, _36486_, _06019_);
  or _86073_ (_36488_, _36487_, _36482_);
  and _86074_ (_36489_, _36488_, _36435_);
  or _86075_ (_36490_, _36489_, _06112_);
  and _86076_ (_36491_, _14086_, _07705_);
  or _86077_ (_36492_, _36491_, _36430_);
  or _86078_ (_36493_, _36492_, _08751_);
  and _86079_ (_36495_, _36493_, _08756_);
  and _86080_ (_36496_, _36495_, _36490_);
  nor _86081_ (_36497_, _12302_, _13745_);
  or _86082_ (_36498_, _36497_, _36430_);
  and _86083_ (_36499_, _36429_, _06284_);
  and _86084_ (_36500_, _36499_, _36498_);
  or _86085_ (_36501_, _36500_, _36496_);
  and _86086_ (_36502_, _36501_, _07032_);
  nand _86087_ (_36503_, _36434_, _06108_);
  nor _86088_ (_36504_, _36503_, _36440_);
  or _86089_ (_36506_, _36504_, _06277_);
  or _86090_ (_36507_, _36506_, _36502_);
  and _86091_ (_36508_, _36507_, _36432_);
  or _86092_ (_36509_, _36508_, _06130_);
  and _86093_ (_36510_, _14083_, _07705_);
  or _86094_ (_36511_, _36430_, _08777_);
  or _86095_ (_36512_, _36511_, _36510_);
  and _86096_ (_36513_, _36512_, _08782_);
  and _86097_ (_36514_, _36513_, _36509_);
  and _86098_ (_36515_, _36498_, _06292_);
  or _86099_ (_36517_, _36515_, _06316_);
  or _86100_ (_36518_, _36517_, _36514_);
  or _86101_ (_36519_, _36441_, _06718_);
  and _86102_ (_36520_, _36519_, _36518_);
  or _86103_ (_36521_, _36520_, _05652_);
  or _86104_ (_36522_, _36430_, _05653_);
  and _86105_ (_36523_, _36522_, _36521_);
  or _86106_ (_36524_, _36523_, _06047_);
  or _86107_ (_36525_, _36441_, _06048_);
  and _86108_ (_36526_, _36525_, _01336_);
  and _86109_ (_36528_, _36526_, _36524_);
  or _86110_ (_36529_, _36528_, _36427_);
  and _86111_ (_43510_, _36529_, _42882_);
  not _86112_ (_36530_, \oc8051_golden_model_1.PSW [1]);
  nor _86113_ (_36531_, _01336_, _36530_);
  nor _86114_ (_36532_, _07705_, _36530_);
  nor _86115_ (_36533_, _10993_, _13745_);
  or _86116_ (_36534_, _36533_, _36532_);
  or _86117_ (_36535_, _36534_, _08782_);
  or _86118_ (_36536_, _14367_, _13745_);
  or _86119_ (_36538_, _07705_, \oc8051_golden_model_1.PSW [1]);
  and _86120_ (_36539_, _36538_, _09833_);
  and _86121_ (_36540_, _36539_, _36536_);
  and _86122_ (_36541_, _09075_, _07705_);
  or _86123_ (_36542_, _36541_, _36532_);
  and _86124_ (_36543_, _36542_, _07011_);
  nor _86125_ (_36544_, _13745_, _07132_);
  or _86126_ (_36545_, _36544_, _36532_);
  and _86127_ (_36546_, _36545_, _06239_);
  nor _86128_ (_36547_, _08355_, _36530_);
  and _86129_ (_36549_, _14266_, _08355_);
  or _86130_ (_36550_, _36549_, _36547_);
  or _86131_ (_36551_, _36550_, _06044_);
  and _86132_ (_36552_, _14284_, _07705_);
  not _86133_ (_36553_, _36552_);
  and _86134_ (_36554_, _36553_, _36538_);
  and _86135_ (_36555_, _36554_, _06102_);
  nor _86136_ (_36556_, _06938_, _36530_);
  and _86137_ (_36557_, _07705_, \oc8051_golden_model_1.ACC [1]);
  or _86138_ (_36558_, _36557_, _36532_);
  and _86139_ (_36560_, _36558_, _06938_);
  or _86140_ (_36561_, _36560_, _36556_);
  and _86141_ (_36562_, _36561_, _06954_);
  or _86142_ (_36563_, _36562_, _06043_);
  or _86143_ (_36564_, _36563_, _36555_);
  and _86144_ (_36565_, _36564_, _36551_);
  and _86145_ (_36566_, _36565_, _06848_);
  or _86146_ (_36567_, _36566_, _36546_);
  or _86147_ (_36568_, _36567_, _06219_);
  or _86148_ (_36569_, _36558_, _06220_);
  and _86149_ (_36571_, _36569_, _06040_);
  and _86150_ (_36572_, _36571_, _36568_);
  and _86151_ (_36573_, _14273_, _08355_);
  or _86152_ (_36574_, _36573_, _36547_);
  and _86153_ (_36575_, _36574_, _06039_);
  or _86154_ (_36576_, _36575_, _06032_);
  or _86155_ (_36577_, _36576_, _36572_);
  or _86156_ (_36578_, _36547_, _14302_);
  and _86157_ (_36579_, _36578_, _36550_);
  or _86158_ (_36580_, _36579_, _06033_);
  and _86159_ (_36582_, _36580_, _06027_);
  and _86160_ (_36583_, _36582_, _36577_);
  or _86161_ (_36584_, _36547_, _14267_);
  and _86162_ (_36585_, _36584_, _06026_);
  and _86163_ (_36586_, _36585_, _36550_);
  or _86164_ (_36587_, _36586_, _09815_);
  or _86165_ (_36588_, _36587_, _36583_);
  or _86166_ (_36589_, _36545_, _09827_);
  and _86167_ (_36590_, _36589_, _07012_);
  and _86168_ (_36591_, _36590_, _36588_);
  or _86169_ (_36593_, _36591_, _36543_);
  and _86170_ (_36594_, _36593_, _05669_);
  or _86171_ (_36595_, _36594_, _36540_);
  and _86172_ (_36596_, _36595_, _06020_);
  nand _86173_ (_36597_, _07705_, _06832_);
  and _86174_ (_36598_, _36538_, _06019_);
  and _86175_ (_36599_, _36598_, _36597_);
  or _86176_ (_36600_, _36599_, _36596_);
  and _86177_ (_36601_, _36600_, _08751_);
  or _86178_ (_36602_, _14263_, _13745_);
  and _86179_ (_36604_, _36538_, _06112_);
  and _86180_ (_36605_, _36604_, _36602_);
  or _86181_ (_36606_, _36605_, _06284_);
  or _86182_ (_36607_, _36606_, _36601_);
  nand _86183_ (_36608_, _10992_, _07705_);
  and _86184_ (_36609_, _36608_, _36534_);
  or _86185_ (_36610_, _36609_, _08756_);
  and _86186_ (_36611_, _36610_, _07032_);
  and _86187_ (_36612_, _36611_, _36607_);
  or _86188_ (_36613_, _14261_, _13745_);
  and _86189_ (_36615_, _36538_, _06108_);
  and _86190_ (_36616_, _36615_, _36613_);
  or _86191_ (_36617_, _36616_, _06277_);
  or _86192_ (_36618_, _36617_, _36612_);
  nor _86193_ (_36619_, _36532_, _06278_);
  nand _86194_ (_36620_, _36619_, _36608_);
  and _86195_ (_36621_, _36620_, _08777_);
  and _86196_ (_36622_, _36621_, _36618_);
  or _86197_ (_36623_, _36597_, _08078_);
  and _86198_ (_36624_, _36538_, _06130_);
  and _86199_ (_36626_, _36624_, _36623_);
  or _86200_ (_36627_, _36626_, _06292_);
  or _86201_ (_36628_, _36627_, _36622_);
  and _86202_ (_36629_, _36628_, _36535_);
  or _86203_ (_36630_, _36629_, _06316_);
  or _86204_ (_36631_, _36554_, _06718_);
  and _86205_ (_36632_, _36631_, _05653_);
  and _86206_ (_36633_, _36632_, _36630_);
  and _86207_ (_36634_, _36574_, _05652_);
  or _86208_ (_36635_, _36634_, _06047_);
  or _86209_ (_36637_, _36635_, _36633_);
  or _86210_ (_36638_, _36532_, _06048_);
  or _86211_ (_36639_, _36638_, _36552_);
  and _86212_ (_36640_, _36639_, _01336_);
  and _86213_ (_36641_, _36640_, _36637_);
  or _86214_ (_36642_, _36641_, _36531_);
  and _86215_ (_43511_, _36642_, _42882_);
  not _86216_ (_36643_, \oc8051_golden_model_1.PSW [2]);
  nor _86217_ (_36644_, _01336_, _36643_);
  not _86218_ (_36645_, _10692_);
  nand _86219_ (_36647_, _10967_, _36645_);
  or _86220_ (_36648_, _10967_, _10691_);
  and _86221_ (_36649_, _36648_, _36647_);
  and _86222_ (_36650_, _36649_, _06692_);
  nor _86223_ (_36651_, _10570_, _13739_);
  not _86224_ (_36652_, _36651_);
  nor _86225_ (_36653_, _10570_, _06053_);
  or _86226_ (_36654_, _36653_, \oc8051_golden_model_1.ACC [7]);
  and _86227_ (_36655_, _36654_, _36652_);
  not _86228_ (_36656_, _36655_);
  or _86229_ (_36658_, _36656_, _14017_);
  and _86230_ (_36659_, _36658_, _10880_);
  or _86231_ (_36660_, _36659_, _36651_);
  or _86232_ (_36661_, _36652_, _10877_);
  and _86233_ (_36662_, _36661_, _10824_);
  and _86234_ (_36663_, _36662_, _36660_);
  and _86235_ (_36664_, _09182_, _07705_);
  nor _86236_ (_36665_, _07705_, _36643_);
  or _86237_ (_36666_, _36665_, _07012_);
  or _86238_ (_36667_, _36666_, _36664_);
  nor _86239_ (_36669_, _13745_, _07530_);
  or _86240_ (_36670_, _36669_, _36665_);
  or _86241_ (_36671_, _36670_, _09827_);
  nor _86242_ (_36672_, _10496_, \oc8051_golden_model_1.ACC [7]);
  nor _86243_ (_36673_, _10495_, _36645_);
  nor _86244_ (_36674_, _36673_, _36672_);
  nor _86245_ (_36675_, _36674_, _10501_);
  nor _86246_ (_36676_, _13934_, _10497_);
  nor _86247_ (_36677_, _36676_, _36675_);
  and _86248_ (_36678_, _36677_, _10556_);
  nor _86249_ (_36680_, _36677_, _10556_);
  or _86250_ (_36681_, _36680_, _36678_);
  and _86251_ (_36682_, _36681_, _12361_);
  nor _86252_ (_36683_, _08355_, _36643_);
  and _86253_ (_36684_, _14479_, _08355_);
  or _86254_ (_36685_, _36684_, _36683_);
  and _86255_ (_36686_, _36685_, _06039_);
  or _86256_ (_36687_, _36670_, _06848_);
  and _86257_ (_36688_, _14493_, _07705_);
  or _86258_ (_36689_, _36688_, _36665_);
  or _86259_ (_36691_, _36689_, _06954_);
  and _86260_ (_36692_, _07705_, \oc8051_golden_model_1.ACC [2]);
  or _86261_ (_36693_, _36692_, _36665_);
  and _86262_ (_36694_, _36693_, _06938_);
  nor _86263_ (_36695_, _06938_, _36643_);
  or _86264_ (_36696_, _36695_, _06102_);
  or _86265_ (_36697_, _36696_, _36694_);
  and _86266_ (_36698_, _36697_, _06044_);
  and _86267_ (_36699_, _36698_, _36691_);
  and _86268_ (_36700_, _14497_, _08355_);
  or _86269_ (_36702_, _36700_, _36683_);
  and _86270_ (_36703_, _36702_, _06043_);
  or _86271_ (_36704_, _36703_, _06239_);
  or _86272_ (_36705_, _36704_, _36699_);
  and _86273_ (_36706_, _36705_, _36687_);
  or _86274_ (_36707_, _36706_, _06219_);
  or _86275_ (_36708_, _36693_, _06220_);
  and _86276_ (_36709_, _36708_, _06040_);
  and _86277_ (_36710_, _36709_, _36707_);
  or _86278_ (_36711_, _36710_, _36686_);
  and _86279_ (_36713_, _36711_, _06033_);
  and _86280_ (_36714_, _36700_, _14512_);
  or _86281_ (_36715_, _36714_, _36683_);
  and _86282_ (_36716_, _36715_, _06032_);
  or _86283_ (_36717_, _36716_, _36713_);
  and _86284_ (_36718_, _36717_, _09800_);
  or _86285_ (_36719_, _16187_, _09803_);
  or _86286_ (_36720_, _36719_, _16295_);
  or _86287_ (_36721_, _36720_, _16411_);
  or _86288_ (_36722_, _36721_, _16527_);
  or _86289_ (_36724_, _36722_, _16643_);
  or _86290_ (_36725_, _36724_, _16757_);
  or _86291_ (_36726_, _36725_, _16877_);
  and _86292_ (_36727_, _36726_, _09269_);
  or _86293_ (_36728_, _36727_, _10468_);
  or _86294_ (_36729_, _36728_, _36718_);
  nor _86295_ (_36730_, _10719_, _10240_);
  or _86296_ (_36731_, _10240_, _07785_);
  and _86297_ (_36732_, _36731_, _08393_);
  or _86298_ (_36733_, _36732_, _36730_);
  and _86299_ (_36735_, _36733_, _13925_);
  nor _86300_ (_36736_, _36733_, _13925_);
  nor _86301_ (_36737_, _36736_, _36735_);
  not _86302_ (_36738_, _36737_);
  nor _86303_ (_36739_, _36738_, _10490_);
  and _86304_ (_36740_, _36738_, _10490_);
  or _86305_ (_36741_, _36740_, _36739_);
  or _86306_ (_36742_, _36741_, _10469_);
  and _86307_ (_36743_, _36742_, _13935_);
  and _86308_ (_36744_, _36743_, _36729_);
  or _86309_ (_36746_, _36744_, _36682_);
  and _86310_ (_36747_, _36746_, _06267_);
  nor _86311_ (_36748_, _10314_, _14043_);
  nor _86312_ (_36749_, _10315_, \oc8051_golden_model_1.ACC [7]);
  nor _86313_ (_36750_, _36749_, _36748_);
  nor _86314_ (_36751_, _36750_, _10320_);
  nor _86315_ (_36752_, _13761_, _10316_);
  or _86316_ (_36753_, _36752_, _36751_);
  nand _86317_ (_36754_, _36753_, _10370_);
  or _86318_ (_36755_, _36753_, _10370_);
  and _86319_ (_36757_, _36755_, _06261_);
  and _86320_ (_36758_, _36757_, _36754_);
  or _86321_ (_36759_, _36758_, _10306_);
  or _86322_ (_36760_, _36759_, _36747_);
  nor _86323_ (_36761_, _36655_, _13947_);
  and _86324_ (_36762_, _36655_, _13947_);
  nor _86325_ (_36763_, _36762_, _36761_);
  and _86326_ (_36764_, _36763_, _10631_);
  nor _86327_ (_36765_, _36763_, _10631_);
  or _86328_ (_36766_, _36765_, _36764_);
  or _86329_ (_36768_, _36766_, _10307_);
  and _86330_ (_36769_, _36768_, _06027_);
  and _86331_ (_36770_, _36769_, _36760_);
  or _86332_ (_36771_, _36683_, _14525_);
  and _86333_ (_36772_, _36771_, _06026_);
  and _86334_ (_36773_, _36772_, _36702_);
  or _86335_ (_36774_, _36773_, _09815_);
  or _86336_ (_36775_, _36774_, _36770_);
  and _86337_ (_36776_, _36775_, _36671_);
  or _86338_ (_36777_, _36776_, _07011_);
  and _86339_ (_36779_, _36777_, _36667_);
  or _86340_ (_36780_, _36779_, _09833_);
  and _86341_ (_36781_, _14580_, _07705_);
  or _86342_ (_36782_, _36665_, _05669_);
  or _86343_ (_36783_, _36782_, _36781_);
  and _86344_ (_36784_, _36783_, _09839_);
  and _86345_ (_36785_, _36784_, _36780_);
  nor _86346_ (_36786_, \oc8051_golden_model_1.B [1], \oc8051_golden_model_1.B [0]);
  and _86347_ (_36787_, _36786_, _09832_);
  and _86348_ (_36788_, _36787_, _09860_);
  or _86349_ (_36790_, _36788_, _06019_);
  or _86350_ (_36791_, _36790_, _36785_);
  and _86351_ (_36792_, _07705_, _08730_);
  or _86352_ (_36793_, _36792_, _36665_);
  or _86353_ (_36794_, _36793_, _06020_);
  and _86354_ (_36795_, _36794_, _36791_);
  or _86355_ (_36796_, _36795_, _06112_);
  and _86356_ (_36797_, _14596_, _07705_);
  or _86357_ (_36798_, _36797_, _36665_);
  or _86358_ (_36799_, _36798_, _08751_);
  and _86359_ (_36801_, _36799_, _08756_);
  and _86360_ (_36802_, _36801_, _36796_);
  and _86361_ (_36803_, _10991_, _07705_);
  or _86362_ (_36804_, _36803_, _36665_);
  and _86363_ (_36805_, _36804_, _06284_);
  or _86364_ (_36806_, _36805_, _36802_);
  and _86365_ (_36807_, _36806_, _07032_);
  or _86366_ (_36808_, _36665_, _08177_);
  and _86367_ (_36809_, _36793_, _06108_);
  and _86368_ (_36810_, _36809_, _36808_);
  or _86369_ (_36812_, _36810_, _36807_);
  and _86370_ (_36813_, _36812_, _06278_);
  and _86371_ (_36814_, _36693_, _06277_);
  and _86372_ (_36815_, _36814_, _36808_);
  or _86373_ (_36816_, _36815_, _06130_);
  or _86374_ (_36817_, _36816_, _36813_);
  and _86375_ (_36818_, _14593_, _07705_);
  or _86376_ (_36819_, _36665_, _08777_);
  or _86377_ (_36820_, _36819_, _36818_);
  and _86378_ (_36821_, _36820_, _08782_);
  and _86379_ (_36823_, _36821_, _36817_);
  nor _86380_ (_36824_, _10990_, _13745_);
  or _86381_ (_36825_, _36824_, _36665_);
  and _86382_ (_36826_, _36825_, _06292_);
  or _86383_ (_36827_, _36826_, _10303_);
  or _86384_ (_36828_, _36827_, _36823_);
  nor _86385_ (_36829_, _36733_, _13999_);
  nor _86386_ (_36830_, _36829_, _36730_);
  and _86387_ (_36831_, _36830_, _10302_);
  and _86388_ (_36832_, _36730_, _10299_);
  or _86389_ (_36834_, _36832_, _10304_);
  or _86390_ (_36835_, _36834_, _36831_);
  and _86391_ (_36836_, _36835_, _17410_);
  and _86392_ (_36837_, _36836_, _36828_);
  not _86393_ (_36838_, _36674_);
  nor _86394_ (_36839_, _36838_, _14006_);
  nor _86395_ (_36840_, _36839_, _36673_);
  and _86396_ (_36841_, _36840_, _10820_);
  and _86397_ (_36842_, _36673_, _10817_);
  or _86398_ (_36843_, _36842_, _36841_);
  and _86399_ (_36845_, _36843_, _17409_);
  or _86400_ (_36846_, _36845_, _36837_);
  and _86401_ (_36847_, _36846_, _17423_);
  nand _86402_ (_36848_, _36843_, _17416_);
  nand _86403_ (_36849_, _36848_, _06289_);
  or _86404_ (_36850_, _36849_, _36847_);
  nor _86405_ (_36851_, _36749_, _14011_);
  nor _86406_ (_36852_, _36851_, _36748_);
  and _86407_ (_36853_, _36852_, _10850_);
  and _86408_ (_36854_, _36748_, _10847_);
  or _86409_ (_36856_, _36854_, _36853_);
  or _86410_ (_36857_, _36856_, _06289_);
  and _86411_ (_36858_, _36857_, _10856_);
  and _86412_ (_36859_, _36858_, _36850_);
  or _86413_ (_36860_, _36859_, _36663_);
  and _86414_ (_36861_, _36860_, _10890_);
  nand _86415_ (_36862_, _10926_, _10719_);
  and _86416_ (_36863_, _36862_, _16956_);
  and _86417_ (_36864_, _36863_, _14027_);
  or _86418_ (_36865_, _36864_, _17437_);
  or _86419_ (_36867_, _36865_, _36861_);
  and _86420_ (_36868_, _36649_, _17443_);
  or _86421_ (_36869_, _36868_, _10934_);
  and _86422_ (_36870_, _36869_, _36867_);
  or _86423_ (_36871_, _36870_, _36650_);
  and _86424_ (_36872_, _36871_, _10975_);
  or _86425_ (_36873_, _11008_, _08767_);
  and _86426_ (_36874_, _14045_, _36873_);
  nand _86427_ (_36875_, _11048_, _13739_);
  and _86428_ (_36876_, _36875_, _13741_);
  or _86429_ (_36878_, _36876_, _06316_);
  or _86430_ (_36879_, _36878_, _36874_);
  or _86431_ (_36880_, _36879_, _36872_);
  or _86432_ (_36881_, _36689_, _06718_);
  and _86433_ (_36882_, _36881_, _05653_);
  and _86434_ (_36883_, _36882_, _36880_);
  and _86435_ (_36884_, _36685_, _05652_);
  or _86436_ (_36885_, _36884_, _06047_);
  or _86437_ (_36886_, _36885_, _36883_);
  and _86438_ (_36887_, _14657_, _07705_);
  or _86439_ (_36889_, _36665_, _06048_);
  or _86440_ (_36890_, _36889_, _36887_);
  and _86441_ (_36891_, _36890_, _01336_);
  and _86442_ (_36892_, _36891_, _36886_);
  or _86443_ (_36893_, _36892_, _36644_);
  and _86444_ (_43512_, _36893_, _42882_);
  nor _86445_ (_36894_, _01336_, _07369_);
  nor _86446_ (_36895_, _07705_, _07369_);
  nor _86447_ (_36896_, _13745_, _07353_);
  or _86448_ (_36897_, _36896_, _36895_);
  or _86449_ (_36899_, _36897_, _09827_);
  nor _86450_ (_36900_, _08355_, _07369_);
  and _86451_ (_36901_, _14681_, _08355_);
  or _86452_ (_36902_, _36901_, _36900_);
  and _86453_ (_36903_, _36902_, _06039_);
  and _86454_ (_36904_, _14672_, _07705_);
  or _86455_ (_36905_, _36904_, _36895_);
  or _86456_ (_36906_, _36905_, _06954_);
  and _86457_ (_36907_, _07705_, \oc8051_golden_model_1.ACC [3]);
  or _86458_ (_36908_, _36907_, _36895_);
  and _86459_ (_36910_, _36908_, _06938_);
  nor _86460_ (_36911_, _06938_, _07369_);
  or _86461_ (_36912_, _36911_, _06102_);
  or _86462_ (_36913_, _36912_, _36910_);
  and _86463_ (_36914_, _36913_, _06044_);
  and _86464_ (_36915_, _36914_, _36906_);
  and _86465_ (_36916_, _14683_, _08355_);
  or _86466_ (_36917_, _36916_, _36900_);
  and _86467_ (_36918_, _36917_, _06043_);
  or _86468_ (_36919_, _36918_, _06239_);
  or _86469_ (_36921_, _36919_, _36915_);
  or _86470_ (_36922_, _36897_, _06848_);
  and _86471_ (_36923_, _36922_, _36921_);
  or _86472_ (_36924_, _36923_, _06219_);
  or _86473_ (_36925_, _36908_, _06220_);
  and _86474_ (_36926_, _36925_, _06040_);
  and _86475_ (_36927_, _36926_, _36924_);
  or _86476_ (_36928_, _36927_, _36903_);
  and _86477_ (_36929_, _36928_, _06033_);
  and _86478_ (_36930_, _14709_, _08355_);
  or _86479_ (_36932_, _36930_, _36900_);
  and _86480_ (_36933_, _36932_, _06032_);
  or _86481_ (_36934_, _36933_, _36929_);
  and _86482_ (_36935_, _36934_, _06027_);
  and _86483_ (_36936_, _14724_, _08355_);
  or _86484_ (_36937_, _36936_, _36900_);
  and _86485_ (_36938_, _36937_, _06026_);
  or _86486_ (_36939_, _36938_, _09815_);
  or _86487_ (_36940_, _36939_, _36935_);
  and _86488_ (_36941_, _36940_, _36899_);
  or _86489_ (_36943_, _36941_, _07011_);
  and _86490_ (_36944_, _09181_, _07705_);
  or _86491_ (_36945_, _36895_, _07012_);
  or _86492_ (_36946_, _36945_, _36944_);
  and _86493_ (_36947_, _36946_, _36943_);
  or _86494_ (_36948_, _36947_, _09833_);
  and _86495_ (_36949_, _14778_, _07705_);
  or _86496_ (_36950_, _36949_, _36895_);
  or _86497_ (_36951_, _36950_, _05669_);
  and _86498_ (_36952_, _36951_, _06020_);
  and _86499_ (_36954_, _36952_, _36948_);
  and _86500_ (_36955_, _07705_, _08662_);
  or _86501_ (_36956_, _36955_, _36895_);
  and _86502_ (_36957_, _36956_, _06019_);
  or _86503_ (_36958_, _36957_, _06112_);
  or _86504_ (_36959_, _36958_, _36954_);
  and _86505_ (_36960_, _14793_, _07705_);
  or _86506_ (_36961_, _36960_, _36895_);
  or _86507_ (_36962_, _36961_, _08751_);
  and _86508_ (_36963_, _36962_, _08756_);
  and _86509_ (_36965_, _36963_, _36959_);
  and _86510_ (_36966_, _12299_, _07705_);
  or _86511_ (_36967_, _36966_, _36895_);
  and _86512_ (_36968_, _36967_, _06284_);
  or _86513_ (_36969_, _36968_, _36965_);
  and _86514_ (_36970_, _36969_, _07032_);
  or _86515_ (_36971_, _36895_, _08029_);
  and _86516_ (_36972_, _36956_, _06108_);
  and _86517_ (_36973_, _36972_, _36971_);
  or _86518_ (_36974_, _36973_, _36970_);
  and _86519_ (_36976_, _36974_, _06278_);
  and _86520_ (_36977_, _36908_, _06277_);
  and _86521_ (_36978_, _36977_, _36971_);
  or _86522_ (_36979_, _36978_, _06130_);
  or _86523_ (_36980_, _36979_, _36976_);
  and _86524_ (_36981_, _14792_, _07705_);
  or _86525_ (_36982_, _36895_, _08777_);
  or _86526_ (_36983_, _36982_, _36981_);
  and _86527_ (_36984_, _36983_, _08782_);
  and _86528_ (_36985_, _36984_, _36980_);
  nor _86529_ (_36987_, _10988_, _13745_);
  or _86530_ (_36988_, _36987_, _36895_);
  and _86531_ (_36989_, _36988_, _06292_);
  or _86532_ (_36990_, _36989_, _06316_);
  or _86533_ (_36991_, _36990_, _36985_);
  or _86534_ (_36992_, _36905_, _06718_);
  and _86535_ (_36993_, _36992_, _05653_);
  and _86536_ (_36994_, _36993_, _36991_);
  and _86537_ (_36995_, _36902_, _05652_);
  or _86538_ (_36996_, _36995_, _06047_);
  or _86539_ (_36998_, _36996_, _36994_);
  and _86540_ (_36999_, _14849_, _07705_);
  or _86541_ (_37000_, _36895_, _06048_);
  or _86542_ (_37001_, _37000_, _36999_);
  and _86543_ (_37002_, _37001_, _01336_);
  and _86544_ (_37003_, _37002_, _36998_);
  or _86545_ (_37004_, _37003_, _36894_);
  and _86546_ (_43513_, _37004_, _42882_);
  not _86547_ (_37005_, \oc8051_golden_model_1.PSW [4]);
  nor _86548_ (_37006_, _01336_, _37005_);
  nor _86549_ (_37008_, _07705_, _37005_);
  nor _86550_ (_37009_, _08270_, _13745_);
  or _86551_ (_37010_, _37009_, _37008_);
  or _86552_ (_37011_, _37010_, _09827_);
  nor _86553_ (_37012_, _08355_, _37005_);
  and _86554_ (_37013_, _14882_, _08355_);
  or _86555_ (_37014_, _37013_, _37012_);
  and _86556_ (_37015_, _37014_, _06039_);
  and _86557_ (_37016_, _14887_, _07705_);
  or _86558_ (_37017_, _37016_, _37008_);
  or _86559_ (_37019_, _37017_, _06954_);
  and _86560_ (_37020_, _07705_, \oc8051_golden_model_1.ACC [4]);
  or _86561_ (_37021_, _37020_, _37008_);
  and _86562_ (_37022_, _37021_, _06938_);
  nor _86563_ (_37023_, _06938_, _37005_);
  or _86564_ (_37024_, _37023_, _06102_);
  or _86565_ (_37025_, _37024_, _37022_);
  and _86566_ (_37026_, _37025_, _06044_);
  and _86567_ (_37027_, _37026_, _37019_);
  and _86568_ (_37028_, _14878_, _08355_);
  or _86569_ (_37030_, _37028_, _37012_);
  and _86570_ (_37031_, _37030_, _06043_);
  or _86571_ (_37032_, _37031_, _06239_);
  or _86572_ (_37033_, _37032_, _37027_);
  or _86573_ (_37034_, _37010_, _06848_);
  and _86574_ (_37035_, _37034_, _37033_);
  or _86575_ (_37036_, _37035_, _06219_);
  or _86576_ (_37037_, _37021_, _06220_);
  and _86577_ (_37038_, _37037_, _06040_);
  and _86578_ (_37039_, _37038_, _37036_);
  or _86579_ (_37041_, _37039_, _37015_);
  and _86580_ (_37042_, _37041_, _06033_);
  and _86581_ (_37043_, _14915_, _08355_);
  or _86582_ (_37044_, _37043_, _37012_);
  and _86583_ (_37045_, _37044_, _06032_);
  or _86584_ (_37046_, _37045_, _37042_);
  and _86585_ (_37047_, _37046_, _06027_);
  or _86586_ (_37048_, _37012_, _14879_);
  and _86587_ (_37049_, _37048_, _06026_);
  and _86588_ (_37050_, _37049_, _37030_);
  or _86589_ (_37052_, _37050_, _09815_);
  or _86590_ (_37053_, _37052_, _37047_);
  and _86591_ (_37054_, _37053_, _37011_);
  or _86592_ (_37055_, _37054_, _07011_);
  and _86593_ (_37056_, _09180_, _07705_);
  or _86594_ (_37057_, _37008_, _07012_);
  or _86595_ (_37058_, _37057_, _37056_);
  and _86596_ (_37059_, _37058_, _37055_);
  or _86597_ (_37060_, _37059_, _09833_);
  and _86598_ (_37061_, _14983_, _07705_);
  or _86599_ (_37063_, _37061_, _37008_);
  or _86600_ (_37064_, _37063_, _05669_);
  and _86601_ (_37065_, _37064_, _06020_);
  and _86602_ (_37066_, _37065_, _37060_);
  and _86603_ (_37067_, _08665_, _07705_);
  or _86604_ (_37068_, _37067_, _37008_);
  and _86605_ (_37069_, _37068_, _06019_);
  or _86606_ (_37070_, _37069_, _06112_);
  or _86607_ (_37071_, _37070_, _37066_);
  and _86608_ (_37072_, _14876_, _07705_);
  or _86609_ (_37074_, _37008_, _08751_);
  or _86610_ (_37075_, _37074_, _37072_);
  and _86611_ (_37076_, _37075_, _08756_);
  and _86612_ (_37077_, _37076_, _37071_);
  and _86613_ (_37078_, _10986_, _07705_);
  or _86614_ (_37079_, _37078_, _37008_);
  and _86615_ (_37080_, _37079_, _06284_);
  or _86616_ (_37081_, _37080_, _37077_);
  and _86617_ (_37082_, _37081_, _07032_);
  or _86618_ (_37083_, _37008_, _08273_);
  and _86619_ (_37085_, _37068_, _06108_);
  and _86620_ (_37086_, _37085_, _37083_);
  or _86621_ (_37087_, _37086_, _37082_);
  and _86622_ (_37088_, _37087_, _06278_);
  and _86623_ (_37089_, _37021_, _06277_);
  and _86624_ (_37090_, _37089_, _37083_);
  or _86625_ (_37091_, _37090_, _06130_);
  or _86626_ (_37092_, _37091_, _37088_);
  and _86627_ (_37093_, _14873_, _07705_);
  or _86628_ (_37094_, _37008_, _08777_);
  or _86629_ (_37096_, _37094_, _37093_);
  and _86630_ (_37097_, _37096_, _08782_);
  and _86631_ (_37098_, _37097_, _37092_);
  nor _86632_ (_37099_, _10985_, _13745_);
  or _86633_ (_37100_, _37099_, _37008_);
  and _86634_ (_37101_, _37100_, _06292_);
  or _86635_ (_37102_, _37101_, _06316_);
  or _86636_ (_37103_, _37102_, _37098_);
  or _86637_ (_37104_, _37017_, _06718_);
  and _86638_ (_37105_, _37104_, _05653_);
  and _86639_ (_37107_, _37105_, _37103_);
  and _86640_ (_37108_, _37014_, _05652_);
  or _86641_ (_37109_, _37108_, _06047_);
  or _86642_ (_37110_, _37109_, _37107_);
  and _86643_ (_37111_, _15055_, _07705_);
  or _86644_ (_37112_, _37008_, _06048_);
  or _86645_ (_37113_, _37112_, _37111_);
  and _86646_ (_37114_, _37113_, _01336_);
  and _86647_ (_37115_, _37114_, _37110_);
  or _86648_ (_37116_, _37115_, _37006_);
  and _86649_ (_43514_, _37116_, _42882_);
  not _86650_ (_37118_, \oc8051_golden_model_1.PSW [5]);
  nor _86651_ (_37119_, _01336_, _37118_);
  nor _86652_ (_37120_, _07705_, _37118_);
  nor _86653_ (_37121_, _07977_, _13745_);
  or _86654_ (_37122_, _37121_, _37120_);
  or _86655_ (_37123_, _37122_, _09827_);
  and _86656_ (_37124_, _15093_, _07705_);
  or _86657_ (_37125_, _37124_, _37120_);
  or _86658_ (_37126_, _37125_, _06954_);
  and _86659_ (_37128_, _07705_, \oc8051_golden_model_1.ACC [5]);
  or _86660_ (_37129_, _37128_, _37120_);
  and _86661_ (_37130_, _37129_, _06938_);
  nor _86662_ (_37131_, _06938_, _37118_);
  or _86663_ (_37132_, _37131_, _06102_);
  or _86664_ (_37133_, _37132_, _37130_);
  and _86665_ (_37134_, _37133_, _06044_);
  and _86666_ (_37135_, _37134_, _37126_);
  nor _86667_ (_37136_, _08355_, _37118_);
  and _86668_ (_37137_, _15073_, _08355_);
  or _86669_ (_37139_, _37137_, _37136_);
  and _86670_ (_37140_, _37139_, _06043_);
  or _86671_ (_37141_, _37140_, _06239_);
  or _86672_ (_37142_, _37141_, _37135_);
  or _86673_ (_37143_, _37122_, _06848_);
  and _86674_ (_37144_, _37143_, _37142_);
  or _86675_ (_37145_, _37144_, _06219_);
  or _86676_ (_37146_, _37129_, _06220_);
  and _86677_ (_37147_, _37146_, _06040_);
  and _86678_ (_37148_, _37147_, _37145_);
  and _86679_ (_37150_, _15077_, _08355_);
  or _86680_ (_37151_, _37150_, _37136_);
  and _86681_ (_37152_, _37151_, _06039_);
  or _86682_ (_37153_, _37152_, _06032_);
  or _86683_ (_37154_, _37153_, _37148_);
  or _86684_ (_37155_, _37136_, _15110_);
  and _86685_ (_37156_, _37155_, _37139_);
  or _86686_ (_37157_, _37156_, _06033_);
  and _86687_ (_37158_, _37157_, _06027_);
  and _86688_ (_37159_, _37158_, _37154_);
  or _86689_ (_37161_, _37136_, _15074_);
  and _86690_ (_37162_, _37161_, _06026_);
  and _86691_ (_37163_, _37162_, _37139_);
  or _86692_ (_37164_, _37163_, _09815_);
  or _86693_ (_37165_, _37164_, _37159_);
  and _86694_ (_37166_, _37165_, _37123_);
  or _86695_ (_37167_, _37166_, _07011_);
  and _86696_ (_37168_, _09179_, _07705_);
  or _86697_ (_37169_, _37120_, _07012_);
  or _86698_ (_37170_, _37169_, _37168_);
  and _86699_ (_37172_, _37170_, _05669_);
  and _86700_ (_37173_, _37172_, _37167_);
  and _86701_ (_37174_, _15179_, _07705_);
  or _86702_ (_37175_, _37174_, _37120_);
  and _86703_ (_37176_, _37175_, _09833_);
  or _86704_ (_37177_, _37176_, _06019_);
  or _86705_ (_37178_, _37177_, _37173_);
  and _86706_ (_37179_, _08652_, _07705_);
  or _86707_ (_37180_, _37179_, _37120_);
  or _86708_ (_37181_, _37180_, _06020_);
  and _86709_ (_37183_, _37181_, _37178_);
  or _86710_ (_37184_, _37183_, _06112_);
  and _86711_ (_37185_, _15195_, _07705_);
  or _86712_ (_37186_, _37185_, _37120_);
  or _86713_ (_37187_, _37186_, _08751_);
  and _86714_ (_37188_, _37187_, _08756_);
  and _86715_ (_37189_, _37188_, _37184_);
  and _86716_ (_37190_, _12306_, _07705_);
  or _86717_ (_37191_, _37190_, _37120_);
  and _86718_ (_37192_, _37191_, _06284_);
  or _86719_ (_37194_, _37192_, _37189_);
  and _86720_ (_37195_, _37194_, _07032_);
  or _86721_ (_37196_, _37120_, _07980_);
  and _86722_ (_37197_, _37180_, _06108_);
  and _86723_ (_37198_, _37197_, _37196_);
  or _86724_ (_37199_, _37198_, _37195_);
  and _86725_ (_37200_, _37199_, _06278_);
  and _86726_ (_37201_, _37129_, _06277_);
  and _86727_ (_37202_, _37201_, _37196_);
  or _86728_ (_37203_, _37202_, _06130_);
  or _86729_ (_37205_, _37203_, _37200_);
  and _86730_ (_37206_, _15194_, _07705_);
  or _86731_ (_37207_, _37120_, _08777_);
  or _86732_ (_37208_, _37207_, _37206_);
  and _86733_ (_37209_, _37208_, _08782_);
  and _86734_ (_37210_, _37209_, _37205_);
  nor _86735_ (_37211_, _10982_, _13745_);
  or _86736_ (_37212_, _37211_, _37120_);
  and _86737_ (_37213_, _37212_, _06292_);
  or _86738_ (_37214_, _37213_, _06316_);
  or _86739_ (_37216_, _37214_, _37210_);
  or _86740_ (_37217_, _37125_, _06718_);
  and _86741_ (_37218_, _37217_, _05653_);
  and _86742_ (_37219_, _37218_, _37216_);
  and _86743_ (_37220_, _37151_, _05652_);
  or _86744_ (_37221_, _37220_, _06047_);
  or _86745_ (_37222_, _37221_, _37219_);
  and _86746_ (_37223_, _15253_, _07705_);
  or _86747_ (_37224_, _37120_, _06048_);
  or _86748_ (_37225_, _37224_, _37223_);
  and _86749_ (_37227_, _37225_, _01336_);
  and _86750_ (_37228_, _37227_, _37222_);
  or _86751_ (_37229_, _37228_, _37119_);
  and _86752_ (_43515_, _37229_, _42882_);
  nor _86753_ (_37230_, _01336_, _17846_);
  or _86754_ (_37231_, _10871_, _10567_);
  and _86755_ (_37232_, _37231_, _10824_);
  or _86756_ (_37233_, _10796_, _10512_);
  or _86757_ (_37234_, _37233_, _10811_);
  and _86758_ (_37235_, _06229_, _05731_);
  and _86759_ (_37237_, _06136_, _05731_);
  and _86760_ (_37238_, _07005_, _05731_);
  or _86761_ (_37239_, _10293_, _10237_);
  and _86762_ (_37240_, _37239_, _37238_);
  and _86763_ (_37241_, _15396_, _07705_);
  nor _86764_ (_37242_, _07705_, _17846_);
  or _86765_ (_37243_, _37242_, _08777_);
  or _86766_ (_37244_, _37243_, _37241_);
  nor _86767_ (_37245_, _07883_, _13745_);
  or _86768_ (_37246_, _37245_, _37242_);
  or _86769_ (_37248_, _37246_, _09827_);
  and _86770_ (_37249_, _15293_, _07705_);
  or _86771_ (_37250_, _37249_, _37242_);
  or _86772_ (_37251_, _37250_, _06954_);
  and _86773_ (_37252_, _07705_, \oc8051_golden_model_1.ACC [6]);
  or _86774_ (_37253_, _37252_, _37242_);
  and _86775_ (_37254_, _37253_, _06938_);
  nor _86776_ (_37255_, _06938_, _17846_);
  or _86777_ (_37256_, _37255_, _06102_);
  or _86778_ (_37257_, _37256_, _37254_);
  and _86779_ (_37259_, _37257_, _06044_);
  and _86780_ (_37260_, _37259_, _37251_);
  nor _86781_ (_37261_, _08355_, _17846_);
  and _86782_ (_37262_, _15280_, _08355_);
  or _86783_ (_37263_, _37262_, _37261_);
  and _86784_ (_37264_, _37263_, _06043_);
  or _86785_ (_37265_, _37264_, _06239_);
  or _86786_ (_37266_, _37265_, _37260_);
  or _86787_ (_37267_, _37246_, _06848_);
  and _86788_ (_37268_, _37267_, _37266_);
  or _86789_ (_37270_, _37268_, _06219_);
  or _86790_ (_37271_, _37253_, _06220_);
  and _86791_ (_37272_, _37271_, _06040_);
  and _86792_ (_37273_, _37272_, _37270_);
  and _86793_ (_37274_, _15278_, _08355_);
  or _86794_ (_37275_, _37274_, _37261_);
  and _86795_ (_37276_, _37275_, _06039_);
  or _86796_ (_37277_, _37276_, _06032_);
  or _86797_ (_37278_, _37277_, _37273_);
  or _86798_ (_37279_, _37261_, _15310_);
  and _86799_ (_37281_, _37279_, _37263_);
  or _86800_ (_37282_, _37281_, _06033_);
  and _86801_ (_37283_, _37282_, _10469_);
  and _86802_ (_37284_, _37283_, _37278_);
  or _86803_ (_37285_, _12361_, _10237_);
  or _86804_ (_37286_, _37285_, _10483_);
  and _86805_ (_37287_, _37286_, _12368_);
  or _86806_ (_37288_, _37287_, _37284_);
  or _86807_ (_37289_, _10512_, _13935_);
  or _86808_ (_37290_, _37289_, _10549_);
  and _86809_ (_37292_, _37290_, _37288_);
  or _86810_ (_37293_, _37292_, _12367_);
  or _86811_ (_37294_, _10311_, _06267_);
  or _86812_ (_37295_, _37294_, _10360_);
  or _86813_ (_37296_, _10567_, _10307_);
  or _86814_ (_37297_, _37296_, _10621_);
  and _86815_ (_37298_, _37297_, _06027_);
  and _86816_ (_37299_, _37298_, _37295_);
  and _86817_ (_37300_, _37299_, _37293_);
  or _86818_ (_37301_, _37261_, _15326_);
  and _86819_ (_37303_, _37301_, _06026_);
  and _86820_ (_37304_, _37303_, _37263_);
  or _86821_ (_37305_, _37304_, _09815_);
  or _86822_ (_37306_, _37305_, _37300_);
  and _86823_ (_37307_, _37306_, _37248_);
  or _86824_ (_37308_, _37307_, _07011_);
  and _86825_ (_37309_, _09178_, _07705_);
  or _86826_ (_37310_, _37242_, _07012_);
  or _86827_ (_37311_, _37310_, _37309_);
  and _86828_ (_37312_, _37311_, _05669_);
  and _86829_ (_37314_, _37312_, _37308_);
  and _86830_ (_37315_, _15382_, _07705_);
  or _86831_ (_37316_, _37315_, _37242_);
  and _86832_ (_37317_, _37316_, _09833_);
  or _86833_ (_37318_, _37317_, _06019_);
  or _86834_ (_37319_, _37318_, _37314_);
  and _86835_ (_37320_, _15389_, _07705_);
  or _86836_ (_37321_, _37320_, _37242_);
  or _86837_ (_37322_, _37321_, _06020_);
  and _86838_ (_37323_, _37322_, _37319_);
  or _86839_ (_37325_, _37323_, _06112_);
  and _86840_ (_37326_, _15399_, _07705_);
  or _86841_ (_37327_, _37326_, _37242_);
  or _86842_ (_37328_, _37327_, _08751_);
  and _86843_ (_37329_, _37328_, _08756_);
  and _86844_ (_37330_, _37329_, _37325_);
  and _86845_ (_37331_, _10980_, _07705_);
  or _86846_ (_37332_, _37331_, _37242_);
  and _86847_ (_37333_, _37332_, _06284_);
  or _86848_ (_37334_, _37333_, _37330_);
  and _86849_ (_37336_, _37334_, _07032_);
  or _86850_ (_37337_, _37242_, _07886_);
  and _86851_ (_37338_, _37321_, _06108_);
  and _86852_ (_37339_, _37338_, _37337_);
  or _86853_ (_37340_, _37339_, _37336_);
  and _86854_ (_37341_, _37340_, _06278_);
  and _86855_ (_37342_, _37253_, _06277_);
  and _86856_ (_37343_, _37342_, _37337_);
  or _86857_ (_37344_, _37343_, _06130_);
  or _86858_ (_37345_, _37344_, _37341_);
  and _86859_ (_37347_, _37345_, _37244_);
  or _86860_ (_37348_, _37347_, _06292_);
  nor _86861_ (_37349_, _10979_, _13745_);
  or _86862_ (_37350_, _37349_, _37242_);
  nor _86863_ (_37351_, _37350_, _08782_);
  nor _86864_ (_37352_, _37351_, _37238_);
  and _86865_ (_37353_, _37352_, _37348_);
  nor _86866_ (_37354_, _37353_, _37240_);
  nor _86867_ (_37355_, _37354_, _37237_);
  and _86868_ (_37356_, _37239_, _37237_);
  nor _86869_ (_37358_, _37356_, _37355_);
  nor _86870_ (_37359_, _37358_, _37235_);
  and _86871_ (_37360_, _06227_, _05731_);
  and _86872_ (_37361_, _37239_, _37235_);
  or _86873_ (_37362_, _37361_, _37360_);
  or _86874_ (_37363_, _37362_, _37359_);
  and _86875_ (_37364_, _07002_, _05731_);
  not _86876_ (_37365_, _37360_);
  nor _86877_ (_37366_, _37239_, _37365_);
  nor _86878_ (_37367_, _37366_, _37364_);
  and _86879_ (_37369_, _37367_, _37363_);
  and _86880_ (_37370_, _37239_, _37364_);
  or _86881_ (_37371_, _37370_, _10794_);
  or _86882_ (_37372_, _37371_, _37369_);
  and _86883_ (_37373_, _37372_, _37234_);
  or _86884_ (_37374_, _37373_, _06288_);
  or _86885_ (_37375_, _10311_, _06289_);
  or _86886_ (_37376_, _37375_, _10841_);
  and _86887_ (_37377_, _37376_, _10856_);
  and _86888_ (_37378_, _37377_, _37374_);
  or _86889_ (_37380_, _37378_, _37232_);
  and _86890_ (_37381_, _37380_, _10890_);
  and _86891_ (_37382_, _10920_, _16956_);
  or _86892_ (_37383_, _37382_, _10932_);
  or _86893_ (_37384_, _37383_, _37381_);
  or _86894_ (_37385_, _10961_, _10934_);
  and _86895_ (_37386_, _37385_, _06052_);
  and _86896_ (_37387_, _37386_, _37384_);
  or _86897_ (_37388_, _11002_, _10974_);
  and _86898_ (_37389_, _37388_, _10976_);
  or _86899_ (_37391_, _37389_, _37387_);
  or _86900_ (_37392_, _11042_, _11050_);
  and _86901_ (_37393_, _37392_, _37391_);
  or _86902_ (_37394_, _37393_, _06316_);
  or _86903_ (_37395_, _37250_, _06718_);
  and _86904_ (_37396_, _37395_, _05653_);
  and _86905_ (_37397_, _37396_, _37394_);
  and _86906_ (_37398_, _37275_, _05652_);
  or _86907_ (_37399_, _37398_, _06047_);
  or _86908_ (_37400_, _37399_, _37397_);
  and _86909_ (_37402_, _15451_, _07705_);
  or _86910_ (_37403_, _37242_, _06048_);
  or _86911_ (_37404_, _37403_, _37402_);
  and _86912_ (_37405_, _37404_, _01336_);
  and _86913_ (_37406_, _37405_, _37400_);
  or _86914_ (_37407_, _37406_, _37230_);
  and _86915_ (_43516_, _37407_, _42882_);
  and _86916_ (_37408_, _05750_, op0_cnst);
  or _86917_ (_00001_, _37408_, rst);
  and _86918_ (_37409_, inst_finished_r, op0_cnst);
  nor _86919_ (_37411_, word_in[3], word_in[2]);
  not _86920_ (_37412_, _37411_);
  not _86921_ (_37413_, word_in[1]);
  and _86922_ (_37414_, _37413_, word_in[0]);
  and _86923_ (_37415_, _37414_, \oc8051_golden_model_1.IRAM[1] [1]);
  nor _86924_ (_37416_, _37413_, word_in[0]);
  and _86925_ (_37417_, _37416_, \oc8051_golden_model_1.IRAM[2] [1]);
  nor _86926_ (_37418_, _37417_, _37415_);
  nor _86927_ (_37419_, word_in[1], word_in[0]);
  and _86928_ (_37420_, _37419_, \oc8051_golden_model_1.IRAM[0] [1]);
  and _86929_ (_37422_, word_in[1], word_in[0]);
  and _86930_ (_37423_, _37422_, \oc8051_golden_model_1.IRAM[3] [1]);
  nor _86931_ (_37424_, _37423_, _37420_);
  and _86932_ (_37425_, _37424_, _37418_);
  nor _86933_ (_37426_, _37425_, _37412_);
  and _86934_ (_37427_, word_in[3], word_in[2]);
  not _86935_ (_37428_, _37427_);
  and _86936_ (_37429_, _37414_, \oc8051_golden_model_1.IRAM[13] [1]);
  and _86937_ (_37430_, _37416_, \oc8051_golden_model_1.IRAM[14] [1]);
  nor _86938_ (_37431_, _37430_, _37429_);
  and _86939_ (_37433_, _37419_, \oc8051_golden_model_1.IRAM[12] [1]);
  and _86940_ (_37434_, _37422_, \oc8051_golden_model_1.IRAM[15] [1]);
  nor _86941_ (_37435_, _37434_, _37433_);
  and _86942_ (_37436_, _37435_, _37431_);
  nor _86943_ (_37437_, _37436_, _37428_);
  nor _86944_ (_37438_, _37437_, _37426_);
  not _86945_ (_37439_, word_in[3]);
  and _86946_ (_37440_, _37439_, word_in[2]);
  not _86947_ (_37441_, _37440_);
  and _86948_ (_37442_, _37414_, \oc8051_golden_model_1.IRAM[5] [1]);
  and _86949_ (_37444_, _37416_, \oc8051_golden_model_1.IRAM[6] [1]);
  nor _86950_ (_37445_, _37444_, _37442_);
  and _86951_ (_37446_, _37419_, \oc8051_golden_model_1.IRAM[4] [1]);
  and _86952_ (_37447_, _37422_, \oc8051_golden_model_1.IRAM[7] [1]);
  nor _86953_ (_37448_, _37447_, _37446_);
  and _86954_ (_37449_, _37448_, _37445_);
  nor _86955_ (_37450_, _37449_, _37441_);
  nor _86956_ (_37451_, _37439_, word_in[2]);
  not _86957_ (_37452_, _37451_);
  and _86958_ (_37453_, _37414_, \oc8051_golden_model_1.IRAM[9] [1]);
  and _86959_ (_37455_, _37416_, \oc8051_golden_model_1.IRAM[10] [1]);
  nor _86960_ (_37456_, _37455_, _37453_);
  and _86961_ (_37457_, _37419_, \oc8051_golden_model_1.IRAM[8] [1]);
  and _86962_ (_37458_, _37422_, \oc8051_golden_model_1.IRAM[11] [1]);
  nor _86963_ (_37459_, _37458_, _37457_);
  and _86964_ (_37460_, _37459_, _37456_);
  nor _86965_ (_37461_, _37460_, _37452_);
  nor _86966_ (_37462_, _37461_, _37450_);
  and _86967_ (_37463_, _37462_, _37438_);
  and _86968_ (_37464_, _37440_, _37422_);
  and _86969_ (_37466_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  and _86970_ (_37467_, _37440_, _37416_);
  and _86971_ (_37468_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nor _86972_ (_37469_, _37468_, _37466_);
  and _86973_ (_37470_, _37427_, _37414_);
  and _86974_ (_37471_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  and _86975_ (_37472_, _37427_, _37419_);
  and _86976_ (_37473_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor _86977_ (_37474_, _37473_, _37471_);
  and _86978_ (_37475_, _37474_, _37469_);
  and _86979_ (_37477_, _37416_, _37411_);
  and _86980_ (_37478_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  and _86981_ (_37479_, _37414_, _37411_);
  and _86982_ (_37480_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor _86983_ (_37481_, _37480_, _37478_);
  and _86984_ (_37482_, _37427_, _37416_);
  and _86985_ (_37483_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  and _86986_ (_37484_, _37451_, _37419_);
  and _86987_ (_37485_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nor _86988_ (_37486_, _37485_, _37483_);
  and _86989_ (_37488_, _37486_, _37481_);
  and _86990_ (_37489_, _37488_, _37475_);
  and _86991_ (_37490_, _37451_, _37414_);
  and _86992_ (_37491_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  and _86993_ (_37492_, _37419_, _37411_);
  and _86994_ (_37493_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor _86995_ (_37494_, _37493_, _37491_);
  and _86996_ (_37495_, _37451_, _37416_);
  and _86997_ (_37496_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  and _86998_ (_37497_, _37440_, _37414_);
  and _86999_ (_37499_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor _87000_ (_37500_, _37499_, _37496_);
  and _87001_ (_37501_, _37500_, _37494_);
  and _87002_ (_37502_, _37427_, _37422_);
  and _87003_ (_37503_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  and _87004_ (_37504_, _37440_, _37419_);
  and _87005_ (_37505_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor _87006_ (_37506_, _37505_, _37503_);
  and _87007_ (_37507_, _37451_, _37422_);
  and _87008_ (_37508_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  and _87009_ (_37510_, _37422_, _37411_);
  and _87010_ (_37511_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor _87011_ (_37512_, _37511_, _37508_);
  and _87012_ (_37513_, _37512_, _37506_);
  and _87013_ (_37514_, _37513_, _37501_);
  and _87014_ (_37515_, _37514_, _37489_);
  nand _87015_ (_37516_, _37515_, _37463_);
  or _87016_ (_37517_, _37515_, _37463_);
  and _87017_ (_37518_, _37517_, _37516_);
  and _87018_ (_37519_, _37414_, \oc8051_golden_model_1.IRAM[1] [0]);
  and _87019_ (_37521_, _37416_, \oc8051_golden_model_1.IRAM[2] [0]);
  nor _87020_ (_37522_, _37521_, _37519_);
  and _87021_ (_37523_, _37419_, \oc8051_golden_model_1.IRAM[0] [0]);
  and _87022_ (_37524_, _37422_, \oc8051_golden_model_1.IRAM[3] [0]);
  nor _87023_ (_37525_, _37524_, _37523_);
  and _87024_ (_37526_, _37525_, _37522_);
  nor _87025_ (_37527_, _37526_, _37412_);
  and _87026_ (_37528_, _37414_, \oc8051_golden_model_1.IRAM[9] [0]);
  and _87027_ (_37529_, _37416_, \oc8051_golden_model_1.IRAM[10] [0]);
  nor _87028_ (_37530_, _37529_, _37528_);
  and _87029_ (_37532_, _37419_, \oc8051_golden_model_1.IRAM[8] [0]);
  and _87030_ (_37533_, _37422_, \oc8051_golden_model_1.IRAM[11] [0]);
  nor _87031_ (_37534_, _37533_, _37532_);
  and _87032_ (_37535_, _37534_, _37530_);
  nor _87033_ (_37536_, _37535_, _37452_);
  nor _87034_ (_37537_, _37536_, _37527_);
  and _87035_ (_37538_, _37414_, \oc8051_golden_model_1.IRAM[5] [0]);
  and _87036_ (_37539_, _37416_, \oc8051_golden_model_1.IRAM[6] [0]);
  nor _87037_ (_37540_, _37539_, _37538_);
  and _87038_ (_37541_, _37419_, \oc8051_golden_model_1.IRAM[4] [0]);
  and _87039_ (_37543_, _37422_, \oc8051_golden_model_1.IRAM[7] [0]);
  nor _87040_ (_37544_, _37543_, _37541_);
  and _87041_ (_37545_, _37544_, _37540_);
  nor _87042_ (_37546_, _37545_, _37441_);
  and _87043_ (_37547_, _37414_, \oc8051_golden_model_1.IRAM[13] [0]);
  and _87044_ (_37548_, _37416_, \oc8051_golden_model_1.IRAM[14] [0]);
  nor _87045_ (_37549_, _37548_, _37547_);
  and _87046_ (_37550_, _37419_, \oc8051_golden_model_1.IRAM[12] [0]);
  and _87047_ (_37551_, _37422_, \oc8051_golden_model_1.IRAM[15] [0]);
  nor _87048_ (_37552_, _37551_, _37550_);
  and _87049_ (_37554_, _37552_, _37549_);
  nor _87050_ (_37555_, _37554_, _37428_);
  nor _87051_ (_37556_, _37555_, _37546_);
  and _87052_ (_37557_, _37556_, _37537_);
  and _87053_ (_37558_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  and _87054_ (_37559_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor _87055_ (_37560_, _37559_, _37558_);
  and _87056_ (_37561_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  and _87057_ (_37562_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor _87058_ (_37563_, _37562_, _37561_);
  and _87059_ (_37565_, _37563_, _37560_);
  and _87060_ (_37566_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  and _87061_ (_37567_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor _87062_ (_37568_, _37567_, _37566_);
  and _87063_ (_37569_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  and _87064_ (_37570_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor _87065_ (_37571_, _37570_, _37569_);
  and _87066_ (_37572_, _37571_, _37568_);
  and _87067_ (_37573_, _37572_, _37565_);
  and _87068_ (_37574_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  and _87069_ (_37576_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor _87070_ (_37577_, _37576_, _37574_);
  and _87071_ (_37578_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  and _87072_ (_37579_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor _87073_ (_37580_, _37579_, _37578_);
  and _87074_ (_37581_, _37580_, _37577_);
  and _87075_ (_37582_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  and _87076_ (_37583_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor _87077_ (_37584_, _37583_, _37582_);
  and _87078_ (_37585_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  and _87079_ (_37587_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor _87080_ (_37588_, _37587_, _37585_);
  and _87081_ (_37589_, _37588_, _37584_);
  and _87082_ (_37590_, _37589_, _37581_);
  and _87083_ (_37591_, _37590_, _37573_);
  not _87084_ (_37592_, _37591_);
  nor _87085_ (_37593_, _37592_, _37557_);
  and _87086_ (_37594_, _37592_, _37557_);
  or _87087_ (_37595_, _37594_, _37593_);
  or _87088_ (_37596_, _37595_, _37518_);
  and _87089_ (_37598_, _37414_, \oc8051_golden_model_1.IRAM[1] [3]);
  and _87090_ (_37599_, _37416_, \oc8051_golden_model_1.IRAM[2] [3]);
  nor _87091_ (_37600_, _37599_, _37598_);
  and _87092_ (_37601_, _37419_, \oc8051_golden_model_1.IRAM[0] [3]);
  and _87093_ (_37602_, _37422_, \oc8051_golden_model_1.IRAM[3] [3]);
  nor _87094_ (_37603_, _37602_, _37601_);
  and _87095_ (_37604_, _37603_, _37600_);
  nor _87096_ (_37605_, _37604_, _37412_);
  and _87097_ (_37606_, _37414_, \oc8051_golden_model_1.IRAM[13] [3]);
  and _87098_ (_37607_, _37416_, \oc8051_golden_model_1.IRAM[14] [3]);
  nor _87099_ (_37609_, _37607_, _37606_);
  and _87100_ (_37610_, _37419_, \oc8051_golden_model_1.IRAM[12] [3]);
  and _87101_ (_37611_, _37422_, \oc8051_golden_model_1.IRAM[15] [3]);
  nor _87102_ (_37612_, _37611_, _37610_);
  and _87103_ (_37613_, _37612_, _37609_);
  nor _87104_ (_37614_, _37613_, _37428_);
  nor _87105_ (_37615_, _37614_, _37605_);
  and _87106_ (_37616_, _37414_, \oc8051_golden_model_1.IRAM[5] [3]);
  and _87107_ (_37617_, _37416_, \oc8051_golden_model_1.IRAM[6] [3]);
  nor _87108_ (_37618_, _37617_, _37616_);
  and _87109_ (_37620_, _37419_, \oc8051_golden_model_1.IRAM[4] [3]);
  and _87110_ (_37621_, _37422_, \oc8051_golden_model_1.IRAM[7] [3]);
  nor _87111_ (_37622_, _37621_, _37620_);
  and _87112_ (_37623_, _37622_, _37618_);
  nor _87113_ (_37624_, _37623_, _37441_);
  and _87114_ (_37625_, _37414_, \oc8051_golden_model_1.IRAM[9] [3]);
  and _87115_ (_37626_, _37416_, \oc8051_golden_model_1.IRAM[10] [3]);
  nor _87116_ (_37627_, _37626_, _37625_);
  and _87117_ (_37628_, _37419_, \oc8051_golden_model_1.IRAM[8] [3]);
  and _87118_ (_37629_, _37422_, \oc8051_golden_model_1.IRAM[11] [3]);
  nor _87119_ (_37631_, _37629_, _37628_);
  and _87120_ (_37632_, _37631_, _37627_);
  nor _87121_ (_37633_, _37632_, _37452_);
  nor _87122_ (_37634_, _37633_, _37624_);
  and _87123_ (_37635_, _37634_, _37615_);
  and _87124_ (_37636_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  and _87125_ (_37637_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor _87126_ (_37638_, _37637_, _37636_);
  and _87127_ (_37639_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  and _87128_ (_37640_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor _87129_ (_37642_, _37640_, _37639_);
  and _87130_ (_37643_, _37642_, _37638_);
  and _87131_ (_37644_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  and _87132_ (_37645_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor _87133_ (_37646_, _37645_, _37644_);
  and _87134_ (_37647_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  and _87135_ (_37648_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor _87136_ (_37649_, _37648_, _37647_);
  and _87137_ (_37650_, _37649_, _37646_);
  and _87138_ (_37651_, _37650_, _37643_);
  and _87139_ (_37653_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  and _87140_ (_37654_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor _87141_ (_37655_, _37654_, _37653_);
  and _87142_ (_37656_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  and _87143_ (_37657_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nor _87144_ (_37658_, _37657_, _37656_);
  and _87145_ (_37659_, _37658_, _37655_);
  and _87146_ (_37660_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  and _87147_ (_37661_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor _87148_ (_37662_, _37661_, _37660_);
  and _87149_ (_37664_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  and _87150_ (_37665_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor _87151_ (_37666_, _37665_, _37664_);
  and _87152_ (_37667_, _37666_, _37662_);
  and _87153_ (_37668_, _37667_, _37659_);
  and _87154_ (_37669_, _37668_, _37651_);
  nand _87155_ (_37670_, _37669_, _37635_);
  or _87156_ (_37671_, _37669_, _37635_);
  and _87157_ (_37672_, _37671_, _37670_);
  and _87158_ (_37673_, _37414_, \oc8051_golden_model_1.IRAM[1] [2]);
  and _87159_ (_37675_, _37416_, \oc8051_golden_model_1.IRAM[2] [2]);
  nor _87160_ (_37676_, _37675_, _37673_);
  and _87161_ (_37677_, _37419_, \oc8051_golden_model_1.IRAM[0] [2]);
  and _87162_ (_37678_, _37422_, \oc8051_golden_model_1.IRAM[3] [2]);
  nor _87163_ (_37679_, _37678_, _37677_);
  and _87164_ (_37680_, _37679_, _37676_);
  nor _87165_ (_37681_, _37680_, _37412_);
  and _87166_ (_37682_, _37414_, \oc8051_golden_model_1.IRAM[9] [2]);
  and _87167_ (_37683_, _37416_, \oc8051_golden_model_1.IRAM[10] [2]);
  nor _87168_ (_37684_, _37683_, _37682_);
  and _87169_ (_37686_, _37419_, \oc8051_golden_model_1.IRAM[8] [2]);
  and _87170_ (_37687_, _37422_, \oc8051_golden_model_1.IRAM[11] [2]);
  nor _87171_ (_37688_, _37687_, _37686_);
  and _87172_ (_37689_, _37688_, _37684_);
  nor _87173_ (_37690_, _37689_, _37452_);
  nor _87174_ (_37691_, _37690_, _37681_);
  and _87175_ (_37692_, _37414_, \oc8051_golden_model_1.IRAM[5] [2]);
  and _87176_ (_37693_, _37416_, \oc8051_golden_model_1.IRAM[6] [2]);
  nor _87177_ (_37694_, _37693_, _37692_);
  and _87178_ (_37695_, _37419_, \oc8051_golden_model_1.IRAM[4] [2]);
  and _87179_ (_37697_, _37422_, \oc8051_golden_model_1.IRAM[7] [2]);
  nor _87180_ (_37698_, _37697_, _37695_);
  and _87181_ (_37699_, _37698_, _37694_);
  nor _87182_ (_37700_, _37699_, _37441_);
  and _87183_ (_37701_, _37414_, \oc8051_golden_model_1.IRAM[13] [2]);
  and _87184_ (_37702_, _37416_, \oc8051_golden_model_1.IRAM[14] [2]);
  nor _87185_ (_37703_, _37702_, _37701_);
  and _87186_ (_37704_, _37419_, \oc8051_golden_model_1.IRAM[12] [2]);
  and _87187_ (_37705_, _37422_, \oc8051_golden_model_1.IRAM[15] [2]);
  nor _87188_ (_37706_, _37705_, _37704_);
  and _87189_ (_37708_, _37706_, _37703_);
  nor _87190_ (_37709_, _37708_, _37428_);
  nor _87191_ (_37710_, _37709_, _37700_);
  and _87192_ (_37711_, _37710_, _37691_);
  and _87193_ (_37712_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  and _87194_ (_37713_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor _87195_ (_37714_, _37713_, _37712_);
  and _87196_ (_37715_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  and _87197_ (_37716_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor _87198_ (_37717_, _37716_, _37715_);
  and _87199_ (_37719_, _37717_, _37714_);
  and _87200_ (_37720_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  and _87201_ (_37721_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor _87202_ (_37722_, _37721_, _37720_);
  and _87203_ (_37723_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  and _87204_ (_37724_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor _87205_ (_37725_, _37724_, _37723_);
  and _87206_ (_37726_, _37725_, _37722_);
  and _87207_ (_37727_, _37726_, _37719_);
  and _87208_ (_37728_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  and _87209_ (_37730_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor _87210_ (_37731_, _37730_, _37728_);
  and _87211_ (_37732_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  and _87212_ (_37733_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor _87213_ (_37734_, _37733_, _37732_);
  and _87214_ (_37735_, _37734_, _37731_);
  and _87215_ (_37736_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  and _87216_ (_37737_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor _87217_ (_37738_, _37737_, _37736_);
  and _87218_ (_37739_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  and _87219_ (_37741_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor _87220_ (_37742_, _37741_, _37739_);
  and _87221_ (_37743_, _37742_, _37738_);
  and _87222_ (_37744_, _37743_, _37735_);
  and _87223_ (_37745_, _37744_, _37727_);
  nand _87224_ (_37746_, _37745_, _37711_);
  or _87225_ (_37747_, _37745_, _37711_);
  and _87226_ (_37748_, _37747_, _37746_);
  or _87227_ (_37749_, _37748_, _37672_);
  or _87228_ (_37750_, _37749_, _37596_);
  and _87229_ (_37752_, _37414_, \oc8051_golden_model_1.IRAM[5] [4]);
  and _87230_ (_37753_, _37416_, \oc8051_golden_model_1.IRAM[6] [4]);
  nor _87231_ (_37754_, _37753_, _37752_);
  and _87232_ (_37755_, _37419_, \oc8051_golden_model_1.IRAM[4] [4]);
  and _87233_ (_37756_, _37422_, \oc8051_golden_model_1.IRAM[7] [4]);
  nor _87234_ (_37757_, _37756_, _37755_);
  and _87235_ (_37758_, _37757_, _37754_);
  nor _87236_ (_37759_, _37758_, _37441_);
  and _87237_ (_37760_, _37414_, \oc8051_golden_model_1.IRAM[9] [4]);
  and _87238_ (_37761_, _37416_, \oc8051_golden_model_1.IRAM[10] [4]);
  nor _87239_ (_37763_, _37761_, _37760_);
  and _87240_ (_37764_, _37419_, \oc8051_golden_model_1.IRAM[8] [4]);
  and _87241_ (_37765_, _37422_, \oc8051_golden_model_1.IRAM[11] [4]);
  nor _87242_ (_37766_, _37765_, _37764_);
  and _87243_ (_37767_, _37766_, _37763_);
  nor _87244_ (_37768_, _37767_, _37452_);
  nor _87245_ (_37769_, _37768_, _37759_);
  and _87246_ (_37770_, _37414_, \oc8051_golden_model_1.IRAM[1] [4]);
  and _87247_ (_37771_, _37416_, \oc8051_golden_model_1.IRAM[2] [4]);
  nor _87248_ (_37772_, _37771_, _37770_);
  and _87249_ (_37774_, _37419_, \oc8051_golden_model_1.IRAM[0] [4]);
  and _87250_ (_37775_, _37422_, \oc8051_golden_model_1.IRAM[3] [4]);
  nor _87251_ (_37776_, _37775_, _37774_);
  and _87252_ (_37777_, _37776_, _37772_);
  nor _87253_ (_37778_, _37777_, _37412_);
  and _87254_ (_37779_, _37414_, \oc8051_golden_model_1.IRAM[13] [4]);
  and _87255_ (_37780_, _37416_, \oc8051_golden_model_1.IRAM[14] [4]);
  nor _87256_ (_37781_, _37780_, _37779_);
  and _87257_ (_37782_, _37419_, \oc8051_golden_model_1.IRAM[12] [4]);
  and _87258_ (_37783_, _37422_, \oc8051_golden_model_1.IRAM[15] [4]);
  nor _87259_ (_37785_, _37783_, _37782_);
  and _87260_ (_37786_, _37785_, _37781_);
  nor _87261_ (_37787_, _37786_, _37428_);
  nor _87262_ (_37788_, _37787_, _37778_);
  and _87263_ (_37789_, _37788_, _37769_);
  not _87264_ (_37790_, _37789_);
  and _87265_ (_37791_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  and _87266_ (_37792_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor _87267_ (_37793_, _37792_, _37791_);
  and _87268_ (_37794_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  and _87269_ (_37796_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor _87270_ (_37797_, _37796_, _37794_);
  and _87271_ (_37798_, _37797_, _37793_);
  and _87272_ (_37799_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  and _87273_ (_37800_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor _87274_ (_37801_, _37800_, _37799_);
  and _87275_ (_37802_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  and _87276_ (_37803_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor _87277_ (_37804_, _37803_, _37802_);
  and _87278_ (_37805_, _37804_, _37801_);
  and _87279_ (_37807_, _37805_, _37798_);
  and _87280_ (_37808_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  and _87281_ (_37809_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor _87282_ (_37810_, _37809_, _37808_);
  and _87283_ (_37811_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  and _87284_ (_37812_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor _87285_ (_37813_, _37812_, _37811_);
  and _87286_ (_37814_, _37813_, _37810_);
  and _87287_ (_37815_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  and _87288_ (_37816_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor _87289_ (_37818_, _37816_, _37815_);
  and _87290_ (_37819_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  and _87291_ (_37820_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor _87292_ (_37821_, _37820_, _37819_);
  and _87293_ (_37822_, _37821_, _37818_);
  and _87294_ (_37823_, _37822_, _37814_);
  and _87295_ (_37824_, _37823_, _37807_);
  nor _87296_ (_37825_, _37824_, _37790_);
  and _87297_ (_37826_, _37824_, _37790_);
  or _87298_ (_37827_, _37826_, _37825_);
  and _87299_ (_37829_, _37414_, \oc8051_golden_model_1.IRAM[1] [5]);
  and _87300_ (_37830_, _37416_, \oc8051_golden_model_1.IRAM[2] [5]);
  nor _87301_ (_37831_, _37830_, _37829_);
  and _87302_ (_37832_, _37419_, \oc8051_golden_model_1.IRAM[0] [5]);
  and _87303_ (_37833_, _37422_, \oc8051_golden_model_1.IRAM[3] [5]);
  nor _87304_ (_37834_, _37833_, _37832_);
  and _87305_ (_37835_, _37834_, _37831_);
  nor _87306_ (_37836_, _37835_, _37412_);
  and _87307_ (_37837_, _37414_, \oc8051_golden_model_1.IRAM[13] [5]);
  and _87308_ (_37838_, _37416_, \oc8051_golden_model_1.IRAM[14] [5]);
  nor _87309_ (_37840_, _37838_, _37837_);
  and _87310_ (_37841_, _37419_, \oc8051_golden_model_1.IRAM[12] [5]);
  and _87311_ (_37842_, _37422_, \oc8051_golden_model_1.IRAM[15] [5]);
  nor _87312_ (_37843_, _37842_, _37841_);
  and _87313_ (_37844_, _37843_, _37840_);
  nor _87314_ (_37845_, _37844_, _37428_);
  nor _87315_ (_37846_, _37845_, _37836_);
  and _87316_ (_37847_, _37414_, \oc8051_golden_model_1.IRAM[5] [5]);
  and _87317_ (_37848_, _37416_, \oc8051_golden_model_1.IRAM[6] [5]);
  nor _87318_ (_37849_, _37848_, _37847_);
  and _87319_ (_37851_, _37419_, \oc8051_golden_model_1.IRAM[4] [5]);
  and _87320_ (_37852_, _37422_, \oc8051_golden_model_1.IRAM[7] [5]);
  nor _87321_ (_37853_, _37852_, _37851_);
  and _87322_ (_37854_, _37853_, _37849_);
  nor _87323_ (_37855_, _37854_, _37441_);
  and _87324_ (_37856_, _37414_, \oc8051_golden_model_1.IRAM[9] [5]);
  and _87325_ (_37857_, _37416_, \oc8051_golden_model_1.IRAM[10] [5]);
  nor _87326_ (_37858_, _37857_, _37856_);
  and _87327_ (_37859_, _37419_, \oc8051_golden_model_1.IRAM[8] [5]);
  and _87328_ (_37860_, _37422_, \oc8051_golden_model_1.IRAM[11] [5]);
  nor _87329_ (_37862_, _37860_, _37859_);
  and _87330_ (_37863_, _37862_, _37858_);
  nor _87331_ (_37864_, _37863_, _37452_);
  nor _87332_ (_37865_, _37864_, _37855_);
  and _87333_ (_37866_, _37865_, _37846_);
  and _87334_ (_37867_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  and _87335_ (_37868_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor _87336_ (_37869_, _37868_, _37867_);
  and _87337_ (_37870_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  and _87338_ (_37871_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor _87339_ (_37873_, _37871_, _37870_);
  and _87340_ (_37874_, _37873_, _37869_);
  and _87341_ (_37875_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  and _87342_ (_37876_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor _87343_ (_37877_, _37876_, _37875_);
  and _87344_ (_37878_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  and _87345_ (_37879_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor _87346_ (_37880_, _37879_, _37878_);
  and _87347_ (_37881_, _37880_, _37877_);
  and _87348_ (_37882_, _37881_, _37874_);
  and _87349_ (_37884_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  and _87350_ (_37885_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor _87351_ (_37886_, _37885_, _37884_);
  and _87352_ (_37887_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  and _87353_ (_37888_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor _87354_ (_37889_, _37888_, _37887_);
  and _87355_ (_37890_, _37889_, _37886_);
  and _87356_ (_37891_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  and _87357_ (_37892_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor _87358_ (_37893_, _37892_, _37891_);
  and _87359_ (_37895_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  and _87360_ (_37896_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor _87361_ (_37897_, _37896_, _37895_);
  and _87362_ (_37898_, _37897_, _37893_);
  and _87363_ (_37899_, _37898_, _37890_);
  and _87364_ (_37900_, _37899_, _37882_);
  nand _87365_ (_37901_, _37900_, _37866_);
  or _87366_ (_37902_, _37900_, _37866_);
  and _87367_ (_37903_, _37902_, _37901_);
  or _87368_ (_37904_, _37903_, _37827_);
  and _87369_ (_37906_, _37414_, \oc8051_golden_model_1.IRAM[1] [6]);
  and _87370_ (_37907_, _37416_, \oc8051_golden_model_1.IRAM[2] [6]);
  nor _87371_ (_37908_, _37907_, _37906_);
  and _87372_ (_37909_, _37419_, \oc8051_golden_model_1.IRAM[0] [6]);
  and _87373_ (_37910_, _37422_, \oc8051_golden_model_1.IRAM[3] [6]);
  nor _87374_ (_37911_, _37910_, _37909_);
  and _87375_ (_37912_, _37911_, _37908_);
  nor _87376_ (_37913_, _37912_, _37412_);
  and _87377_ (_37914_, _37414_, \oc8051_golden_model_1.IRAM[9] [6]);
  and _87378_ (_37915_, _37416_, \oc8051_golden_model_1.IRAM[10] [6]);
  nor _87379_ (_37917_, _37915_, _37914_);
  and _87380_ (_37918_, _37419_, \oc8051_golden_model_1.IRAM[8] [6]);
  and _87381_ (_37919_, _37422_, \oc8051_golden_model_1.IRAM[11] [6]);
  nor _87382_ (_37920_, _37919_, _37918_);
  and _87383_ (_37921_, _37920_, _37917_);
  nor _87384_ (_37922_, _37921_, _37452_);
  nor _87385_ (_37923_, _37922_, _37913_);
  and _87386_ (_37924_, _37414_, \oc8051_golden_model_1.IRAM[5] [6]);
  and _87387_ (_37925_, _37416_, \oc8051_golden_model_1.IRAM[6] [6]);
  nor _87388_ (_37926_, _37925_, _37924_);
  and _87389_ (_37928_, _37419_, \oc8051_golden_model_1.IRAM[4] [6]);
  and _87390_ (_37929_, _37422_, \oc8051_golden_model_1.IRAM[7] [6]);
  nor _87391_ (_37930_, _37929_, _37928_);
  and _87392_ (_37931_, _37930_, _37926_);
  nor _87393_ (_37932_, _37931_, _37441_);
  and _87394_ (_37933_, _37414_, \oc8051_golden_model_1.IRAM[13] [6]);
  and _87395_ (_37934_, _37416_, \oc8051_golden_model_1.IRAM[14] [6]);
  nor _87396_ (_37935_, _37934_, _37933_);
  and _87397_ (_37936_, _37419_, \oc8051_golden_model_1.IRAM[12] [6]);
  and _87398_ (_37937_, _37422_, \oc8051_golden_model_1.IRAM[15] [6]);
  nor _87399_ (_37939_, _37937_, _37936_);
  and _87400_ (_37940_, _37939_, _37935_);
  nor _87401_ (_37941_, _37940_, _37428_);
  nor _87402_ (_37942_, _37941_, _37932_);
  and _87403_ (_37943_, _37942_, _37923_);
  and _87404_ (_37944_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  and _87405_ (_37945_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor _87406_ (_37946_, _37945_, _37944_);
  and _87407_ (_37947_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  and _87408_ (_37948_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor _87409_ (_37950_, _37948_, _37947_);
  and _87410_ (_37951_, _37950_, _37946_);
  and _87411_ (_37952_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  and _87412_ (_37953_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor _87413_ (_37954_, _37953_, _37952_);
  and _87414_ (_37955_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  and _87415_ (_37956_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor _87416_ (_37957_, _37956_, _37955_);
  and _87417_ (_37958_, _37957_, _37954_);
  and _87418_ (_37959_, _37958_, _37951_);
  and _87419_ (_37961_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  and _87420_ (_37962_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor _87421_ (_37963_, _37962_, _37961_);
  and _87422_ (_37964_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  and _87423_ (_37965_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor _87424_ (_37966_, _37965_, _37964_);
  and _87425_ (_37967_, _37966_, _37963_);
  and _87426_ (_37968_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  and _87427_ (_37969_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor _87428_ (_37970_, _37969_, _37968_);
  and _87429_ (_37972_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  and _87430_ (_37973_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor _87431_ (_37974_, _37973_, _37972_);
  and _87432_ (_37975_, _37974_, _37970_);
  and _87433_ (_37976_, _37975_, _37967_);
  and _87434_ (_37977_, _37976_, _37959_);
  nand _87435_ (_37978_, _37977_, _37943_);
  or _87436_ (_37979_, _37977_, _37943_);
  and _87437_ (_37980_, _37979_, _37978_);
  and _87438_ (_37981_, _37414_, \oc8051_golden_model_1.IRAM[5] [7]);
  and _87439_ (_37983_, _37416_, \oc8051_golden_model_1.IRAM[6] [7]);
  nor _87440_ (_37984_, _37983_, _37981_);
  and _87441_ (_37985_, _37419_, \oc8051_golden_model_1.IRAM[4] [7]);
  and _87442_ (_37986_, _37422_, \oc8051_golden_model_1.IRAM[7] [7]);
  nor _87443_ (_37987_, _37986_, _37985_);
  and _87444_ (_37988_, _37987_, _37984_);
  nor _87445_ (_37989_, _37988_, _37441_);
  and _87446_ (_37990_, _37414_, \oc8051_golden_model_1.IRAM[13] [7]);
  and _87447_ (_37991_, _37416_, \oc8051_golden_model_1.IRAM[14] [7]);
  nor _87448_ (_37992_, _37991_, _37990_);
  and _87449_ (_37994_, _37419_, \oc8051_golden_model_1.IRAM[12] [7]);
  and _87450_ (_37995_, _37422_, \oc8051_golden_model_1.IRAM[15] [7]);
  nor _87451_ (_37996_, _37995_, _37994_);
  and _87452_ (_37997_, _37996_, _37992_);
  nor _87453_ (_37998_, _37997_, _37428_);
  nor _87454_ (_37999_, _37998_, _37989_);
  and _87455_ (_38000_, _37414_, \oc8051_golden_model_1.IRAM[1] [7]);
  and _87456_ (_38001_, _37416_, \oc8051_golden_model_1.IRAM[2] [7]);
  nor _87457_ (_38002_, _38001_, _38000_);
  and _87458_ (_38003_, _37419_, \oc8051_golden_model_1.IRAM[0] [7]);
  and _87459_ (_38005_, _37422_, \oc8051_golden_model_1.IRAM[3] [7]);
  nor _87460_ (_38006_, _38005_, _38003_);
  and _87461_ (_38007_, _38006_, _38002_);
  nor _87462_ (_38008_, _38007_, _37412_);
  and _87463_ (_38009_, _37414_, \oc8051_golden_model_1.IRAM[9] [7]);
  and _87464_ (_38010_, _37416_, \oc8051_golden_model_1.IRAM[10] [7]);
  nor _87465_ (_38011_, _38010_, _38009_);
  and _87466_ (_38012_, _37419_, \oc8051_golden_model_1.IRAM[8] [7]);
  and _87467_ (_38013_, _37422_, \oc8051_golden_model_1.IRAM[11] [7]);
  nor _87468_ (_38014_, _38013_, _38012_);
  and _87469_ (_38016_, _38014_, _38011_);
  nor _87470_ (_38017_, _38016_, _37452_);
  nor _87471_ (_38018_, _38017_, _38008_);
  and _87472_ (_38019_, _38018_, _37999_);
  and _87473_ (_38020_, _37484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  and _87474_ (_38021_, _37477_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor _87475_ (_38022_, _38021_, _38020_);
  and _87476_ (_38023_, _37497_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  and _87477_ (_38024_, _37504_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nor _87478_ (_38025_, _38024_, _38023_);
  and _87479_ (_38027_, _38025_, _38022_);
  and _87480_ (_38028_, _37507_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  and _87481_ (_38029_, _37490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nor _87482_ (_38030_, _38029_, _38028_);
  and _87483_ (_38031_, _37472_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  and _87484_ (_38032_, _37510_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor _87485_ (_38033_, _38032_, _38031_);
  and _87486_ (_38034_, _38033_, _38030_);
  and _87487_ (_38035_, _38034_, _38027_);
  and _87488_ (_38036_, _37482_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  and _87489_ (_38038_, _37470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nor _87490_ (_38039_, _38038_, _38036_);
  and _87491_ (_38040_, _37464_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  and _87492_ (_38041_, _37467_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor _87493_ (_38042_, _38041_, _38040_);
  and _87494_ (_38043_, _38042_, _38039_);
  and _87495_ (_38044_, _37495_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  and _87496_ (_38045_, _37492_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor _87497_ (_38046_, _38045_, _38044_);
  and _87498_ (_38047_, _37502_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  and _87499_ (_38049_, _37479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nor _87500_ (_38050_, _38049_, _38047_);
  and _87501_ (_38051_, _38050_, _38046_);
  and _87502_ (_38052_, _38051_, _38043_);
  and _87503_ (_38053_, _38052_, _38035_);
  nand _87504_ (_38054_, _38053_, _38019_);
  or _87505_ (_38055_, _38053_, _38019_);
  and _87506_ (_38056_, _38055_, _38054_);
  or _87507_ (_38057_, _38056_, _37980_);
  or _87508_ (_38058_, _38057_, _37904_);
  or _87509_ (_38060_, _38058_, _37750_);
  and _87510_ (property_invalid_iram, _38060_, _37409_);
  nor _87511_ (_38061_, _09956_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _87512_ (_38062_, _09956_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _87513_ (_38063_, _38062_, _38061_);
  nand _87514_ (_38064_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _87515_ (_38065_, \oc8051_golden_model_1.ACC [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _87516_ (_38066_, _38065_, _38064_);
  or _87517_ (_38067_, _38066_, _38063_);
  and _87518_ (_38068_, _05784_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor _87519_ (_38070_, _05784_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _87520_ (_38071_, _38070_, _38068_);
  and _87521_ (_38072_, _05758_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _87522_ (_38073_, \oc8051_golden_model_1.ACC [0], _39048_);
  or _87523_ (_38074_, _38073_, _38072_);
  or _87524_ (_38075_, _38074_, _38071_);
  or _87525_ (_38076_, _38075_, _38067_);
  or _87526_ (_38077_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand _87527_ (_38078_, \oc8051_golden_model_1.ACC [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _87528_ (_38079_, _38078_, _38077_);
  or _87529_ (_38081_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _87530_ (_38082_, \oc8051_golden_model_1.ACC [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and _87531_ (_38083_, _38082_, _38081_);
  or _87532_ (_38084_, _38083_, _38079_);
  nand _87533_ (_38085_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _87534_ (_38086_, \oc8051_golden_model_1.ACC [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _87535_ (_38087_, _38086_, _38085_);
  and _87536_ (_38088_, _08393_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor _87537_ (_38089_, _08393_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or _87538_ (_38090_, _38089_, _38088_);
  or _87539_ (_38092_, _38090_, _38087_);
  or _87540_ (_38093_, _38092_, _38084_);
  or _87541_ (_38094_, _38093_, _38076_);
  and _87542_ (property_invalid_acc, _38094_, _37409_);
  and _87543_ (_38095_, _37408_, _01336_);
  nor _87544_ (_38096_, _25378_, _01937_);
  and _87545_ (_38097_, _25378_, _01937_);
  or _87546_ (_38098_, _38097_, _38096_);
  nor _87547_ (_38099_, _25728_, _01941_);
  nor _87548_ (_38100_, _26416_, _01949_);
  or _87549_ (_38102_, _38100_, _38099_);
  nor _87550_ (_38103_, _26769_, _01953_);
  and _87551_ (_38104_, _26416_, _01949_);
  or _87552_ (_38105_, _38104_, _38103_);
  or _87553_ (_38106_, _38105_, _38102_);
  nor _87554_ (_38107_, _26067_, _01945_);
  and _87555_ (_38108_, _28118_, _38558_);
  nor _87556_ (_38109_, _28118_, _38558_);
  and _87557_ (_38110_, _12796_, _38536_);
  nor _87558_ (_38111_, _12796_, _38536_);
  or _87559_ (_38113_, _38111_, _38110_);
  and _87560_ (_38114_, _27796_, _38552_);
  nor _87561_ (_38115_, _29339_, _38544_);
  or _87562_ (_38116_, _38115_, _38114_);
  or _87563_ (_38117_, _38116_, _38113_);
  nand _87564_ (_38118_, _25007_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or _87565_ (_38119_, _25007_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _87566_ (_38120_, _38119_, _38118_);
  nor _87567_ (_38121_, _29649_, _38540_);
  or _87568_ (_38122_, _38121_, _38120_);
  nor _87569_ (_38124_, _28728_, _38548_);
  and _87570_ (_38125_, _28728_, _38548_);
  and _87571_ (_38126_, _29649_, _38540_);
  or _87572_ (_38127_, _38126_, _38125_);
  or _87573_ (_38128_, _38127_, _38124_);
  or _87574_ (_38129_, _38128_, _38122_);
  nor _87575_ (_38130_, _27796_, _38552_);
  and _87576_ (_38131_, _29339_, _38544_);
  or _87577_ (_38132_, _38131_, _38130_);
  or _87578_ (_38133_, _38132_, _38129_);
  or _87579_ (_38135_, _38133_, _38117_);
  and _87580_ (_38136_, _28426_, _38563_);
  nor _87581_ (_38137_, _28426_, _38563_);
  or _87582_ (_38138_, _38137_, _38136_);
  and _87583_ (_38139_, _29035_, _38569_);
  nor _87584_ (_38140_, _29035_, _38569_);
  or _87585_ (_38141_, _38140_, _38139_);
  or _87586_ (_38142_, _38141_, _38138_);
  or _87587_ (_38143_, _38142_, _38135_);
  or _87588_ (_38144_, _38143_, _38109_);
  or _87589_ (_38146_, _38144_, _38108_);
  or _87590_ (_38147_, _38146_, _38107_);
  nor _87591_ (_38148_, _27474_, _01960_);
  and _87592_ (_38149_, _27474_, _01960_);
  or _87593_ (_38150_, _38149_, _38148_);
  and _87594_ (_38151_, _26067_, _01945_);
  nand _87595_ (_38152_, _27119_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _87596_ (_38153_, _27119_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _87597_ (_38154_, _38153_, _38152_);
  or _87598_ (_38155_, _38154_, _38151_);
  or _87599_ (_38157_, _38155_, _38150_);
  or _87600_ (_38158_, _38157_, _38147_);
  and _87601_ (_38159_, _25728_, _01941_);
  and _87602_ (_38160_, _26769_, _01953_);
  or _87603_ (_38161_, _38160_, _38159_);
  or _87604_ (_38162_, _38161_, _38158_);
  or _87605_ (_38163_, _38162_, _38106_);
  or _87606_ (_38164_, _38163_, _38098_);
  and _87607_ (property_invalid_pc, _38164_, _38095_);
  buf _87608_ (_00543_, _42885_);
  buf _87609_ (_05103_, _42882_);
  buf _87610_ (_05155_, _42882_);
  buf _87611_ (_05206_, _42882_);
  buf _87612_ (_05258_, _42882_);
  buf _87613_ (_05309_, _42882_);
  buf _87614_ (_05362_, _42882_);
  buf _87615_ (_05415_, _42882_);
  buf _87616_ (_05468_, _42882_);
  buf _87617_ (_05521_, _42882_);
  buf _87618_ (_05574_, _42882_);
  buf _87619_ (_05627_, _42882_);
  buf _87620_ (_05680_, _42882_);
  buf _87621_ (_05733_, _42882_);
  buf _87622_ (_05786_, _42882_);
  buf _87623_ (_05839_, _42882_);
  buf _87624_ (_05892_, _42882_);
  buf _87625_ (_39058_, _38956_);
  buf _87626_ (_39060_, _38958_);
  buf _87627_ (_39073_, _38956_);
  buf _87628_ (_39074_, _38958_);
  buf _87629_ (_39386_, _38975_);
  buf _87630_ (_39387_, _38976_);
  buf _87631_ (_39388_, _38978_);
  buf _87632_ (_39389_, _38979_);
  buf _87633_ (_39390_, _38980_);
  buf _87634_ (_39391_, _38981_);
  buf _87635_ (_39392_, _38982_);
  buf _87636_ (_39393_, _38984_);
  buf _87637_ (_39394_, _38985_);
  buf _87638_ (_39396_, _38986_);
  buf _87639_ (_39397_, _38987_);
  buf _87640_ (_39398_, _38988_);
  buf _87641_ (_39399_, _38990_);
  buf _87642_ (_39400_, _38991_);
  buf _87643_ (_39451_, _38975_);
  buf _87644_ (_39452_, _38976_);
  buf _87645_ (_39453_, _38978_);
  buf _87646_ (_39454_, _38979_);
  buf _87647_ (_39455_, _38980_);
  buf _87648_ (_39456_, _38981_);
  buf _87649_ (_39457_, _38982_);
  buf _87650_ (_39458_, _38984_);
  buf _87651_ (_39459_, _38985_);
  buf _87652_ (_39461_, _38986_);
  buf _87653_ (_39462_, _38987_);
  buf _87654_ (_39463_, _38988_);
  buf _87655_ (_39464_, _38990_);
  buf _87656_ (_39465_, _38991_);
  buf _87657_ (_39855_, _39760_);
  buf _87658_ (_40018_, _39760_);
  dff _87659_ (op0_cnst, _00001_, clk);
  dff _87660_ (inst_finished_r, _00000_, clk);
  dff _87661_ (\oc8051_gm_cxrom_1.cell0.data [0], _05107_, clk);
  dff _87662_ (\oc8051_gm_cxrom_1.cell0.data [1], _05111_, clk);
  dff _87663_ (\oc8051_gm_cxrom_1.cell0.data [2], _05115_, clk);
  dff _87664_ (\oc8051_gm_cxrom_1.cell0.data [3], _05119_, clk);
  dff _87665_ (\oc8051_gm_cxrom_1.cell0.data [4], _05123_, clk);
  dff _87666_ (\oc8051_gm_cxrom_1.cell0.data [5], _05126_, clk);
  dff _87667_ (\oc8051_gm_cxrom_1.cell0.data [6], _05130_, clk);
  dff _87668_ (\oc8051_gm_cxrom_1.cell0.data [7], _05100_, clk);
  dff _87669_ (\oc8051_gm_cxrom_1.cell0.valid , _05103_, clk);
  dff _87670_ (\oc8051_gm_cxrom_1.cell1.data [0], _05159_, clk);
  dff _87671_ (\oc8051_gm_cxrom_1.cell1.data [1], _05162_, clk);
  dff _87672_ (\oc8051_gm_cxrom_1.cell1.data [2], _05166_, clk);
  dff _87673_ (\oc8051_gm_cxrom_1.cell1.data [3], _05170_, clk);
  dff _87674_ (\oc8051_gm_cxrom_1.cell1.data [4], _05174_, clk);
  dff _87675_ (\oc8051_gm_cxrom_1.cell1.data [5], _05178_, clk);
  dff _87676_ (\oc8051_gm_cxrom_1.cell1.data [6], _05182_, clk);
  dff _87677_ (\oc8051_gm_cxrom_1.cell1.data [7], _05152_, clk);
  dff _87678_ (\oc8051_gm_cxrom_1.cell1.valid , _05155_, clk);
  dff _87679_ (\oc8051_gm_cxrom_1.cell10.data [0], _05631_, clk);
  dff _87680_ (\oc8051_gm_cxrom_1.cell10.data [1], _05635_, clk);
  dff _87681_ (\oc8051_gm_cxrom_1.cell10.data [2], _05639_, clk);
  dff _87682_ (\oc8051_gm_cxrom_1.cell10.data [3], _05643_, clk);
  dff _87683_ (\oc8051_gm_cxrom_1.cell10.data [4], _05647_, clk);
  dff _87684_ (\oc8051_gm_cxrom_1.cell10.data [5], _05651_, clk);
  dff _87685_ (\oc8051_gm_cxrom_1.cell10.data [6], _05655_, clk);
  dff _87686_ (\oc8051_gm_cxrom_1.cell10.data [7], _05624_, clk);
  dff _87687_ (\oc8051_gm_cxrom_1.cell10.valid , _05627_, clk);
  dff _87688_ (\oc8051_gm_cxrom_1.cell11.data [0], _05684_, clk);
  dff _87689_ (\oc8051_gm_cxrom_1.cell11.data [1], _05688_, clk);
  dff _87690_ (\oc8051_gm_cxrom_1.cell11.data [2], _05692_, clk);
  dff _87691_ (\oc8051_gm_cxrom_1.cell11.data [3], _05696_, clk);
  dff _87692_ (\oc8051_gm_cxrom_1.cell11.data [4], _05700_, clk);
  dff _87693_ (\oc8051_gm_cxrom_1.cell11.data [5], _05704_, clk);
  dff _87694_ (\oc8051_gm_cxrom_1.cell11.data [6], _05708_, clk);
  dff _87695_ (\oc8051_gm_cxrom_1.cell11.data [7], _05677_, clk);
  dff _87696_ (\oc8051_gm_cxrom_1.cell11.valid , _05680_, clk);
  dff _87697_ (\oc8051_gm_cxrom_1.cell12.data [0], _05737_, clk);
  dff _87698_ (\oc8051_gm_cxrom_1.cell12.data [1], _05741_, clk);
  dff _87699_ (\oc8051_gm_cxrom_1.cell12.data [2], _05745_, clk);
  dff _87700_ (\oc8051_gm_cxrom_1.cell12.data [3], _05749_, clk);
  dff _87701_ (\oc8051_gm_cxrom_1.cell12.data [4], _05753_, clk);
  dff _87702_ (\oc8051_gm_cxrom_1.cell12.data [5], _05757_, clk);
  dff _87703_ (\oc8051_gm_cxrom_1.cell12.data [6], _05761_, clk);
  dff _87704_ (\oc8051_gm_cxrom_1.cell12.data [7], _05730_, clk);
  dff _87705_ (\oc8051_gm_cxrom_1.cell12.valid , _05733_, clk);
  dff _87706_ (\oc8051_gm_cxrom_1.cell13.data [0], _05790_, clk);
  dff _87707_ (\oc8051_gm_cxrom_1.cell13.data [1], _05794_, clk);
  dff _87708_ (\oc8051_gm_cxrom_1.cell13.data [2], _05798_, clk);
  dff _87709_ (\oc8051_gm_cxrom_1.cell13.data [3], _05802_, clk);
  dff _87710_ (\oc8051_gm_cxrom_1.cell13.data [4], _05806_, clk);
  dff _87711_ (\oc8051_gm_cxrom_1.cell13.data [5], _05810_, clk);
  dff _87712_ (\oc8051_gm_cxrom_1.cell13.data [6], _05814_, clk);
  dff _87713_ (\oc8051_gm_cxrom_1.cell13.data [7], _05783_, clk);
  dff _87714_ (\oc8051_gm_cxrom_1.cell13.valid , _05786_, clk);
  dff _87715_ (\oc8051_gm_cxrom_1.cell14.data [0], _05843_, clk);
  dff _87716_ (\oc8051_gm_cxrom_1.cell14.data [1], _05847_, clk);
  dff _87717_ (\oc8051_gm_cxrom_1.cell14.data [2], _05851_, clk);
  dff _87718_ (\oc8051_gm_cxrom_1.cell14.data [3], _05855_, clk);
  dff _87719_ (\oc8051_gm_cxrom_1.cell14.data [4], _05859_, clk);
  dff _87720_ (\oc8051_gm_cxrom_1.cell14.data [5], _05863_, clk);
  dff _87721_ (\oc8051_gm_cxrom_1.cell14.data [6], _05867_, clk);
  dff _87722_ (\oc8051_gm_cxrom_1.cell14.data [7], _05836_, clk);
  dff _87723_ (\oc8051_gm_cxrom_1.cell14.valid , _05839_, clk);
  dff _87724_ (\oc8051_gm_cxrom_1.cell15.data [0], _05896_, clk);
  dff _87725_ (\oc8051_gm_cxrom_1.cell15.data [1], _05900_, clk);
  dff _87726_ (\oc8051_gm_cxrom_1.cell15.data [2], _05904_, clk);
  dff _87727_ (\oc8051_gm_cxrom_1.cell15.data [3], _05908_, clk);
  dff _87728_ (\oc8051_gm_cxrom_1.cell15.data [4], _05912_, clk);
  dff _87729_ (\oc8051_gm_cxrom_1.cell15.data [5], _05916_, clk);
  dff _87730_ (\oc8051_gm_cxrom_1.cell15.data [6], _05920_, clk);
  dff _87731_ (\oc8051_gm_cxrom_1.cell15.data [7], _05889_, clk);
  dff _87732_ (\oc8051_gm_cxrom_1.cell15.valid , _05892_, clk);
  dff _87733_ (\oc8051_gm_cxrom_1.cell2.data [0], _05210_, clk);
  dff _87734_ (\oc8051_gm_cxrom_1.cell2.data [1], _05214_, clk);
  dff _87735_ (\oc8051_gm_cxrom_1.cell2.data [2], _05218_, clk);
  dff _87736_ (\oc8051_gm_cxrom_1.cell2.data [3], _05222_, clk);
  dff _87737_ (\oc8051_gm_cxrom_1.cell2.data [4], _05226_, clk);
  dff _87738_ (\oc8051_gm_cxrom_1.cell2.data [5], _05230_, clk);
  dff _87739_ (\oc8051_gm_cxrom_1.cell2.data [6], _05234_, clk);
  dff _87740_ (\oc8051_gm_cxrom_1.cell2.data [7], _05203_, clk);
  dff _87741_ (\oc8051_gm_cxrom_1.cell2.valid , _05206_, clk);
  dff _87742_ (\oc8051_gm_cxrom_1.cell3.data [0], _05262_, clk);
  dff _87743_ (\oc8051_gm_cxrom_1.cell3.data [1], _05266_, clk);
  dff _87744_ (\oc8051_gm_cxrom_1.cell3.data [2], _05270_, clk);
  dff _87745_ (\oc8051_gm_cxrom_1.cell3.data [3], _05273_, clk);
  dff _87746_ (\oc8051_gm_cxrom_1.cell3.data [4], _05277_, clk);
  dff _87747_ (\oc8051_gm_cxrom_1.cell3.data [5], _05281_, clk);
  dff _87748_ (\oc8051_gm_cxrom_1.cell3.data [6], _05285_, clk);
  dff _87749_ (\oc8051_gm_cxrom_1.cell3.data [7], _05255_, clk);
  dff _87750_ (\oc8051_gm_cxrom_1.cell3.valid , _05258_, clk);
  dff _87751_ (\oc8051_gm_cxrom_1.cell4.data [0], _05313_, clk);
  dff _87752_ (\oc8051_gm_cxrom_1.cell4.data [1], _05317_, clk);
  dff _87753_ (\oc8051_gm_cxrom_1.cell4.data [2], _05321_, clk);
  dff _87754_ (\oc8051_gm_cxrom_1.cell4.data [3], _05325_, clk);
  dff _87755_ (\oc8051_gm_cxrom_1.cell4.data [4], _05329_, clk);
  dff _87756_ (\oc8051_gm_cxrom_1.cell4.data [5], _05333_, clk);
  dff _87757_ (\oc8051_gm_cxrom_1.cell4.data [6], _05337_, clk);
  dff _87758_ (\oc8051_gm_cxrom_1.cell4.data [7], _05306_, clk);
  dff _87759_ (\oc8051_gm_cxrom_1.cell4.valid , _05309_, clk);
  dff _87760_ (\oc8051_gm_cxrom_1.cell5.data [0], _05366_, clk);
  dff _87761_ (\oc8051_gm_cxrom_1.cell5.data [1], _05370_, clk);
  dff _87762_ (\oc8051_gm_cxrom_1.cell5.data [2], _05374_, clk);
  dff _87763_ (\oc8051_gm_cxrom_1.cell5.data [3], _05378_, clk);
  dff _87764_ (\oc8051_gm_cxrom_1.cell5.data [4], _05382_, clk);
  dff _87765_ (\oc8051_gm_cxrom_1.cell5.data [5], _05386_, clk);
  dff _87766_ (\oc8051_gm_cxrom_1.cell5.data [6], _05390_, clk);
  dff _87767_ (\oc8051_gm_cxrom_1.cell5.data [7], _05359_, clk);
  dff _87768_ (\oc8051_gm_cxrom_1.cell5.valid , _05362_, clk);
  dff _87769_ (\oc8051_gm_cxrom_1.cell6.data [0], _05419_, clk);
  dff _87770_ (\oc8051_gm_cxrom_1.cell6.data [1], _05423_, clk);
  dff _87771_ (\oc8051_gm_cxrom_1.cell6.data [2], _05427_, clk);
  dff _87772_ (\oc8051_gm_cxrom_1.cell6.data [3], _05431_, clk);
  dff _87773_ (\oc8051_gm_cxrom_1.cell6.data [4], _05435_, clk);
  dff _87774_ (\oc8051_gm_cxrom_1.cell6.data [5], _05439_, clk);
  dff _87775_ (\oc8051_gm_cxrom_1.cell6.data [6], _05443_, clk);
  dff _87776_ (\oc8051_gm_cxrom_1.cell6.data [7], _05412_, clk);
  dff _87777_ (\oc8051_gm_cxrom_1.cell6.valid , _05415_, clk);
  dff _87778_ (\oc8051_gm_cxrom_1.cell7.data [0], _05472_, clk);
  dff _87779_ (\oc8051_gm_cxrom_1.cell7.data [1], _05476_, clk);
  dff _87780_ (\oc8051_gm_cxrom_1.cell7.data [2], _05480_, clk);
  dff _87781_ (\oc8051_gm_cxrom_1.cell7.data [3], _05484_, clk);
  dff _87782_ (\oc8051_gm_cxrom_1.cell7.data [4], _05488_, clk);
  dff _87783_ (\oc8051_gm_cxrom_1.cell7.data [5], _05492_, clk);
  dff _87784_ (\oc8051_gm_cxrom_1.cell7.data [6], _05496_, clk);
  dff _87785_ (\oc8051_gm_cxrom_1.cell7.data [7], _05465_, clk);
  dff _87786_ (\oc8051_gm_cxrom_1.cell7.valid , _05468_, clk);
  dff _87787_ (\oc8051_gm_cxrom_1.cell8.data [0], _05525_, clk);
  dff _87788_ (\oc8051_gm_cxrom_1.cell8.data [1], _05529_, clk);
  dff _87789_ (\oc8051_gm_cxrom_1.cell8.data [2], _05533_, clk);
  dff _87790_ (\oc8051_gm_cxrom_1.cell8.data [3], _05537_, clk);
  dff _87791_ (\oc8051_gm_cxrom_1.cell8.data [4], _05541_, clk);
  dff _87792_ (\oc8051_gm_cxrom_1.cell8.data [5], _05545_, clk);
  dff _87793_ (\oc8051_gm_cxrom_1.cell8.data [6], _05549_, clk);
  dff _87794_ (\oc8051_gm_cxrom_1.cell8.data [7], _05518_, clk);
  dff _87795_ (\oc8051_gm_cxrom_1.cell8.valid , _05521_, clk);
  dff _87796_ (\oc8051_gm_cxrom_1.cell9.data [0], _05578_, clk);
  dff _87797_ (\oc8051_gm_cxrom_1.cell9.data [1], _05582_, clk);
  dff _87798_ (\oc8051_gm_cxrom_1.cell9.data [2], _05586_, clk);
  dff _87799_ (\oc8051_gm_cxrom_1.cell9.data [3], _05590_, clk);
  dff _87800_ (\oc8051_gm_cxrom_1.cell9.data [4], _05594_, clk);
  dff _87801_ (\oc8051_gm_cxrom_1.cell9.data [5], _05598_, clk);
  dff _87802_ (\oc8051_gm_cxrom_1.cell9.data [6], _05602_, clk);
  dff _87803_ (\oc8051_gm_cxrom_1.cell9.data [7], _05571_, clk);
  dff _87804_ (\oc8051_gm_cxrom_1.cell9.valid , _05574_, clk);
  dff _87805_ (\oc8051_golden_model_1.IRAM[15] [0], _40967_, clk);
  dff _87806_ (\oc8051_golden_model_1.IRAM[15] [1], _40968_, clk);
  dff _87807_ (\oc8051_golden_model_1.IRAM[15] [2], _40969_, clk);
  dff _87808_ (\oc8051_golden_model_1.IRAM[15] [3], _40970_, clk);
  dff _87809_ (\oc8051_golden_model_1.IRAM[15] [4], _40971_, clk);
  dff _87810_ (\oc8051_golden_model_1.IRAM[15] [5], _40972_, clk);
  dff _87811_ (\oc8051_golden_model_1.IRAM[15] [6], _40973_, clk);
  dff _87812_ (\oc8051_golden_model_1.IRAM[15] [7], _40751_, clk);
  dff _87813_ (\oc8051_golden_model_1.IRAM[14] [0], _40956_, clk);
  dff _87814_ (\oc8051_golden_model_1.IRAM[14] [1], _40957_, clk);
  dff _87815_ (\oc8051_golden_model_1.IRAM[14] [2], _40958_, clk);
  dff _87816_ (\oc8051_golden_model_1.IRAM[14] [3], _40959_, clk);
  dff _87817_ (\oc8051_golden_model_1.IRAM[14] [4], _40960_, clk);
  dff _87818_ (\oc8051_golden_model_1.IRAM[14] [5], _40962_, clk);
  dff _87819_ (\oc8051_golden_model_1.IRAM[14] [6], _40963_, clk);
  dff _87820_ (\oc8051_golden_model_1.IRAM[14] [7], _40964_, clk);
  dff _87821_ (\oc8051_golden_model_1.IRAM[13] [0], _40943_, clk);
  dff _87822_ (\oc8051_golden_model_1.IRAM[13] [1], _40945_, clk);
  dff _87823_ (\oc8051_golden_model_1.IRAM[13] [2], _40946_, clk);
  dff _87824_ (\oc8051_golden_model_1.IRAM[13] [3], _40947_, clk);
  dff _87825_ (\oc8051_golden_model_1.IRAM[13] [4], _40948_, clk);
  dff _87826_ (\oc8051_golden_model_1.IRAM[13] [5], _40949_, clk);
  dff _87827_ (\oc8051_golden_model_1.IRAM[13] [6], _40951_, clk);
  dff _87828_ (\oc8051_golden_model_1.IRAM[13] [7], _40952_, clk);
  dff _87829_ (\oc8051_golden_model_1.IRAM[12] [0], _40932_, clk);
  dff _87830_ (\oc8051_golden_model_1.IRAM[12] [1], _40933_, clk);
  dff _87831_ (\oc8051_golden_model_1.IRAM[12] [2], _40934_, clk);
  dff _87832_ (\oc8051_golden_model_1.IRAM[12] [3], _40935_, clk);
  dff _87833_ (\oc8051_golden_model_1.IRAM[12] [4], _40936_, clk);
  dff _87834_ (\oc8051_golden_model_1.IRAM[12] [5], _40937_, clk);
  dff _87835_ (\oc8051_golden_model_1.IRAM[12] [6], _40939_, clk);
  dff _87836_ (\oc8051_golden_model_1.IRAM[12] [7], _40940_, clk);
  dff _87837_ (\oc8051_golden_model_1.IRAM[11] [0], _40919_, clk);
  dff _87838_ (\oc8051_golden_model_1.IRAM[11] [1], _40920_, clk);
  dff _87839_ (\oc8051_golden_model_1.IRAM[11] [2], _40921_, clk);
  dff _87840_ (\oc8051_golden_model_1.IRAM[11] [3], _40924_, clk);
  dff _87841_ (\oc8051_golden_model_1.IRAM[11] [4], _40925_, clk);
  dff _87842_ (\oc8051_golden_model_1.IRAM[11] [5], _40926_, clk);
  dff _87843_ (\oc8051_golden_model_1.IRAM[11] [6], _40927_, clk);
  dff _87844_ (\oc8051_golden_model_1.IRAM[11] [7], _40928_, clk);
  dff _87845_ (\oc8051_golden_model_1.IRAM[10] [0], _40908_, clk);
  dff _87846_ (\oc8051_golden_model_1.IRAM[10] [1], _40909_, clk);
  dff _87847_ (\oc8051_golden_model_1.IRAM[10] [2], _40910_, clk);
  dff _87848_ (\oc8051_golden_model_1.IRAM[10] [3], _40912_, clk);
  dff _87849_ (\oc8051_golden_model_1.IRAM[10] [4], _40913_, clk);
  dff _87850_ (\oc8051_golden_model_1.IRAM[10] [5], _40914_, clk);
  dff _87851_ (\oc8051_golden_model_1.IRAM[10] [6], _40915_, clk);
  dff _87852_ (\oc8051_golden_model_1.IRAM[10] [7], _40916_, clk);
  dff _87853_ (\oc8051_golden_model_1.IRAM[9] [0], _40896_, clk);
  dff _87854_ (\oc8051_golden_model_1.IRAM[9] [1], _40897_, clk);
  dff _87855_ (\oc8051_golden_model_1.IRAM[9] [2], _40898_, clk);
  dff _87856_ (\oc8051_golden_model_1.IRAM[9] [3], _40899_, clk);
  dff _87857_ (\oc8051_golden_model_1.IRAM[9] [4], _40901_, clk);
  dff _87858_ (\oc8051_golden_model_1.IRAM[9] [5], _40902_, clk);
  dff _87859_ (\oc8051_golden_model_1.IRAM[9] [6], _40903_, clk);
  dff _87860_ (\oc8051_golden_model_1.IRAM[9] [7], _40904_, clk);
  dff _87861_ (\oc8051_golden_model_1.IRAM[8] [0], _40884_, clk);
  dff _87862_ (\oc8051_golden_model_1.IRAM[8] [1], _40885_, clk);
  dff _87863_ (\oc8051_golden_model_1.IRAM[8] [2], _40886_, clk);
  dff _87864_ (\oc8051_golden_model_1.IRAM[8] [3], _40887_, clk);
  dff _87865_ (\oc8051_golden_model_1.IRAM[8] [4], _40889_, clk);
  dff _87866_ (\oc8051_golden_model_1.IRAM[8] [5], _40890_, clk);
  dff _87867_ (\oc8051_golden_model_1.IRAM[8] [6], _40891_, clk);
  dff _87868_ (\oc8051_golden_model_1.IRAM[8] [7], _40892_, clk);
  dff _87869_ (\oc8051_golden_model_1.IRAM[7] [0], _40872_, clk);
  dff _87870_ (\oc8051_golden_model_1.IRAM[7] [1], _40873_, clk);
  dff _87871_ (\oc8051_golden_model_1.IRAM[7] [2], _40874_, clk);
  dff _87872_ (\oc8051_golden_model_1.IRAM[7] [3], _40876_, clk);
  dff _87873_ (\oc8051_golden_model_1.IRAM[7] [4], _40877_, clk);
  dff _87874_ (\oc8051_golden_model_1.IRAM[7] [5], _40878_, clk);
  dff _87875_ (\oc8051_golden_model_1.IRAM[7] [6], _40879_, clk);
  dff _87876_ (\oc8051_golden_model_1.IRAM[7] [7], _40880_, clk);
  dff _87877_ (\oc8051_golden_model_1.IRAM[6] [0], _40860_, clk);
  dff _87878_ (\oc8051_golden_model_1.IRAM[6] [1], _40861_, clk);
  dff _87879_ (\oc8051_golden_model_1.IRAM[6] [2], _40862_, clk);
  dff _87880_ (\oc8051_golden_model_1.IRAM[6] [3], _40863_, clk);
  dff _87881_ (\oc8051_golden_model_1.IRAM[6] [4], _40864_, clk);
  dff _87882_ (\oc8051_golden_model_1.IRAM[6] [5], _40865_, clk);
  dff _87883_ (\oc8051_golden_model_1.IRAM[6] [6], _40866_, clk);
  dff _87884_ (\oc8051_golden_model_1.IRAM[6] [7], _40867_, clk);
  dff _87885_ (\oc8051_golden_model_1.IRAM[5] [0], _40848_, clk);
  dff _87886_ (\oc8051_golden_model_1.IRAM[5] [1], _40849_, clk);
  dff _87887_ (\oc8051_golden_model_1.IRAM[5] [2], _40850_, clk);
  dff _87888_ (\oc8051_golden_model_1.IRAM[5] [3], _40851_, clk);
  dff _87889_ (\oc8051_golden_model_1.IRAM[5] [4], _40853_, clk);
  dff _87890_ (\oc8051_golden_model_1.IRAM[5] [5], _40854_, clk);
  dff _87891_ (\oc8051_golden_model_1.IRAM[5] [6], _40855_, clk);
  dff _87892_ (\oc8051_golden_model_1.IRAM[5] [7], _40856_, clk);
  dff _87893_ (\oc8051_golden_model_1.IRAM[4] [0], _40835_, clk);
  dff _87894_ (\oc8051_golden_model_1.IRAM[4] [1], _40836_, clk);
  dff _87895_ (\oc8051_golden_model_1.IRAM[4] [2], _40837_, clk);
  dff _87896_ (\oc8051_golden_model_1.IRAM[4] [3], _40838_, clk);
  dff _87897_ (\oc8051_golden_model_1.IRAM[4] [4], _40841_, clk);
  dff _87898_ (\oc8051_golden_model_1.IRAM[4] [5], _40842_, clk);
  dff _87899_ (\oc8051_golden_model_1.IRAM[4] [6], _40843_, clk);
  dff _87900_ (\oc8051_golden_model_1.IRAM[4] [7], _40844_, clk);
  dff _87901_ (\oc8051_golden_model_1.IRAM[3] [0], _40823_, clk);
  dff _87902_ (\oc8051_golden_model_1.IRAM[3] [1], _40824_, clk);
  dff _87903_ (\oc8051_golden_model_1.IRAM[3] [2], _40825_, clk);
  dff _87904_ (\oc8051_golden_model_1.IRAM[3] [3], _40827_, clk);
  dff _87905_ (\oc8051_golden_model_1.IRAM[3] [4], _40828_, clk);
  dff _87906_ (\oc8051_golden_model_1.IRAM[3] [5], _40829_, clk);
  dff _87907_ (\oc8051_golden_model_1.IRAM[3] [6], _40830_, clk);
  dff _87908_ (\oc8051_golden_model_1.IRAM[3] [7], _40831_, clk);
  dff _87909_ (\oc8051_golden_model_1.IRAM[2] [0], _40813_, clk);
  dff _87910_ (\oc8051_golden_model_1.IRAM[2] [1], _40814_, clk);
  dff _87911_ (\oc8051_golden_model_1.IRAM[2] [2], _40815_, clk);
  dff _87912_ (\oc8051_golden_model_1.IRAM[2] [3], _40816_, clk);
  dff _87913_ (\oc8051_golden_model_1.IRAM[2] [4], _40818_, clk);
  dff _87914_ (\oc8051_golden_model_1.IRAM[2] [5], _40819_, clk);
  dff _87915_ (\oc8051_golden_model_1.IRAM[2] [6], _40820_, clk);
  dff _87916_ (\oc8051_golden_model_1.IRAM[2] [7], _40821_, clk);
  dff _87917_ (\oc8051_golden_model_1.IRAM[1] [0], _40801_, clk);
  dff _87918_ (\oc8051_golden_model_1.IRAM[1] [1], _40802_, clk);
  dff _87919_ (\oc8051_golden_model_1.IRAM[1] [2], _40803_, clk);
  dff _87920_ (\oc8051_golden_model_1.IRAM[1] [3], _40805_, clk);
  dff _87921_ (\oc8051_golden_model_1.IRAM[1] [4], _40806_, clk);
  dff _87922_ (\oc8051_golden_model_1.IRAM[1] [5], _40807_, clk);
  dff _87923_ (\oc8051_golden_model_1.IRAM[1] [6], _40808_, clk);
  dff _87924_ (\oc8051_golden_model_1.IRAM[1] [7], _40809_, clk);
  dff _87925_ (\oc8051_golden_model_1.IRAM[0] [0], _40792_, clk);
  dff _87926_ (\oc8051_golden_model_1.IRAM[0] [1], _40793_, clk);
  dff _87927_ (\oc8051_golden_model_1.IRAM[0] [2], _40794_, clk);
  dff _87928_ (\oc8051_golden_model_1.IRAM[0] [3], _40795_, clk);
  dff _87929_ (\oc8051_golden_model_1.IRAM[0] [4], _40797_, clk);
  dff _87930_ (\oc8051_golden_model_1.IRAM[0] [5], _40798_, clk);
  dff _87931_ (\oc8051_golden_model_1.IRAM[0] [6], _40799_, clk);
  dff _87932_ (\oc8051_golden_model_1.IRAM[0] [7], _40800_, clk);
  dff _87933_ (\oc8051_golden_model_1.B [0], _43324_, clk);
  dff _87934_ (\oc8051_golden_model_1.B [1], _43325_, clk);
  dff _87935_ (\oc8051_golden_model_1.B [2], _43326_, clk);
  dff _87936_ (\oc8051_golden_model_1.B [3], _43327_, clk);
  dff _87937_ (\oc8051_golden_model_1.B [4], _43328_, clk);
  dff _87938_ (\oc8051_golden_model_1.B [5], _43329_, clk);
  dff _87939_ (\oc8051_golden_model_1.B [6], _43330_, clk);
  dff _87940_ (\oc8051_golden_model_1.B [7], _40752_, clk);
  dff _87941_ (\oc8051_golden_model_1.ACC [0], _43332_, clk);
  dff _87942_ (\oc8051_golden_model_1.ACC [1], _43333_, clk);
  dff _87943_ (\oc8051_golden_model_1.ACC [2], _43334_, clk);
  dff _87944_ (\oc8051_golden_model_1.ACC [3], _43335_, clk);
  dff _87945_ (\oc8051_golden_model_1.ACC [4], _43336_, clk);
  dff _87946_ (\oc8051_golden_model_1.ACC [5], _43338_, clk);
  dff _87947_ (\oc8051_golden_model_1.ACC [6], _43339_, clk);
  dff _87948_ (\oc8051_golden_model_1.ACC [7], _40753_, clk);
  dff _87949_ (\oc8051_golden_model_1.PCON [0], _43340_, clk);
  dff _87950_ (\oc8051_golden_model_1.PCON [1], _43342_, clk);
  dff _87951_ (\oc8051_golden_model_1.PCON [2], _43343_, clk);
  dff _87952_ (\oc8051_golden_model_1.PCON [3], _43344_, clk);
  dff _87953_ (\oc8051_golden_model_1.PCON [4], _43345_, clk);
  dff _87954_ (\oc8051_golden_model_1.PCON [5], _43346_, clk);
  dff _87955_ (\oc8051_golden_model_1.PCON [6], _43347_, clk);
  dff _87956_ (\oc8051_golden_model_1.PCON [7], _40756_, clk);
  dff _87957_ (\oc8051_golden_model_1.TMOD [0], _43349_, clk);
  dff _87958_ (\oc8051_golden_model_1.TMOD [1], _43350_, clk);
  dff _87959_ (\oc8051_golden_model_1.TMOD [2], _43351_, clk);
  dff _87960_ (\oc8051_golden_model_1.TMOD [3], _43352_, clk);
  dff _87961_ (\oc8051_golden_model_1.TMOD [4], _43353_, clk);
  dff _87962_ (\oc8051_golden_model_1.TMOD [5], _43354_, clk);
  dff _87963_ (\oc8051_golden_model_1.TMOD [6], _43355_, clk);
  dff _87964_ (\oc8051_golden_model_1.TMOD [7], _40757_, clk);
  dff _87965_ (\oc8051_golden_model_1.DPL [0], _43357_, clk);
  dff _87966_ (\oc8051_golden_model_1.DPL [1], _43358_, clk);
  dff _87967_ (\oc8051_golden_model_1.DPL [2], _43359_, clk);
  dff _87968_ (\oc8051_golden_model_1.DPL [3], _43361_, clk);
  dff _87969_ (\oc8051_golden_model_1.DPL [4], _43362_, clk);
  dff _87970_ (\oc8051_golden_model_1.DPL [5], _43363_, clk);
  dff _87971_ (\oc8051_golden_model_1.DPL [6], _43364_, clk);
  dff _87972_ (\oc8051_golden_model_1.DPL [7], _40758_, clk);
  dff _87973_ (\oc8051_golden_model_1.DPH [0], _43366_, clk);
  dff _87974_ (\oc8051_golden_model_1.DPH [1], _43367_, clk);
  dff _87975_ (\oc8051_golden_model_1.DPH [2], _43368_, clk);
  dff _87976_ (\oc8051_golden_model_1.DPH [3], _43369_, clk);
  dff _87977_ (\oc8051_golden_model_1.DPH [4], _43370_, clk);
  dff _87978_ (\oc8051_golden_model_1.DPH [5], _43371_, clk);
  dff _87979_ (\oc8051_golden_model_1.DPH [6], _43372_, clk);
  dff _87980_ (\oc8051_golden_model_1.DPH [7], _40759_, clk);
  dff _87981_ (\oc8051_golden_model_1.TL1 [0], _43374_, clk);
  dff _87982_ (\oc8051_golden_model_1.TL1 [1], _43375_, clk);
  dff _87983_ (\oc8051_golden_model_1.TL1 [2], _43376_, clk);
  dff _87984_ (\oc8051_golden_model_1.TL1 [3], _43377_, clk);
  dff _87985_ (\oc8051_golden_model_1.TL1 [4], _43378_, clk);
  dff _87986_ (\oc8051_golden_model_1.TL1 [5], _43380_, clk);
  dff _87987_ (\oc8051_golden_model_1.TL1 [6], _43381_, clk);
  dff _87988_ (\oc8051_golden_model_1.TL1 [7], _40760_, clk);
  dff _87989_ (\oc8051_golden_model_1.TL0 [0], _43382_, clk);
  dff _87990_ (\oc8051_golden_model_1.TL0 [1], _43384_, clk);
  dff _87991_ (\oc8051_golden_model_1.TL0 [2], _43385_, clk);
  dff _87992_ (\oc8051_golden_model_1.TL0 [3], _43386_, clk);
  dff _87993_ (\oc8051_golden_model_1.TL0 [4], _43387_, clk);
  dff _87994_ (\oc8051_golden_model_1.TL0 [5], _43388_, clk);
  dff _87995_ (\oc8051_golden_model_1.TL0 [6], _43389_, clk);
  dff _87996_ (\oc8051_golden_model_1.TL0 [7], _40762_, clk);
  dff _87997_ (\oc8051_golden_model_1.TCON [0], _43391_, clk);
  dff _87998_ (\oc8051_golden_model_1.TCON [1], _43392_, clk);
  dff _87999_ (\oc8051_golden_model_1.TCON [2], _43393_, clk);
  dff _88000_ (\oc8051_golden_model_1.TCON [3], _43394_, clk);
  dff _88001_ (\oc8051_golden_model_1.TCON [4], _43395_, clk);
  dff _88002_ (\oc8051_golden_model_1.TCON [5], _43396_, clk);
  dff _88003_ (\oc8051_golden_model_1.TCON [6], _43397_, clk);
  dff _88004_ (\oc8051_golden_model_1.TCON [7], _40763_, clk);
  dff _88005_ (\oc8051_golden_model_1.TH1 [0], _43399_, clk);
  dff _88006_ (\oc8051_golden_model_1.TH1 [1], _43400_, clk);
  dff _88007_ (\oc8051_golden_model_1.TH1 [2], _43401_, clk);
  dff _88008_ (\oc8051_golden_model_1.TH1 [3], _43403_, clk);
  dff _88009_ (\oc8051_golden_model_1.TH1 [4], _43404_, clk);
  dff _88010_ (\oc8051_golden_model_1.TH1 [5], _43405_, clk);
  dff _88011_ (\oc8051_golden_model_1.TH1 [6], _43406_, clk);
  dff _88012_ (\oc8051_golden_model_1.TH1 [7], _40764_, clk);
  dff _88013_ (\oc8051_golden_model_1.TH0 [0], _43408_, clk);
  dff _88014_ (\oc8051_golden_model_1.TH0 [1], _43409_, clk);
  dff _88015_ (\oc8051_golden_model_1.TH0 [2], _43410_, clk);
  dff _88016_ (\oc8051_golden_model_1.TH0 [3], _43411_, clk);
  dff _88017_ (\oc8051_golden_model_1.TH0 [4], _43412_, clk);
  dff _88018_ (\oc8051_golden_model_1.TH0 [5], _43413_, clk);
  dff _88019_ (\oc8051_golden_model_1.TH0 [6], _43414_, clk);
  dff _88020_ (\oc8051_golden_model_1.TH0 [7], _40765_, clk);
  dff _88021_ (\oc8051_golden_model_1.PC [0], _43417_, clk);
  dff _88022_ (\oc8051_golden_model_1.PC [1], _43418_, clk);
  dff _88023_ (\oc8051_golden_model_1.PC [2], _43419_, clk);
  dff _88024_ (\oc8051_golden_model_1.PC [3], _43420_, clk);
  dff _88025_ (\oc8051_golden_model_1.PC [4], _43421_, clk);
  dff _88026_ (\oc8051_golden_model_1.PC [5], _43422_, clk);
  dff _88027_ (\oc8051_golden_model_1.PC [6], _43423_, clk);
  dff _88028_ (\oc8051_golden_model_1.PC [7], _43425_, clk);
  dff _88029_ (\oc8051_golden_model_1.PC [8], _43426_, clk);
  dff _88030_ (\oc8051_golden_model_1.PC [9], _43427_, clk);
  dff _88031_ (\oc8051_golden_model_1.PC [10], _43428_, clk);
  dff _88032_ (\oc8051_golden_model_1.PC [11], _43429_, clk);
  dff _88033_ (\oc8051_golden_model_1.PC [12], _43430_, clk);
  dff _88034_ (\oc8051_golden_model_1.PC [13], _43431_, clk);
  dff _88035_ (\oc8051_golden_model_1.PC [14], _43432_, clk);
  dff _88036_ (\oc8051_golden_model_1.PC [15], _40766_, clk);
  dff _88037_ (\oc8051_golden_model_1.P2 [0], _43434_, clk);
  dff _88038_ (\oc8051_golden_model_1.P2 [1], _43435_, clk);
  dff _88039_ (\oc8051_golden_model_1.P2 [2], _43436_, clk);
  dff _88040_ (\oc8051_golden_model_1.P2 [3], _43437_, clk);
  dff _88041_ (\oc8051_golden_model_1.P2 [4], _43438_, clk);
  dff _88042_ (\oc8051_golden_model_1.P2 [5], _43440_, clk);
  dff _88043_ (\oc8051_golden_model_1.P2 [6], _43441_, clk);
  dff _88044_ (\oc8051_golden_model_1.P2 [7], _40768_, clk);
  dff _88045_ (\oc8051_golden_model_1.P3 [0], _43442_, clk);
  dff _88046_ (\oc8051_golden_model_1.P3 [1], _43444_, clk);
  dff _88047_ (\oc8051_golden_model_1.P3 [2], _43445_, clk);
  dff _88048_ (\oc8051_golden_model_1.P3 [3], _43446_, clk);
  dff _88049_ (\oc8051_golden_model_1.P3 [4], _43447_, clk);
  dff _88050_ (\oc8051_golden_model_1.P3 [5], _43448_, clk);
  dff _88051_ (\oc8051_golden_model_1.P3 [6], _43449_, clk);
  dff _88052_ (\oc8051_golden_model_1.P3 [7], _40769_, clk);
  dff _88053_ (\oc8051_golden_model_1.P0 [0], _43451_, clk);
  dff _88054_ (\oc8051_golden_model_1.P0 [1], _43452_, clk);
  dff _88055_ (\oc8051_golden_model_1.P0 [2], _43453_, clk);
  dff _88056_ (\oc8051_golden_model_1.P0 [3], _43454_, clk);
  dff _88057_ (\oc8051_golden_model_1.P0 [4], _43455_, clk);
  dff _88058_ (\oc8051_golden_model_1.P0 [5], _43456_, clk);
  dff _88059_ (\oc8051_golden_model_1.P0 [6], _43457_, clk);
  dff _88060_ (\oc8051_golden_model_1.P0 [7], _40770_, clk);
  dff _88061_ (\oc8051_golden_model_1.P1 [0], _43459_, clk);
  dff _88062_ (\oc8051_golden_model_1.P1 [1], _43460_, clk);
  dff _88063_ (\oc8051_golden_model_1.P1 [2], _43461_, clk);
  dff _88064_ (\oc8051_golden_model_1.P1 [3], _43463_, clk);
  dff _88065_ (\oc8051_golden_model_1.P1 [4], _43464_, clk);
  dff _88066_ (\oc8051_golden_model_1.P1 [5], _43465_, clk);
  dff _88067_ (\oc8051_golden_model_1.P1 [6], _43466_, clk);
  dff _88068_ (\oc8051_golden_model_1.P1 [7], _40771_, clk);
  dff _88069_ (\oc8051_golden_model_1.IP [0], _43468_, clk);
  dff _88070_ (\oc8051_golden_model_1.IP [1], _43469_, clk);
  dff _88071_ (\oc8051_golden_model_1.IP [2], _43470_, clk);
  dff _88072_ (\oc8051_golden_model_1.IP [3], _43471_, clk);
  dff _88073_ (\oc8051_golden_model_1.IP [4], _43472_, clk);
  dff _88074_ (\oc8051_golden_model_1.IP [5], _43473_, clk);
  dff _88075_ (\oc8051_golden_model_1.IP [6], _43474_, clk);
  dff _88076_ (\oc8051_golden_model_1.IP [7], _40772_, clk);
  dff _88077_ (\oc8051_golden_model_1.IE [0], _43476_, clk);
  dff _88078_ (\oc8051_golden_model_1.IE [1], _43477_, clk);
  dff _88079_ (\oc8051_golden_model_1.IE [2], _43478_, clk);
  dff _88080_ (\oc8051_golden_model_1.IE [3], _43479_, clk);
  dff _88081_ (\oc8051_golden_model_1.IE [4], _43480_, clk);
  dff _88082_ (\oc8051_golden_model_1.IE [5], _43482_, clk);
  dff _88083_ (\oc8051_golden_model_1.IE [6], _43483_, clk);
  dff _88084_ (\oc8051_golden_model_1.IE [7], _40774_, clk);
  dff _88085_ (\oc8051_golden_model_1.SCON [0], _43484_, clk);
  dff _88086_ (\oc8051_golden_model_1.SCON [1], _43486_, clk);
  dff _88087_ (\oc8051_golden_model_1.SCON [2], _43487_, clk);
  dff _88088_ (\oc8051_golden_model_1.SCON [3], _43488_, clk);
  dff _88089_ (\oc8051_golden_model_1.SCON [4], _43489_, clk);
  dff _88090_ (\oc8051_golden_model_1.SCON [5], _43490_, clk);
  dff _88091_ (\oc8051_golden_model_1.SCON [6], _43491_, clk);
  dff _88092_ (\oc8051_golden_model_1.SCON [7], _40775_, clk);
  dff _88093_ (\oc8051_golden_model_1.SP [0], _43493_, clk);
  dff _88094_ (\oc8051_golden_model_1.SP [1], _43494_, clk);
  dff _88095_ (\oc8051_golden_model_1.SP [2], _43495_, clk);
  dff _88096_ (\oc8051_golden_model_1.SP [3], _43496_, clk);
  dff _88097_ (\oc8051_golden_model_1.SP [4], _43497_, clk);
  dff _88098_ (\oc8051_golden_model_1.SP [5], _43498_, clk);
  dff _88099_ (\oc8051_golden_model_1.SP [6], _43499_, clk);
  dff _88100_ (\oc8051_golden_model_1.SP [7], _40776_, clk);
  dff _88101_ (\oc8051_golden_model_1.SBUF [0], _43501_, clk);
  dff _88102_ (\oc8051_golden_model_1.SBUF [1], _43502_, clk);
  dff _88103_ (\oc8051_golden_model_1.SBUF [2], _43503_, clk);
  dff _88104_ (\oc8051_golden_model_1.SBUF [3], _43505_, clk);
  dff _88105_ (\oc8051_golden_model_1.SBUF [4], _43506_, clk);
  dff _88106_ (\oc8051_golden_model_1.SBUF [5], _43507_, clk);
  dff _88107_ (\oc8051_golden_model_1.SBUF [6], _43508_, clk);
  dff _88108_ (\oc8051_golden_model_1.SBUF [7], _40777_, clk);
  dff _88109_ (\oc8051_golden_model_1.PSW [0], _43510_, clk);
  dff _88110_ (\oc8051_golden_model_1.PSW [1], _43511_, clk);
  dff _88111_ (\oc8051_golden_model_1.PSW [2], _43512_, clk);
  dff _88112_ (\oc8051_golden_model_1.PSW [3], _43513_, clk);
  dff _88113_ (\oc8051_golden_model_1.PSW [4], _43514_, clk);
  dff _88114_ (\oc8051_golden_model_1.PSW [5], _43515_, clk);
  dff _88115_ (\oc8051_golden_model_1.PSW [6], _43516_, clk);
  dff _88116_ (\oc8051_golden_model_1.PSW [7], _40778_, clk);
  dff _88117_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _02832_, clk);
  dff _88118_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _02844_, clk);
  dff _88119_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _02866_, clk);
  dff _88120_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _02890_, clk);
  dff _88121_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _02914_, clk);
  dff _88122_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _00956_, clk);
  dff _88123_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _02924_, clk);
  dff _88124_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _00925_, clk);
  dff _88125_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _02936_, clk);
  dff _88126_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _02948_, clk);
  dff _88127_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _02960_, clk);
  dff _88128_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _02971_, clk);
  dff _88129_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _02984_, clk);
  dff _88130_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _02997_, clk);
  dff _88131_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _03011_, clk);
  dff _88132_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _00976_, clk);
  dff _88133_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _02356_, clk);
  dff _88134_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _22216_, clk);
  dff _88135_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _02542_, clk);
  dff _88136_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _02695_, clk);
  dff _88137_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _02877_, clk);
  dff _88138_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _03117_, clk);
  dff _88139_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _03361_, clk);
  dff _88140_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _03562_, clk);
  dff _88141_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _03757_, clk);
  dff _88142_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _03954_, clk);
  dff _88143_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _04054_, clk);
  dff _88144_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _04147_, clk);
  dff _88145_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _04246_, clk);
  dff _88146_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _04345_, clk);
  dff _88147_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _04444_, clk);
  dff _88148_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _04542_, clk);
  dff _88149_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [14], _04641_, clk);
  dff _88150_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [15], _24374_, clk);
  dff _88151_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _38968_, clk);
  dff _88152_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _38969_, clk);
  dff _88153_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _38970_, clk);
  dff _88154_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _38971_, clk);
  dff _88155_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _38972_, clk);
  dff _88156_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _38973_, clk);
  dff _88157_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _38974_, clk);
  dff _88158_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _38955_, clk);
  dff _88159_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _38975_, clk);
  dff _88160_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _38976_, clk);
  dff _88161_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _38978_, clk);
  dff _88162_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], _38979_, clk);
  dff _88163_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _38980_, clk);
  dff _88164_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _38981_, clk);
  dff _88165_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _38982_, clk);
  dff _88166_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _38956_, clk);
  dff _88167_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _38984_, clk);
  dff _88168_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], _38985_, clk);
  dff _88169_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], _38986_, clk);
  dff _88170_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _38987_, clk);
  dff _88171_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _38988_, clk);
  dff _88172_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _38990_, clk);
  dff _88173_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _38991_, clk);
  dff _88174_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _38958_, clk);
  dff _88175_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _34275_, clk);
  dff _88176_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _34278_, clk);
  dff _88177_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _09716_, clk);
  dff _88178_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _34280_, clk);
  dff _88179_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _34282_, clk);
  dff _88180_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _09719_, clk);
  dff _88181_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _34284_, clk);
  dff _88182_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _09722_, clk);
  dff _88183_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _34286_, clk);
  dff _88184_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _34288_, clk);
  dff _88185_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _34290_, clk);
  dff _88186_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _09725_, clk);
  dff _88187_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _34292_, clk);
  dff _88188_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _09728_, clk);
  dff _88189_ (\oc8051_top_1.oc8051_decoder1.wr , _09731_, clk);
  dff _88190_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _09790_, clk);
  dff _88191_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _09792_, clk);
  dff _88192_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _09695_, clk);
  dff _88193_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _09795_, clk);
  dff _88194_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _09798_, clk);
  dff _88195_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _09698_, clk);
  dff _88196_ (\oc8051_top_1.oc8051_decoder1.state [0], _09801_, clk);
  dff _88197_ (\oc8051_top_1.oc8051_decoder1.state [1], _09701_, clk);
  dff _88198_ (\oc8051_top_1.oc8051_decoder1.op [0], _09804_, clk);
  dff _88199_ (\oc8051_top_1.oc8051_decoder1.op [1], _09807_, clk);
  dff _88200_ (\oc8051_top_1.oc8051_decoder1.op [2], _09810_, clk);
  dff _88201_ (\oc8051_top_1.oc8051_decoder1.op [3], _09813_, clk);
  dff _88202_ (\oc8051_top_1.oc8051_decoder1.op [4], _09816_, clk);
  dff _88203_ (\oc8051_top_1.oc8051_decoder1.op [5], _09819_, clk);
  dff _88204_ (\oc8051_top_1.oc8051_decoder1.op [6], _09822_, clk);
  dff _88205_ (\oc8051_top_1.oc8051_decoder1.op [7], _09704_, clk);
  dff _88206_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _09707_, clk);
  dff _88207_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _34273_, clk);
  dff _88208_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _09713_, clk);
  dff _88209_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _09825_, clk);
  dff _88210_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _09710_, clk);
  dff _88211_ (\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , _39760_, clk);
  dff _88212_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _39792_, clk);
  dff _88213_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _39793_, clk);
  dff _88214_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _39794_, clk);
  dff _88215_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _39795_, clk);
  dff _88216_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _39796_, clk);
  dff _88217_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _39797_, clk);
  dff _88218_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _39798_, clk);
  dff _88219_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _39762_, clk);
  dff _88220_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _39799_, clk);
  dff _88221_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _39800_, clk);
  dff _88222_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _39801_, clk);
  dff _88223_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _39803_, clk);
  dff _88224_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _39804_, clk);
  dff _88225_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _39805_, clk);
  dff _88226_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _39806_, clk);
  dff _88227_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _39763_, clk);
  dff _88228_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _39807_, clk);
  dff _88229_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _39808_, clk);
  dff _88230_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _39809_, clk);
  dff _88231_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _39810_, clk);
  dff _88232_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _39811_, clk);
  dff _88233_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _39812_, clk);
  dff _88234_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _39814_, clk);
  dff _88235_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _39764_, clk);
  dff _88236_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _39815_, clk);
  dff _88237_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _39816_, clk);
  dff _88238_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _39817_, clk);
  dff _88239_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _39818_, clk);
  dff _88240_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _39819_, clk);
  dff _88241_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _39820_, clk);
  dff _88242_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _39821_, clk);
  dff _88243_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _39765_, clk);
  dff _88244_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _39339_, clk);
  dff _88245_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _39340_, clk);
  dff _88246_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _39341_, clk);
  dff _88247_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _39342_, clk);
  dff _88248_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _39056_, clk);
  dff _88249_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _39128_, clk);
  dff _88250_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _39129_, clk);
  dff _88251_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _39130_, clk);
  dff _88252_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _39131_, clk);
  dff _88253_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _39132_, clk);
  dff _88254_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _39134_, clk);
  dff _88255_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _39135_, clk);
  dff _88256_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _39136_, clk);
  dff _88257_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _39137_, clk);
  dff _88258_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _39138_, clk);
  dff _88259_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _39139_, clk);
  dff _88260_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _39140_, clk);
  dff _88261_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _39141_, clk);
  dff _88262_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _39142_, clk);
  dff _88263_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _39143_, clk);
  dff _88264_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _39015_, clk);
  dff _88265_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _39148_, clk);
  dff _88266_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _39149_, clk);
  dff _88267_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _39150_, clk);
  dff _88268_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _39151_, clk);
  dff _88269_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _39152_, clk);
  dff _88270_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _39153_, clk);
  dff _88271_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _39154_, clk);
  dff _88272_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _39155_, clk);
  dff _88273_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _39156_, clk);
  dff _88274_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _39157_, clk);
  dff _88275_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _39159_, clk);
  dff _88276_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _39160_, clk);
  dff _88277_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _39161_, clk);
  dff _88278_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _39162_, clk);
  dff _88279_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _39163_, clk);
  dff _88280_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _39016_, clk);
  dff _88281_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _39343_, clk);
  dff _88282_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _39344_, clk);
  dff _88283_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _39345_, clk);
  dff _88284_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _39346_, clk);
  dff _88285_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _39348_, clk);
  dff _88286_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _39349_, clk);
  dff _88287_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _39350_, clk);
  dff _88288_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _39351_, clk);
  dff _88289_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _39352_, clk);
  dff _88290_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _39353_, clk);
  dff _88291_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _39354_, clk);
  dff _88292_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _39355_, clk);
  dff _88293_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _39356_, clk);
  dff _88294_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _39357_, clk);
  dff _88295_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _39359_, clk);
  dff _88296_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _39360_, clk);
  dff _88297_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _39361_, clk);
  dff _88298_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _39362_, clk);
  dff _88299_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _39363_, clk);
  dff _88300_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _39364_, clk);
  dff _88301_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _39365_, clk);
  dff _88302_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _39366_, clk);
  dff _88303_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _39367_, clk);
  dff _88304_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _39368_, clk);
  dff _88305_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _39370_, clk);
  dff _88306_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _39371_, clk);
  dff _88307_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _39372_, clk);
  dff _88308_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _39373_, clk);
  dff _88309_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _39374_, clk);
  dff _88310_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _39375_, clk);
  dff _88311_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _39376_, clk);
  dff _88312_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _39081_, clk);
  dff _88313_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _39054_, clk);
  dff _88314_ (\oc8051_top_1.oc8051_memory_interface1.dack_ir , 1'b0, clk);
  dff _88315_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _39377_, clk);
  dff _88316_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _39379_, clk);
  dff _88317_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _39380_, clk);
  dff _88318_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _39381_, clk);
  dff _88319_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _39382_, clk);
  dff _88320_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _39383_, clk);
  dff _88321_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _39385_, clk);
  dff _88322_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _39057_, clk);
  dff _88323_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _39386_, clk);
  dff _88324_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _39387_, clk);
  dff _88325_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _39388_, clk);
  dff _88326_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _39389_, clk);
  dff _88327_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _39390_, clk);
  dff _88328_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _39391_, clk);
  dff _88329_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _39392_, clk);
  dff _88330_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _39058_, clk);
  dff _88331_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _39393_, clk);
  dff _88332_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _39394_, clk);
  dff _88333_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _39396_, clk);
  dff _88334_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _39397_, clk);
  dff _88335_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _39398_, clk);
  dff _88336_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _39399_, clk);
  dff _88337_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _39400_, clk);
  dff _88338_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], _39060_, clk);
  dff _88339_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _39061_, clk);
  dff _88340_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _39062_, clk);
  dff _88341_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [0], _39401_, clk);
  dff _88342_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [1], _39402_, clk);
  dff _88343_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [2], _39403_, clk);
  dff _88344_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [3], _39404_, clk);
  dff _88345_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [4], _39405_, clk);
  dff _88346_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [5], _39407_, clk);
  dff _88347_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [6], _39408_, clk);
  dff _88348_ (\oc8051_top_1.oc8051_memory_interface1.ddat_ir [7], _39063_, clk);
  dff _88349_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _39409_, clk);
  dff _88350_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _39410_, clk);
  dff _88351_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _39411_, clk);
  dff _88352_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _39412_, clk);
  dff _88353_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _39413_, clk);
  dff _88354_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _39414_, clk);
  dff _88355_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _39415_, clk);
  dff _88356_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _39416_, clk);
  dff _88357_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _39418_, clk);
  dff _88358_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _39419_, clk);
  dff _88359_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _39420_, clk);
  dff _88360_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _39421_, clk);
  dff _88361_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _39422_, clk);
  dff _88362_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _39423_, clk);
  dff _88363_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _39424_, clk);
  dff _88364_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _39064_, clk);
  dff _88365_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _39425_, clk);
  dff _88366_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _39426_, clk);
  dff _88367_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _39427_, clk);
  dff _88368_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _39429_, clk);
  dff _88369_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _39430_, clk);
  dff _88370_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _39431_, clk);
  dff _88371_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _39432_, clk);
  dff _88372_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _39433_, clk);
  dff _88373_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _39434_, clk);
  dff _88374_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _39435_, clk);
  dff _88375_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _39436_, clk);
  dff _88376_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _39437_, clk);
  dff _88377_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _39438_, clk);
  dff _88378_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _39440_, clk);
  dff _88379_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _39441_, clk);
  dff _88380_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _39066_, clk);
  dff _88381_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _39067_, clk);
  dff _88382_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _39069_, clk);
  dff _88383_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _39068_, clk);
  dff _88384_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _39442_, clk);
  dff _88385_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _39443_, clk);
  dff _88386_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _39444_, clk);
  dff _88387_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _39445_, clk);
  dff _88388_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _39446_, clk);
  dff _88389_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _39447_, clk);
  dff _88390_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _39448_, clk);
  dff _88391_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _39071_, clk);
  dff _88392_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _39449_, clk);
  dff _88393_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _39450_, clk);
  dff _88394_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _39072_, clk);
  dff _88395_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], _39451_, clk);
  dff _88396_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], _39452_, clk);
  dff _88397_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], _39453_, clk);
  dff _88398_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], _39454_, clk);
  dff _88399_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], _39455_, clk);
  dff _88400_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], _39456_, clk);
  dff _88401_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], _39457_, clk);
  dff _88402_ (\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], _39073_, clk);
  dff _88403_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], _39458_, clk);
  dff _88404_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _39459_, clk);
  dff _88405_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _39461_, clk);
  dff _88406_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], _39462_, clk);
  dff _88407_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], _39463_, clk);
  dff _88408_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], _39464_, clk);
  dff _88409_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], _39465_, clk);
  dff _88410_ (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _39074_, clk);
  dff _88411_ (\oc8051_top_1.oc8051_memory_interface1.reti , _39075_, clk);
  dff _88412_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _39466_, clk);
  dff _88413_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _39467_, clk);
  dff _88414_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _39468_, clk);
  dff _88415_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _39469_, clk);
  dff _88416_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _39470_, clk);
  dff _88417_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _39472_, clk);
  dff _88418_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _39473_, clk);
  dff _88419_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _39076_, clk);
  dff _88420_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _39078_, clk);
  dff _88421_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _39079_, clk);
  dff _88422_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _39474_, clk);
  dff _88423_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _39475_, clk);
  dff _88424_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _39476_, clk);
  dff _88425_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _39080_, clk);
  dff _88426_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _39477_, clk);
  dff _88427_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _39478_, clk);
  dff _88428_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _39479_, clk);
  dff _88429_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _39480_, clk);
  dff _88430_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _39481_, clk);
  dff _88431_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _39483_, clk);
  dff _88432_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _39484_, clk);
  dff _88433_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _39485_, clk);
  dff _88434_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _39486_, clk);
  dff _88435_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _39487_, clk);
  dff _88436_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _39488_, clk);
  dff _88437_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _39489_, clk);
  dff _88438_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _39490_, clk);
  dff _88439_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _39491_, clk);
  dff _88440_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _39492_, clk);
  dff _88441_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _39494_, clk);
  dff _88442_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _39495_, clk);
  dff _88443_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _39496_, clk);
  dff _88444_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _39497_, clk);
  dff _88445_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _39498_, clk);
  dff _88446_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _39499_, clk);
  dff _88447_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _39500_, clk);
  dff _88448_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _39501_, clk);
  dff _88449_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _39502_, clk);
  dff _88450_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _39503_, clk);
  dff _88451_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _39505_, clk);
  dff _88452_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _39506_, clk);
  dff _88453_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _39507_, clk);
  dff _88454_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _39508_, clk);
  dff _88455_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _39509_, clk);
  dff _88456_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _39510_, clk);
  dff _88457_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _39082_, clk);
  dff _88458_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [0], _39511_, clk);
  dff _88459_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [1], _39512_, clk);
  dff _88460_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [2], _39513_, clk);
  dff _88461_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [3], _39514_, clk);
  dff _88462_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [4], _39516_, clk);
  dff _88463_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [5], _39517_, clk);
  dff _88464_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [6], _39518_, clk);
  dff _88465_ (\oc8051_top_1.oc8051_memory_interface1.ddat_o [7], _39083_, clk);
  dff _88466_ (\oc8051_top_1.oc8051_memory_interface1.dwe_o , _39084_, clk);
  dff _88467_ (\oc8051_top_1.oc8051_memory_interface1.dstb_o , _39086_, clk);
  dff _88468_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [0], _39519_, clk);
  dff _88469_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [1], _39520_, clk);
  dff _88470_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [2], _39521_, clk);
  dff _88471_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [3], _39522_, clk);
  dff _88472_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [4], _39523_, clk);
  dff _88473_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [5], _39524_, clk);
  dff _88474_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [6], _39525_, clk);
  dff _88475_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [7], _39527_, clk);
  dff _88476_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [8], _39528_, clk);
  dff _88477_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [9], _39529_, clk);
  dff _88478_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [10], _39530_, clk);
  dff _88479_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [11], _39531_, clk);
  dff _88480_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [12], _39532_, clk);
  dff _88481_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [13], _39533_, clk);
  dff _88482_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [14], _39534_, clk);
  dff _88483_ (\oc8051_top_1.oc8051_memory_interface1.dadr_ot [15], _39087_, clk);
  dff _88484_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _39088_, clk);
  dff _88485_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _39089_, clk);
  dff _88486_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _39090_, clk);
  dff _88487_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _39535_, clk);
  dff _88488_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _39536_, clk);
  dff _88489_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _39538_, clk);
  dff _88490_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _39539_, clk);
  dff _88491_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [4], _39540_, clk);
  dff _88492_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [5], _39541_, clk);
  dff _88493_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [6], _39542_, clk);
  dff _88494_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [7], _39543_, clk);
  dff _88495_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [8], _39544_, clk);
  dff _88496_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [9], _39545_, clk);
  dff _88497_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [10], _39546_, clk);
  dff _88498_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [11], _39547_, clk);
  dff _88499_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [12], _39549_, clk);
  dff _88500_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [13], _39550_, clk);
  dff _88501_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [14], _39551_, clk);
  dff _88502_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [15], _39091_, clk);
  dff _88503_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _39092_, clk);
  dff _88504_ (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _40015_, clk);
  dff _88505_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _40036_, clk);
  dff _88506_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _40037_, clk);
  dff _88507_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _40039_, clk);
  dff _88508_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _40040_, clk);
  dff _88509_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _40041_, clk);
  dff _88510_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _40042_, clk);
  dff _88511_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _40043_, clk);
  dff _88512_ (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _40016_, clk);
  dff _88513_ (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _40018_, clk);
  dff _88514_ (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _40044_, clk);
  dff _88515_ (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _40045_, clk);
  dff _88516_ (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _40019_, clk);
  dff _88517_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _03167_, clk);
  dff _88518_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _03171_, clk);
  dff _88519_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _03175_, clk);
  dff _88520_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03179_, clk);
  dff _88521_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03183_, clk);
  dff _88522_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03187_, clk);
  dff _88523_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03191_, clk);
  dff _88524_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _03194_, clk);
  dff _88525_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _03134_, clk);
  dff _88526_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _03138_, clk);
  dff _88527_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _03142_, clk);
  dff _88528_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _03146_, clk);
  dff _88529_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _03150_, clk);
  dff _88530_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03154_, clk);
  dff _88531_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03158_, clk);
  dff _88532_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _03161_, clk);
  dff _88533_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _02796_, clk);
  dff _88534_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _02801_, clk);
  dff _88535_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _02806_, clk);
  dff _88536_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _02811_, clk);
  dff _88537_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _02815_, clk);
  dff _88538_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _02820_, clk);
  dff _88539_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _02825_, clk);
  dff _88540_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _02827_, clk);
  dff _88541_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _02835_, clk);
  dff _88542_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _02838_, clk);
  dff _88543_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _02841_, clk);
  dff _88544_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _02845_, clk);
  dff _88545_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _02849_, clk);
  dff _88546_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _02852_, clk);
  dff _88547_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _02855_, clk);
  dff _88548_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _02858_, clk);
  dff _88549_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _02864_, clk);
  dff _88550_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _02868_, clk);
  dff _88551_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _02871_, clk);
  dff _88552_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _02875_, clk);
  dff _88553_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _02878_, clk);
  dff _88554_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _02882_, clk);
  dff _88555_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _02885_, clk);
  dff _88556_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _02888_, clk);
  dff _88557_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _02926_, clk);
  dff _88558_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _02929_, clk);
  dff _88559_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _02933_, clk);
  dff _88560_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _02937_, clk);
  dff _88561_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _02940_, clk);
  dff _88562_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _02943_, clk);
  dff _88563_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _02947_, clk);
  dff _88564_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _02950_, clk);
  dff _88565_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _02894_, clk);
  dff _88566_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _02898_, clk);
  dff _88567_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _02902_, clk);
  dff _88568_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _02905_, clk);
  dff _88569_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _02909_, clk);
  dff _88570_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _02912_, clk);
  dff _88571_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _02916_, clk);
  dff _88572_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _02919_, clk);
  dff _88573_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _03071_, clk);
  dff _88574_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _03074_, clk);
  dff _88575_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _03078_, clk);
  dff _88576_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _03081_, clk);
  dff _88577_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _03085_, clk);
  dff _88578_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _03089_, clk);
  dff _88579_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _03093_, clk);
  dff _88580_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _03096_, clk);
  dff _88581_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _03045_, clk);
  dff _88582_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _03048_, clk);
  dff _88583_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _03051_, clk);
  dff _88584_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _03054_, clk);
  dff _88585_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _03058_, clk);
  dff _88586_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _03061_, clk);
  dff _88587_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _03064_, clk);
  dff _88588_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _03067_, clk);
  dff _88589_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _03014_, clk);
  dff _88590_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _03018_, clk);
  dff _88591_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _03021_, clk);
  dff _88592_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _03025_, clk);
  dff _88593_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _03028_, clk);
  dff _88594_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _03032_, clk);
  dff _88595_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _03036_, clk);
  dff _88596_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _03038_, clk);
  dff _88597_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _02983_, clk);
  dff _88598_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _02987_, clk);
  dff _88599_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _02991_, clk);
  dff _88600_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _02994_, clk);
  dff _88601_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _02999_, clk);
  dff _88602_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _03002_, clk);
  dff _88603_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _03006_, clk);
  dff _88604_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _03009_, clk);
  dff _88605_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _02954_, clk);
  dff _88606_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _02957_, clk);
  dff _88607_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _02962_, clk);
  dff _88608_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _02965_, clk);
  dff _88609_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _02968_, clk);
  dff _88610_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _02972_, clk);
  dff _88611_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _02976_, clk);
  dff _88612_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _02978_, clk);
  dff _88613_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _03101_, clk);
  dff _88614_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _03105_, clk);
  dff _88615_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _03109_, clk);
  dff _88616_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _03113_, clk);
  dff _88617_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _03118_, clk);
  dff _88618_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _03122_, clk);
  dff _88619_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _03126_, clk);
  dff _88620_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _03129_, clk);
  dff _88621_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _03263_, clk);
  dff _88622_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _03267_, clk);
  dff _88623_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03271_, clk);
  dff _88624_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03275_, clk);
  dff _88625_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _03279_, clk);
  dff _88626_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03283_, clk);
  dff _88627_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03287_, clk);
  dff _88628_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _02573_, clk);
  dff _88629_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03231_, clk);
  dff _88630_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03235_, clk);
  dff _88631_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _03239_, clk);
  dff _88632_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03243_, clk);
  dff _88633_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _03247_, clk);
  dff _88634_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03251_, clk);
  dff _88635_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03255_, clk);
  dff _88636_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _03258_, clk);
  dff _88637_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03199_, clk);
  dff _88638_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _03203_, clk);
  dff _88639_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03207_, clk);
  dff _88640_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03211_, clk);
  dff _88641_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _03215_, clk);
  dff _88642_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03219_, clk);
  dff _88643_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _03223_, clk);
  dff _88644_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _03226_, clk);
  dff _88645_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _05081_, clk);
  dff _88646_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _05083_, clk);
  dff _88647_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _05084_, clk);
  dff _88648_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _05086_, clk);
  dff _88649_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _05088_, clk);
  dff _88650_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _05090_, clk);
  dff _88651_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _05092_, clk);
  dff _88652_ (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _02563_, clk);
  dff _88653_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0], clk);
  dff _88654_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1], clk);
  dff _88655_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2], clk);
  dff _88656_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3], clk);
  dff _88657_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4], clk);
  dff _88658_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5], clk);
  dff _88659_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6], clk);
  dff _88660_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7], clk);
  dff _88661_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8], clk);
  dff _88662_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9], clk);
  dff _88663_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10], clk);
  dff _88664_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11], clk);
  dff _88665_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12], clk);
  dff _88666_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13], clk);
  dff _88667_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14], clk);
  dff _88668_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15], clk);
  dff _88669_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16], clk);
  dff _88670_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17], clk);
  dff _88671_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18], clk);
  dff _88672_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19], clk);
  dff _88673_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20], clk);
  dff _88674_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21], clk);
  dff _88675_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22], clk);
  dff _88676_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23], clk);
  dff _88677_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24], clk);
  dff _88678_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25], clk);
  dff _88679_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26], clk);
  dff _88680_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27], clk);
  dff _88681_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28], clk);
  dff _88682_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29], clk);
  dff _88683_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30], clk);
  dff _88684_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31], clk);
  dff _88685_ (\oc8051_top_1.oc8051_rom1.ea_int , 1'b1, clk);
  dff _88686_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _39849_, clk);
  dff _88687_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _39935_, clk);
  dff _88688_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _39936_, clk);
  dff _88689_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _39937_, clk);
  dff _88690_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _39850_, clk);
  dff _88691_ (\oc8051_top_1.oc8051_sfr1.bit_out , _39851_, clk);
  dff _88692_ (\oc8051_top_1.oc8051_sfr1.wait_data , _39853_, clk);
  dff _88693_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _39938_, clk);
  dff _88694_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _39939_, clk);
  dff _88695_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _39940_, clk);
  dff _88696_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _39941_, clk);
  dff _88697_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _39943_, clk);
  dff _88698_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _39944_, clk);
  dff _88699_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _39945_, clk);
  dff _88700_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _39854_, clk);
  dff _88701_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _39855_, clk);
  dff _88702_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _19849_, clk);
  dff _88703_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _19860_, clk);
  dff _88704_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _19872_, clk);
  dff _88705_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _19884_, clk);
  dff _88706_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _19896_, clk);
  dff _88707_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _19908_, clk);
  dff _88708_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _19920_, clk);
  dff _88709_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _17998_, clk);
  dff _88710_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _08903_, clk);
  dff _88711_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _08914_, clk);
  dff _88712_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _08925_, clk);
  dff _88713_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _08936_, clk);
  dff _88714_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _08947_, clk);
  dff _88715_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _08958_, clk);
  dff _88716_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _08969_, clk);
  dff _88717_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _06662_, clk);
  dff _88718_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _13647_, clk);
  dff _88719_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _13657_, clk);
  dff _88720_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _13668_, clk);
  dff _88721_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _13679_, clk);
  dff _88722_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _13690_, clk);
  dff _88723_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _13701_, clk);
  dff _88724_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _13712_, clk);
  dff _88725_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _12713_, clk);
  dff _88726_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13723_, clk);
  dff _88727_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _13733_, clk);
  dff _88728_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _13744_, clk);
  dff _88729_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _13755_, clk);
  dff _88730_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _13766_, clk);
  dff _88731_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _13777_, clk);
  dff _88732_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _13788_, clk);
  dff _88733_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _12734_, clk);
  dff _88734_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _42886_, clk);
  dff _88735_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , _42885_, clk);
  dff _88736_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie0_buff , 1'b0, clk);
  dff _88737_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie1_buff , _42882_, clk);
  dff _88738_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00130_, clk);
  dff _88739_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00132_, clk);
  dff _88740_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00134_, clk);
  dff _88741_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00136_, clk);
  dff _88742_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00138_, clk);
  dff _88743_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00140_, clk);
  dff _88744_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00141_, clk);
  dff _88745_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _42880_, clk);
  dff _88746_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00143_, clk);
  dff _88747_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _42879_, clk);
  dff _88748_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _42877_, clk);
  dff _88749_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00145_, clk);
  dff _88750_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00147_, clk);
  dff _88751_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _42875_, clk);
  dff _88752_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00149_, clk);
  dff _88753_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00151_, clk);
  dff _88754_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _42873_, clk);
  dff _88755_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00152_, clk);
  dff _88756_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [1], _42872_, clk);
  dff _88757_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00154_, clk);
  dff _88758_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [1], _42870_, clk);
  dff _88759_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _42840_, clk);
  dff _88760_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _42838_, clk);
  dff _88761_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _42836_, clk);
  dff _88762_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _42834_, clk);
  dff _88763_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00156_, clk);
  dff _88764_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00158_, clk);
  dff _88765_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00160_, clk);
  dff _88766_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _42832_, clk);
  dff _88767_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00162_, clk);
  dff _88768_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00163_, clk);
  dff _88769_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00165_, clk);
  dff _88770_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00167_, clk);
  dff _88771_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00169_, clk);
  dff _88772_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00171_, clk);
  dff _88773_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00173_, clk);
  dff _88774_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _42830_, clk);
  dff _88775_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00174_, clk);
  dff _88776_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00176_, clk);
  dff _88777_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00178_, clk);
  dff _88778_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00180_, clk);
  dff _88779_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00182_, clk);
  dff _88780_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00184_, clk);
  dff _88781_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00185_, clk);
  dff _88782_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _42827_, clk);
  dff _88783_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _40589_, clk);
  dff _88784_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _40591_, clk);
  dff _88785_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _40593_, clk);
  dff _88786_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _40595_, clk);
  dff _88787_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _40597_, clk);
  dff _88788_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _40599_, clk);
  dff _88789_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _40601_, clk);
  dff _88790_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _31126_, clk);
  dff _88791_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _40603_, clk);
  dff _88792_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _40605_, clk);
  dff _88793_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _40607_, clk);
  dff _88794_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _40609_, clk);
  dff _88795_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _40611_, clk);
  dff _88796_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _40612_, clk);
  dff _88797_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _40614_, clk);
  dff _88798_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _31149_, clk);
  dff _88799_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _40616_, clk);
  dff _88800_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _40618_, clk);
  dff _88801_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _40620_, clk);
  dff _88802_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _40622_, clk);
  dff _88803_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _40624_, clk);
  dff _88804_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _40626_, clk);
  dff _88805_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _40628_, clk);
  dff _88806_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _31172_, clk);
  dff _88807_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _40630_, clk);
  dff _88808_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _40632_, clk);
  dff _88809_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _40634_, clk);
  dff _88810_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _40636_, clk);
  dff _88811_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _40638_, clk);
  dff _88812_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _40640_, clk);
  dff _88813_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _40642_, clk);
  dff _88814_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _31194_, clk);
  dff _88815_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _17374_, clk);
  dff _88816_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _17385_, clk);
  dff _88817_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _17396_, clk);
  dff _88818_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _17407_, clk);
  dff _88819_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _17418_, clk);
  dff _88820_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _17429_, clk);
  dff _88821_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _15193_, clk);
  dff _88822_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _09519_, clk);
  dff _88823_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _10696_, clk);
  dff _88824_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _10707_, clk);
  dff _88825_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _10718_, clk);
  dff _88826_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _10729_, clk);
  dff _88827_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _10740_, clk);
  dff _88828_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _10751_, clk);
  dff _88829_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _10762_, clk);
  dff _88830_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _09540_, clk);
  dff _88831_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _41092_, clk);
  dff _88832_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _41095_, clk);
  dff _88833_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _41601_, clk);
  dff _88834_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _41603_, clk);
  dff _88835_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _41605_, clk);
  dff _88836_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _41606_, clk);
  dff _88837_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _41608_, clk);
  dff _88838_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _41610_, clk);
  dff _88839_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _41612_, clk);
  dff _88840_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _41098_, clk);
  dff _88841_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _41614_, clk);
  dff _88842_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _41616_, clk);
  dff _88843_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _41618_, clk);
  dff _88844_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _41620_, clk);
  dff _88845_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _41622_, clk);
  dff _88846_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _41623_, clk);
  dff _88847_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _41625_, clk);
  dff _88848_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _41101_, clk);
  dff _88849_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _41104_, clk);
  dff _88850_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _41107_, clk);
  dff _88851_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _41627_, clk);
  dff _88852_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _41629_, clk);
  dff _88853_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _41631_, clk);
  dff _88854_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _41633_, clk);
  dff _88855_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _41635_, clk);
  dff _88856_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _41637_, clk);
  dff _88857_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _41638_, clk);
  dff _88858_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _41110_, clk);
  dff _88859_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _41640_, clk);
  dff _88860_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _41642_, clk);
  dff _88861_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _41644_, clk);
  dff _88862_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _41646_, clk);
  dff _88863_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _41648_, clk);
  dff _88864_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _41650_, clk);
  dff _88865_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _41652_, clk);
  dff _88866_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _41113_, clk);
  dff _88867_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _41116_, clk);
  dff _88868_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _41653_, clk);
  dff _88869_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _41655_, clk);
  dff _88870_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _41657_, clk);
  dff _88871_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _41659_, clk);
  dff _88872_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _41660_, clk);
  dff _88873_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _41662_, clk);
  dff _88874_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _41664_, clk);
  dff _88875_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _41119_, clk);
  dff _88876_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01628_, clk);
  dff _88877_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01631_, clk);
  dff _88878_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01634_, clk);
  dff _88879_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01637_, clk);
  dff _88880_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _02108_, clk);
  dff _88881_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _02109_, clk);
  dff _88882_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _02111_, clk);
  dff _88883_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _02113_, clk);
  dff _88884_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _02115_, clk);
  dff _88885_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _02116_, clk);
  dff _88886_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _02118_, clk);
  dff _88887_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01640_, clk);
  dff _88888_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _02120_, clk);
  dff _88889_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _02122_, clk);
  dff _88890_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _02123_, clk);
  dff _88891_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _02125_, clk);
  dff _88892_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _02127_, clk);
  dff _88893_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _02129_, clk);
  dff _88894_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _02130_, clk);
  dff _88895_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01643_, clk);
  dff _88896_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01646_, clk);
  dff _88897_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _02132_, clk);
  dff _88898_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _02134_, clk);
  dff _88899_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _02136_, clk);
  dff _88900_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _02137_, clk);
  dff _88901_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _02139_, clk);
  dff _88902_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _02141_, clk);
  dff _88903_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _02143_, clk);
  dff _88904_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01649_, clk);
  dff _88905_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _02144_, clk);
  dff _88906_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _02145_, clk);
  dff _88907_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _02146_, clk);
  dff _88908_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _02147_, clk);
  dff _88909_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _02148_, clk);
  dff _88910_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _02149_, clk);
  dff _88911_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _02150_, clk);
  dff _88912_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01652_, clk);
  dff _88913_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01655_, clk);
  dff _88914_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _02151_, clk);
  dff _88915_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _02152_, clk);
  dff _88916_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _02153_, clk);
  dff _88917_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _02154_, clk);
  dff _88918_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _02155_, clk);
  dff _88919_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _02156_, clk);
  dff _88920_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _02157_, clk);
  dff _88921_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01658_, clk);
  dff _88922_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _01210_, clk);
  dff _88923_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _01212_, clk);
  dff _88924_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _01214_, clk);
  dff _88925_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _01216_, clk);
  dff _88926_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01218_, clk);
  dff _88927_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01220_, clk);
  dff _88928_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _01222_, clk);
  dff _88929_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _01224_, clk);
  dff _88930_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _01226_, clk);
  dff _88931_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _01228_, clk);
  dff _88932_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _01229_, clk);
  dff _88933_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00567_, clk);
  dff _88934_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _00543_, clk);
  dff _88935_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _00546_, clk);
  dff _88936_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00548_, clk);
  dff _88937_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _00551_, clk);
  dff _88938_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _00554_, clk);
  dff _88939_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _00556_, clk);
  dff _88940_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _01231_, clk);
  dff _88941_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _00559_, clk);
  dff _88942_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01233_, clk);
  dff _88943_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _01235_, clk);
  dff _88944_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01237_, clk);
  dff _88945_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _00562_, clk);
  dff _88946_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _01239_, clk);
  dff _88947_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01241_, clk);
  dff _88948_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01243_, clk);
  dff _88949_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01245_, clk);
  dff _88950_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01247_, clk);
  dff _88951_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01249_, clk);
  dff _88952_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01251_, clk);
  dff _88953_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00564_, clk);
  dff _88954_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _00570_, clk);
  dff _88955_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _00572_, clk);
  dff _88956_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd , _00575_, clk);
  dff _88957_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _00578_, clk);
  dff _88958_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _00580_, clk);
  dff _88959_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01253_, clk);
  dff _88960_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _01255_, clk);
  dff _88961_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01257_, clk);
  dff _88962_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _00583_, clk);
  dff _88963_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _01259_, clk);
  dff _88964_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _01261_, clk);
  dff _88965_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _01263_, clk);
  dff _88966_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _01264_, clk);
  dff _88967_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _01266_, clk);
  dff _88968_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _01268_, clk);
  dff _88969_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _01270_, clk);
  dff _88970_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _01272_, clk);
  dff _88971_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _01274_, clk);
  dff _88972_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _01276_, clk);
  dff _88973_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00586_, clk);
  dff _88974_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _01278_, clk);
  dff _88975_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _01280_, clk);
  dff _88976_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _01282_, clk);
  dff _88977_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _01284_, clk);
  dff _88978_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _01286_, clk);
  dff _88979_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _01288_, clk);
  dff _88980_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _01290_, clk);
  dff _88981_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _00588_, clk);
  dff _88982_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01292_, clk);
  dff _88983_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01294_, clk);
  dff _88984_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _01296_, clk);
  dff _88985_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01298_, clk);
  dff _88986_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _01299_, clk);
  dff _88987_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _01301_, clk);
  dff _88988_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _01303_, clk);
  dff _88989_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _00591_, clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell0.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell0.word [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.cell0.word [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.cell0.word [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.cell0.word [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.cell0.word [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.cell0.word [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.cell0.word [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.cell0.word [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.cell1.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell1.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell1.word [0], word_in[8]);
  buf(\oc8051_gm_cxrom_1.cell1.word [1], word_in[9]);
  buf(\oc8051_gm_cxrom_1.cell1.word [2], word_in[10]);
  buf(\oc8051_gm_cxrom_1.cell1.word [3], word_in[11]);
  buf(\oc8051_gm_cxrom_1.cell1.word [4], word_in[12]);
  buf(\oc8051_gm_cxrom_1.cell1.word [5], word_in[13]);
  buf(\oc8051_gm_cxrom_1.cell1.word [6], word_in[14]);
  buf(\oc8051_gm_cxrom_1.cell1.word [7], word_in[15]);
  buf(\oc8051_gm_cxrom_1.cell2.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell2.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell2.word [0], word_in[16]);
  buf(\oc8051_gm_cxrom_1.cell2.word [1], word_in[17]);
  buf(\oc8051_gm_cxrom_1.cell2.word [2], word_in[18]);
  buf(\oc8051_gm_cxrom_1.cell2.word [3], word_in[19]);
  buf(\oc8051_gm_cxrom_1.cell2.word [4], word_in[20]);
  buf(\oc8051_gm_cxrom_1.cell2.word [5], word_in[21]);
  buf(\oc8051_gm_cxrom_1.cell2.word [6], word_in[22]);
  buf(\oc8051_gm_cxrom_1.cell2.word [7], word_in[23]);
  buf(\oc8051_gm_cxrom_1.cell3.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell3.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell3.word [0], word_in[24]);
  buf(\oc8051_gm_cxrom_1.cell3.word [1], word_in[25]);
  buf(\oc8051_gm_cxrom_1.cell3.word [2], word_in[26]);
  buf(\oc8051_gm_cxrom_1.cell3.word [3], word_in[27]);
  buf(\oc8051_gm_cxrom_1.cell3.word [4], word_in[28]);
  buf(\oc8051_gm_cxrom_1.cell3.word [5], word_in[29]);
  buf(\oc8051_gm_cxrom_1.cell3.word [6], word_in[30]);
  buf(\oc8051_gm_cxrom_1.cell3.word [7], word_in[31]);
  buf(\oc8051_gm_cxrom_1.cell4.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell4.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell4.word [0], word_in[32]);
  buf(\oc8051_gm_cxrom_1.cell4.word [1], word_in[33]);
  buf(\oc8051_gm_cxrom_1.cell4.word [2], word_in[34]);
  buf(\oc8051_gm_cxrom_1.cell4.word [3], word_in[35]);
  buf(\oc8051_gm_cxrom_1.cell4.word [4], word_in[36]);
  buf(\oc8051_gm_cxrom_1.cell4.word [5], word_in[37]);
  buf(\oc8051_gm_cxrom_1.cell4.word [6], word_in[38]);
  buf(\oc8051_gm_cxrom_1.cell4.word [7], word_in[39]);
  buf(\oc8051_gm_cxrom_1.cell5.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell5.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell5.word [0], word_in[40]);
  buf(\oc8051_gm_cxrom_1.cell5.word [1], word_in[41]);
  buf(\oc8051_gm_cxrom_1.cell5.word [2], word_in[42]);
  buf(\oc8051_gm_cxrom_1.cell5.word [3], word_in[43]);
  buf(\oc8051_gm_cxrom_1.cell5.word [4], word_in[44]);
  buf(\oc8051_gm_cxrom_1.cell5.word [5], word_in[45]);
  buf(\oc8051_gm_cxrom_1.cell5.word [6], word_in[46]);
  buf(\oc8051_gm_cxrom_1.cell5.word [7], word_in[47]);
  buf(\oc8051_gm_cxrom_1.cell6.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell6.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell6.word [0], word_in[48]);
  buf(\oc8051_gm_cxrom_1.cell6.word [1], word_in[49]);
  buf(\oc8051_gm_cxrom_1.cell6.word [2], word_in[50]);
  buf(\oc8051_gm_cxrom_1.cell6.word [3], word_in[51]);
  buf(\oc8051_gm_cxrom_1.cell6.word [4], word_in[52]);
  buf(\oc8051_gm_cxrom_1.cell6.word [5], word_in[53]);
  buf(\oc8051_gm_cxrom_1.cell6.word [6], word_in[54]);
  buf(\oc8051_gm_cxrom_1.cell6.word [7], word_in[55]);
  buf(\oc8051_gm_cxrom_1.cell7.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell7.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell7.word [0], word_in[56]);
  buf(\oc8051_gm_cxrom_1.cell7.word [1], word_in[57]);
  buf(\oc8051_gm_cxrom_1.cell7.word [2], word_in[58]);
  buf(\oc8051_gm_cxrom_1.cell7.word [3], word_in[59]);
  buf(\oc8051_gm_cxrom_1.cell7.word [4], word_in[60]);
  buf(\oc8051_gm_cxrom_1.cell7.word [5], word_in[61]);
  buf(\oc8051_gm_cxrom_1.cell7.word [6], word_in[62]);
  buf(\oc8051_gm_cxrom_1.cell7.word [7], word_in[63]);
  buf(\oc8051_gm_cxrom_1.cell8.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell8.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell8.word [0], word_in[64]);
  buf(\oc8051_gm_cxrom_1.cell8.word [1], word_in[65]);
  buf(\oc8051_gm_cxrom_1.cell8.word [2], word_in[66]);
  buf(\oc8051_gm_cxrom_1.cell8.word [3], word_in[67]);
  buf(\oc8051_gm_cxrom_1.cell8.word [4], word_in[68]);
  buf(\oc8051_gm_cxrom_1.cell8.word [5], word_in[69]);
  buf(\oc8051_gm_cxrom_1.cell8.word [6], word_in[70]);
  buf(\oc8051_gm_cxrom_1.cell8.word [7], word_in[71]);
  buf(\oc8051_gm_cxrom_1.cell9.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell9.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell9.word [0], word_in[72]);
  buf(\oc8051_gm_cxrom_1.cell9.word [1], word_in[73]);
  buf(\oc8051_gm_cxrom_1.cell9.word [2], word_in[74]);
  buf(\oc8051_gm_cxrom_1.cell9.word [3], word_in[75]);
  buf(\oc8051_gm_cxrom_1.cell9.word [4], word_in[76]);
  buf(\oc8051_gm_cxrom_1.cell9.word [5], word_in[77]);
  buf(\oc8051_gm_cxrom_1.cell9.word [6], word_in[78]);
  buf(\oc8051_gm_cxrom_1.cell9.word [7], word_in[79]);
  buf(\oc8051_gm_cxrom_1.cell10.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell10.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell10.word [0], word_in[80]);
  buf(\oc8051_gm_cxrom_1.cell10.word [1], word_in[81]);
  buf(\oc8051_gm_cxrom_1.cell10.word [2], word_in[82]);
  buf(\oc8051_gm_cxrom_1.cell10.word [3], word_in[83]);
  buf(\oc8051_gm_cxrom_1.cell10.word [4], word_in[84]);
  buf(\oc8051_gm_cxrom_1.cell10.word [5], word_in[85]);
  buf(\oc8051_gm_cxrom_1.cell10.word [6], word_in[86]);
  buf(\oc8051_gm_cxrom_1.cell10.word [7], word_in[87]);
  buf(\oc8051_gm_cxrom_1.cell11.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell11.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell11.word [0], word_in[88]);
  buf(\oc8051_gm_cxrom_1.cell11.word [1], word_in[89]);
  buf(\oc8051_gm_cxrom_1.cell11.word [2], word_in[90]);
  buf(\oc8051_gm_cxrom_1.cell11.word [3], word_in[91]);
  buf(\oc8051_gm_cxrom_1.cell11.word [4], word_in[92]);
  buf(\oc8051_gm_cxrom_1.cell11.word [5], word_in[93]);
  buf(\oc8051_gm_cxrom_1.cell11.word [6], word_in[94]);
  buf(\oc8051_gm_cxrom_1.cell11.word [7], word_in[95]);
  buf(\oc8051_gm_cxrom_1.cell12.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell12.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell12.word [0], word_in[96]);
  buf(\oc8051_gm_cxrom_1.cell12.word [1], word_in[97]);
  buf(\oc8051_gm_cxrom_1.cell12.word [2], word_in[98]);
  buf(\oc8051_gm_cxrom_1.cell12.word [3], word_in[99]);
  buf(\oc8051_gm_cxrom_1.cell12.word [4], word_in[100]);
  buf(\oc8051_gm_cxrom_1.cell12.word [5], word_in[101]);
  buf(\oc8051_gm_cxrom_1.cell12.word [6], word_in[102]);
  buf(\oc8051_gm_cxrom_1.cell12.word [7], word_in[103]);
  buf(\oc8051_gm_cxrom_1.cell13.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell13.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell13.word [0], word_in[104]);
  buf(\oc8051_gm_cxrom_1.cell13.word [1], word_in[105]);
  buf(\oc8051_gm_cxrom_1.cell13.word [2], word_in[106]);
  buf(\oc8051_gm_cxrom_1.cell13.word [3], word_in[107]);
  buf(\oc8051_gm_cxrom_1.cell13.word [4], word_in[108]);
  buf(\oc8051_gm_cxrom_1.cell13.word [5], word_in[109]);
  buf(\oc8051_gm_cxrom_1.cell13.word [6], word_in[110]);
  buf(\oc8051_gm_cxrom_1.cell13.word [7], word_in[111]);
  buf(\oc8051_gm_cxrom_1.cell14.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell14.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell14.word [0], word_in[112]);
  buf(\oc8051_gm_cxrom_1.cell14.word [1], word_in[113]);
  buf(\oc8051_gm_cxrom_1.cell14.word [2], word_in[114]);
  buf(\oc8051_gm_cxrom_1.cell14.word [3], word_in[115]);
  buf(\oc8051_gm_cxrom_1.cell14.word [4], word_in[116]);
  buf(\oc8051_gm_cxrom_1.cell14.word [5], word_in[117]);
  buf(\oc8051_gm_cxrom_1.cell14.word [6], word_in[118]);
  buf(\oc8051_gm_cxrom_1.cell14.word [7], word_in[119]);
  buf(\oc8051_gm_cxrom_1.cell15.clk , clk);
  buf(\oc8051_gm_cxrom_1.cell15.rst , rst);
  buf(\oc8051_gm_cxrom_1.cell15.word [0], word_in[120]);
  buf(\oc8051_gm_cxrom_1.cell15.word [1], word_in[121]);
  buf(\oc8051_gm_cxrom_1.cell15.word [2], word_in[122]);
  buf(\oc8051_gm_cxrom_1.cell15.word [3], word_in[123]);
  buf(\oc8051_gm_cxrom_1.cell15.word [4], word_in[124]);
  buf(\oc8051_gm_cxrom_1.cell15.word [5], word_in[125]);
  buf(\oc8051_gm_cxrom_1.cell15.word [6], word_in[126]);
  buf(\oc8051_gm_cxrom_1.cell15.word [7], word_in[127]);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dadr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [0], \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [1], \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [2], \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [3], \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [4], \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [5], \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [6], \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff0 [7], \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [0], \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [1], \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [2], \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [3], \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [4], \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [5], \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [6], \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff1 [7], \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [0], \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [1], \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [2], \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [3], \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [4], \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [5], \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [6], \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff2 [7], \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [0], \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [1], \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [2], \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [3], \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [4], \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [5], \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [6], \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.buff3 [7], \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [0], psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.txd , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.p , psw[0]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_gm_cxrom_1.clk , clk);
  buf(\oc8051_gm_cxrom_1.rst , rst);
  buf(\oc8051_gm_cxrom_1.word_in [0], word_in[0]);
  buf(\oc8051_gm_cxrom_1.word_in [1], word_in[1]);
  buf(\oc8051_gm_cxrom_1.word_in [2], word_in[2]);
  buf(\oc8051_gm_cxrom_1.word_in [3], word_in[3]);
  buf(\oc8051_gm_cxrom_1.word_in [4], word_in[4]);
  buf(\oc8051_gm_cxrom_1.word_in [5], word_in[5]);
  buf(\oc8051_gm_cxrom_1.word_in [6], word_in[6]);
  buf(\oc8051_gm_cxrom_1.word_in [7], word_in[7]);
  buf(\oc8051_gm_cxrom_1.word_in [8], word_in[8]);
  buf(\oc8051_gm_cxrom_1.word_in [9], word_in[9]);
  buf(\oc8051_gm_cxrom_1.word_in [10], word_in[10]);
  buf(\oc8051_gm_cxrom_1.word_in [11], word_in[11]);
  buf(\oc8051_gm_cxrom_1.word_in [12], word_in[12]);
  buf(\oc8051_gm_cxrom_1.word_in [13], word_in[13]);
  buf(\oc8051_gm_cxrom_1.word_in [14], word_in[14]);
  buf(\oc8051_gm_cxrom_1.word_in [15], word_in[15]);
  buf(\oc8051_gm_cxrom_1.word_in [16], word_in[16]);
  buf(\oc8051_gm_cxrom_1.word_in [17], word_in[17]);
  buf(\oc8051_gm_cxrom_1.word_in [18], word_in[18]);
  buf(\oc8051_gm_cxrom_1.word_in [19], word_in[19]);
  buf(\oc8051_gm_cxrom_1.word_in [20], word_in[20]);
  buf(\oc8051_gm_cxrom_1.word_in [21], word_in[21]);
  buf(\oc8051_gm_cxrom_1.word_in [22], word_in[22]);
  buf(\oc8051_gm_cxrom_1.word_in [23], word_in[23]);
  buf(\oc8051_gm_cxrom_1.word_in [24], word_in[24]);
  buf(\oc8051_gm_cxrom_1.word_in [25], word_in[25]);
  buf(\oc8051_gm_cxrom_1.word_in [26], word_in[26]);
  buf(\oc8051_gm_cxrom_1.word_in [27], word_in[27]);
  buf(\oc8051_gm_cxrom_1.word_in [28], word_in[28]);
  buf(\oc8051_gm_cxrom_1.word_in [29], word_in[29]);
  buf(\oc8051_gm_cxrom_1.word_in [30], word_in[30]);
  buf(\oc8051_gm_cxrom_1.word_in [31], word_in[31]);
  buf(\oc8051_gm_cxrom_1.word_in [32], word_in[32]);
  buf(\oc8051_gm_cxrom_1.word_in [33], word_in[33]);
  buf(\oc8051_gm_cxrom_1.word_in [34], word_in[34]);
  buf(\oc8051_gm_cxrom_1.word_in [35], word_in[35]);
  buf(\oc8051_gm_cxrom_1.word_in [36], word_in[36]);
  buf(\oc8051_gm_cxrom_1.word_in [37], word_in[37]);
  buf(\oc8051_gm_cxrom_1.word_in [38], word_in[38]);
  buf(\oc8051_gm_cxrom_1.word_in [39], word_in[39]);
  buf(\oc8051_gm_cxrom_1.word_in [40], word_in[40]);
  buf(\oc8051_gm_cxrom_1.word_in [41], word_in[41]);
  buf(\oc8051_gm_cxrom_1.word_in [42], word_in[42]);
  buf(\oc8051_gm_cxrom_1.word_in [43], word_in[43]);
  buf(\oc8051_gm_cxrom_1.word_in [44], word_in[44]);
  buf(\oc8051_gm_cxrom_1.word_in [45], word_in[45]);
  buf(\oc8051_gm_cxrom_1.word_in [46], word_in[46]);
  buf(\oc8051_gm_cxrom_1.word_in [47], word_in[47]);
  buf(\oc8051_gm_cxrom_1.word_in [48], word_in[48]);
  buf(\oc8051_gm_cxrom_1.word_in [49], word_in[49]);
  buf(\oc8051_gm_cxrom_1.word_in [50], word_in[50]);
  buf(\oc8051_gm_cxrom_1.word_in [51], word_in[51]);
  buf(\oc8051_gm_cxrom_1.word_in [52], word_in[52]);
  buf(\oc8051_gm_cxrom_1.word_in [53], word_in[53]);
  buf(\oc8051_gm_cxrom_1.word_in [54], word_in[54]);
  buf(\oc8051_gm_cxrom_1.word_in [55], word_in[55]);
  buf(\oc8051_gm_cxrom_1.word_in [56], word_in[56]);
  buf(\oc8051_gm_cxrom_1.word_in [57], word_in[57]);
  buf(\oc8051_gm_cxrom_1.word_in [58], word_in[58]);
  buf(\oc8051_gm_cxrom_1.word_in [59], word_in[59]);
  buf(\oc8051_gm_cxrom_1.word_in [60], word_in[60]);
  buf(\oc8051_gm_cxrom_1.word_in [61], word_in[61]);
  buf(\oc8051_gm_cxrom_1.word_in [62], word_in[62]);
  buf(\oc8051_gm_cxrom_1.word_in [63], word_in[63]);
  buf(\oc8051_gm_cxrom_1.word_in [64], word_in[64]);
  buf(\oc8051_gm_cxrom_1.word_in [65], word_in[65]);
  buf(\oc8051_gm_cxrom_1.word_in [66], word_in[66]);
  buf(\oc8051_gm_cxrom_1.word_in [67], word_in[67]);
  buf(\oc8051_gm_cxrom_1.word_in [68], word_in[68]);
  buf(\oc8051_gm_cxrom_1.word_in [69], word_in[69]);
  buf(\oc8051_gm_cxrom_1.word_in [70], word_in[70]);
  buf(\oc8051_gm_cxrom_1.word_in [71], word_in[71]);
  buf(\oc8051_gm_cxrom_1.word_in [72], word_in[72]);
  buf(\oc8051_gm_cxrom_1.word_in [73], word_in[73]);
  buf(\oc8051_gm_cxrom_1.word_in [74], word_in[74]);
  buf(\oc8051_gm_cxrom_1.word_in [75], word_in[75]);
  buf(\oc8051_gm_cxrom_1.word_in [76], word_in[76]);
  buf(\oc8051_gm_cxrom_1.word_in [77], word_in[77]);
  buf(\oc8051_gm_cxrom_1.word_in [78], word_in[78]);
  buf(\oc8051_gm_cxrom_1.word_in [79], word_in[79]);
  buf(\oc8051_gm_cxrom_1.word_in [80], word_in[80]);
  buf(\oc8051_gm_cxrom_1.word_in [81], word_in[81]);
  buf(\oc8051_gm_cxrom_1.word_in [82], word_in[82]);
  buf(\oc8051_gm_cxrom_1.word_in [83], word_in[83]);
  buf(\oc8051_gm_cxrom_1.word_in [84], word_in[84]);
  buf(\oc8051_gm_cxrom_1.word_in [85], word_in[85]);
  buf(\oc8051_gm_cxrom_1.word_in [86], word_in[86]);
  buf(\oc8051_gm_cxrom_1.word_in [87], word_in[87]);
  buf(\oc8051_gm_cxrom_1.word_in [88], word_in[88]);
  buf(\oc8051_gm_cxrom_1.word_in [89], word_in[89]);
  buf(\oc8051_gm_cxrom_1.word_in [90], word_in[90]);
  buf(\oc8051_gm_cxrom_1.word_in [91], word_in[91]);
  buf(\oc8051_gm_cxrom_1.word_in [92], word_in[92]);
  buf(\oc8051_gm_cxrom_1.word_in [93], word_in[93]);
  buf(\oc8051_gm_cxrom_1.word_in [94], word_in[94]);
  buf(\oc8051_gm_cxrom_1.word_in [95], word_in[95]);
  buf(\oc8051_gm_cxrom_1.word_in [96], word_in[96]);
  buf(\oc8051_gm_cxrom_1.word_in [97], word_in[97]);
  buf(\oc8051_gm_cxrom_1.word_in [98], word_in[98]);
  buf(\oc8051_gm_cxrom_1.word_in [99], word_in[99]);
  buf(\oc8051_gm_cxrom_1.word_in [100], word_in[100]);
  buf(\oc8051_gm_cxrom_1.word_in [101], word_in[101]);
  buf(\oc8051_gm_cxrom_1.word_in [102], word_in[102]);
  buf(\oc8051_gm_cxrom_1.word_in [103], word_in[103]);
  buf(\oc8051_gm_cxrom_1.word_in [104], word_in[104]);
  buf(\oc8051_gm_cxrom_1.word_in [105], word_in[105]);
  buf(\oc8051_gm_cxrom_1.word_in [106], word_in[106]);
  buf(\oc8051_gm_cxrom_1.word_in [107], word_in[107]);
  buf(\oc8051_gm_cxrom_1.word_in [108], word_in[108]);
  buf(\oc8051_gm_cxrom_1.word_in [109], word_in[109]);
  buf(\oc8051_gm_cxrom_1.word_in [110], word_in[110]);
  buf(\oc8051_gm_cxrom_1.word_in [111], word_in[111]);
  buf(\oc8051_gm_cxrom_1.word_in [112], word_in[112]);
  buf(\oc8051_gm_cxrom_1.word_in [113], word_in[113]);
  buf(\oc8051_gm_cxrom_1.word_in [114], word_in[114]);
  buf(\oc8051_gm_cxrom_1.word_in [115], word_in[115]);
  buf(\oc8051_gm_cxrom_1.word_in [116], word_in[116]);
  buf(\oc8051_gm_cxrom_1.word_in [117], word_in[117]);
  buf(\oc8051_gm_cxrom_1.word_in [118], word_in[118]);
  buf(\oc8051_gm_cxrom_1.word_in [119], word_in[119]);
  buf(\oc8051_gm_cxrom_1.word_in [120], word_in[120]);
  buf(\oc8051_gm_cxrom_1.word_in [121], word_in[121]);
  buf(\oc8051_gm_cxrom_1.word_in [122], word_in[122]);
  buf(\oc8051_gm_cxrom_1.word_in [123], word_in[123]);
  buf(\oc8051_gm_cxrom_1.word_in [124], word_in[124]);
  buf(\oc8051_gm_cxrom_1.word_in [125], word_in[125]);
  buf(\oc8051_gm_cxrom_1.word_in [126], word_in[126]);
  buf(\oc8051_gm_cxrom_1.word_in [127], word_in[127]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_gm_cxrom_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_gm_cxrom_1.rd_addr_0 [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [0], \oc8051_golden_model_1.PC [0]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [1], \oc8051_golden_model_1.PC [1]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [2], \oc8051_golden_model_1.PC [2]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [3], \oc8051_golden_model_1.PC [3]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [4], \oc8051_golden_model_1.PC [4]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [5], \oc8051_golden_model_1.PC [5]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [6], \oc8051_golden_model_1.PC [6]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [7], \oc8051_golden_model_1.PC [7]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [8], \oc8051_golden_model_1.PC [8]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [9], \oc8051_golden_model_1.PC [9]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [10], \oc8051_golden_model_1.PC [10]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [11], \oc8051_golden_model_1.PC [11]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [12], \oc8051_golden_model_1.PC [12]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [13], \oc8051_golden_model_1.PC [13]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [14], \oc8051_golden_model_1.PC [14]);
  buf(\oc8051_golden_model_1.RD_ROM_0_ADDR [15], \oc8051_golden_model_1.PC [15]);
  buf(\oc8051_golden_model_1.clk , clk);
  buf(\oc8051_golden_model_1.rst , rst);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [0], word_in[0]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [1], word_in[1]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [2], word_in[2]);
  buf(\oc8051_golden_model_1.RD_IRAM_ADDR [3], word_in[3]);
  buf(\oc8051_golden_model_1.ACC_03 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_03 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_03 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_03 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_03 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_03 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_03 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_03 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_13 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_13 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_13 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_13 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_13 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_13 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_13 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_13 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_23 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_23 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_23 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_23 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_23 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_23 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_23 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_23 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_33 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.ACC_33 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_33 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_33 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_33 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_33 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_33 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_33 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_c4 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_c4 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_c4 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_c4 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.ACC_c4 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.ACC_c4 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.ACC_c4 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d6 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d6 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d6 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d6 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d6 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d6 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d6 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_d7 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_d7 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_d7 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_d7 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_d7 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.ACC_d7 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.ACC_d7 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.ACC_d7 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.ACC_e4 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.ACC_e4 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.ACC_e4 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.ACC_e4 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.ACC_e4 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.ACC_e4 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.ACC_e4 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.ACC_e4 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_22 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_22 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_22 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_22 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_22 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_22 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_22 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_22 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_22 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_22 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_22 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_22 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_22 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_22 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_22 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PC_32 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.PC_32 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.PC_32 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.PC_32 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.PC_32 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.PC_32 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.PC_32 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.PC_32 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.PC_32 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.PC_32 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.PC_32 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.PC_32 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.PC_32 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.PC_32 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.PC_32 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.PC_32 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.PSW_13 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_13 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_13 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_13 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_13 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_13 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_13 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_13 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.PSW_24 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_24 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_24 [2], \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.PSW_24 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_24 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_24 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_24 [6], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.PSW_24 [7], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.PSW_25 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_25 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_25 [2], \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.PSW_25 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_25 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_25 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_25 [6], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.PSW_25 [7], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.PSW_26 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_26 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_26 [2], \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.PSW_26 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_26 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_26 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_26 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_26 [7], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.PSW_27 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_27 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_27 [2], \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.PSW_27 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_27 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_27 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_27 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.PSW_27 [7], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.PSW_28 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_28 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_28 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_28 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_28 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_28 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_28 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_28 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_29 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_29 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_29 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_29 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_29 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_29 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_29 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_29 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2a [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2a [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2a [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2b [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2b [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2b [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2c [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2c [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.PSW_2c [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2d [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.PSW_2d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2d [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2d [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.PSW_2e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2e [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2e [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2e [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_2f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_2f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_2f [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.PSW_2f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_2f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_2f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_2f [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.PSW_2f [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.PSW_33 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_33 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_33 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_33 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_33 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_33 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_33 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_33 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.PSW_34 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_34 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_34 [2], \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.PSW_34 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_34 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_34 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_34 [6], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.PSW_34 [7], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.PSW_35 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_35 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_35 [2], \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.PSW_35 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_35 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_35 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_35 [6], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.PSW_35 [7], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.PSW_36 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_36 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_36 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_36 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_36 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_36 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_36 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_36 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_37 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_37 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_37 [2], \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.PSW_37 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_37 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_37 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_37 [6], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.PSW_37 [7], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.PSW_38 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_38 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_38 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_38 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_38 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_38 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_38 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_38 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_39 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_39 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_39 [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_39 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_39 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_39 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_39 [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_39 [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3a [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3a [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3a [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3b [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3b [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3b [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3c [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3c [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3c [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3d [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3d [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3d [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3e [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3e [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3e [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_3f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_3f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_3f [2], \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.PSW_3f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_3f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_3f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_3f [6], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.PSW_3f [7], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.PSW_72 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_72 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_72 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_72 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_72 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_72 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_72 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_72 [7], \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.PSW_82 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_82 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_82 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_82 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_82 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_82 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_82 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_82 [7], \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.PSW_84 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_84 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_84 [2], \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.PSW_84 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_84 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_84 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_84 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_84 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_94 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_94 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_94 [2], \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.PSW_94 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_94 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_94 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_94 [6], \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.PSW_94 [7], \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.PSW_95 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_95 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_95 [2], \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.PSW_95 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_95 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_95 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_95 [6], \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.PSW_95 [7], \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.PSW_96 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_96 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_96 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_96 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_96 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_96 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_96 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_96 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_97 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_97 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_97 [2], \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.PSW_97 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_97 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_97 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_97 [6], \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.PSW_97 [7], \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.PSW_98 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_98 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_98 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_98 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_98 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_98 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_98 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_98 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_99 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_99 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_99 [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_99 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_99 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_99 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_99 [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_99 [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9a [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9a [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9a [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9a [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9a [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9a [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9a [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9a [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9b [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9b [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9b [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9b [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9b [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9b [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9b [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9b [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9c [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9c [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9c [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9c [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9c [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9c [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9c [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9c [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9d [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9d [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9d [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9d [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9d [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9d [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9d [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9d [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9e [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9e [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9e [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9e [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9e [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9e [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9e [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9e [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_9f [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_9f [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_9f [2], \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.PSW_9f [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_9f [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_9f [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_9f [6], \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.PSW_9f [7], \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.PSW_a0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a0 [7], \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.PSW_a2 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a2 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a2 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_a2 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a2 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a2 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a2 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a2 [7], \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.PSW_a4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_a4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_a4 [2], \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.PSW_a4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_a4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_a4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_a4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_a4 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_b0 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b0 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b0 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b0 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b0 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b0 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b0 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b0 [7], \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.PSW_b3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b3 [7], \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.PSW_b4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b4 [7], \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.PSW_b5 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b5 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b5 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b5 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b5 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b5 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b5 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b5 [7], \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.PSW_b6 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b6 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b6 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b6 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b6 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b6 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b6 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b6 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b7 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b7 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b7 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b7 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b7 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b7 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b7 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b7 [7], \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.PSW_b8 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b8 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b8 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b8 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b8 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b8 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b8 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b8 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_b9 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_b9 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_b9 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_b9 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_b9 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_b9 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_b9 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_b9 [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_ba [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_ba [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_ba [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_ba [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_ba [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_ba [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_ba [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_ba [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bb [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bb [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bb [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bb [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bb [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bb [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bb [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bb [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bc [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bc [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bc [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bc [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bc [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bc [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bc [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bc [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bd [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bd [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bd [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bd [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bd [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bd [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bd [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bd [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_be [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_be [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_be [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_be [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_be [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_be [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_be [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_be [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_bf [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_bf [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_bf [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_bf [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_bf [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_bf [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_bf [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_bf [7], \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.PSW_c3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_c3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_c3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_c3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_c3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_c3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_c3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_c3 [7], 1'b0);
  buf(\oc8051_golden_model_1.PSW_d3 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d3 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d3 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d3 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d3 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d3 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d3 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d3 [7], 1'b1);
  buf(\oc8051_golden_model_1.PSW_d4 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.PSW_d4 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.PSW_d4 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.PSW_d4 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.PSW_d4 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.PSW_d4 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.PSW_d4 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.PSW_d4 [7], \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_0 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.RD_IRAM_1 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0006 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0006 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0007 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0007 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0007 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0011 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0011 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0011 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0011 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0019 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0019 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0019 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0019 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0023 [2], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0023 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0023 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0023 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0027 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0027 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0027 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0027 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [1], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0031 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0031 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0031 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0031 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [0], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0035 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0035 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0035 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0035 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [0], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [1], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [2], 1'b1);
  buf(\oc8051_golden_model_1.n0039 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n0039 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n0039 [5], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [6], 1'b0);
  buf(\oc8051_golden_model_1.n0039 [7], 1'b0);
  buf(\oc8051_golden_model_1.n0561 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n0561 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n0561 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n0561 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n0561 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n0561 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n0561 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n0561 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n0594 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n0594 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n0594 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n0594 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n0594 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n0594 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n0594 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n0594 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n0701 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n0701 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0701 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0701 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0701 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0701 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0701 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0701 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0701 [8], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [9], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [10], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [11], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [12], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [13], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [14], 1'b0);
  buf(\oc8051_golden_model_1.n0701 [15], 1'b0);
  buf(\oc8051_golden_model_1.n0733 [0], \oc8051_golden_model_1.DPL [0]);
  buf(\oc8051_golden_model_1.n0733 [1], \oc8051_golden_model_1.DPL [1]);
  buf(\oc8051_golden_model_1.n0733 [2], \oc8051_golden_model_1.DPL [2]);
  buf(\oc8051_golden_model_1.n0733 [3], \oc8051_golden_model_1.DPL [3]);
  buf(\oc8051_golden_model_1.n0733 [4], \oc8051_golden_model_1.DPL [4]);
  buf(\oc8051_golden_model_1.n0733 [5], \oc8051_golden_model_1.DPL [5]);
  buf(\oc8051_golden_model_1.n0733 [6], \oc8051_golden_model_1.DPL [6]);
  buf(\oc8051_golden_model_1.n0733 [7], \oc8051_golden_model_1.DPL [7]);
  buf(\oc8051_golden_model_1.n0733 [8], \oc8051_golden_model_1.DPH [0]);
  buf(\oc8051_golden_model_1.n0733 [9], \oc8051_golden_model_1.DPH [1]);
  buf(\oc8051_golden_model_1.n0733 [10], \oc8051_golden_model_1.DPH [2]);
  buf(\oc8051_golden_model_1.n0733 [11], \oc8051_golden_model_1.DPH [3]);
  buf(\oc8051_golden_model_1.n0733 [12], \oc8051_golden_model_1.DPH [4]);
  buf(\oc8051_golden_model_1.n0733 [13], \oc8051_golden_model_1.DPH [5]);
  buf(\oc8051_golden_model_1.n0733 [14], \oc8051_golden_model_1.DPH [6]);
  buf(\oc8051_golden_model_1.n0733 [15], \oc8051_golden_model_1.DPH [7]);
  buf(\oc8051_golden_model_1.n0994 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n0994 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n0994 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n0994 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n0994 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n0994 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n0994 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n0994 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1071 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1071 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1071 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1071 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1073 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1073 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1075 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1075 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1075 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1076 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1076 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1076 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1077 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1077 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1077 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1078 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1078 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1078 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1079 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1079 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1079 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1080 [0], 1'b0);
  buf(\oc8051_golden_model_1.n1080 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1080 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1081 [0], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [1], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [2], 1'b1);
  buf(\oc8051_golden_model_1.n1081 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1118 , \oc8051_golden_model_1.n1735 [7]);
  buf(\oc8051_golden_model_1.n1146 , \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1147 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1147 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1147 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1147 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1147 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1147 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1147 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1147 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1148 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1148 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1148 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1148 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1148 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1148 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1148 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1148 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1149 [0], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1149 [1], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1149 [2], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1149 [3], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1149 [4], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1149 [5], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1149 [6], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1149 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1150 , \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1151 , \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1152 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1152 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1152 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1153 , \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1154 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1154 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1155 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1155 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1155 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1155 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1155 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1155 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1155 [7], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1181 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1181 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1181 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1181 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1181 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1181 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1181 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1181 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1181 [8], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1181 [9], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1181 [10], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1181 [11], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1181 [12], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1181 [13], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1181 [14], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1181 [15], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1183 [0], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1183 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1183 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1183 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1183 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1183 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1183 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1183 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1185 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1185 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1185 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1185 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1185 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1185 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1185 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1185 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1189 [8], \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1190 , \oc8051_golden_model_1.n1207 [7]);
  buf(\oc8051_golden_model_1.n1191 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1191 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1191 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1191 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1192 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1192 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1192 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1192 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1196 [4], \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1197 , \oc8051_golden_model_1.n1207 [6]);
  buf(\oc8051_golden_model_1.n1198 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1198 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1198 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1198 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1198 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1198 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1198 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1198 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1198 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1206 , \oc8051_golden_model_1.n1207 [2]);
  buf(\oc8051_golden_model_1.n1207 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1207 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1207 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1207 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1207 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1211 [8], \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1212 , \oc8051_golden_model_1.n1227 [7]);
  buf(\oc8051_golden_model_1.n1217 [4], \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1218 , \oc8051_golden_model_1.n1227 [6]);
  buf(\oc8051_golden_model_1.n1226 , \oc8051_golden_model_1.n1227 [2]);
  buf(\oc8051_golden_model_1.n1227 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1227 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1227 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1227 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1227 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1229 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1229 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1229 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1229 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1229 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1229 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1229 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1229 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1229 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1231 [8], \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1232 , \oc8051_golden_model_1.n1246 [7]);
  buf(\oc8051_golden_model_1.n1233 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1233 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1233 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1233 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1234 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1234 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1234 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1234 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1236 [4], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1237 , \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1238 [0], \oc8051_golden_model_1.n1852 [0]);
  buf(\oc8051_golden_model_1.n1238 [1], \oc8051_golden_model_1.n1852 [1]);
  buf(\oc8051_golden_model_1.n1238 [2], \oc8051_golden_model_1.n1852 [2]);
  buf(\oc8051_golden_model_1.n1238 [3], \oc8051_golden_model_1.n1852 [3]);
  buf(\oc8051_golden_model_1.n1238 [4], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1238 [5], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1238 [6], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1238 [7], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1238 [8], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1245 , \oc8051_golden_model_1.n1246 [2]);
  buf(\oc8051_golden_model_1.n1246 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1246 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1246 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1246 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1246 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1246 [6], \oc8051_golden_model_1.n1258 [6]);
  buf(\oc8051_golden_model_1.n1249 [8], \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1250 , \oc8051_golden_model_1.n1258 [7]);
  buf(\oc8051_golden_model_1.n1257 , \oc8051_golden_model_1.n1258 [2]);
  buf(\oc8051_golden_model_1.n1258 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1258 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1258 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1258 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1258 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1260 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1260 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1260 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1260 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1260 [4], \oc8051_golden_model_1.n1268 [4]);
  buf(\oc8051_golden_model_1.n1260 [5], \oc8051_golden_model_1.n1268 [5]);
  buf(\oc8051_golden_model_1.n1260 [6], \oc8051_golden_model_1.n1268 [6]);
  buf(\oc8051_golden_model_1.n1260 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1260 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1262 [8], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1263 , \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1264 [0], \oc8051_golden_model_1.n1268 [0]);
  buf(\oc8051_golden_model_1.n1264 [1], \oc8051_golden_model_1.n1268 [1]);
  buf(\oc8051_golden_model_1.n1264 [2], \oc8051_golden_model_1.n1268 [2]);
  buf(\oc8051_golden_model_1.n1264 [3], \oc8051_golden_model_1.n1268 [3]);
  buf(\oc8051_golden_model_1.n1264 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1266 [4], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1267 , \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1268 [7], \oc8051_golden_model_1.n1268 [8]);
  buf(\oc8051_golden_model_1.n1275 , \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1276 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1276 [2], \oc8051_golden_model_1.n1280 [2]);
  buf(\oc8051_golden_model_1.n1276 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1276 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1276 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1276 [6], \oc8051_golden_model_1.n1292 [6]);
  buf(\oc8051_golden_model_1.n1276 [7], \oc8051_golden_model_1.n1280 [7]);
  buf(\oc8051_golden_model_1.n1278 [4], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1279 , \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1280 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1280 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1280 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1280 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1280 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1280 [6], \oc8051_golden_model_1.n1291 [6]);
  buf(\oc8051_golden_model_1.n1282 [8], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1283 , \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1290 , \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1291 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1291 [2], \oc8051_golden_model_1.n1292 [2]);
  buf(\oc8051_golden_model_1.n1291 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1291 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1291 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1291 [7], \oc8051_golden_model_1.n1292 [7]);
  buf(\oc8051_golden_model_1.n1292 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1292 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1292 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1292 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1292 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1295 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1295 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1295 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1295 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1295 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1295 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1295 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1295 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1295 [8], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1296 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1296 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1296 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1296 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1296 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1296 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1296 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1296 [8], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1297 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1297 [1], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1297 [2], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1297 [3], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1297 [4], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1297 [5], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1297 [6], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1297 [7], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1298 , \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1299 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1299 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1299 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1299 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1299 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1299 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1299 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1299 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1300 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1300 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1300 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1303 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [5], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [6], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1303 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1305 [8], \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1306 , \oc8051_golden_model_1.n1318 [7]);
  buf(\oc8051_golden_model_1.n1307 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1307 [1], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [2], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [3], 1'b0);
  buf(\oc8051_golden_model_1.n1307 [4], 1'b0);
  buf(\oc8051_golden_model_1.n1309 [4], \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1310 , \oc8051_golden_model_1.n1318 [6]);
  buf(\oc8051_golden_model_1.n1317 , \oc8051_golden_model_1.n1318 [2]);
  buf(\oc8051_golden_model_1.n1318 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1318 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1318 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1318 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1318 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1322 [8], \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1323 , \oc8051_golden_model_1.n1334 [7]);
  buf(\oc8051_golden_model_1.n1325 [4], \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1326 , \oc8051_golden_model_1.n1334 [6]);
  buf(\oc8051_golden_model_1.n1333 , \oc8051_golden_model_1.n1334 [2]);
  buf(\oc8051_golden_model_1.n1334 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1334 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1334 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1334 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1334 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1338 [8], \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1339 , \oc8051_golden_model_1.n1350 [7]);
  buf(\oc8051_golden_model_1.n1341 [4], \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1342 , \oc8051_golden_model_1.n1350 [6]);
  buf(\oc8051_golden_model_1.n1349 , \oc8051_golden_model_1.n1350 [2]);
  buf(\oc8051_golden_model_1.n1350 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1350 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1350 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1350 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1350 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1354 [8], \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1355 , \oc8051_golden_model_1.n1366 [7]);
  buf(\oc8051_golden_model_1.n1357 [4], \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1358 , \oc8051_golden_model_1.n1366 [6]);
  buf(\oc8051_golden_model_1.n1365 , \oc8051_golden_model_1.n1366 [2]);
  buf(\oc8051_golden_model_1.n1366 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1366 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1366 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1366 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1366 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1520 , \oc8051_golden_model_1.n1522 [7]);
  buf(\oc8051_golden_model_1.n1521 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1521 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1521 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1521 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1521 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1521 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1521 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1522 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1522 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1522 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1522 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1522 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1522 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1522 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1545 , \oc8051_golden_model_1.n1546 [7]);
  buf(\oc8051_golden_model_1.n1546 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1546 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1546 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1546 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1546 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1546 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1546 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1553 [0], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1553 [1], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1553 [2], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1553 [3], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1554 , \oc8051_golden_model_1.n1555 [2]);
  buf(\oc8051_golden_model_1.n1555 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1555 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1555 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1555 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1555 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1555 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1555 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1680 [0], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [1], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [2], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [3], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [4], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [5], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [6], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1680 [7], \oc8051_golden_model_1.PSW [7]);
  buf(\oc8051_golden_model_1.n1683 , \oc8051_golden_model_1.n1692 [7]);
  buf(\oc8051_golden_model_1.n1685 , \oc8051_golden_model_1.n1692 [6]);
  buf(\oc8051_golden_model_1.n1691 , \oc8051_golden_model_1.n1692 [2]);
  buf(\oc8051_golden_model_1.n1692 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1692 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1692 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1692 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1692 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1696 , \oc8051_golden_model_1.n1705 [7]);
  buf(\oc8051_golden_model_1.n1698 , \oc8051_golden_model_1.n1705 [6]);
  buf(\oc8051_golden_model_1.n1704 , \oc8051_golden_model_1.n1705 [2]);
  buf(\oc8051_golden_model_1.n1705 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1705 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1705 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1705 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1705 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1709 , \oc8051_golden_model_1.n1718 [7]);
  buf(\oc8051_golden_model_1.n1711 , \oc8051_golden_model_1.n1718 [6]);
  buf(\oc8051_golden_model_1.n1717 , \oc8051_golden_model_1.n1718 [2]);
  buf(\oc8051_golden_model_1.n1718 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1718 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1718 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1718 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1718 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1722 , \oc8051_golden_model_1.n1731 [7]);
  buf(\oc8051_golden_model_1.n1724 , \oc8051_golden_model_1.n1731 [6]);
  buf(\oc8051_golden_model_1.n1730 , \oc8051_golden_model_1.n1731 [2]);
  buf(\oc8051_golden_model_1.n1731 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1731 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1731 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1731 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1731 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1733 , \oc8051_golden_model_1.n1734 [7]);
  buf(\oc8051_golden_model_1.n1734 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1734 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1734 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1734 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1734 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1734 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1734 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1735 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1735 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1735 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1735 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1735 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1735 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1735 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1739 [0], \oc8051_golden_model_1.B [0]);
  buf(\oc8051_golden_model_1.n1739 [1], \oc8051_golden_model_1.B [1]);
  buf(\oc8051_golden_model_1.n1739 [2], \oc8051_golden_model_1.B [2]);
  buf(\oc8051_golden_model_1.n1739 [3], \oc8051_golden_model_1.B [3]);
  buf(\oc8051_golden_model_1.n1739 [4], \oc8051_golden_model_1.B [4]);
  buf(\oc8051_golden_model_1.n1739 [5], \oc8051_golden_model_1.B [5]);
  buf(\oc8051_golden_model_1.n1739 [6], \oc8051_golden_model_1.B [6]);
  buf(\oc8051_golden_model_1.n1739 [7], \oc8051_golden_model_1.B [7]);
  buf(\oc8051_golden_model_1.n1739 [8], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [9], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [10], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [11], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [12], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [13], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [14], 1'b0);
  buf(\oc8051_golden_model_1.n1739 [15], 1'b0);
  buf(\oc8051_golden_model_1.n1745 , \oc8051_golden_model_1.n1746 [2]);
  buf(\oc8051_golden_model_1.n1746 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1746 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1746 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1746 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1746 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1746 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1746 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1749 , \oc8051_golden_model_1.n1750 [7]);
  buf(\oc8051_golden_model_1.n1750 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1750 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1750 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1750 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1750 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1750 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1750 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1765 , \oc8051_golden_model_1.n1766 [7]);
  buf(\oc8051_golden_model_1.n1766 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1766 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1766 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1766 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1766 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1766 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1766 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1771 , \oc8051_golden_model_1.n1772 [7]);
  buf(\oc8051_golden_model_1.n1772 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1772 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1772 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1772 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1772 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1772 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1772 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1777 , \oc8051_golden_model_1.n1778 [7]);
  buf(\oc8051_golden_model_1.n1778 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1778 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1778 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1778 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1778 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1778 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1778 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1783 , \oc8051_golden_model_1.n1784 [7]);
  buf(\oc8051_golden_model_1.n1784 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1784 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1784 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1784 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1784 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1784 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1784 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1789 , \oc8051_golden_model_1.n1790 [7]);
  buf(\oc8051_golden_model_1.n1790 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1790 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1790 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1790 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1790 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1790 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1790 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1791 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1791 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1791 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1791 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1791 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1791 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1791 [7], 1'b0);
  buf(\oc8051_golden_model_1.n1792 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1792 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1792 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1792 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [0], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1793 [1], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1793 [2], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1793 [3], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1793 [4], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1793 [5], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1793 [6], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1793 [7], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_golden_model_1.n1828 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1828 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1828 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1828 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1828 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1828 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1828 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1828 [7], 1'b1);
  buf(\oc8051_golden_model_1.n1847 , \oc8051_golden_model_1.n1848 [7]);
  buf(\oc8051_golden_model_1.n1848 [0], \oc8051_golden_model_1.PSW [0]);
  buf(\oc8051_golden_model_1.n1848 [1], \oc8051_golden_model_1.PSW [1]);
  buf(\oc8051_golden_model_1.n1848 [2], \oc8051_golden_model_1.PSW [2]);
  buf(\oc8051_golden_model_1.n1848 [3], \oc8051_golden_model_1.PSW [3]);
  buf(\oc8051_golden_model_1.n1848 [4], \oc8051_golden_model_1.PSW [4]);
  buf(\oc8051_golden_model_1.n1848 [5], \oc8051_golden_model_1.PSW [5]);
  buf(\oc8051_golden_model_1.n1848 [6], \oc8051_golden_model_1.PSW [6]);
  buf(\oc8051_golden_model_1.n1852 [4], \oc8051_golden_model_1.ACC [4]);
  buf(\oc8051_golden_model_1.n1852 [5], \oc8051_golden_model_1.ACC [5]);
  buf(\oc8051_golden_model_1.n1852 [6], \oc8051_golden_model_1.ACC [6]);
  buf(\oc8051_golden_model_1.n1852 [7], \oc8051_golden_model_1.ACC [7]);
  buf(\oc8051_golden_model_1.n1853 [0], \oc8051_golden_model_1.n1854 [4]);
  buf(\oc8051_golden_model_1.n1853 [1], \oc8051_golden_model_1.n1854 [5]);
  buf(\oc8051_golden_model_1.n1853 [2], \oc8051_golden_model_1.n1854 [6]);
  buf(\oc8051_golden_model_1.n1853 [3], \oc8051_golden_model_1.n1854 [7]);
  buf(\oc8051_golden_model_1.n1854 [0], \oc8051_golden_model_1.ACC [0]);
  buf(\oc8051_golden_model_1.n1854 [1], \oc8051_golden_model_1.ACC [1]);
  buf(\oc8051_golden_model_1.n1854 [2], \oc8051_golden_model_1.ACC [2]);
  buf(\oc8051_golden_model_1.n1854 [3], \oc8051_golden_model_1.ACC [3]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.psw [0], psw[0]);
  buf(\oc8051_top_1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.wbd_we_o , \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(\oc8051_top_1.wbd_stb_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_cyc_o , \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(\oc8051_top_1.wbd_dat_o [0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(\oc8051_top_1.wbd_dat_o [1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(\oc8051_top_1.wbd_dat_o [2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(\oc8051_top_1.wbd_dat_o [3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(\oc8051_top_1.wbd_dat_o [4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(\oc8051_top_1.wbd_dat_o [5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(\oc8051_top_1.wbd_dat_o [6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(\oc8051_top_1.wbd_dat_o [7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(\oc8051_top_1.wbd_adr_o [0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(\oc8051_top_1.wbd_adr_o [1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(\oc8051_top_1.wbd_adr_o [2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(\oc8051_top_1.wbd_adr_o [3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(\oc8051_top_1.wbd_adr_o [4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(\oc8051_top_1.wbd_adr_o [5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(\oc8051_top_1.wbd_adr_o [6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(\oc8051_top_1.wbd_adr_o [7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(\oc8051_top_1.wbd_adr_o [8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(\oc8051_top_1.wbd_adr_o [9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(\oc8051_top_1.wbd_adr_o [10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(\oc8051_top_1.wbd_adr_o [11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(\oc8051_top_1.wbd_adr_o [12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(\oc8051_top_1.wbd_adr_o [13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(\oc8051_top_1.wbd_adr_o [14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(\oc8051_top_1.wbd_adr_o [15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.txd_o , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.ea_int , \oc8051_top_1.oc8051_rom1.ea_int );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(rd_iram_addr[0], word_in[0]);
  buf(rd_iram_addr[1], word_in[1]);
  buf(rd_iram_addr[2], word_in[2]);
  buf(rd_iram_addr[3], word_in[3]);
  buf(rd_rom_0_addr[0], \oc8051_golden_model_1.PC [0]);
  buf(rd_rom_0_addr[1], \oc8051_golden_model_1.PC [1]);
  buf(rd_rom_0_addr[2], \oc8051_golden_model_1.PC [2]);
  buf(rd_rom_0_addr[3], \oc8051_golden_model_1.PC [3]);
  buf(rd_rom_0_addr[4], \oc8051_golden_model_1.PC [4]);
  buf(rd_rom_0_addr[5], \oc8051_golden_model_1.PC [5]);
  buf(rd_rom_0_addr[6], \oc8051_golden_model_1.PC [6]);
  buf(rd_rom_0_addr[7], \oc8051_golden_model_1.PC [7]);
  buf(rd_rom_0_addr[8], \oc8051_golden_model_1.PC [8]);
  buf(rd_rom_0_addr[9], \oc8051_golden_model_1.PC [9]);
  buf(rd_rom_0_addr[10], \oc8051_golden_model_1.PC [10]);
  buf(rd_rom_0_addr[11], \oc8051_golden_model_1.PC [11]);
  buf(rd_rom_0_addr[12], \oc8051_golden_model_1.PC [12]);
  buf(rd_rom_0_addr[13], \oc8051_golden_model_1.PC [13]);
  buf(rd_rom_0_addr[14], \oc8051_golden_model_1.PC [14]);
  buf(rd_rom_0_addr[15], \oc8051_golden_model_1.PC [15]);
  buf(ACC_gm[0], \oc8051_golden_model_1.ACC [0]);
  buf(ACC_gm[1], \oc8051_golden_model_1.ACC [1]);
  buf(ACC_gm[2], \oc8051_golden_model_1.ACC [2]);
  buf(ACC_gm[3], \oc8051_golden_model_1.ACC [3]);
  buf(ACC_gm[4], \oc8051_golden_model_1.ACC [4]);
  buf(ACC_gm[5], \oc8051_golden_model_1.ACC [5]);
  buf(ACC_gm[6], \oc8051_golden_model_1.ACC [6]);
  buf(ACC_gm[7], \oc8051_golden_model_1.ACC [7]);
  buf(acc[0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(acc[1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(acc[2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(acc[3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(acc[4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(acc[5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(acc[6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(acc[7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(psw[1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(psw[2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(psw[3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(psw[4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(psw[5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(psw[6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(psw[7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(cxrom_data_out[0], \oc8051_top_1.oc8051_rom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_top_1.oc8051_rom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_top_1.oc8051_rom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_top_1.oc8051_rom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_top_1.oc8051_rom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_top_1.oc8051_rom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_top_1.oc8051_rom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_top_1.oc8051_rom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_top_1.oc8051_rom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_top_1.oc8051_rom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_top_1.oc8051_rom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_top_1.oc8051_rom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_top_1.oc8051_rom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_top_1.oc8051_rom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_top_1.oc8051_rom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_top_1.oc8051_rom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_top_1.oc8051_rom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_top_1.oc8051_rom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_top_1.oc8051_rom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_top_1.oc8051_rom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_top_1.oc8051_rom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_top_1.oc8051_rom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_top_1.oc8051_rom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_top_1.oc8051_rom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_top_1.oc8051_rom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_top_1.oc8051_rom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_top_1.oc8051_rom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_top_1.oc8051_rom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_top_1.oc8051_rom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_top_1.oc8051_rom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_top_1.oc8051_rom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_top_1.oc8051_rom1.cxrom_data_out [31]);
  buf(wbd_adr_o[0], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [0]);
  buf(wbd_adr_o[1], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [1]);
  buf(wbd_adr_o[2], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [2]);
  buf(wbd_adr_o[3], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [3]);
  buf(wbd_adr_o[4], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [4]);
  buf(wbd_adr_o[5], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [5]);
  buf(wbd_adr_o[6], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [6]);
  buf(wbd_adr_o[7], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [7]);
  buf(wbd_adr_o[8], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [8]);
  buf(wbd_adr_o[9], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [9]);
  buf(wbd_adr_o[10], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [10]);
  buf(wbd_adr_o[11], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [11]);
  buf(wbd_adr_o[12], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [12]);
  buf(wbd_adr_o[13], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [13]);
  buf(wbd_adr_o[14], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [14]);
  buf(wbd_adr_o[15], \oc8051_top_1.oc8051_memory_interface1.dadr_ot [15]);
  buf(wbd_dat_o[0], \oc8051_top_1.oc8051_memory_interface1.ddat_o [0]);
  buf(wbd_dat_o[1], \oc8051_top_1.oc8051_memory_interface1.ddat_o [1]);
  buf(wbd_dat_o[2], \oc8051_top_1.oc8051_memory_interface1.ddat_o [2]);
  buf(wbd_dat_o[3], \oc8051_top_1.oc8051_memory_interface1.ddat_o [3]);
  buf(wbd_dat_o[4], \oc8051_top_1.oc8051_memory_interface1.ddat_o [4]);
  buf(wbd_dat_o[5], \oc8051_top_1.oc8051_memory_interface1.ddat_o [5]);
  buf(wbd_dat_o[6], \oc8051_top_1.oc8051_memory_interface1.ddat_o [6]);
  buf(wbd_dat_o[7], \oc8051_top_1.oc8051_memory_interface1.ddat_o [7]);
  buf(wbd_cyc_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_stb_o, \oc8051_top_1.oc8051_memory_interface1.dstb_o );
  buf(wbd_we_o, \oc8051_top_1.oc8051_memory_interface1.dwe_o );
  buf(txd_o, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.txd );
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
