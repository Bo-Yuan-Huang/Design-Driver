
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid, ABINPUT);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  wire _14711_;
  wire _14712_;
  wire _14713_;
  wire _14714_;
  wire _14715_;
  wire _14716_;
  wire _14717_;
  wire _14718_;
  wire _14719_;
  wire _14720_;
  wire _14721_;
  wire _14722_;
  wire _14723_;
  wire _14724_;
  wire _14725_;
  wire _14726_;
  wire _14727_;
  wire _14728_;
  wire _14729_;
  wire _14730_;
  wire _14731_;
  wire _14732_;
  wire _14733_;
  wire _14734_;
  wire _14735_;
  wire _14736_;
  wire _14737_;
  wire _14738_;
  wire _14739_;
  wire _14740_;
  wire _14741_;
  wire _14742_;
  wire _14743_;
  wire _14744_;
  wire _14745_;
  wire _14746_;
  wire _14747_;
  wire _14748_;
  wire _14749_;
  wire _14750_;
  wire _14751_;
  wire _14752_;
  wire _14753_;
  wire _14754_;
  wire _14755_;
  wire _14756_;
  wire _14757_;
  wire _14758_;
  wire _14759_;
  wire _14760_;
  wire _14761_;
  wire _14762_;
  wire _14763_;
  wire _14764_;
  wire _14765_;
  wire _14766_;
  wire _14767_;
  wire _14768_;
  wire _14769_;
  wire _14770_;
  wire _14771_;
  wire _14772_;
  wire _14773_;
  wire _14774_;
  wire _14775_;
  wire _14776_;
  wire _14777_;
  wire _14778_;
  wire _14779_;
  wire _14780_;
  wire _14781_;
  wire _14782_;
  wire _14783_;
  wire _14784_;
  wire _14785_;
  wire _14786_;
  wire _14787_;
  wire _14788_;
  wire _14789_;
  wire _14790_;
  wire _14791_;
  wire _14792_;
  wire _14793_;
  wire _14794_;
  wire _14795_;
  wire _14796_;
  wire _14797_;
  wire _14798_;
  wire _14799_;
  wire _14800_;
  wire _14801_;
  wire _14802_;
  wire _14803_;
  wire _14804_;
  wire _14805_;
  wire _14806_;
  wire _14807_;
  wire _14808_;
  wire _14809_;
  wire _14810_;
  wire _14811_;
  wire _14812_;
  wire _14813_;
  wire _14814_;
  wire _14815_;
  wire _14816_;
  wire _14817_;
  wire _14818_;
  wire _14819_;
  wire _14820_;
  wire _14821_;
  wire _14822_;
  wire _14823_;
  wire _14824_;
  wire _14825_;
  wire _14826_;
  wire _14827_;
  wire _14828_;
  wire _14829_;
  wire _14830_;
  wire _14831_;
  wire _14832_;
  wire _14833_;
  wire _14834_;
  wire _14835_;
  wire _14836_;
  wire _14837_;
  wire _14838_;
  wire _14839_;
  wire _14840_;
  wire _14841_;
  wire _14842_;
  wire _14843_;
  wire _14844_;
  wire _14845_;
  wire _14846_;
  wire _14847_;
  wire _14848_;
  wire _14849_;
  wire _14850_;
  wire _14851_;
  wire _14852_;
  wire _14853_;
  wire _14854_;
  wire _14855_;
  wire _14856_;
  wire _14857_;
  wire _14858_;
  wire _14859_;
  wire _14860_;
  wire _14861_;
  wire _14862_;
  wire _14863_;
  wire _14864_;
  wire _14865_;
  wire _14866_;
  wire _14867_;
  wire _14868_;
  wire _14869_;
  wire _14870_;
  wire _14871_;
  wire _14872_;
  wire _14873_;
  wire _14874_;
  wire _14875_;
  wire _14876_;
  wire _14877_;
  wire _14878_;
  wire _14879_;
  wire _14880_;
  wire _14881_;
  wire _14882_;
  wire _14883_;
  wire _14884_;
  wire _14885_;
  wire _14886_;
  wire _14887_;
  wire _14888_;
  wire _14889_;
  wire _14890_;
  wire _14891_;
  wire _14892_;
  wire _14893_;
  wire _14894_;
  wire _14895_;
  wire _14896_;
  wire _14897_;
  wire _14898_;
  wire _14899_;
  wire _14900_;
  wire _14901_;
  wire _14902_;
  wire _14903_;
  wire _14904_;
  wire _14905_;
  wire _14906_;
  wire _14907_;
  wire _14908_;
  wire _14909_;
  wire _14910_;
  wire _14911_;
  wire _14912_;
  wire _14913_;
  wire _14914_;
  wire _14915_;
  wire _14916_;
  wire _14917_;
  wire _14918_;
  wire _14919_;
  wire _14920_;
  wire _14921_;
  wire _14922_;
  wire _14923_;
  wire _14924_;
  wire _14925_;
  wire _14926_;
  wire _14927_;
  wire _14928_;
  wire _14929_;
  wire _14930_;
  wire _14931_;
  wire _14932_;
  wire _14933_;
  wire _14934_;
  wire _14935_;
  wire _14936_;
  wire _14937_;
  wire _14938_;
  wire _14939_;
  wire _14940_;
  wire _14941_;
  wire _14942_;
  wire _14943_;
  wire _14944_;
  wire _14945_;
  wire _14946_;
  wire _14947_;
  wire _14948_;
  wire _14949_;
  wire _14950_;
  wire _14951_;
  wire _14952_;
  wire _14953_;
  wire _14954_;
  wire _14955_;
  wire _14956_;
  wire _14957_;
  wire _14958_;
  wire _14959_;
  wire _14960_;
  wire _14961_;
  wire _14962_;
  wire _14963_;
  wire _14964_;
  wire _14965_;
  wire _14966_;
  wire _14967_;
  wire _14968_;
  wire _14969_;
  wire _14970_;
  wire _14971_;
  wire _14972_;
  wire _14973_;
  wire _14974_;
  wire _14975_;
  wire _14976_;
  wire _14977_;
  wire _14978_;
  wire _14979_;
  wire _14980_;
  wire _14981_;
  wire _14982_;
  wire _14983_;
  wire _14984_;
  wire _14985_;
  wire _14986_;
  wire _14987_;
  wire _14988_;
  wire _14989_;
  wire _14990_;
  wire _14991_;
  wire _14992_;
  wire _14993_;
  wire _14994_;
  wire _14995_;
  wire _14996_;
  wire _14997_;
  wire _14998_;
  wire _14999_;
  wire _15000_;
  wire _15001_;
  wire _15002_;
  wire _15003_;
  wire _15004_;
  wire _15005_;
  wire _15006_;
  wire _15007_;
  wire _15008_;
  wire _15009_;
  wire _15010_;
  wire _15011_;
  wire _15012_;
  wire _15013_;
  wire _15014_;
  wire _15015_;
  wire _15016_;
  wire _15017_;
  wire _15018_;
  wire _15019_;
  wire _15020_;
  wire _15021_;
  wire _15022_;
  wire _15023_;
  wire _15024_;
  wire _15025_;
  wire _15026_;
  wire _15027_;
  wire _15028_;
  wire _15029_;
  wire _15030_;
  wire _15031_;
  wire _15032_;
  wire _15033_;
  wire _15034_;
  wire _15035_;
  wire _15036_;
  wire _15037_;
  wire _15038_;
  wire _15039_;
  wire _15040_;
  wire _15041_;
  wire _15042_;
  wire _15043_;
  wire _15044_;
  wire _15045_;
  wire _15046_;
  wire _15047_;
  wire _15048_;
  wire _15049_;
  wire _15050_;
  wire _15051_;
  wire _15052_;
  wire _15053_;
  wire _15054_;
  wire _15055_;
  wire _15056_;
  wire _15057_;
  wire _15058_;
  wire _15059_;
  wire _15060_;
  wire _15061_;
  wire _15062_;
  wire _15063_;
  wire _15064_;
  wire _15065_;
  wire _15066_;
  wire _15067_;
  wire _15068_;
  wire _15069_;
  wire _15070_;
  wire _15071_;
  wire _15072_;
  wire _15073_;
  wire _15074_;
  wire _15075_;
  wire _15076_;
  wire _15077_;
  wire _15078_;
  wire _15079_;
  wire _15080_;
  wire _15081_;
  wire _15082_;
  wire _15083_;
  wire _15084_;
  wire _15085_;
  wire _15086_;
  wire _15087_;
  wire _15088_;
  wire _15089_;
  wire _15090_;
  wire _15091_;
  wire _15092_;
  wire _15093_;
  wire _15094_;
  wire _15095_;
  wire _15096_;
  wire _15097_;
  wire _15098_;
  wire _15099_;
  wire _15100_;
  wire _15101_;
  wire _15102_;
  wire _15103_;
  wire _15104_;
  wire _15105_;
  wire _15106_;
  wire _15107_;
  wire _15108_;
  wire _15109_;
  wire _15110_;
  wire _15111_;
  wire _15112_;
  wire _15113_;
  wire _15114_;
  wire _15115_;
  wire _15116_;
  wire _15117_;
  wire _15118_;
  wire _15119_;
  wire _15120_;
  wire _15121_;
  wire _15122_;
  wire _15123_;
  wire _15124_;
  wire _15125_;
  wire _15126_;
  wire _15127_;
  wire _15128_;
  wire _15129_;
  wire _15130_;
  wire _15131_;
  wire _15132_;
  wire _15133_;
  wire _15134_;
  wire _15135_;
  wire _15136_;
  wire _15137_;
  wire _15138_;
  wire _15139_;
  wire _15140_;
  wire _15141_;
  wire _15142_;
  wire _15143_;
  wire _15144_;
  wire _15145_;
  wire _15146_;
  wire _15147_;
  wire _15148_;
  wire _15149_;
  wire _15150_;
  wire _15151_;
  wire _15152_;
  wire _15153_;
  wire _15154_;
  wire _15155_;
  wire _15156_;
  wire _15157_;
  wire _15158_;
  wire _15159_;
  wire _15160_;
  wire _15161_;
  wire _15162_;
  wire _15163_;
  wire _15164_;
  wire _15165_;
  wire _15166_;
  wire _15167_;
  wire _15168_;
  wire _15169_;
  wire _15170_;
  wire _15171_;
  wire _15172_;
  wire _15173_;
  wire _15174_;
  wire _15175_;
  wire _15176_;
  wire _15177_;
  wire _15178_;
  wire _15179_;
  wire _15180_;
  wire _15181_;
  wire _15182_;
  wire _15183_;
  wire _15184_;
  wire _15185_;
  wire _15186_;
  wire _15187_;
  wire _15188_;
  wire _15189_;
  wire _15190_;
  wire _15191_;
  wire _15192_;
  wire _15193_;
  wire _15194_;
  wire _15195_;
  wire _15196_;
  wire _15197_;
  wire _15198_;
  wire _15199_;
  wire _15200_;
  wire _15201_;
  wire _15202_;
  wire _15203_;
  wire _15204_;
  wire _15205_;
  wire _15206_;
  wire _15207_;
  wire _15208_;
  wire _15209_;
  wire _15210_;
  wire _15211_;
  wire _15212_;
  wire _15213_;
  wire _15214_;
  wire _15215_;
  wire _15216_;
  wire _15217_;
  wire _15218_;
  wire _15219_;
  wire _15220_;
  wire _15221_;
  wire _15222_;
  wire _15223_;
  wire _15224_;
  wire _15225_;
  wire _15226_;
  wire _15227_;
  wire _15228_;
  wire _15229_;
  wire _15230_;
  wire _15231_;
  wire _15232_;
  wire _15233_;
  wire _15234_;
  wire _15235_;
  wire _15236_;
  wire _15237_;
  wire _15238_;
  wire _15239_;
  wire _15240_;
  wire _15241_;
  wire _15242_;
  wire _15243_;
  wire _15244_;
  wire _15245_;
  wire _15246_;
  wire _15247_;
  wire _15248_;
  wire _15249_;
  wire _15250_;
  wire _15251_;
  wire _15252_;
  wire _15253_;
  wire _15254_;
  wire _15255_;
  wire _15256_;
  wire _15257_;
  wire _15258_;
  wire _15259_;
  wire _15260_;
  wire _15261_;
  wire _15262_;
  wire _15263_;
  wire _15264_;
  wire _15265_;
  wire _15266_;
  wire _15267_;
  wire _15268_;
  wire _15269_;
  wire _15270_;
  wire _15271_;
  wire _15272_;
  wire _15273_;
  wire _15274_;
  wire _15275_;
  wire _15276_;
  wire _15277_;
  wire _15278_;
  wire _15279_;
  wire _15280_;
  wire _15281_;
  wire _15282_;
  wire _15283_;
  wire _15284_;
  wire _15285_;
  wire _15286_;
  wire _15287_;
  wire _15288_;
  wire _15289_;
  wire _15290_;
  wire _15291_;
  wire _15292_;
  wire _15293_;
  wire _15294_;
  wire _15295_;
  wire _15296_;
  wire _15297_;
  wire _15298_;
  wire _15299_;
  wire _15300_;
  wire _15301_;
  wire _15302_;
  wire _15303_;
  wire _15304_;
  wire _15305_;
  wire _15306_;
  wire _15307_;
  wire _15308_;
  wire _15309_;
  wire _15310_;
  wire _15311_;
  wire _15312_;
  wire _15313_;
  wire _15314_;
  wire _15315_;
  wire _15316_;
  wire _15317_;
  wire _15318_;
  wire _15319_;
  wire _15320_;
  wire _15321_;
  wire _15322_;
  wire _15323_;
  wire _15324_;
  wire _15325_;
  wire _15326_;
  wire _15327_;
  wire _15328_;
  wire _15329_;
  wire _15330_;
  wire _15331_;
  wire _15332_;
  wire _15333_;
  wire _15334_;
  wire _15335_;
  wire _15336_;
  wire _15337_;
  wire _15338_;
  wire _15339_;
  wire _15340_;
  wire _15341_;
  wire _15342_;
  wire _15343_;
  wire _15344_;
  wire _15345_;
  wire _15346_;
  wire _15347_;
  wire _15348_;
  wire _15349_;
  wire _15350_;
  wire _15351_;
  wire _15352_;
  wire _15353_;
  wire _15354_;
  wire _15355_;
  wire _15356_;
  wire _15357_;
  wire _15358_;
  wire _15359_;
  wire _15360_;
  wire _15361_;
  wire _15362_;
  wire _15363_;
  wire _15364_;
  wire _15365_;
  wire _15366_;
  wire _15367_;
  wire _15368_;
  wire _15369_;
  wire _15370_;
  wire _15371_;
  wire _15372_;
  wire _15373_;
  wire _15374_;
  wire _15375_;
  wire _15376_;
  wire _15377_;
  wire _15378_;
  wire _15379_;
  wire _15380_;
  wire _15381_;
  wire _15382_;
  wire _15383_;
  wire _15384_;
  wire _15385_;
  wire _15386_;
  wire _15387_;
  wire _15388_;
  wire _15389_;
  wire _15390_;
  wire _15391_;
  wire _15392_;
  wire _15393_;
  wire _15394_;
  wire _15395_;
  wire _15396_;
  wire _15397_;
  wire _15398_;
  wire _15399_;
  wire _15400_;
  wire _15401_;
  wire _15402_;
  wire _15403_;
  wire _15404_;
  wire _15405_;
  wire _15406_;
  wire _15407_;
  wire _15408_;
  wire _15409_;
  wire _15410_;
  wire _15411_;
  wire _15412_;
  wire _15413_;
  wire _15414_;
  wire _15415_;
  wire _15416_;
  wire _15417_;
  wire _15418_;
  wire _15419_;
  wire _15420_;
  wire _15421_;
  wire _15422_;
  wire _15423_;
  wire _15424_;
  wire _15425_;
  wire _15426_;
  wire _15427_;
  wire _15428_;
  wire _15429_;
  wire _15430_;
  wire _15431_;
  wire _15432_;
  wire _15433_;
  wire _15434_;
  wire _15435_;
  wire _15436_;
  wire _15437_;
  wire _15438_;
  wire _15439_;
  wire _15440_;
  wire _15441_;
  wire _15442_;
  wire _15443_;
  wire _15444_;
  wire _15445_;
  wire _15446_;
  wire _15447_;
  wire _15448_;
  wire _15449_;
  wire _15450_;
  wire _15451_;
  wire _15452_;
  wire _15453_;
  wire _15454_;
  wire _15455_;
  wire _15456_;
  wire _15457_;
  wire _15458_;
  wire _15459_;
  wire _15460_;
  wire _15461_;
  wire _15462_;
  wire _15463_;
  wire _15464_;
  wire _15465_;
  wire _15466_;
  wire _15467_;
  wire _15468_;
  wire _15469_;
  wire _15470_;
  wire _15471_;
  wire _15472_;
  wire _15473_;
  wire _15474_;
  wire _15475_;
  wire _15476_;
  wire _15477_;
  wire _15478_;
  wire _15479_;
  wire _15480_;
  wire _15481_;
  wire _15482_;
  wire _15483_;
  wire _15484_;
  wire _15485_;
  wire _15486_;
  wire _15487_;
  wire _15488_;
  wire _15489_;
  wire _15490_;
  wire _15491_;
  wire _15492_;
  wire _15493_;
  wire _15494_;
  wire _15495_;
  wire _15496_;
  wire _15497_;
  wire _15498_;
  wire _15499_;
  wire _15500_;
  wire _15501_;
  wire _15502_;
  wire _15503_;
  wire _15504_;
  wire _15505_;
  wire _15506_;
  wire _15507_;
  wire _15508_;
  wire _15509_;
  wire _15510_;
  wire _15511_;
  wire _15512_;
  wire _15513_;
  wire _15514_;
  wire _15515_;
  wire _15516_;
  wire _15517_;
  wire _15518_;
  wire _15519_;
  wire _15520_;
  wire _15521_;
  wire _15522_;
  wire _15523_;
  wire _15524_;
  wire _15525_;
  wire _15526_;
  wire _15527_;
  wire _15528_;
  wire _15529_;
  wire _15530_;
  wire _15531_;
  wire _15532_;
  wire _15533_;
  wire _15534_;
  wire _15535_;
  wire _15536_;
  wire _15537_;
  wire _15538_;
  wire _15539_;
  wire _15540_;
  wire _15541_;
  wire _15542_;
  wire _15543_;
  wire _15544_;
  wire _15545_;
  wire _15546_;
  wire _15547_;
  wire _15548_;
  wire _15549_;
  wire _15550_;
  wire _15551_;
  wire _15552_;
  wire _15553_;
  wire _15554_;
  wire _15555_;
  wire _15556_;
  wire _15557_;
  wire _15558_;
  wire _15559_;
  wire _15560_;
  wire _15561_;
  wire _15562_;
  wire _15563_;
  wire _15564_;
  wire _15565_;
  wire _15566_;
  wire _15567_;
  wire _15568_;
  wire _15569_;
  wire _15570_;
  wire _15571_;
  wire _15572_;
  wire _15573_;
  wire _15574_;
  wire _15575_;
  wire _15576_;
  wire _15577_;
  wire _15578_;
  wire _15579_;
  wire _15580_;
  wire _15581_;
  wire _15582_;
  wire _15583_;
  wire _15584_;
  wire _15585_;
  wire _15586_;
  wire _15587_;
  wire _15588_;
  wire _15589_;
  wire _15590_;
  wire _15591_;
  wire _15592_;
  wire _15593_;
  wire _15594_;
  wire _15595_;
  wire _15596_;
  wire _15597_;
  wire _15598_;
  wire _15599_;
  wire _15600_;
  wire _15601_;
  wire _15602_;
  wire _15603_;
  wire _15604_;
  wire _15605_;
  wire _15606_;
  wire _15607_;
  wire _15608_;
  wire _15609_;
  wire _15610_;
  wire _15611_;
  wire _15612_;
  wire _15613_;
  wire _15614_;
  wire _15615_;
  wire _15616_;
  wire _15617_;
  wire _15618_;
  wire _15619_;
  wire _15620_;
  wire _15621_;
  wire _15622_;
  wire _15623_;
  wire _15624_;
  wire _15625_;
  wire _15626_;
  wire _15627_;
  wire _15628_;
  wire _15629_;
  wire _15630_;
  wire _15631_;
  wire _15632_;
  wire _15633_;
  wire _15634_;
  wire _15635_;
  wire _15636_;
  wire _15637_;
  wire _15638_;
  wire _15639_;
  wire _15640_;
  wire _15641_;
  wire _15642_;
  wire _15643_;
  wire _15644_;
  wire _15645_;
  wire _15646_;
  wire _15647_;
  wire _15648_;
  wire _15649_;
  wire _15650_;
  wire _15651_;
  wire _15652_;
  wire _15653_;
  wire _15654_;
  wire _15655_;
  wire _15656_;
  wire _15657_;
  wire _15658_;
  wire _15659_;
  wire _15660_;
  wire _15661_;
  wire _15662_;
  wire _15663_;
  wire _15664_;
  wire _15665_;
  wire _15666_;
  wire _15667_;
  wire _15668_;
  wire _15669_;
  wire _15670_;
  wire _15671_;
  wire _15672_;
  wire _15673_;
  wire _15674_;
  wire _15675_;
  wire _15676_;
  wire _15677_;
  wire _15678_;
  wire _15679_;
  wire _15680_;
  wire _15681_;
  wire _15682_;
  wire _15683_;
  wire _15684_;
  wire _15685_;
  wire _15686_;
  wire _15687_;
  wire _15688_;
  wire _15689_;
  wire _15690_;
  wire _15691_;
  wire _15692_;
  wire _15693_;
  wire _15694_;
  wire _15695_;
  wire _15696_;
  wire _15697_;
  wire _15698_;
  wire _15699_;
  wire _15700_;
  wire _15701_;
  wire _15702_;
  wire _15703_;
  wire _15704_;
  wire _15705_;
  wire _15706_;
  wire _15707_;
  wire _15708_;
  wire _15709_;
  wire _15710_;
  wire _15711_;
  wire _15712_;
  wire _15713_;
  wire _15714_;
  wire _15715_;
  wire _15716_;
  wire _15717_;
  wire _15718_;
  wire _15719_;
  wire _15720_;
  wire _15721_;
  wire _15722_;
  wire _15723_;
  wire _15724_;
  wire _15725_;
  wire _15726_;
  wire _15727_;
  wire _15728_;
  wire _15729_;
  wire _15730_;
  wire _15731_;
  wire _15732_;
  wire _15733_;
  wire _15734_;
  wire _15735_;
  wire _15736_;
  wire _15737_;
  wire _15738_;
  wire _15739_;
  wire _15740_;
  wire _15741_;
  wire _15742_;
  wire _15743_;
  wire _15744_;
  wire _15745_;
  wire _15746_;
  wire _15747_;
  wire _15748_;
  wire _15749_;
  wire _15750_;
  wire _15751_;
  wire _15752_;
  wire _15753_;
  wire _15754_;
  wire _15755_;
  wire _15756_;
  wire _15757_;
  wire _15758_;
  wire _15759_;
  wire _15760_;
  wire _15761_;
  wire _15762_;
  wire _15763_;
  wire _15764_;
  wire _15765_;
  wire _15766_;
  wire _15767_;
  wire _15768_;
  wire _15769_;
  wire _15770_;
  wire _15771_;
  wire _15772_;
  wire _15773_;
  wire _15774_;
  wire _15775_;
  wire _15776_;
  wire _15777_;
  wire _15778_;
  wire _15779_;
  wire _15780_;
  wire _15781_;
  wire _15782_;
  wire _15783_;
  wire _15784_;
  wire _15785_;
  wire _15786_;
  wire _15787_;
  wire _15788_;
  wire _15789_;
  wire _15790_;
  wire _15791_;
  wire _15792_;
  wire _15793_;
  wire _15794_;
  wire _15795_;
  wire _15796_;
  wire _15797_;
  wire _15798_;
  wire _15799_;
  wire _15800_;
  wire _15801_;
  wire _15802_;
  wire _15803_;
  wire _15804_;
  wire _15805_;
  wire _15806_;
  wire _15807_;
  wire _15808_;
  wire _15809_;
  wire _15810_;
  wire _15811_;
  wire _15812_;
  wire _15813_;
  wire _15814_;
  wire _15815_;
  wire _15816_;
  wire _15817_;
  wire _15818_;
  wire _15819_;
  wire _15820_;
  wire _15821_;
  wire _15822_;
  wire _15823_;
  wire _15824_;
  wire _15825_;
  wire _15826_;
  wire _15827_;
  wire _15828_;
  wire _15829_;
  wire _15830_;
  wire _15831_;
  wire _15832_;
  wire _15833_;
  wire _15834_;
  wire _15835_;
  wire _15836_;
  wire _15837_;
  wire _15838_;
  wire _15839_;
  wire _15840_;
  wire _15841_;
  wire _15842_;
  wire _15843_;
  wire _15844_;
  wire _15845_;
  wire _15846_;
  wire _15847_;
  wire _15848_;
  wire _15849_;
  wire _15850_;
  wire _15851_;
  wire _15852_;
  wire _15853_;
  wire _15854_;
  wire _15855_;
  wire _15856_;
  wire _15857_;
  wire _15858_;
  wire _15859_;
  wire _15860_;
  wire _15861_;
  wire _15862_;
  wire _15863_;
  wire _15864_;
  wire _15865_;
  wire _15866_;
  wire _15867_;
  wire _15868_;
  wire _15869_;
  wire _15870_;
  wire _15871_;
  wire _15872_;
  wire _15873_;
  wire _15874_;
  wire _15875_;
  wire _15876_;
  wire _15877_;
  wire _15878_;
  wire _15879_;
  wire _15880_;
  wire _15881_;
  wire _15882_;
  wire _15883_;
  wire _15884_;
  wire _15885_;
  wire _15886_;
  wire _15887_;
  wire _15888_;
  wire _15889_;
  wire _15890_;
  wire _15891_;
  wire _15892_;
  wire _15893_;
  wire _15894_;
  wire _15895_;
  wire _15896_;
  wire _15897_;
  wire _15898_;
  wire _15899_;
  wire _15900_;
  wire _15901_;
  wire _15902_;
  wire _15903_;
  wire _15904_;
  wire _15905_;
  wire _15906_;
  wire _15907_;
  wire _15908_;
  wire _15909_;
  wire _15910_;
  wire _15911_;
  wire _15912_;
  wire _15913_;
  wire _15914_;
  wire _15915_;
  wire _15916_;
  wire _15917_;
  wire _15918_;
  wire _15919_;
  wire _15920_;
  wire _15921_;
  wire _15922_;
  wire _15923_;
  wire _15924_;
  wire _15925_;
  wire _15926_;
  wire _15927_;
  wire _15928_;
  wire _15929_;
  wire _15930_;
  wire _15931_;
  wire _15932_;
  wire _15933_;
  wire _15934_;
  wire _15935_;
  wire _15936_;
  wire _15937_;
  wire _15938_;
  wire _15939_;
  wire _15940_;
  wire _15941_;
  wire _15942_;
  wire _15943_;
  wire _15944_;
  wire _15945_;
  wire _15946_;
  wire _15947_;
  wire _15948_;
  wire _15949_;
  wire _15950_;
  wire _15951_;
  wire _15952_;
  wire _15953_;
  wire _15954_;
  wire _15955_;
  wire _15956_;
  wire _15957_;
  wire _15958_;
  wire _15959_;
  wire _15960_;
  wire _15961_;
  wire _15962_;
  wire _15963_;
  wire _15964_;
  wire _15965_;
  wire _15966_;
  wire _15967_;
  wire _15968_;
  wire _15969_;
  wire _15970_;
  wire _15971_;
  wire _15972_;
  wire _15973_;
  wire _15974_;
  wire _15975_;
  wire _15976_;
  wire _15977_;
  wire _15978_;
  wire _15979_;
  wire _15980_;
  wire _15981_;
  wire _15982_;
  wire _15983_;
  wire _15984_;
  wire _15985_;
  wire _15986_;
  wire _15987_;
  wire _15988_;
  wire _15989_;
  wire _15990_;
  wire _15991_;
  wire _15992_;
  wire _15993_;
  wire _15994_;
  wire _15995_;
  wire _15996_;
  wire _15997_;
  wire _15998_;
  wire _15999_;
  wire _16000_;
  wire _16001_;
  wire _16002_;
  wire _16003_;
  wire _16004_;
  wire _16005_;
  wire _16006_;
  wire _16007_;
  wire _16008_;
  wire _16009_;
  wire _16010_;
  wire _16011_;
  wire _16012_;
  wire _16013_;
  wire _16014_;
  wire _16015_;
  wire _16016_;
  wire _16017_;
  wire _16018_;
  wire _16019_;
  wire _16020_;
  wire _16021_;
  wire _16022_;
  wire _16023_;
  wire _16024_;
  wire _16025_;
  wire _16026_;
  wire _16027_;
  wire _16028_;
  wire _16029_;
  wire _16030_;
  wire _16031_;
  wire _16032_;
  wire _16033_;
  wire _16034_;
  wire _16035_;
  wire _16036_;
  wire _16037_;
  wire _16038_;
  wire _16039_;
  wire _16040_;
  wire _16041_;
  wire _16042_;
  wire _16043_;
  wire _16044_;
  wire _16045_;
  wire _16046_;
  wire _16047_;
  wire _16048_;
  wire _16049_;
  wire _16050_;
  wire _16051_;
  wire _16052_;
  wire _16053_;
  wire _16054_;
  wire _16055_;
  wire _16056_;
  wire _16057_;
  wire _16058_;
  wire _16059_;
  wire _16060_;
  wire _16061_;
  wire _16062_;
  wire _16063_;
  wire _16064_;
  wire _16065_;
  wire _16066_;
  wire _16067_;
  wire _16068_;
  wire _16069_;
  wire _16070_;
  wire _16071_;
  wire _16072_;
  wire _16073_;
  wire _16074_;
  wire _16075_;
  wire _16076_;
  wire _16077_;
  wire _16078_;
  wire _16079_;
  wire _16080_;
  wire _16081_;
  wire _16082_;
  wire _16083_;
  wire _16084_;
  wire _16085_;
  wire _16086_;
  wire _16087_;
  wire _16088_;
  wire _16089_;
  wire _16090_;
  wire _16091_;
  wire _16092_;
  wire _16093_;
  wire _16094_;
  wire _16095_;
  wire _16096_;
  wire _16097_;
  wire _16098_;
  wire _16099_;
  wire _16100_;
  wire _16101_;
  wire _16102_;
  wire _16103_;
  wire _16104_;
  wire _16105_;
  wire _16106_;
  wire _16107_;
  wire _16108_;
  wire _16109_;
  wire _16110_;
  wire _16111_;
  wire _16112_;
  wire _16113_;
  wire _16114_;
  wire _16115_;
  wire _16116_;
  wire _16117_;
  wire _16118_;
  wire _16119_;
  wire _16120_;
  wire _16121_;
  wire _16122_;
  wire _16123_;
  wire _16124_;
  wire _16125_;
  wire _16126_;
  wire _16127_;
  wire _16128_;
  wire _16129_;
  wire _16130_;
  wire _16131_;
  wire _16132_;
  wire _16133_;
  wire _16134_;
  wire _16135_;
  wire _16136_;
  wire _16137_;
  wire _16138_;
  wire _16139_;
  wire _16140_;
  wire _16141_;
  wire _16142_;
  wire _16143_;
  wire _16144_;
  wire _16145_;
  wire _16146_;
  wire _16147_;
  wire _16148_;
  wire _16149_;
  wire _16150_;
  wire _16151_;
  wire _16152_;
  wire _16153_;
  wire _16154_;
  wire _16155_;
  wire _16156_;
  wire _16157_;
  wire _16158_;
  wire _16159_;
  wire _16160_;
  wire _16161_;
  wire _16162_;
  wire _16163_;
  wire _16164_;
  wire _16165_;
  wire _16166_;
  wire _16167_;
  wire _16168_;
  wire _16169_;
  wire _16170_;
  wire _16171_;
  wire _16172_;
  wire _16173_;
  wire _16174_;
  wire _16175_;
  wire _16176_;
  wire _16177_;
  wire _16178_;
  wire _16179_;
  wire _16180_;
  wire _16181_;
  wire _16182_;
  wire _16183_;
  wire _16184_;
  wire _16185_;
  wire _16186_;
  wire _16187_;
  wire _16188_;
  wire _16189_;
  wire _16190_;
  wire _16191_;
  wire _16192_;
  wire _16193_;
  wire _16194_;
  wire _16195_;
  wire _16196_;
  wire _16197_;
  wire _16198_;
  wire _16199_;
  wire _16200_;
  wire _16201_;
  wire _16202_;
  wire _16203_;
  wire _16204_;
  wire _16205_;
  wire _16206_;
  wire _16207_;
  wire _16208_;
  wire _16209_;
  wire _16210_;
  wire _16211_;
  wire _16212_;
  wire _16213_;
  wire _16214_;
  wire _16215_;
  wire _16216_;
  wire _16217_;
  wire _16218_;
  wire _16219_;
  wire _16220_;
  wire _16221_;
  wire _16222_;
  wire _16223_;
  wire _16224_;
  wire _16225_;
  wire _16226_;
  wire _16227_;
  wire _16228_;
  wire _16229_;
  wire _16230_;
  wire _16231_;
  wire _16232_;
  wire _16233_;
  wire _16234_;
  wire _16235_;
  wire _16236_;
  wire _16237_;
  wire _16238_;
  wire _16239_;
  wire _16240_;
  wire _16241_;
  wire _16242_;
  wire _16243_;
  wire _16244_;
  wire _16245_;
  wire _16246_;
  wire _16247_;
  wire _16248_;
  wire _16249_;
  wire _16250_;
  wire _16251_;
  wire _16252_;
  wire _16253_;
  wire _16254_;
  wire _16255_;
  wire _16256_;
  wire _16257_;
  wire _16258_;
  wire _16259_;
  wire _16260_;
  wire _16261_;
  wire _16262_;
  wire _16263_;
  wire _16264_;
  wire _16265_;
  wire _16266_;
  wire _16267_;
  wire _16268_;
  wire _16269_;
  wire _16270_;
  wire _16271_;
  wire _16272_;
  wire _16273_;
  wire _16274_;
  wire _16275_;
  wire _16276_;
  wire _16277_;
  wire _16278_;
  wire _16279_;
  wire _16280_;
  wire _16281_;
  wire _16282_;
  wire _16283_;
  wire _16284_;
  wire _16285_;
  wire _16286_;
  wire _16287_;
  wire _16288_;
  wire _16289_;
  wire _16290_;
  wire _16291_;
  wire _16292_;
  wire _16293_;
  wire _16294_;
  wire _16295_;
  wire _16296_;
  wire _16297_;
  wire _16298_;
  wire _16299_;
  wire _16300_;
  wire _16301_;
  wire _16302_;
  wire _16303_;
  wire _16304_;
  wire _16305_;
  wire _16306_;
  wire _16307_;
  wire _16308_;
  wire _16309_;
  wire _16310_;
  wire _16311_;
  wire _16312_;
  wire _16313_;
  wire _16314_;
  wire _16315_;
  wire _16316_;
  wire _16317_;
  wire _16318_;
  wire _16319_;
  wire _16320_;
  wire _16321_;
  wire _16322_;
  wire _16323_;
  wire _16324_;
  wire _16325_;
  wire _16326_;
  wire _16327_;
  wire _16328_;
  wire _16329_;
  wire _16330_;
  wire _16331_;
  wire _16332_;
  wire _16333_;
  wire _16334_;
  wire _16335_;
  wire _16336_;
  wire _16337_;
  wire _16338_;
  wire _16339_;
  wire _16340_;
  wire _16341_;
  wire _16342_;
  wire _16343_;
  wire _16344_;
  wire _16345_;
  wire _16346_;
  wire _16347_;
  wire _16348_;
  wire _16349_;
  wire _16350_;
  wire _16351_;
  wire _16352_;
  wire _16353_;
  wire _16354_;
  wire _16355_;
  wire _16356_;
  wire _16357_;
  wire _16358_;
  wire _16359_;
  wire _16360_;
  wire _16361_;
  wire _16362_;
  wire _16363_;
  wire _16364_;
  wire _16365_;
  wire _16366_;
  wire _16367_;
  wire _16368_;
  wire _16369_;
  wire _16370_;
  wire _16371_;
  wire _16372_;
  wire _16373_;
  wire _16374_;
  wire _16375_;
  wire _16376_;
  wire _16377_;
  wire _16378_;
  wire _16379_;
  wire _16380_;
  wire _16381_;
  wire _16382_;
  wire _16383_;
  wire _16384_;
  wire _16385_;
  wire _16386_;
  wire _16387_;
  wire _16388_;
  wire _16389_;
  wire _16390_;
  wire _16391_;
  wire _16392_;
  wire _16393_;
  wire _16394_;
  wire _16395_;
  wire _16396_;
  wire _16397_;
  wire _16398_;
  wire _16399_;
  wire _16400_;
  wire _16401_;
  wire _16402_;
  wire _16403_;
  wire _16404_;
  wire _16405_;
  wire _16406_;
  wire _16407_;
  wire _16408_;
  wire _16409_;
  wire _16410_;
  wire _16411_;
  wire _16412_;
  wire _16413_;
  wire _16414_;
  wire _16415_;
  wire _16416_;
  wire _16417_;
  wire _16418_;
  wire _16419_;
  wire _16420_;
  wire _16421_;
  wire _16422_;
  wire _16423_;
  wire _16424_;
  wire _16425_;
  wire _16426_;
  wire _16427_;
  wire _16428_;
  wire _16429_;
  wire _16430_;
  wire _16431_;
  wire _16432_;
  wire _16433_;
  wire _16434_;
  wire _16435_;
  wire _16436_;
  wire _16437_;
  wire _16438_;
  wire _16439_;
  wire _16440_;
  wire _16441_;
  wire _16442_;
  wire _16443_;
  wire _16444_;
  wire _16445_;
  wire _16446_;
  wire _16447_;
  wire _16448_;
  wire _16449_;
  wire _16450_;
  wire _16451_;
  wire _16452_;
  wire _16453_;
  wire _16454_;
  wire _16455_;
  wire _16456_;
  wire _16457_;
  wire _16458_;
  wire _16459_;
  wire _16460_;
  wire _16461_;
  wire _16462_;
  wire _16463_;
  wire _16464_;
  wire _16465_;
  wire _16466_;
  wire _16467_;
  wire _16468_;
  wire _16469_;
  wire _16470_;
  wire _16471_;
  wire _16472_;
  wire _16473_;
  wire _16474_;
  wire _16475_;
  wire _16476_;
  wire _16477_;
  wire _16478_;
  wire _16479_;
  wire _16480_;
  wire _16481_;
  wire _16482_;
  wire _16483_;
  wire _16484_;
  wire _16485_;
  wire _16486_;
  wire _16487_;
  wire _16488_;
  wire _16489_;
  wire _16490_;
  wire _16491_;
  wire _16492_;
  wire _16493_;
  wire _16494_;
  wire _16495_;
  wire _16496_;
  wire _16497_;
  wire _16498_;
  wire _16499_;
  wire _16500_;
  wire _16501_;
  wire _16502_;
  wire _16503_;
  wire _16504_;
  wire _16505_;
  wire _16506_;
  wire _16507_;
  wire _16508_;
  wire _16509_;
  wire _16510_;
  wire _16511_;
  wire _16512_;
  wire _16513_;
  wire _16514_;
  wire _16515_;
  wire _16516_;
  wire _16517_;
  wire _16518_;
  wire _16519_;
  wire _16520_;
  wire _16521_;
  wire _16522_;
  wire _16523_;
  wire _16524_;
  wire _16525_;
  wire _16526_;
  wire _16527_;
  wire _16528_;
  wire _16529_;
  wire _16530_;
  wire _16531_;
  wire _16532_;
  wire _16533_;
  wire _16534_;
  wire _16535_;
  wire _16536_;
  wire _16537_;
  wire _16538_;
  wire _16539_;
  wire _16540_;
  wire _16541_;
  wire _16542_;
  wire _16543_;
  wire _16544_;
  wire _16545_;
  wire _16546_;
  wire _16547_;
  wire _16548_;
  wire _16549_;
  wire _16550_;
  wire _16551_;
  wire _16552_;
  wire _16553_;
  wire _16554_;
  wire _16555_;
  wire _16556_;
  wire _16557_;
  wire _16558_;
  wire _16559_;
  wire _16560_;
  wire _16561_;
  wire _16562_;
  wire _16563_;
  wire _16564_;
  wire _16565_;
  wire _16566_;
  wire _16567_;
  wire _16568_;
  wire _16569_;
  wire _16570_;
  wire _16571_;
  wire _16572_;
  wire _16573_;
  wire _16574_;
  wire _16575_;
  wire _16576_;
  wire _16577_;
  wire _16578_;
  wire _16579_;
  wire _16580_;
  wire _16581_;
  wire _16582_;
  wire _16583_;
  wire _16584_;
  wire _16585_;
  wire _16586_;
  wire _16587_;
  wire _16588_;
  wire _16589_;
  wire _16590_;
  wire _16591_;
  wire _16592_;
  wire _16593_;
  wire _16594_;
  wire _16595_;
  wire _16596_;
  wire _16597_;
  wire _16598_;
  wire _16599_;
  wire _16600_;
  wire _16601_;
  wire _16602_;
  wire _16603_;
  wire _16604_;
  wire _16605_;
  wire _16606_;
  wire _16607_;
  wire _16608_;
  wire _16609_;
  wire _16610_;
  wire _16611_;
  wire _16612_;
  wire _16613_;
  wire _16614_;
  wire _16615_;
  wire _16616_;
  wire _16617_;
  wire _16618_;
  wire _16619_;
  wire _16620_;
  wire _16621_;
  wire _16622_;
  wire _16623_;
  wire _16624_;
  wire _16625_;
  wire _16626_;
  wire _16627_;
  wire _16628_;
  wire _16629_;
  wire _16630_;
  wire _16631_;
  wire _16632_;
  wire _16633_;
  wire _16634_;
  wire _16635_;
  wire _16636_;
  wire _16637_;
  wire _16638_;
  wire _16639_;
  wire _16640_;
  wire _16641_;
  wire _16642_;
  wire _16643_;
  wire _16644_;
  wire _16645_;
  wire _16646_;
  wire _16647_;
  wire _16648_;
  wire _16649_;
  wire _16650_;
  wire _16651_;
  wire _16652_;
  wire _16653_;
  wire _16654_;
  wire _16655_;
  wire _16656_;
  wire _16657_;
  wire _16658_;
  wire _16659_;
  wire _16660_;
  wire _16661_;
  wire _16662_;
  wire _16663_;
  wire _16664_;
  wire _16665_;
  wire _16666_;
  wire _16667_;
  wire _16668_;
  wire _16669_;
  wire _16670_;
  wire _16671_;
  wire _16672_;
  wire _16673_;
  wire _16674_;
  wire _16675_;
  wire _16676_;
  wire _16677_;
  wire _16678_;
  wire _16679_;
  wire _16680_;
  wire _16681_;
  wire _16682_;
  wire _16683_;
  wire _16684_;
  wire _16685_;
  wire _16686_;
  wire _16687_;
  wire _16688_;
  wire _16689_;
  wire _16690_;
  wire _16691_;
  wire _16692_;
  wire _16693_;
  wire _16694_;
  wire _16695_;
  wire _16696_;
  wire _16697_;
  wire _16698_;
  wire _16699_;
  wire _16700_;
  wire _16701_;
  wire _16702_;
  wire _16703_;
  wire _16704_;
  wire _16705_;
  wire _16706_;
  wire _16707_;
  wire _16708_;
  wire _16709_;
  wire _16710_;
  wire _16711_;
  wire _16712_;
  wire _16713_;
  wire _16714_;
  wire _16715_;
  wire _16716_;
  wire _16717_;
  wire _16718_;
  wire _16719_;
  wire _16720_;
  wire _16721_;
  wire _16722_;
  wire _16723_;
  wire _16724_;
  wire _16725_;
  wire _16726_;
  wire _16727_;
  wire _16728_;
  wire _16729_;
  wire _16730_;
  wire _16731_;
  wire _16732_;
  wire _16733_;
  wire _16734_;
  wire _16735_;
  wire _16736_;
  wire _16737_;
  wire _16738_;
  wire _16739_;
  wire _16740_;
  wire _16741_;
  wire _16742_;
  wire _16743_;
  wire _16744_;
  wire _16745_;
  wire _16746_;
  wire _16747_;
  wire _16748_;
  wire _16749_;
  wire _16750_;
  wire _16751_;
  wire _16752_;
  wire _16753_;
  wire _16754_;
  wire _16755_;
  wire _16756_;
  wire _16757_;
  wire _16758_;
  wire _16759_;
  wire _16760_;
  wire _16761_;
  wire _16762_;
  wire _16763_;
  wire _16764_;
  wire _16765_;
  wire _16766_;
  wire _16767_;
  wire _16768_;
  wire _16769_;
  wire _16770_;
  wire _16771_;
  wire _16772_;
  wire _16773_;
  wire _16774_;
  wire _16775_;
  wire _16776_;
  wire _16777_;
  wire _16778_;
  wire _16779_;
  wire _16780_;
  wire _16781_;
  wire _16782_;
  wire _16783_;
  wire _16784_;
  wire _16785_;
  wire _16786_;
  wire _16787_;
  wire _16788_;
  wire _16789_;
  wire _16790_;
  wire _16791_;
  wire _16792_;
  wire _16793_;
  wire _16794_;
  wire _16795_;
  wire _16796_;
  wire _16797_;
  wire _16798_;
  wire _16799_;
  wire _16800_;
  wire _16801_;
  wire _16802_;
  wire _16803_;
  wire _16804_;
  wire _16805_;
  wire _16806_;
  wire _16807_;
  wire _16808_;
  wire _16809_;
  wire _16810_;
  wire _16811_;
  wire _16812_;
  wire _16813_;
  wire _16814_;
  wire _16815_;
  wire _16816_;
  wire _16817_;
  wire _16818_;
  wire _16819_;
  wire _16820_;
  wire _16821_;
  wire _16822_;
  wire _16823_;
  wire _16824_;
  wire _16825_;
  wire _16826_;
  wire _16827_;
  wire _16828_;
  wire _16829_;
  wire _16830_;
  wire _16831_;
  wire _16832_;
  wire _16833_;
  wire _16834_;
  wire _16835_;
  wire _16836_;
  wire _16837_;
  wire _16838_;
  wire _16839_;
  wire _16840_;
  wire _16841_;
  wire _16842_;
  wire _16843_;
  wire _16844_;
  wire _16845_;
  wire _16846_;
  wire _16847_;
  wire _16848_;
  wire _16849_;
  wire _16850_;
  wire _16851_;
  wire _16852_;
  wire _16853_;
  wire _16854_;
  wire _16855_;
  wire _16856_;
  wire _16857_;
  wire _16858_;
  wire _16859_;
  wire _16860_;
  wire _16861_;
  wire _16862_;
  wire _16863_;
  wire _16864_;
  wire _16865_;
  wire _16866_;
  wire _16867_;
  wire _16868_;
  wire _16869_;
  wire _16870_;
  wire _16871_;
  wire _16872_;
  wire _16873_;
  wire _16874_;
  wire _16875_;
  wire _16876_;
  wire _16877_;
  wire _16878_;
  wire _16879_;
  wire _16880_;
  wire _16881_;
  wire _16882_;
  wire _16883_;
  wire _16884_;
  wire _16885_;
  wire _16886_;
  wire _16887_;
  wire _16888_;
  wire _16889_;
  wire _16890_;
  wire _16891_;
  wire _16892_;
  wire _16893_;
  wire _16894_;
  wire _16895_;
  wire _16896_;
  wire _16897_;
  wire _16898_;
  wire _16899_;
  wire _16900_;
  wire _16901_;
  wire _16902_;
  wire _16903_;
  wire _16904_;
  wire _16905_;
  wire _16906_;
  wire _16907_;
  wire _16908_;
  wire _16909_;
  wire _16910_;
  wire _16911_;
  wire _16912_;
  wire _16913_;
  wire _16914_;
  wire _16915_;
  wire _16916_;
  wire _16917_;
  wire _16918_;
  wire _16919_;
  wire _16920_;
  wire _16921_;
  wire _16922_;
  wire _16923_;
  wire _16924_;
  wire _16925_;
  wire _16926_;
  wire _16927_;
  wire _16928_;
  wire _16929_;
  wire _16930_;
  wire _16931_;
  wire _16932_;
  wire _16933_;
  wire _16934_;
  wire _16935_;
  wire _16936_;
  wire _16937_;
  wire _16938_;
  wire _16939_;
  wire _16940_;
  wire _16941_;
  wire _16942_;
  wire _16943_;
  wire _16944_;
  wire _16945_;
  wire _16946_;
  wire _16947_;
  wire _16948_;
  wire _16949_;
  wire _16950_;
  wire _16951_;
  wire _16952_;
  wire _16953_;
  wire _16954_;
  wire _16955_;
  wire _16956_;
  wire _16957_;
  wire _16958_;
  wire _16959_;
  wire _16960_;
  wire _16961_;
  wire _16962_;
  wire _16963_;
  wire _16964_;
  wire _16965_;
  wire _16966_;
  wire _16967_;
  wire _16968_;
  wire _16969_;
  wire _16970_;
  wire _16971_;
  wire _16972_;
  wire _16973_;
  wire _16974_;
  wire _16975_;
  wire _16976_;
  wire _16977_;
  wire _16978_;
  wire _16979_;
  wire _16980_;
  wire _16981_;
  wire _16982_;
  wire _16983_;
  wire _16984_;
  wire _16985_;
  wire _16986_;
  wire _16987_;
  wire _16988_;
  wire _16989_;
  wire _16990_;
  wire _16991_;
  wire _16992_;
  wire _16993_;
  wire _16994_;
  wire _16995_;
  wire _16996_;
  wire _16997_;
  wire _16998_;
  wire _16999_;
  wire _17000_;
  wire _17001_;
  wire _17002_;
  wire _17003_;
  wire _17004_;
  wire _17005_;
  wire _17006_;
  wire _17007_;
  wire _17008_;
  wire _17009_;
  wire _17010_;
  wire _17011_;
  wire _17012_;
  wire _17013_;
  wire _17014_;
  wire _17015_;
  wire _17016_;
  wire _17017_;
  wire _17018_;
  wire _17019_;
  wire _17020_;
  wire _17021_;
  wire _17022_;
  wire _17023_;
  wire _17024_;
  wire _17025_;
  wire _17026_;
  wire _17027_;
  wire _17028_;
  wire _17029_;
  wire _17030_;
  wire _17031_;
  wire _17032_;
  wire _17033_;
  wire _17034_;
  wire _17035_;
  wire _17036_;
  wire _17037_;
  wire _17038_;
  wire _17039_;
  wire _17040_;
  wire _17041_;
  wire _17042_;
  wire _17043_;
  wire _17044_;
  wire _17045_;
  wire _17046_;
  wire _17047_;
  wire _17048_;
  wire _17049_;
  wire _17050_;
  wire _17051_;
  wire _17052_;
  wire _17053_;
  wire _17054_;
  wire _17055_;
  wire _17056_;
  wire _17057_;
  wire _17058_;
  wire _17059_;
  wire _17060_;
  wire _17061_;
  wire _17062_;
  wire _17063_;
  wire _17064_;
  wire _17065_;
  wire _17066_;
  wire _17067_;
  wire _17068_;
  wire _17069_;
  wire _17070_;
  wire _17071_;
  wire _17072_;
  wire _17073_;
  wire _17074_;
  wire _17075_;
  wire _17076_;
  wire _17077_;
  wire _17078_;
  wire _17079_;
  wire _17080_;
  wire _17081_;
  wire _17082_;
  wire _17083_;
  wire _17084_;
  wire _17085_;
  wire _17086_;
  wire _17087_;
  wire _17088_;
  wire _17089_;
  wire _17090_;
  wire _17091_;
  wire _17092_;
  wire _17093_;
  wire _17094_;
  wire _17095_;
  wire _17096_;
  wire _17097_;
  wire _17098_;
  wire _17099_;
  wire _17100_;
  wire _17101_;
  wire _17102_;
  wire _17103_;
  wire _17104_;
  wire _17105_;
  wire _17106_;
  wire _17107_;
  wire _17108_;
  wire _17109_;
  wire _17110_;
  wire _17111_;
  wire _17112_;
  wire _17113_;
  wire _17114_;
  wire _17115_;
  wire _17116_;
  wire _17117_;
  wire _17118_;
  wire _17119_;
  wire _17120_;
  wire _17121_;
  wire _17122_;
  wire _17123_;
  wire _17124_;
  wire _17125_;
  wire _17126_;
  wire _17127_;
  wire _17128_;
  wire _17129_;
  wire _17130_;
  wire _17131_;
  wire _17132_;
  wire _17133_;
  wire _17134_;
  wire _17135_;
  wire _17136_;
  wire _17137_;
  wire _17138_;
  wire _17139_;
  wire _17140_;
  wire _17141_;
  wire _17142_;
  wire _17143_;
  wire _17144_;
  wire _17145_;
  wire _17146_;
  wire _17147_;
  wire _17148_;
  wire _17149_;
  wire _17150_;
  wire _17151_;
  wire _17152_;
  wire _17153_;
  wire _17154_;
  wire _17155_;
  wire _17156_;
  wire _17157_;
  wire _17158_;
  wire _17159_;
  wire _17160_;
  wire _17161_;
  wire _17162_;
  wire _17163_;
  wire _17164_;
  wire _17165_;
  wire _17166_;
  wire _17167_;
  wire _17168_;
  wire _17169_;
  wire _17170_;
  wire _17171_;
  wire _17172_;
  wire _17173_;
  wire _17174_;
  wire _17175_;
  wire _17176_;
  wire _17177_;
  wire _17178_;
  wire _17179_;
  wire _17180_;
  wire _17181_;
  wire _17182_;
  wire _17183_;
  wire _17184_;
  wire _17185_;
  wire _17186_;
  wire _17187_;
  wire _17188_;
  wire _17189_;
  wire _17190_;
  wire _17191_;
  wire _17192_;
  wire _17193_;
  wire _17194_;
  wire _17195_;
  wire _17196_;
  wire _17197_;
  wire _17198_;
  wire _17199_;
  wire _17200_;
  wire _17201_;
  wire _17202_;
  wire _17203_;
  wire _17204_;
  wire _17205_;
  wire _17206_;
  wire _17207_;
  wire _17208_;
  wire _17209_;
  wire _17210_;
  wire _17211_;
  wire _17212_;
  wire _17213_;
  wire _17214_;
  wire _17215_;
  wire _17216_;
  wire _17217_;
  wire _17218_;
  wire _17219_;
  wire _17220_;
  wire _17221_;
  wire _17222_;
  wire _17223_;
  wire _17224_;
  wire _17225_;
  wire _17226_;
  wire _17227_;
  wire _17228_;
  wire _17229_;
  wire _17230_;
  wire _17231_;
  wire _17232_;
  wire _17233_;
  wire _17234_;
  wire _17235_;
  wire _17236_;
  wire _17237_;
  wire _17238_;
  wire _17239_;
  wire _17240_;
  wire _17241_;
  wire _17242_;
  wire _17243_;
  wire _17244_;
  wire _17245_;
  wire _17246_;
  wire _17247_;
  wire _17248_;
  wire _17249_;
  wire _17250_;
  wire _17251_;
  wire _17252_;
  wire _17253_;
  wire _17254_;
  wire _17255_;
  wire _17256_;
  wire _17257_;
  wire _17258_;
  wire _17259_;
  wire _17260_;
  wire _17261_;
  wire _17262_;
  wire _17263_;
  wire _17264_;
  wire _17265_;
  wire _17266_;
  wire _17267_;
  wire _17268_;
  wire _17269_;
  wire _17270_;
  wire _17271_;
  wire _17272_;
  wire _17273_;
  wire _17274_;
  wire _17275_;
  wire _17276_;
  wire _17277_;
  wire _17278_;
  wire _17279_;
  wire _17280_;
  wire _17281_;
  wire _17282_;
  wire _17283_;
  wire _17284_;
  wire _17285_;
  wire _17286_;
  wire _17287_;
  wire _17288_;
  wire _17289_;
  wire _17290_;
  wire _17291_;
  wire _17292_;
  wire _17293_;
  wire _17294_;
  wire _17295_;
  wire _17296_;
  wire _17297_;
  wire _17298_;
  wire _17299_;
  wire _17300_;
  wire _17301_;
  wire _17302_;
  wire _17303_;
  wire _17304_;
  wire _17305_;
  wire _17306_;
  wire _17307_;
  wire _17308_;
  wire _17309_;
  wire _17310_;
  wire _17311_;
  wire _17312_;
  wire _17313_;
  wire _17314_;
  wire _17315_;
  wire _17316_;
  wire _17317_;
  wire _17318_;
  wire _17319_;
  wire _17320_;
  wire _17321_;
  wire _17322_;
  wire _17323_;
  wire _17324_;
  wire _17325_;
  wire _17326_;
  wire _17327_;
  wire _17328_;
  wire _17329_;
  wire _17330_;
  wire _17331_;
  wire _17332_;
  wire _17333_;
  wire _17334_;
  wire _17335_;
  wire _17336_;
  wire _17337_;
  wire _17338_;
  wire _17339_;
  wire _17340_;
  wire _17341_;
  wire _17342_;
  wire _17343_;
  wire _17344_;
  wire _17345_;
  wire _17346_;
  wire _17347_;
  wire _17348_;
  wire _17349_;
  wire _17350_;
  wire _17351_;
  wire _17352_;
  wire _17353_;
  wire _17354_;
  wire _17355_;
  wire _17356_;
  wire _17357_;
  wire _17358_;
  wire _17359_;
  wire _17360_;
  wire _17361_;
  wire _17362_;
  wire _17363_;
  wire _17364_;
  wire _17365_;
  wire _17366_;
  wire _17367_;
  wire _17368_;
  wire _17369_;
  wire _17370_;
  wire _17371_;
  wire _17372_;
  wire _17373_;
  wire _17374_;
  wire _17375_;
  wire _17376_;
  wire _17377_;
  wire _17378_;
  wire _17379_;
  wire _17380_;
  wire _17381_;
  wire _17382_;
  wire _17383_;
  wire _17384_;
  wire _17385_;
  wire _17386_;
  wire _17387_;
  wire _17388_;
  wire _17389_;
  wire _17390_;
  wire _17391_;
  wire _17392_;
  wire _17393_;
  wire _17394_;
  wire _17395_;
  wire _17396_;
  wire _17397_;
  wire _17398_;
  wire _17399_;
  wire _17400_;
  wire _17401_;
  wire _17402_;
  wire _17403_;
  wire _17404_;
  wire _17405_;
  wire _17406_;
  wire _17407_;
  wire _17408_;
  wire _17409_;
  wire _17410_;
  wire _17411_;
  wire _17412_;
  wire _17413_;
  wire _17414_;
  wire _17415_;
  wire _17416_;
  wire _17417_;
  wire _17418_;
  wire _17419_;
  wire _17420_;
  wire _17421_;
  wire _17422_;
  wire _17423_;
  wire _17424_;
  wire _17425_;
  wire _17426_;
  wire _17427_;
  wire _17428_;
  wire _17429_;
  wire _17430_;
  wire _17431_;
  wire _17432_;
  wire _17433_;
  wire _17434_;
  wire _17435_;
  wire _17436_;
  wire _17437_;
  wire _17438_;
  wire _17439_;
  wire _17440_;
  wire _17441_;
  wire _17442_;
  wire _17443_;
  wire _17444_;
  wire _17445_;
  wire _17446_;
  wire _17447_;
  wire _17448_;
  wire _17449_;
  wire _17450_;
  wire _17451_;
  wire _17452_;
  wire _17453_;
  wire _17454_;
  wire _17455_;
  wire _17456_;
  wire _17457_;
  wire _17458_;
  wire _17459_;
  wire _17460_;
  wire _17461_;
  wire _17462_;
  wire _17463_;
  wire _17464_;
  wire _17465_;
  wire _17466_;
  wire _17467_;
  wire _17468_;
  wire _17469_;
  wire _17470_;
  wire _17471_;
  wire _17472_;
  wire _17473_;
  wire _17474_;
  wire _17475_;
  wire _17476_;
  wire _17477_;
  wire _17478_;
  wire _17479_;
  wire _17480_;
  wire _17481_;
  wire _17482_;
  wire _17483_;
  wire _17484_;
  wire _17485_;
  wire _17486_;
  wire _17487_;
  wire _17488_;
  wire _17489_;
  wire _17490_;
  wire _17491_;
  wire _17492_;
  wire _17493_;
  wire _17494_;
  wire _17495_;
  wire _17496_;
  wire _17497_;
  wire _17498_;
  wire _17499_;
  wire _17500_;
  wire _17501_;
  wire _17502_;
  wire _17503_;
  wire _17504_;
  wire _17505_;
  wire _17506_;
  wire _17507_;
  wire _17508_;
  wire _17509_;
  wire _17510_;
  wire _17511_;
  wire _17512_;
  wire _17513_;
  wire _17514_;
  wire _17515_;
  wire _17516_;
  wire _17517_;
  wire _17518_;
  wire _17519_;
  wire _17520_;
  wire _17521_;
  wire _17522_;
  wire _17523_;
  wire _17524_;
  wire _17525_;
  wire _17526_;
  wire _17527_;
  wire _17528_;
  wire _17529_;
  wire _17530_;
  wire _17531_;
  wire _17532_;
  wire _17533_;
  wire _17534_;
  wire _17535_;
  wire _17536_;
  wire _17537_;
  wire _17538_;
  wire _17539_;
  wire _17540_;
  wire _17541_;
  wire _17542_;
  wire _17543_;
  wire _17544_;
  wire _17545_;
  wire _17546_;
  wire _17547_;
  wire _17548_;
  wire _17549_;
  wire _17550_;
  wire _17551_;
  wire _17552_;
  wire _17553_;
  wire _17554_;
  wire _17555_;
  wire _17556_;
  wire _17557_;
  wire _17558_;
  wire _17559_;
  wire _17560_;
  wire _17561_;
  wire _17562_;
  wire _17563_;
  wire _17564_;
  wire _17565_;
  wire _17566_;
  wire _17567_;
  wire _17568_;
  wire _17569_;
  wire _17570_;
  wire _17571_;
  wire _17572_;
  wire _17573_;
  wire _17574_;
  wire _17575_;
  wire _17576_;
  wire _17577_;
  wire _17578_;
  wire _17579_;
  wire _17580_;
  wire _17581_;
  wire _17582_;
  wire _17583_;
  wire _17584_;
  wire _17585_;
  wire _17586_;
  wire _17587_;
  wire _17588_;
  wire _17589_;
  wire _17590_;
  wire _17591_;
  wire _17592_;
  wire _17593_;
  wire _17594_;
  wire _17595_;
  wire _17596_;
  wire _17597_;
  wire _17598_;
  wire _17599_;
  wire _17600_;
  wire _17601_;
  wire _17602_;
  wire _17603_;
  wire _17604_;
  wire _17605_;
  wire _17606_;
  wire _17607_;
  wire _17608_;
  wire _17609_;
  wire _17610_;
  wire _17611_;
  wire _17612_;
  wire _17613_;
  wire _17614_;
  wire _17615_;
  wire _17616_;
  wire _17617_;
  wire _17618_;
  wire _17619_;
  wire _17620_;
  wire _17621_;
  wire _17622_;
  wire _17623_;
  wire _17624_;
  wire _17625_;
  wire _17626_;
  wire _17627_;
  wire _17628_;
  wire _17629_;
  wire _17630_;
  wire _17631_;
  wire _17632_;
  wire _17633_;
  wire _17634_;
  wire _17635_;
  wire _17636_;
  wire _17637_;
  wire _17638_;
  wire _17639_;
  wire _17640_;
  wire _17641_;
  wire _17642_;
  wire _17643_;
  wire _17644_;
  wire _17645_;
  wire _17646_;
  wire _17647_;
  wire _17648_;
  wire _17649_;
  wire _17650_;
  wire _17651_;
  wire _17652_;
  wire _17653_;
  wire _17654_;
  wire _17655_;
  wire _17656_;
  wire _17657_;
  wire _17658_;
  wire _17659_;
  wire _17660_;
  wire _17661_;
  wire _17662_;
  wire _17663_;
  wire _17664_;
  wire _17665_;
  wire _17666_;
  wire _17667_;
  wire _17668_;
  wire _17669_;
  wire _17670_;
  wire _17671_;
  wire _17672_;
  wire _17673_;
  wire _17674_;
  wire _17675_;
  wire _17676_;
  wire _17677_;
  wire _17678_;
  wire _17679_;
  wire _17680_;
  wire _17681_;
  wire _17682_;
  wire _17683_;
  wire _17684_;
  wire _17685_;
  wire _17686_;
  wire _17687_;
  wire _17688_;
  wire _17689_;
  wire _17690_;
  wire _17691_;
  wire _17692_;
  wire _17693_;
  wire _17694_;
  wire _17695_;
  wire _17696_;
  wire _17697_;
  wire _17698_;
  wire _17699_;
  wire _17700_;
  wire _17701_;
  wire _17702_;
  wire _17703_;
  wire _17704_;
  wire _17705_;
  wire _17706_;
  wire _17707_;
  wire _17708_;
  wire _17709_;
  wire _17710_;
  wire _17711_;
  wire _17712_;
  wire _17713_;
  wire _17714_;
  wire _17715_;
  wire _17716_;
  wire _17717_;
  wire _17718_;
  wire _17719_;
  wire _17720_;
  wire _17721_;
  wire _17722_;
  wire _17723_;
  wire _17724_;
  wire _17725_;
  wire _17726_;
  wire _17727_;
  wire _17728_;
  wire _17729_;
  wire _17730_;
  wire _17731_;
  wire _17732_;
  wire _17733_;
  wire _17734_;
  wire _17735_;
  wire _17736_;
  wire _17737_;
  wire _17738_;
  wire _17739_;
  wire _17740_;
  wire _17741_;
  wire _17742_;
  wire _17743_;
  wire _17744_;
  wire _17745_;
  wire _17746_;
  wire _17747_;
  wire _17748_;
  wire _17749_;
  wire _17750_;
  wire _17751_;
  wire _17752_;
  wire _17753_;
  wire _17754_;
  wire _17755_;
  wire _17756_;
  wire _17757_;
  wire _17758_;
  wire _17759_;
  wire _17760_;
  wire _17761_;
  wire _17762_;
  wire _17763_;
  wire _17764_;
  wire _17765_;
  wire _17766_;
  wire _17767_;
  wire _17768_;
  wire _17769_;
  wire _17770_;
  wire _17771_;
  wire _17772_;
  wire _17773_;
  wire _17774_;
  wire _17775_;
  wire _17776_;
  wire _17777_;
  wire _17778_;
  wire _17779_;
  wire _17780_;
  wire _17781_;
  wire _17782_;
  wire _17783_;
  wire _17784_;
  wire _17785_;
  wire _17786_;
  wire _17787_;
  wire _17788_;
  wire _17789_;
  wire _17790_;
  wire _17791_;
  wire _17792_;
  wire _17793_;
  wire _17794_;
  wire _17795_;
  wire _17796_;
  wire _17797_;
  wire _17798_;
  wire _17799_;
  wire _17800_;
  wire _17801_;
  wire _17802_;
  wire _17803_;
  wire _17804_;
  wire _17805_;
  wire _17806_;
  wire _17807_;
  wire _17808_;
  wire _17809_;
  wire _17810_;
  wire _17811_;
  wire _17812_;
  wire _17813_;
  wire _17814_;
  wire _17815_;
  wire _17816_;
  wire _17817_;
  wire _17818_;
  wire _17819_;
  wire _17820_;
  wire _17821_;
  wire _17822_;
  wire _17823_;
  wire _17824_;
  wire _17825_;
  wire _17826_;
  wire _17827_;
  wire _17828_;
  wire _17829_;
  wire _17830_;
  wire _17831_;
  wire _17832_;
  wire _17833_;
  wire _17834_;
  wire _17835_;
  wire _17836_;
  wire _17837_;
  wire _17838_;
  wire _17839_;
  wire _17840_;
  wire _17841_;
  wire _17842_;
  wire _17843_;
  wire _17844_;
  wire _17845_;
  wire _17846_;
  wire _17847_;
  wire _17848_;
  wire _17849_;
  wire _17850_;
  wire _17851_;
  wire _17852_;
  wire _17853_;
  wire _17854_;
  wire _17855_;
  wire _17856_;
  wire _17857_;
  wire _17858_;
  wire _17859_;
  wire _17860_;
  wire _17861_;
  wire _17862_;
  wire _17863_;
  wire _17864_;
  wire _17865_;
  wire _17866_;
  wire _17867_;
  wire _17868_;
  wire _17869_;
  wire _17870_;
  wire _17871_;
  wire _17872_;
  wire _17873_;
  wire _17874_;
  wire _17875_;
  wire _17876_;
  wire _17877_;
  wire _17878_;
  wire _17879_;
  wire _17880_;
  wire _17881_;
  wire _17882_;
  wire _17883_;
  wire _17884_;
  wire _17885_;
  wire _17886_;
  wire _17887_;
  wire _17888_;
  wire _17889_;
  wire _17890_;
  wire _17891_;
  wire _17892_;
  wire _17893_;
  wire _17894_;
  wire _17895_;
  wire _17896_;
  wire _17897_;
  wire _17898_;
  wire _17899_;
  wire _17900_;
  wire _17901_;
  wire _17902_;
  wire _17903_;
  wire _17904_;
  wire _17905_;
  wire _17906_;
  wire _17907_;
  wire _17908_;
  wire _17909_;
  wire _17910_;
  wire _17911_;
  wire _17912_;
  wire _17913_;
  wire _17914_;
  wire _17915_;
  wire _17916_;
  wire _17917_;
  wire _17918_;
  wire _17919_;
  wire _17920_;
  wire _17921_;
  wire _17922_;
  wire _17923_;
  wire _17924_;
  wire _17925_;
  wire _17926_;
  wire _17927_;
  wire _17928_;
  wire _17929_;
  wire _17930_;
  wire _17931_;
  wire _17932_;
  wire _17933_;
  wire _17934_;
  wire _17935_;
  wire _17936_;
  wire _17937_;
  wire _17938_;
  wire _17939_;
  wire _17940_;
  wire _17941_;
  wire _17942_;
  wire _17943_;
  wire _17944_;
  wire _17945_;
  wire _17946_;
  wire _17947_;
  wire _17948_;
  wire _17949_;
  wire _17950_;
  wire _17951_;
  wire _17952_;
  wire _17953_;
  wire _17954_;
  wire _17955_;
  wire _17956_;
  wire _17957_;
  wire _17958_;
  wire _17959_;
  wire _17960_;
  wire _17961_;
  wire _17962_;
  wire _17963_;
  wire _17964_;
  wire _17965_;
  wire _17966_;
  wire _17967_;
  wire _17968_;
  wire _17969_;
  wire _17970_;
  wire _17971_;
  wire _17972_;
  wire _17973_;
  wire _17974_;
  wire _17975_;
  wire _17976_;
  wire _17977_;
  wire _17978_;
  wire _17979_;
  wire _17980_;
  wire _17981_;
  wire _17982_;
  wire _17983_;
  wire _17984_;
  wire _17985_;
  wire _17986_;
  wire _17987_;
  wire _17988_;
  wire _17989_;
  wire _17990_;
  wire _17991_;
  wire _17992_;
  wire _17993_;
  wire _17994_;
  wire _17995_;
  wire _17996_;
  wire _17997_;
  wire _17998_;
  wire _17999_;
  wire _18000_;
  wire _18001_;
  wire _18002_;
  wire _18003_;
  wire _18004_;
  wire _18005_;
  wire _18006_;
  wire _18007_;
  wire _18008_;
  wire _18009_;
  wire _18010_;
  wire _18011_;
  wire _18012_;
  wire _18013_;
  wire _18014_;
  wire _18015_;
  wire _18016_;
  wire _18017_;
  wire _18018_;
  wire _18019_;
  wire _18020_;
  wire _18021_;
  wire _18022_;
  wire _18023_;
  wire _18024_;
  wire _18025_;
  wire _18026_;
  wire _18027_;
  wire _18028_;
  wire _18029_;
  wire _18030_;
  wire _18031_;
  wire _18032_;
  wire _18033_;
  wire _18034_;
  wire _18035_;
  wire _18036_;
  wire _18037_;
  wire _18038_;
  wire _18039_;
  wire _18040_;
  wire _18041_;
  wire _18042_;
  wire _18043_;
  wire _18044_;
  wire _18045_;
  wire _18046_;
  wire _18047_;
  wire _18048_;
  wire _18049_;
  wire _18050_;
  wire _18051_;
  wire _18052_;
  wire _18053_;
  wire _18054_;
  wire _18055_;
  wire _18056_;
  wire _18057_;
  wire _18058_;
  wire _18059_;
  wire _18060_;
  wire _18061_;
  wire _18062_;
  wire _18063_;
  wire _18064_;
  wire _18065_;
  wire _18066_;
  wire _18067_;
  wire _18068_;
  wire _18069_;
  wire _18070_;
  wire _18071_;
  wire _18072_;
  wire _18073_;
  wire _18074_;
  wire _18075_;
  wire _18076_;
  wire _18077_;
  wire _18078_;
  wire _18079_;
  wire _18080_;
  wire _18081_;
  wire _18082_;
  wire _18083_;
  wire _18084_;
  wire _18085_;
  wire _18086_;
  wire _18087_;
  wire _18088_;
  wire _18089_;
  wire _18090_;
  wire _18091_;
  wire _18092_;
  wire _18093_;
  wire _18094_;
  wire _18095_;
  wire _18096_;
  wire _18097_;
  wire _18098_;
  wire _18099_;
  wire _18100_;
  wire _18101_;
  wire _18102_;
  wire _18103_;
  wire _18104_;
  wire _18105_;
  wire _18106_;
  wire _18107_;
  wire _18108_;
  wire _18109_;
  wire _18110_;
  wire _18111_;
  wire _18112_;
  wire _18113_;
  wire _18114_;
  wire _18115_;
  wire _18116_;
  wire _18117_;
  wire _18118_;
  wire _18119_;
  wire _18120_;
  wire _18121_;
  wire _18122_;
  wire _18123_;
  wire _18124_;
  wire _18125_;
  wire _18126_;
  wire _18127_;
  wire _18128_;
  wire _18129_;
  wire _18130_;
  wire _18131_;
  wire _18132_;
  wire _18133_;
  wire _18134_;
  wire _18135_;
  wire _18136_;
  wire _18137_;
  wire _18138_;
  wire _18139_;
  wire _18140_;
  wire _18141_;
  wire _18142_;
  wire _18143_;
  wire _18144_;
  wire _18145_;
  wire _18146_;
  wire _18147_;
  wire _18148_;
  wire _18149_;
  wire _18150_;
  wire _18151_;
  wire _18152_;
  wire _18153_;
  wire _18154_;
  wire _18155_;
  wire _18156_;
  wire _18157_;
  wire _18158_;
  wire _18159_;
  wire _18160_;
  wire _18161_;
  wire _18162_;
  wire _18163_;
  wire _18164_;
  wire _18165_;
  wire _18166_;
  wire _18167_;
  wire _18168_;
  wire _18169_;
  wire _18170_;
  wire _18171_;
  wire _18172_;
  wire _18173_;
  wire _18174_;
  wire _18175_;
  wire _18176_;
  wire _18177_;
  wire _18178_;
  wire _18179_;
  wire _18180_;
  wire _18181_;
  wire _18182_;
  wire _18183_;
  wire _18184_;
  wire _18185_;
  wire _18186_;
  wire _18187_;
  wire _18188_;
  wire _18189_;
  wire _18190_;
  wire _18191_;
  wire _18192_;
  wire _18193_;
  wire _18194_;
  wire _18195_;
  wire _18196_;
  wire _18197_;
  wire _18198_;
  wire _18199_;
  wire _18200_;
  wire _18201_;
  wire _18202_;
  wire _18203_;
  wire _18204_;
  wire _18205_;
  wire _18206_;
  wire _18207_;
  wire _18208_;
  wire _18209_;
  wire _18210_;
  wire _18211_;
  wire _18212_;
  wire _18213_;
  wire _18214_;
  wire _18215_;
  wire _18216_;
  wire _18217_;
  wire _18218_;
  wire _18219_;
  wire _18220_;
  wire _18221_;
  wire _18222_;
  wire _18223_;
  wire _18224_;
  wire _18225_;
  wire _18226_;
  wire _18227_;
  wire _18228_;
  wire _18229_;
  wire _18230_;
  wire _18231_;
  wire _18232_;
  wire _18233_;
  wire _18234_;
  wire _18235_;
  wire _18236_;
  wire _18237_;
  wire _18238_;
  wire _18239_;
  wire _18240_;
  wire _18241_;
  wire _18242_;
  wire _18243_;
  wire _18244_;
  wire _18245_;
  wire _18246_;
  wire _18247_;
  wire _18248_;
  wire _18249_;
  wire _18250_;
  wire _18251_;
  wire _18252_;
  wire _18253_;
  wire _18254_;
  wire _18255_;
  wire _18256_;
  wire _18257_;
  wire _18258_;
  wire _18259_;
  wire _18260_;
  wire _18261_;
  wire _18262_;
  wire _18263_;
  wire _18264_;
  wire _18265_;
  wire _18266_;
  wire _18267_;
  wire _18268_;
  wire _18269_;
  wire _18270_;
  wire _18271_;
  wire _18272_;
  wire _18273_;
  wire _18274_;
  wire _18275_;
  wire _18276_;
  wire _18277_;
  wire _18278_;
  wire _18279_;
  wire _18280_;
  wire _18281_;
  wire _18282_;
  wire _18283_;
  wire _18284_;
  wire _18285_;
  wire _18286_;
  wire _18287_;
  wire _18288_;
  wire _18289_;
  wire _18290_;
  wire _18291_;
  wire _18292_;
  wire _18293_;
  wire _18294_;
  wire _18295_;
  wire _18296_;
  wire _18297_;
  wire _18298_;
  wire _18299_;
  wire _18300_;
  wire _18301_;
  wire _18302_;
  wire _18303_;
  wire _18304_;
  wire _18305_;
  wire _18306_;
  wire _18307_;
  wire _18308_;
  wire _18309_;
  wire _18310_;
  wire _18311_;
  wire _18312_;
  wire _18313_;
  wire _18314_;
  wire _18315_;
  wire _18316_;
  wire _18317_;
  wire _18318_;
  wire _18319_;
  wire _18320_;
  wire _18321_;
  wire _18322_;
  wire _18323_;
  wire _18324_;
  wire _18325_;
  wire _18326_;
  wire _18327_;
  wire _18328_;
  wire _18329_;
  wire _18330_;
  wire _18331_;
  wire _18332_;
  wire _18333_;
  wire _18334_;
  wire _18335_;
  wire _18336_;
  wire _18337_;
  wire _18338_;
  wire _18339_;
  wire _18340_;
  wire _18341_;
  wire _18342_;
  wire _18343_;
  wire _18344_;
  wire _18345_;
  wire _18346_;
  wire _18347_;
  wire _18348_;
  wire _18349_;
  wire _18350_;
  wire _18351_;
  wire _18352_;
  wire _18353_;
  wire _18354_;
  wire _18355_;
  wire _18356_;
  wire _18357_;
  wire _18358_;
  wire _18359_;
  wire _18360_;
  wire _18361_;
  wire _18362_;
  wire _18363_;
  wire _18364_;
  wire _18365_;
  wire _18366_;
  wire _18367_;
  wire _18368_;
  wire _18369_;
  wire _18370_;
  wire _18371_;
  wire _18372_;
  wire _18373_;
  wire _18374_;
  wire _18375_;
  wire _18376_;
  wire _18377_;
  wire _18378_;
  wire _18379_;
  wire _18380_;
  wire _18381_;
  wire _18382_;
  wire _18383_;
  wire _18384_;
  wire _18385_;
  wire _18386_;
  wire _18387_;
  wire _18388_;
  wire _18389_;
  wire _18390_;
  wire _18391_;
  wire _18392_;
  wire _18393_;
  wire _18394_;
  wire _18395_;
  wire _18396_;
  wire _18397_;
  wire _18398_;
  wire _18399_;
  wire _18400_;
  wire _18401_;
  wire _18402_;
  wire _18403_;
  wire _18404_;
  wire _18405_;
  wire _18406_;
  wire _18407_;
  wire _18408_;
  wire _18409_;
  wire _18410_;
  wire _18411_;
  wire _18412_;
  wire _18413_;
  wire _18414_;
  wire _18415_;
  wire _18416_;
  wire _18417_;
  wire _18418_;
  wire _18419_;
  wire _18420_;
  wire _18421_;
  wire _18422_;
  wire _18423_;
  wire _18424_;
  wire _18425_;
  wire _18426_;
  wire _18427_;
  wire _18428_;
  wire _18429_;
  wire _18430_;
  wire _18431_;
  wire _18432_;
  wire _18433_;
  wire _18434_;
  wire _18435_;
  wire _18436_;
  wire _18437_;
  wire _18438_;
  wire _18439_;
  wire _18440_;
  wire _18441_;
  wire _18442_;
  wire _18443_;
  wire _18444_;
  wire _18445_;
  wire _18446_;
  wire _18447_;
  wire _18448_;
  wire _18449_;
  wire _18450_;
  wire _18451_;
  wire _18452_;
  wire _18453_;
  wire _18454_;
  wire _18455_;
  wire _18456_;
  wire _18457_;
  wire _18458_;
  wire _18459_;
  wire _18460_;
  wire _18461_;
  wire _18462_;
  wire _18463_;
  wire _18464_;
  wire _18465_;
  wire _18466_;
  wire _18467_;
  wire _18468_;
  wire _18469_;
  wire _18470_;
  wire _18471_;
  wire _18472_;
  wire _18473_;
  wire _18474_;
  wire _18475_;
  wire _18476_;
  wire _18477_;
  wire _18478_;
  wire _18479_;
  wire _18480_;
  wire _18481_;
  wire _18482_;
  wire _18483_;
  wire _18484_;
  wire _18485_;
  wire _18486_;
  wire _18487_;
  wire _18488_;
  wire _18489_;
  wire _18490_;
  wire _18491_;
  wire _18492_;
  wire _18493_;
  wire _18494_;
  wire _18495_;
  wire _18496_;
  wire _18497_;
  wire _18498_;
  wire _18499_;
  wire _18500_;
  wire _18501_;
  wire _18502_;
  wire _18503_;
  wire _18504_;
  wire _18505_;
  wire _18506_;
  wire _18507_;
  wire _18508_;
  wire _18509_;
  wire _18510_;
  wire _18511_;
  wire _18512_;
  wire _18513_;
  wire _18514_;
  wire _18515_;
  wire _18516_;
  wire _18517_;
  wire _18518_;
  wire _18519_;
  wire _18520_;
  wire _18521_;
  wire _18522_;
  wire _18523_;
  wire _18524_;
  wire _18525_;
  wire _18526_;
  wire _18527_;
  wire _18528_;
  wire _18529_;
  wire _18530_;
  wire _18531_;
  wire _18532_;
  wire _18533_;
  wire _18534_;
  wire _18535_;
  wire _18536_;
  wire _18537_;
  wire _18538_;
  wire _18539_;
  wire _18540_;
  wire _18541_;
  wire _18542_;
  wire _18543_;
  wire _18544_;
  wire _18545_;
  wire _18546_;
  wire _18547_;
  wire _18548_;
  wire _18549_;
  wire _18550_;
  wire _18551_;
  wire _18552_;
  wire _18553_;
  wire _18554_;
  wire _18555_;
  wire _18556_;
  wire _18557_;
  wire _18558_;
  wire _18559_;
  wire _18560_;
  wire _18561_;
  wire _18562_;
  wire _18563_;
  wire _18564_;
  wire _18565_;
  wire _18566_;
  wire _18567_;
  wire _18568_;
  wire _18569_;
  wire _18570_;
  wire _18571_;
  wire _18572_;
  wire _18573_;
  wire _18574_;
  wire _18575_;
  wire _18576_;
  wire _18577_;
  wire _18578_;
  wire _18579_;
  wire _18580_;
  wire _18581_;
  wire _18582_;
  wire _18583_;
  wire _18584_;
  wire _18585_;
  wire _18586_;
  wire _18587_;
  wire _18588_;
  wire _18589_;
  wire _18590_;
  wire _18591_;
  wire _18592_;
  wire _18593_;
  wire _18594_;
  wire _18595_;
  wire _18596_;
  wire _18597_;
  wire _18598_;
  wire _18599_;
  wire _18600_;
  wire _18601_;
  wire _18602_;
  wire _18603_;
  wire _18604_;
  wire _18605_;
  wire _18606_;
  wire _18607_;
  wire _18608_;
  wire _18609_;
  wire _18610_;
  wire _18611_;
  wire _18612_;
  wire _18613_;
  wire _18614_;
  wire _18615_;
  wire _18616_;
  wire _18617_;
  wire _18618_;
  wire _18619_;
  wire _18620_;
  wire _18621_;
  wire _18622_;
  wire _18623_;
  wire _18624_;
  wire _18625_;
  wire _18626_;
  wire _18627_;
  wire _18628_;
  wire _18629_;
  wire _18630_;
  wire _18631_;
  wire _18632_;
  wire _18633_;
  wire _18634_;
  wire _18635_;
  wire _18636_;
  wire _18637_;
  wire _18638_;
  wire _18639_;
  wire _18640_;
  wire _18641_;
  wire _18642_;
  wire _18643_;
  wire _18644_;
  wire _18645_;
  wire _18646_;
  wire _18647_;
  wire _18648_;
  wire _18649_;
  wire _18650_;
  wire _18651_;
  wire _18652_;
  wire _18653_;
  wire _18654_;
  wire _18655_;
  wire _18656_;
  wire _18657_;
  wire _18658_;
  wire _18659_;
  wire _18660_;
  wire _18661_;
  wire _18662_;
  wire _18663_;
  wire _18664_;
  wire _18665_;
  wire _18666_;
  wire _18667_;
  wire _18668_;
  wire _18669_;
  wire _18670_;
  wire _18671_;
  wire _18672_;
  wire _18673_;
  wire _18674_;
  wire _18675_;
  wire _18676_;
  wire _18677_;
  wire _18678_;
  wire _18679_;
  wire _18680_;
  wire _18681_;
  wire _18682_;
  wire _18683_;
  wire _18684_;
  wire _18685_;
  wire _18686_;
  wire _18687_;
  wire _18688_;
  wire _18689_;
  wire _18690_;
  wire _18691_;
  wire _18692_;
  wire _18693_;
  wire _18694_;
  wire _18695_;
  wire _18696_;
  wire _18697_;
  wire _18698_;
  wire _18699_;
  wire _18700_;
  wire _18701_;
  wire _18702_;
  wire _18703_;
  wire _18704_;
  wire _18705_;
  wire _18706_;
  wire _18707_;
  wire _18708_;
  wire _18709_;
  wire _18710_;
  wire _18711_;
  wire _18712_;
  wire _18713_;
  wire _18714_;
  wire _18715_;
  wire _18716_;
  wire _18717_;
  wire _18718_;
  wire _18719_;
  wire _18720_;
  wire _18721_;
  wire _18722_;
  wire _18723_;
  wire _18724_;
  wire _18725_;
  wire _18726_;
  wire _18727_;
  wire _18728_;
  wire _18729_;
  wire _18730_;
  wire _18731_;
  wire _18732_;
  wire _18733_;
  wire _18734_;
  wire _18735_;
  wire _18736_;
  wire _18737_;
  wire _18738_;
  wire _18739_;
  wire _18740_;
  wire _18741_;
  wire _18742_;
  wire _18743_;
  wire _18744_;
  wire _18745_;
  wire _18746_;
  wire _18747_;
  wire _18748_;
  wire _18749_;
  wire _18750_;
  wire _18751_;
  wire _18752_;
  wire _18753_;
  wire _18754_;
  wire _18755_;
  wire _18756_;
  wire _18757_;
  wire _18758_;
  wire _18759_;
  wire _18760_;
  wire _18761_;
  wire _18762_;
  wire _18763_;
  wire _18764_;
  wire _18765_;
  wire _18766_;
  wire _18767_;
  wire _18768_;
  wire _18769_;
  wire _18770_;
  wire _18771_;
  wire _18772_;
  wire _18773_;
  wire _18774_;
  wire _18775_;
  wire _18776_;
  wire _18777_;
  wire _18778_;
  wire _18779_;
  wire _18780_;
  wire _18781_;
  wire _18782_;
  wire _18783_;
  wire _18784_;
  wire _18785_;
  wire _18786_;
  wire _18787_;
  wire _18788_;
  wire _18789_;
  wire _18790_;
  wire _18791_;
  wire _18792_;
  wire _18793_;
  wire _18794_;
  wire _18795_;
  wire _18796_;
  wire _18797_;
  wire _18798_;
  wire _18799_;
  wire _18800_;
  wire _18801_;
  wire _18802_;
  wire _18803_;
  wire _18804_;
  wire _18805_;
  wire _18806_;
  wire _18807_;
  wire _18808_;
  wire _18809_;
  wire _18810_;
  wire _18811_;
  wire _18812_;
  wire _18813_;
  wire _18814_;
  wire _18815_;
  wire _18816_;
  wire _18817_;
  wire _18818_;
  wire _18819_;
  wire _18820_;
  wire _18821_;
  wire _18822_;
  wire _18823_;
  wire _18824_;
  wire _18825_;
  wire _18826_;
  wire _18827_;
  wire _18828_;
  wire _18829_;
  wire _18830_;
  wire _18831_;
  wire _18832_;
  wire _18833_;
  wire _18834_;
  wire _18835_;
  wire _18836_;
  wire _18837_;
  wire _18838_;
  wire _18839_;
  wire _18840_;
  wire _18841_;
  wire _18842_;
  wire _18843_;
  wire _18844_;
  wire _18845_;
  wire _18846_;
  wire _18847_;
  wire _18848_;
  wire _18849_;
  wire _18850_;
  wire _18851_;
  wire _18852_;
  wire _18853_;
  wire _18854_;
  wire _18855_;
  wire _18856_;
  wire _18857_;
  wire _18858_;
  wire _18859_;
  wire _18860_;
  wire _18861_;
  wire _18862_;
  wire _18863_;
  wire _18864_;
  wire _18865_;
  wire _18866_;
  wire _18867_;
  wire _18868_;
  wire _18869_;
  wire _18870_;
  wire _18871_;
  wire _18872_;
  wire _18873_;
  wire _18874_;
  wire _18875_;
  wire _18876_;
  wire _18877_;
  wire _18878_;
  wire _18879_;
  wire _18880_;
  wire _18881_;
  wire _18882_;
  wire _18883_;
  wire _18884_;
  wire _18885_;
  wire _18886_;
  wire _18887_;
  wire _18888_;
  wire _18889_;
  wire _18890_;
  wire _18891_;
  wire _18892_;
  wire _18893_;
  wire _18894_;
  wire _18895_;
  wire _18896_;
  wire _18897_;
  wire _18898_;
  wire _18899_;
  wire _18900_;
  wire _18901_;
  wire _18902_;
  wire _18903_;
  wire _18904_;
  wire _18905_;
  wire _18906_;
  wire _18907_;
  wire _18908_;
  wire _18909_;
  wire _18910_;
  wire _18911_;
  wire _18912_;
  wire _18913_;
  wire _18914_;
  wire _18915_;
  wire _18916_;
  wire _18917_;
  wire _18918_;
  wire _18919_;
  wire _18920_;
  wire _18921_;
  wire _18922_;
  wire _18923_;
  wire _18924_;
  wire _18925_;
  wire _18926_;
  wire _18927_;
  wire _18928_;
  wire _18929_;
  wire _18930_;
  wire _18931_;
  wire _18932_;
  wire _18933_;
  wire _18934_;
  wire _18935_;
  wire _18936_;
  wire _18937_;
  wire _18938_;
  wire _18939_;
  wire _18940_;
  wire _18941_;
  wire _18942_;
  wire _18943_;
  wire _18944_;
  wire _18945_;
  wire _18946_;
  wire _18947_;
  wire _18948_;
  wire _18949_;
  wire _18950_;
  wire _18951_;
  wire _18952_;
  wire _18953_;
  wire _18954_;
  wire _18955_;
  wire _18956_;
  wire _18957_;
  wire _18958_;
  wire _18959_;
  wire _18960_;
  wire _18961_;
  wire _18962_;
  wire _18963_;
  wire _18964_;
  wire _18965_;
  wire _18966_;
  wire _18967_;
  wire _18968_;
  wire _18969_;
  wire _18970_;
  wire _18971_;
  wire _18972_;
  wire _18973_;
  wire _18974_;
  wire _18975_;
  wire _18976_;
  wire _18977_;
  wire _18978_;
  wire _18979_;
  wire _18980_;
  wire _18981_;
  wire _18982_;
  wire _18983_;
  wire _18984_;
  wire _18985_;
  wire _18986_;
  wire _18987_;
  wire _18988_;
  wire _18989_;
  wire _18990_;
  wire _18991_;
  wire _18992_;
  wire _18993_;
  wire _18994_;
  wire _18995_;
  wire _18996_;
  wire _18997_;
  wire _18998_;
  wire _18999_;
  wire _19000_;
  wire _19001_;
  wire _19002_;
  wire _19003_;
  wire _19004_;
  wire _19005_;
  wire _19006_;
  wire _19007_;
  wire _19008_;
  wire _19009_;
  wire _19010_;
  wire _19011_;
  wire _19012_;
  wire _19013_;
  wire _19014_;
  wire _19015_;
  wire _19016_;
  wire _19017_;
  wire _19018_;
  wire _19019_;
  wire _19020_;
  wire _19021_;
  wire _19022_;
  wire _19023_;
  wire _19024_;
  wire _19025_;
  wire _19026_;
  wire _19027_;
  wire _19028_;
  wire _19029_;
  wire _19030_;
  wire _19031_;
  wire _19032_;
  wire _19033_;
  wire _19034_;
  wire _19035_;
  wire _19036_;
  wire _19037_;
  wire _19038_;
  wire _19039_;
  wire _19040_;
  wire _19041_;
  wire _19042_;
  wire _19043_;
  wire _19044_;
  wire _19045_;
  wire _19046_;
  wire _19047_;
  wire _19048_;
  wire _19049_;
  wire _19050_;
  wire _19051_;
  wire _19052_;
  wire _19053_;
  wire _19054_;
  wire _19055_;
  wire _19056_;
  wire _19057_;
  wire _19058_;
  wire _19059_;
  wire _19060_;
  wire _19061_;
  wire _19062_;
  wire _19063_;
  wire _19064_;
  wire _19065_;
  wire _19066_;
  wire _19067_;
  wire _19068_;
  wire _19069_;
  wire _19070_;
  wire _19071_;
  wire _19072_;
  wire _19073_;
  wire _19074_;
  wire _19075_;
  wire _19076_;
  wire _19077_;
  wire _19078_;
  wire _19079_;
  wire _19080_;
  wire _19081_;
  wire _19082_;
  wire _19083_;
  wire _19084_;
  wire _19085_;
  wire _19086_;
  wire _19087_;
  wire _19088_;
  wire _19089_;
  wire _19090_;
  wire _19091_;
  wire _19092_;
  wire _19093_;
  wire _19094_;
  wire _19095_;
  wire _19096_;
  wire _19097_;
  wire _19098_;
  wire _19099_;
  wire _19100_;
  wire _19101_;
  wire _19102_;
  wire _19103_;
  wire _19104_;
  wire _19105_;
  wire _19106_;
  wire _19107_;
  wire _19108_;
  wire _19109_;
  wire _19110_;
  wire _19111_;
  wire _19112_;
  wire _19113_;
  wire _19114_;
  wire _19115_;
  wire _19116_;
  wire _19117_;
  wire _19118_;
  wire _19119_;
  wire _19120_;
  wire _19121_;
  wire _19122_;
  wire _19123_;
  wire _19124_;
  wire _19125_;
  wire _19126_;
  wire _19127_;
  wire _19128_;
  wire _19129_;
  wire _19130_;
  wire _19131_;
  wire _19132_;
  wire _19133_;
  wire _19134_;
  wire _19135_;
  wire _19136_;
  wire _19137_;
  wire _19138_;
  wire _19139_;
  wire _19140_;
  wire _19141_;
  wire _19142_;
  wire _19143_;
  wire _19144_;
  wire _19145_;
  wire _19146_;
  wire _19147_;
  wire _19148_;
  wire _19149_;
  wire _19150_;
  wire _19151_;
  wire _19152_;
  wire _19153_;
  wire _19154_;
  wire _19155_;
  wire _19156_;
  wire _19157_;
  wire _19158_;
  wire _19159_;
  wire _19160_;
  wire _19161_;
  wire _19162_;
  wire _19163_;
  wire _19164_;
  wire _19165_;
  wire _19166_;
  wire _19167_;
  wire _19168_;
  wire _19169_;
  wire _19170_;
  wire _19171_;
  wire _19172_;
  wire _19173_;
  wire _19174_;
  wire _19175_;
  wire _19176_;
  wire _19177_;
  wire _19178_;
  wire _19179_;
  wire _19180_;
  wire _19181_;
  wire _19182_;
  wire _19183_;
  wire _19184_;
  wire _19185_;
  wire _19186_;
  wire _19187_;
  wire _19188_;
  wire _19189_;
  wire _19190_;
  wire _19191_;
  wire _19192_;
  wire _19193_;
  wire _19194_;
  wire _19195_;
  wire _19196_;
  wire _19197_;
  wire _19198_;
  wire _19199_;
  wire _19200_;
  wire _19201_;
  wire _19202_;
  wire _19203_;
  wire _19204_;
  wire _19205_;
  wire _19206_;
  wire _19207_;
  wire _19208_;
  wire _19209_;
  wire _19210_;
  wire _19211_;
  wire _19212_;
  wire _19213_;
  wire _19214_;
  wire _19215_;
  wire _19216_;
  wire _19217_;
  wire _19218_;
  wire _19219_;
  wire _19220_;
  wire _19221_;
  wire _19222_;
  wire _19223_;
  wire _19224_;
  wire _19225_;
  wire _19226_;
  wire _19227_;
  wire _19228_;
  wire _19229_;
  wire _19230_;
  wire _19231_;
  wire _19232_;
  wire _19233_;
  wire _19234_;
  wire _19235_;
  wire _19236_;
  wire _19237_;
  wire _19238_;
  wire _19239_;
  wire _19240_;
  wire _19241_;
  wire _19242_;
  wire _19243_;
  wire _19244_;
  wire _19245_;
  wire _19246_;
  wire _19247_;
  wire _19248_;
  wire _19249_;
  wire _19250_;
  wire _19251_;
  wire _19252_;
  wire _19253_;
  wire _19254_;
  wire _19255_;
  wire _19256_;
  wire _19257_;
  wire _19258_;
  wire _19259_;
  wire _19260_;
  wire _19261_;
  wire _19262_;
  wire _19263_;
  wire _19264_;
  wire _19265_;
  wire _19266_;
  wire _19267_;
  wire _19268_;
  wire _19269_;
  wire _19270_;
  wire _19271_;
  wire _19272_;
  wire _19273_;
  wire _19274_;
  wire _19275_;
  wire _19276_;
  wire _19277_;
  wire _19278_;
  wire _19279_;
  wire _19280_;
  wire _19281_;
  wire _19282_;
  wire _19283_;
  wire _19284_;
  wire _19285_;
  wire _19286_;
  wire _19287_;
  wire _19288_;
  wire _19289_;
  wire _19290_;
  wire _19291_;
  wire _19292_;
  wire _19293_;
  wire _19294_;
  wire _19295_;
  wire _19296_;
  wire _19297_;
  wire _19298_;
  wire _19299_;
  wire _19300_;
  wire _19301_;
  wire _19302_;
  wire _19303_;
  wire _19304_;
  wire _19305_;
  wire _19306_;
  wire _19307_;
  wire _19308_;
  wire _19309_;
  wire _19310_;
  wire _19311_;
  wire _19312_;
  wire _19313_;
  wire _19314_;
  wire _19315_;
  wire _19316_;
  wire _19317_;
  wire _19318_;
  wire _19319_;
  wire _19320_;
  wire _19321_;
  wire _19322_;
  wire _19323_;
  wire _19324_;
  wire _19325_;
  wire _19326_;
  wire _19327_;
  wire _19328_;
  wire _19329_;
  wire _19330_;
  wire _19331_;
  wire _19332_;
  wire _19333_;
  wire _19334_;
  wire _19335_;
  wire _19336_;
  wire _19337_;
  wire _19338_;
  wire _19339_;
  wire _19340_;
  wire _19341_;
  wire _19342_;
  wire _19343_;
  wire _19344_;
  wire _19345_;
  wire _19346_;
  wire _19347_;
  wire _19348_;
  wire _19349_;
  wire _19350_;
  wire _19351_;
  wire _19352_;
  wire _19353_;
  wire _19354_;
  wire _19355_;
  wire _19356_;
  wire _19357_;
  wire _19358_;
  wire _19359_;
  wire _19360_;
  wire _19361_;
  wire _19362_;
  wire _19363_;
  wire _19364_;
  wire _19365_;
  wire _19366_;
  wire _19367_;
  wire _19368_;
  wire _19369_;
  wire _19370_;
  wire _19371_;
  wire _19372_;
  wire _19373_;
  wire _19374_;
  wire _19375_;
  wire _19376_;
  wire _19377_;
  wire _19378_;
  wire _19379_;
  wire _19380_;
  wire _19381_;
  wire _19382_;
  wire _19383_;
  wire _19384_;
  wire _19385_;
  wire _19386_;
  wire _19387_;
  wire _19388_;
  wire _19389_;
  wire _19390_;
  wire _19391_;
  wire _19392_;
  wire _19393_;
  wire _19394_;
  wire _19395_;
  wire _19396_;
  wire _19397_;
  wire _19398_;
  wire _19399_;
  wire _19400_;
  wire _19401_;
  wire _19402_;
  wire _19403_;
  wire _19404_;
  wire _19405_;
  wire _19406_;
  wire _19407_;
  wire _19408_;
  wire _19409_;
  wire _19410_;
  wire _19411_;
  wire _19412_;
  wire _19413_;
  wire _19414_;
  wire _19415_;
  wire _19416_;
  wire _19417_;
  wire _19418_;
  wire _19419_;
  wire _19420_;
  wire _19421_;
  wire _19422_;
  wire _19423_;
  wire _19424_;
  wire _19425_;
  wire _19426_;
  wire _19427_;
  wire _19428_;
  wire _19429_;
  wire _19430_;
  wire _19431_;
  wire _19432_;
  wire _19433_;
  wire _19434_;
  wire _19435_;
  wire _19436_;
  wire _19437_;
  wire _19438_;
  wire _19439_;
  wire _19440_;
  wire _19441_;
  wire _19442_;
  wire _19443_;
  wire _19444_;
  wire _19445_;
  wire _19446_;
  wire _19447_;
  wire _19448_;
  wire _19449_;
  wire _19450_;
  wire _19451_;
  wire _19452_;
  wire _19453_;
  wire _19454_;
  wire _19455_;
  wire _19456_;
  wire _19457_;
  wire _19458_;
  wire _19459_;
  wire _19460_;
  wire _19461_;
  wire _19462_;
  wire _19463_;
  wire _19464_;
  wire _19465_;
  wire _19466_;
  wire _19467_;
  wire _19468_;
  wire _19469_;
  wire _19470_;
  wire _19471_;
  wire _19472_;
  wire _19473_;
  wire _19474_;
  wire _19475_;
  wire _19476_;
  wire _19477_;
  wire _19478_;
  wire _19479_;
  wire _19480_;
  wire _19481_;
  wire _19482_;
  wire _19483_;
  wire _19484_;
  wire _19485_;
  wire _19486_;
  wire _19487_;
  wire _19488_;
  wire _19489_;
  wire _19490_;
  wire _19491_;
  wire _19492_;
  wire _19493_;
  wire _19494_;
  wire _19495_;
  wire _19496_;
  wire _19497_;
  wire _19498_;
  wire _19499_;
  wire _19500_;
  wire _19501_;
  wire _19502_;
  wire _19503_;
  wire _19504_;
  wire _19505_;
  wire _19506_;
  wire _19507_;
  wire _19508_;
  wire _19509_;
  wire _19510_;
  wire _19511_;
  wire _19512_;
  wire _19513_;
  wire _19514_;
  wire _19515_;
  wire _19516_;
  wire _19517_;
  wire _19518_;
  wire _19519_;
  wire _19520_;
  wire _19521_;
  wire _19522_;
  wire _19523_;
  wire _19524_;
  wire _19525_;
  wire _19526_;
  wire _19527_;
  wire _19528_;
  wire _19529_;
  wire _19530_;
  wire _19531_;
  wire _19532_;
  wire _19533_;
  wire _19534_;
  wire _19535_;
  wire _19536_;
  wire _19537_;
  wire _19538_;
  wire _19539_;
  wire _19540_;
  wire _19541_;
  wire _19542_;
  wire _19543_;
  wire _19544_;
  wire _19545_;
  wire _19546_;
  wire _19547_;
  wire _19548_;
  wire _19549_;
  wire _19550_;
  wire _19551_;
  wire _19552_;
  wire _19553_;
  wire _19554_;
  wire _19555_;
  wire _19556_;
  wire _19557_;
  wire _19558_;
  wire _19559_;
  wire _19560_;
  wire _19561_;
  wire _19562_;
  wire _19563_;
  wire _19564_;
  wire _19565_;
  wire _19566_;
  wire _19567_;
  wire _19568_;
  wire _19569_;
  wire _19570_;
  wire _19571_;
  wire _19572_;
  wire _19573_;
  wire _19574_;
  wire _19575_;
  wire _19576_;
  wire _19577_;
  wire _19578_;
  wire _19579_;
  wire _19580_;
  wire _19581_;
  wire _19582_;
  wire _19583_;
  wire _19584_;
  wire _19585_;
  wire _19586_;
  wire _19587_;
  wire _19588_;
  wire _19589_;
  wire _19590_;
  wire _19591_;
  wire _19592_;
  wire _19593_;
  wire _19594_;
  wire _19595_;
  wire _19596_;
  wire _19597_;
  wire _19598_;
  wire _19599_;
  wire _19600_;
  wire _19601_;
  wire _19602_;
  wire _19603_;
  wire _19604_;
  wire _19605_;
  wire _19606_;
  wire _19607_;
  wire _19608_;
  wire _19609_;
  wire _19610_;
  wire _19611_;
  wire _19612_;
  wire _19613_;
  wire _19614_;
  wire _19615_;
  wire _19616_;
  wire _19617_;
  wire _19618_;
  wire _19619_;
  wire _19620_;
  wire _19621_;
  wire _19622_;
  wire _19623_;
  wire _19624_;
  wire _19625_;
  wire _19626_;
  wire _19627_;
  wire _19628_;
  wire _19629_;
  wire _19630_;
  wire _19631_;
  wire _19632_;
  wire _19633_;
  wire _19634_;
  wire _19635_;
  wire _19636_;
  wire _19637_;
  wire _19638_;
  wire _19639_;
  wire _19640_;
  wire _19641_;
  wire _19642_;
  wire _19643_;
  wire _19644_;
  wire _19645_;
  wire _19646_;
  wire _19647_;
  wire _19648_;
  wire _19649_;
  wire _19650_;
  wire _19651_;
  wire _19652_;
  wire _19653_;
  wire _19654_;
  wire _19655_;
  wire _19656_;
  wire _19657_;
  wire _19658_;
  wire _19659_;
  wire _19660_;
  wire _19661_;
  wire _19662_;
  wire _19663_;
  wire _19664_;
  wire _19665_;
  wire _19666_;
  wire _19667_;
  wire _19668_;
  wire _19669_;
  wire _19670_;
  wire _19671_;
  wire _19672_;
  wire _19673_;
  wire _19674_;
  wire _19675_;
  wire _19676_;
  wire _19677_;
  wire _19678_;
  wire _19679_;
  wire _19680_;
  wire _19681_;
  wire _19682_;
  wire _19683_;
  wire _19684_;
  wire _19685_;
  wire _19686_;
  wire _19687_;
  wire _19688_;
  wire _19689_;
  wire _19690_;
  wire _19691_;
  wire _19692_;
  wire _19693_;
  wire _19694_;
  wire _19695_;
  wire _19696_;
  wire _19697_;
  wire _19698_;
  wire _19699_;
  wire _19700_;
  wire _19701_;
  wire _19702_;
  wire _19703_;
  wire _19704_;
  wire _19705_;
  wire _19706_;
  wire _19707_;
  wire _19708_;
  wire _19709_;
  wire _19710_;
  wire _19711_;
  wire _19712_;
  wire _19713_;
  wire _19714_;
  wire _19715_;
  wire _19716_;
  wire _19717_;
  wire _19718_;
  wire _19719_;
  wire _19720_;
  wire _19721_;
  wire _19722_;
  wire _19723_;
  wire _19724_;
  wire _19725_;
  wire _19726_;
  wire _19727_;
  wire _19728_;
  wire _19729_;
  wire _19730_;
  wire _19731_;
  wire _19732_;
  wire _19733_;
  wire _19734_;
  wire _19735_;
  wire _19736_;
  wire _19737_;
  wire _19738_;
  wire _19739_;
  wire _19740_;
  wire _19741_;
  wire _19742_;
  wire _19743_;
  wire _19744_;
  wire _19745_;
  wire _19746_;
  wire _19747_;
  wire _19748_;
  wire _19749_;
  wire _19750_;
  wire _19751_;
  wire _19752_;
  wire _19753_;
  wire _19754_;
  wire _19755_;
  wire _19756_;
  wire _19757_;
  wire _19758_;
  wire _19759_;
  wire _19760_;
  wire _19761_;
  wire _19762_;
  wire _19763_;
  wire _19764_;
  wire _19765_;
  wire _19766_;
  wire _19767_;
  wire _19768_;
  wire _19769_;
  wire _19770_;
  wire _19771_;
  wire _19772_;
  wire _19773_;
  wire _19774_;
  wire _19775_;
  wire _19776_;
  wire _19777_;
  wire _19778_;
  wire _19779_;
  wire _19780_;
  wire _19781_;
  wire _19782_;
  wire _19783_;
  wire _19784_;
  wire _19785_;
  wire _19786_;
  wire _19787_;
  wire _19788_;
  wire _19789_;
  wire _19790_;
  wire _19791_;
  wire _19792_;
  wire _19793_;
  wire _19794_;
  wire _19795_;
  wire _19796_;
  wire _19797_;
  wire _19798_;
  wire _19799_;
  wire _19800_;
  wire _19801_;
  wire _19802_;
  wire _19803_;
  wire _19804_;
  wire _19805_;
  wire _19806_;
  wire _19807_;
  wire _19808_;
  wire _19809_;
  wire _19810_;
  wire _19811_;
  wire _19812_;
  wire _19813_;
  wire _19814_;
  wire _19815_;
  wire _19816_;
  wire _19817_;
  wire _19818_;
  wire _19819_;
  wire _19820_;
  wire _19821_;
  wire _19822_;
  wire _19823_;
  wire _19824_;
  wire _19825_;
  wire _19826_;
  wire _19827_;
  wire _19828_;
  wire _19829_;
  wire _19830_;
  wire _19831_;
  wire _19832_;
  wire _19833_;
  wire _19834_;
  wire _19835_;
  wire _19836_;
  wire _19837_;
  wire _19838_;
  wire _19839_;
  wire _19840_;
  wire _19841_;
  wire _19842_;
  wire _19843_;
  wire _19844_;
  wire _19845_;
  wire _19846_;
  wire _19847_;
  wire _19848_;
  wire _19849_;
  wire _19850_;
  wire _19851_;
  wire _19852_;
  wire _19853_;
  wire _19854_;
  wire _19855_;
  wire _19856_;
  wire _19857_;
  wire _19858_;
  wire _19859_;
  wire _19860_;
  wire _19861_;
  wire _19862_;
  wire _19863_;
  wire _19864_;
  wire _19865_;
  wire _19866_;
  wire _19867_;
  wire _19868_;
  wire _19869_;
  wire _19870_;
  wire _19871_;
  wire _19872_;
  wire _19873_;
  wire _19874_;
  wire _19875_;
  wire _19876_;
  wire _19877_;
  wire _19878_;
  wire _19879_;
  wire _19880_;
  wire _19881_;
  wire _19882_;
  wire _19883_;
  wire _19884_;
  wire _19885_;
  wire _19886_;
  wire _19887_;
  wire _19888_;
  wire _19889_;
  wire _19890_;
  wire _19891_;
  wire _19892_;
  wire _19893_;
  wire _19894_;
  wire _19895_;
  wire _19896_;
  wire _19897_;
  wire _19898_;
  wire _19899_;
  wire _19900_;
  wire _19901_;
  wire _19902_;
  wire _19903_;
  wire _19904_;
  wire _19905_;
  wire _19906_;
  wire _19907_;
  wire _19908_;
  wire _19909_;
  wire _19910_;
  wire _19911_;
  wire _19912_;
  wire _19913_;
  wire _19914_;
  wire _19915_;
  wire _19916_;
  wire _19917_;
  wire _19918_;
  wire _19919_;
  wire _19920_;
  wire _19921_;
  wire _19922_;
  wire _19923_;
  wire _19924_;
  wire _19925_;
  wire _19926_;
  wire _19927_;
  wire _19928_;
  wire _19929_;
  wire _19930_;
  wire _19931_;
  wire _19932_;
  wire _19933_;
  wire _19934_;
  wire _19935_;
  wire _19936_;
  wire _19937_;
  wire _19938_;
  wire _19939_;
  wire _19940_;
  wire _19941_;
  wire _19942_;
  wire _19943_;
  wire _19944_;
  wire _19945_;
  wire _19946_;
  wire _19947_;
  wire _19948_;
  wire _19949_;
  wire _19950_;
  wire _19951_;
  wire _19952_;
  wire _19953_;
  wire _19954_;
  wire _19955_;
  wire _19956_;
  wire _19957_;
  wire _19958_;
  wire _19959_;
  wire _19960_;
  wire _19961_;
  wire _19962_;
  wire _19963_;
  wire _19964_;
  wire _19965_;
  wire _19966_;
  wire _19967_;
  wire _19968_;
  wire _19969_;
  wire _19970_;
  wire _19971_;
  wire _19972_;
  wire _19973_;
  wire _19974_;
  wire _19975_;
  wire _19976_;
  wire _19977_;
  wire _19978_;
  wire _19979_;
  wire _19980_;
  wire _19981_;
  wire _19982_;
  wire _19983_;
  wire _19984_;
  wire _19985_;
  wire _19986_;
  wire _19987_;
  wire _19988_;
  wire _19989_;
  wire _19990_;
  wire _19991_;
  wire _19992_;
  wire _19993_;
  wire _19994_;
  wire _19995_;
  wire _19996_;
  wire _19997_;
  wire _19998_;
  wire _19999_;
  wire _20000_;
  wire _20001_;
  wire _20002_;
  wire _20003_;
  wire _20004_;
  wire _20005_;
  wire _20006_;
  wire _20007_;
  wire _20008_;
  wire _20009_;
  wire _20010_;
  wire _20011_;
  wire _20012_;
  wire _20013_;
  wire _20014_;
  wire _20015_;
  wire _20016_;
  wire _20017_;
  wire _20018_;
  wire _20019_;
  wire _20020_;
  wire _20021_;
  wire _20022_;
  wire _20023_;
  wire _20024_;
  wire _20025_;
  wire _20026_;
  wire _20027_;
  wire _20028_;
  wire _20029_;
  wire _20030_;
  wire _20031_;
  wire _20032_;
  wire _20033_;
  wire _20034_;
  wire _20035_;
  wire _20036_;
  wire _20037_;
  wire _20038_;
  wire _20039_;
  wire _20040_;
  wire _20041_;
  wire _20042_;
  wire _20043_;
  wire _20044_;
  wire _20045_;
  wire _20046_;
  wire _20047_;
  wire _20048_;
  wire _20049_;
  wire _20050_;
  wire _20051_;
  wire _20052_;
  wire _20053_;
  wire _20054_;
  wire _20055_;
  wire _20056_;
  wire _20057_;
  wire _20058_;
  wire _20059_;
  wire _20060_;
  wire _20061_;
  wire _20062_;
  wire _20063_;
  wire _20064_;
  wire _20065_;
  wire _20066_;
  wire _20067_;
  wire _20068_;
  wire _20069_;
  wire _20070_;
  wire _20071_;
  wire _20072_;
  wire _20073_;
  wire _20074_;
  wire _20075_;
  wire _20076_;
  wire _20077_;
  wire _20078_;
  wire _20079_;
  wire _20080_;
  wire _20081_;
  wire _20082_;
  wire _20083_;
  wire _20084_;
  wire _20085_;
  wire _20086_;
  wire _20087_;
  wire _20088_;
  wire _20089_;
  wire _20090_;
  wire _20091_;
  wire _20092_;
  wire _20093_;
  wire _20094_;
  wire _20095_;
  wire _20096_;
  wire _20097_;
  wire _20098_;
  wire _20099_;
  wire _20100_;
  wire _20101_;
  wire _20102_;
  wire _20103_;
  wire _20104_;
  wire _20105_;
  wire _20106_;
  wire _20107_;
  wire _20108_;
  wire _20109_;
  wire _20110_;
  wire _20111_;
  wire _20112_;
  wire _20113_;
  wire _20114_;
  wire _20115_;
  wire _20116_;
  wire _20117_;
  wire _20118_;
  wire _20119_;
  wire _20120_;
  wire _20121_;
  wire _20122_;
  wire _20123_;
  wire _20124_;
  wire _20125_;
  wire _20126_;
  wire _20127_;
  wire _20128_;
  wire _20129_;
  wire _20130_;
  wire _20131_;
  wire _20132_;
  wire _20133_;
  wire _20134_;
  wire _20135_;
  wire _20136_;
  wire _20137_;
  wire _20138_;
  wire _20139_;
  wire _20140_;
  wire _20141_;
  wire _20142_;
  wire _20143_;
  wire _20144_;
  wire _20145_;
  wire _20146_;
  wire _20147_;
  wire _20148_;
  wire _20149_;
  wire _20150_;
  wire _20151_;
  wire _20152_;
  wire _20153_;
  wire _20154_;
  wire _20155_;
  wire _20156_;
  wire _20157_;
  wire _20158_;
  wire _20159_;
  wire _20160_;
  wire _20161_;
  wire _20162_;
  wire _20163_;
  wire _20164_;
  wire _20165_;
  wire _20166_;
  wire _20167_;
  wire _20168_;
  wire _20169_;
  wire _20170_;
  wire _20171_;
  wire _20172_;
  wire _20173_;
  wire _20174_;
  wire _20175_;
  wire _20176_;
  wire _20177_;
  wire _20178_;
  wire _20179_;
  wire _20180_;
  wire _20181_;
  wire _20182_;
  wire _20183_;
  wire _20184_;
  wire _20185_;
  wire _20186_;
  wire _20187_;
  wire _20188_;
  wire _20189_;
  wire _20190_;
  wire _20191_;
  wire _20192_;
  wire _20193_;
  wire _20194_;
  wire _20195_;
  wire _20196_;
  wire _20197_;
  wire _20198_;
  wire _20199_;
  wire _20200_;
  wire _20201_;
  wire _20202_;
  wire _20203_;
  wire _20204_;
  wire _20205_;
  wire _20206_;
  wire _20207_;
  wire _20208_;
  wire _20209_;
  wire _20210_;
  wire _20211_;
  wire _20212_;
  wire _20213_;
  wire _20214_;
  wire _20215_;
  wire _20216_;
  wire _20217_;
  wire _20218_;
  wire _20219_;
  wire _20220_;
  wire _20221_;
  wire _20222_;
  wire _20223_;
  wire _20224_;
  wire _20225_;
  wire _20226_;
  wire _20227_;
  wire _20228_;
  wire _20229_;
  wire _20230_;
  wire _20231_;
  wire _20232_;
  wire _20233_;
  wire _20234_;
  wire _20235_;
  wire _20236_;
  wire _20237_;
  wire _20238_;
  wire _20239_;
  wire _20240_;
  wire _20241_;
  wire _20242_;
  wire _20243_;
  wire _20244_;
  wire _20245_;
  wire _20246_;
  wire _20247_;
  wire _20248_;
  wire _20249_;
  wire _20250_;
  wire _20251_;
  wire _20252_;
  wire _20253_;
  wire _20254_;
  wire _20255_;
  wire _20256_;
  wire _20257_;
  wire _20258_;
  wire _20259_;
  wire _20260_;
  wire _20261_;
  wire _20262_;
  wire _20263_;
  wire _20264_;
  wire _20265_;
  wire _20266_;
  wire _20267_;
  wire _20268_;
  wire _20269_;
  wire _20270_;
  wire _20271_;
  wire _20272_;
  wire _20273_;
  wire _20274_;
  wire _20275_;
  wire _20276_;
  wire _20277_;
  wire _20278_;
  wire _20279_;
  wire _20280_;
  wire _20281_;
  wire _20282_;
  wire _20283_;
  wire _20284_;
  wire _20285_;
  wire _20286_;
  wire _20287_;
  wire _20288_;
  wire _20289_;
  wire _20290_;
  wire _20291_;
  wire _20292_;
  wire _20293_;
  wire _20294_;
  wire _20295_;
  wire _20296_;
  wire _20297_;
  wire _20298_;
  wire _20299_;
  wire _20300_;
  wire _20301_;
  wire _20302_;
  wire _20303_;
  wire _20304_;
  wire _20305_;
  wire _20306_;
  wire _20307_;
  wire _20308_;
  wire _20309_;
  wire _20310_;
  wire _20311_;
  wire _20312_;
  wire _20313_;
  wire _20314_;
  wire _20315_;
  wire _20316_;
  wire _20317_;
  wire _20318_;
  wire _20319_;
  wire _20320_;
  wire _20321_;
  wire _20322_;
  wire _20323_;
  wire _20324_;
  wire _20325_;
  wire _20326_;
  wire _20327_;
  wire _20328_;
  wire _20329_;
  wire _20330_;
  wire _20331_;
  wire _20332_;
  wire _20333_;
  wire _20334_;
  wire _20335_;
  wire _20336_;
  wire _20337_;
  wire _20338_;
  wire _20339_;
  wire _20340_;
  wire _20341_;
  wire _20342_;
  wire _20343_;
  wire _20344_;
  wire _20345_;
  wire _20346_;
  wire _20347_;
  wire _20348_;
  wire _20349_;
  wire _20350_;
  wire _20351_;
  wire _20352_;
  wire _20353_;
  wire _20354_;
  wire _20355_;
  wire _20356_;
  wire _20357_;
  wire _20358_;
  wire _20359_;
  wire _20360_;
  wire _20361_;
  wire _20362_;
  wire _20363_;
  wire _20364_;
  wire _20365_;
  wire _20366_;
  wire _20367_;
  wire _20368_;
  wire _20369_;
  wire _20370_;
  wire _20371_;
  wire _20372_;
  wire _20373_;
  wire _20374_;
  wire _20375_;
  wire _20376_;
  wire _20377_;
  wire _20378_;
  wire _20379_;
  wire _20380_;
  wire _20381_;
  wire _20382_;
  wire _20383_;
  wire _20384_;
  wire _20385_;
  wire _20386_;
  wire _20387_;
  wire _20388_;
  wire _20389_;
  wire _20390_;
  wire _20391_;
  wire _20392_;
  wire _20393_;
  wire _20394_;
  wire _20395_;
  wire _20396_;
  wire _20397_;
  wire _20398_;
  wire _20399_;
  wire _20400_;
  wire _20401_;
  wire _20402_;
  wire _20403_;
  wire _20404_;
  wire _20405_;
  wire _20406_;
  wire _20407_;
  wire _20408_;
  wire _20409_;
  wire _20410_;
  wire _20411_;
  wire _20412_;
  wire _20413_;
  wire _20414_;
  wire _20415_;
  wire _20416_;
  wire _20417_;
  wire _20418_;
  wire _20419_;
  wire _20420_;
  wire _20421_;
  wire _20422_;
  wire _20423_;
  wire _20424_;
  wire _20425_;
  wire _20426_;
  wire _20427_;
  wire _20428_;
  wire _20429_;
  wire _20430_;
  wire _20431_;
  wire _20432_;
  wire _20433_;
  wire _20434_;
  wire _20435_;
  wire _20436_;
  wire _20437_;
  wire _20438_;
  wire _20439_;
  wire _20440_;
  wire _20441_;
  wire _20442_;
  wire _20443_;
  wire _20444_;
  wire _20445_;
  wire _20446_;
  wire _20447_;
  wire _20448_;
  wire _20449_;
  wire _20450_;
  wire _20451_;
  wire _20452_;
  wire _20453_;
  wire _20454_;
  wire _20455_;
  wire _20456_;
  wire _20457_;
  wire _20458_;
  wire _20459_;
  wire _20460_;
  wire _20461_;
  wire _20462_;
  wire _20463_;
  wire _20464_;
  wire _20465_;
  wire _20466_;
  wire _20467_;
  wire _20468_;
  wire _20469_;
  wire _20470_;
  wire _20471_;
  wire _20472_;
  wire _20473_;
  wire _20474_;
  wire _20475_;
  wire _20476_;
  wire _20477_;
  wire _20478_;
  wire _20479_;
  wire _20480_;
  wire _20481_;
  wire _20482_;
  wire _20483_;
  wire _20484_;
  wire _20485_;
  wire _20486_;
  wire _20487_;
  wire _20488_;
  wire _20489_;
  wire _20490_;
  wire _20491_;
  wire _20492_;
  wire _20493_;
  wire _20494_;
  wire _20495_;
  wire _20496_;
  wire _20497_;
  wire _20498_;
  wire _20499_;
  wire _20500_;
  wire _20501_;
  wire _20502_;
  wire _20503_;
  wire _20504_;
  wire _20505_;
  wire _20506_;
  wire _20507_;
  wire _20508_;
  wire _20509_;
  wire _20510_;
  wire _20511_;
  wire _20512_;
  wire _20513_;
  wire _20514_;
  wire _20515_;
  wire _20516_;
  wire _20517_;
  wire _20518_;
  wire _20519_;
  wire _20520_;
  wire _20521_;
  wire _20522_;
  wire _20523_;
  wire _20524_;
  wire _20525_;
  wire _20526_;
  wire _20527_;
  wire _20528_;
  wire _20529_;
  wire _20530_;
  wire _20531_;
  wire _20532_;
  wire _20533_;
  wire _20534_;
  wire _20535_;
  wire _20536_;
  wire _20537_;
  wire _20538_;
  wire _20539_;
  wire _20540_;
  wire _20541_;
  wire _20542_;
  wire _20543_;
  wire _20544_;
  wire _20545_;
  wire _20546_;
  wire _20547_;
  wire _20548_;
  wire _20549_;
  wire _20550_;
  wire _20551_;
  wire _20552_;
  wire _20553_;
  wire _20554_;
  wire _20555_;
  wire _20556_;
  wire _20557_;
  wire _20558_;
  wire _20559_;
  wire _20560_;
  wire _20561_;
  wire _20562_;
  wire _20563_;
  wire _20564_;
  wire _20565_;
  wire _20566_;
  wire _20567_;
  wire _20568_;
  wire _20569_;
  wire _20570_;
  wire _20571_;
  wire _20572_;
  wire _20573_;
  wire _20574_;
  wire _20575_;
  wire _20576_;
  wire _20577_;
  wire _20578_;
  wire _20579_;
  wire _20580_;
  wire _20581_;
  wire _20582_;
  wire _20583_;
  wire _20584_;
  wire _20585_;
  wire _20586_;
  wire _20587_;
  wire _20588_;
  wire _20589_;
  wire _20590_;
  wire _20591_;
  wire _20592_;
  wire _20593_;
  wire _20594_;
  wire _20595_;
  wire _20596_;
  wire _20597_;
  wire _20598_;
  wire _20599_;
  wire _20600_;
  wire _20601_;
  wire _20602_;
  wire _20603_;
  wire _20604_;
  wire _20605_;
  wire _20606_;
  wire _20607_;
  wire _20608_;
  wire _20609_;
  wire _20610_;
  wire _20611_;
  wire _20612_;
  wire _20613_;
  wire _20614_;
  wire _20615_;
  wire _20616_;
  wire _20617_;
  wire _20618_;
  wire _20619_;
  wire _20620_;
  wire _20621_;
  wire _20622_;
  wire _20623_;
  wire _20624_;
  wire _20625_;
  wire _20626_;
  wire _20627_;
  wire _20628_;
  wire _20629_;
  wire _20630_;
  wire _20631_;
  wire _20632_;
  wire _20633_;
  wire _20634_;
  wire _20635_;
  wire _20636_;
  wire _20637_;
  wire _20638_;
  wire _20639_;
  wire _20640_;
  wire _20641_;
  wire _20642_;
  wire _20643_;
  wire _20644_;
  wire _20645_;
  wire _20646_;
  wire _20647_;
  wire _20648_;
  wire _20649_;
  wire _20650_;
  wire _20651_;
  wire _20652_;
  wire _20653_;
  wire _20654_;
  wire _20655_;
  wire _20656_;
  wire _20657_;
  wire _20658_;
  wire _20659_;
  wire _20660_;
  wire _20661_;
  wire _20662_;
  wire _20663_;
  wire _20664_;
  wire _20665_;
  wire _20666_;
  wire _20667_;
  wire _20668_;
  wire _20669_;
  wire _20670_;
  wire _20671_;
  wire _20672_;
  wire _20673_;
  wire _20674_;
  wire _20675_;
  wire _20676_;
  wire _20677_;
  wire _20678_;
  wire _20679_;
  wire _20680_;
  wire _20681_;
  wire _20682_;
  wire _20683_;
  wire _20684_;
  wire _20685_;
  wire _20686_;
  wire _20687_;
  wire _20688_;
  wire _20689_;
  wire _20690_;
  wire _20691_;
  wire _20692_;
  wire _20693_;
  wire _20694_;
  wire _20695_;
  wire _20696_;
  wire _20697_;
  wire _20698_;
  wire _20699_;
  wire _20700_;
  wire _20701_;
  wire _20702_;
  wire _20703_;
  wire _20704_;
  wire _20705_;
  wire _20706_;
  wire _20707_;
  wire _20708_;
  wire _20709_;
  wire _20710_;
  wire _20711_;
  wire _20712_;
  wire _20713_;
  wire _20714_;
  wire _20715_;
  wire _20716_;
  wire _20717_;
  wire _20718_;
  wire _20719_;
  wire _20720_;
  wire _20721_;
  wire _20722_;
  wire _20723_;
  wire _20724_;
  wire _20725_;
  wire _20726_;
  wire _20727_;
  wire _20728_;
  wire _20729_;
  wire _20730_;
  wire _20731_;
  wire _20732_;
  wire _20733_;
  wire _20734_;
  wire _20735_;
  wire _20736_;
  wire _20737_;
  wire _20738_;
  wire _20739_;
  wire _20740_;
  wire _20741_;
  wire _20742_;
  wire _20743_;
  wire _20744_;
  wire _20745_;
  wire _20746_;
  wire _20747_;
  wire _20748_;
  wire _20749_;
  wire _20750_;
  wire _20751_;
  wire _20752_;
  wire _20753_;
  wire _20754_;
  wire _20755_;
  wire _20756_;
  wire _20757_;
  wire _20758_;
  wire _20759_;
  wire _20760_;
  wire _20761_;
  wire _20762_;
  wire _20763_;
  wire _20764_;
  wire _20765_;
  wire _20766_;
  wire _20767_;
  wire _20768_;
  wire _20769_;
  wire _20770_;
  wire _20771_;
  wire _20772_;
  wire _20773_;
  wire _20774_;
  wire _20775_;
  wire _20776_;
  wire _20777_;
  wire _20778_;
  wire _20779_;
  wire _20780_;
  wire _20781_;
  wire _20782_;
  wire _20783_;
  wire _20784_;
  wire _20785_;
  wire _20786_;
  wire _20787_;
  wire _20788_;
  wire _20789_;
  wire _20790_;
  wire _20791_;
  wire _20792_;
  wire _20793_;
  wire _20794_;
  wire _20795_;
  wire _20796_;
  wire _20797_;
  wire _20798_;
  wire _20799_;
  wire _20800_;
  wire _20801_;
  wire _20802_;
  wire _20803_;
  wire _20804_;
  wire _20805_;
  wire _20806_;
  wire _20807_;
  wire _20808_;
  wire _20809_;
  wire _20810_;
  wire _20811_;
  wire _20812_;
  wire _20813_;
  wire _20814_;
  wire _20815_;
  wire _20816_;
  wire _20817_;
  wire _20818_;
  wire _20819_;
  wire _20820_;
  wire _20821_;
  wire _20822_;
  wire _20823_;
  wire _20824_;
  wire _20825_;
  wire _20826_;
  wire _20827_;
  wire _20828_;
  wire _20829_;
  wire _20830_;
  wire _20831_;
  wire _20832_;
  wire _20833_;
  wire _20834_;
  wire _20835_;
  wire _20836_;
  wire _20837_;
  wire _20838_;
  wire _20839_;
  wire _20840_;
  wire _20841_;
  wire _20842_;
  wire _20843_;
  wire _20844_;
  wire _20845_;
  wire _20846_;
  wire _20847_;
  wire _20848_;
  wire _20849_;
  wire _20850_;
  wire _20851_;
  wire _20852_;
  wire _20853_;
  wire _20854_;
  wire _20855_;
  wire _20856_;
  wire _20857_;
  wire _20858_;
  wire _20859_;
  wire _20860_;
  wire _20861_;
  wire _20862_;
  wire _20863_;
  wire _20864_;
  wire _20865_;
  wire _20866_;
  wire _20867_;
  wire _20868_;
  wire _20869_;
  wire _20870_;
  wire _20871_;
  wire _20872_;
  wire _20873_;
  wire _20874_;
  wire _20875_;
  wire _20876_;
  wire _20877_;
  wire _20878_;
  wire _20879_;
  wire _20880_;
  wire _20881_;
  wire _20882_;
  wire _20883_;
  wire _20884_;
  wire _20885_;
  wire _20886_;
  wire _20887_;
  wire _20888_;
  wire _20889_;
  wire _20890_;
  wire _20891_;
  wire _20892_;
  wire _20893_;
  wire _20894_;
  wire _20895_;
  wire _20896_;
  wire _20897_;
  wire _20898_;
  wire _20899_;
  wire _20900_;
  wire _20901_;
  wire _20902_;
  wire _20903_;
  wire _20904_;
  wire _20905_;
  wire _20906_;
  wire _20907_;
  wire _20908_;
  wire _20909_;
  wire _20910_;
  wire _20911_;
  wire _20912_;
  wire _20913_;
  wire _20914_;
  wire _20915_;
  wire _20916_;
  wire _20917_;
  wire _20918_;
  wire _20919_;
  wire _20920_;
  wire _20921_;
  wire _20922_;
  wire _20923_;
  wire _20924_;
  wire _20925_;
  wire _20926_;
  wire _20927_;
  wire _20928_;
  wire _20929_;
  wire _20930_;
  wire _20931_;
  wire _20932_;
  wire _20933_;
  wire _20934_;
  wire _20935_;
  wire _20936_;
  wire _20937_;
  wire _20938_;
  wire _20939_;
  wire _20940_;
  wire _20941_;
  wire _20942_;
  wire _20943_;
  wire _20944_;
  wire _20945_;
  wire _20946_;
  wire _20947_;
  wire _20948_;
  wire _20949_;
  wire _20950_;
  wire _20951_;
  wire _20952_;
  wire _20953_;
  wire _20954_;
  wire _20955_;
  wire _20956_;
  wire _20957_;
  wire _20958_;
  wire _20959_;
  wire _20960_;
  wire _20961_;
  wire _20962_;
  wire _20963_;
  wire _20964_;
  wire _20965_;
  wire _20966_;
  wire _20967_;
  wire _20968_;
  wire _20969_;
  wire _20970_;
  wire _20971_;
  wire _20972_;
  wire _20973_;
  wire _20974_;
  wire _20975_;
  wire _20976_;
  wire _20977_;
  wire _20978_;
  wire _20979_;
  wire _20980_;
  wire _20981_;
  wire _20982_;
  wire _20983_;
  wire _20984_;
  wire _20985_;
  wire _20986_;
  wire _20987_;
  wire _20988_;
  wire _20989_;
  wire _20990_;
  wire _20991_;
  wire _20992_;
  wire _20993_;
  wire _20994_;
  wire _20995_;
  wire _20996_;
  wire _20997_;
  wire _20998_;
  wire _20999_;
  wire _21000_;
  wire _21001_;
  wire _21002_;
  wire _21003_;
  wire _21004_;
  wire _21005_;
  wire _21006_;
  wire _21007_;
  wire _21008_;
  wire _21009_;
  wire _21010_;
  wire _21011_;
  wire _21012_;
  wire _21013_;
  wire _21014_;
  wire _21015_;
  wire _21016_;
  wire _21017_;
  wire _21018_;
  wire _21019_;
  wire _21020_;
  wire _21021_;
  wire _21022_;
  wire _21023_;
  wire _21024_;
  wire _21025_;
  wire _21026_;
  wire _21027_;
  wire _21028_;
  wire _21029_;
  wire _21030_;
  wire _21031_;
  wire _21032_;
  wire _21033_;
  wire _21034_;
  wire _21035_;
  wire _21036_;
  wire _21037_;
  wire _21038_;
  wire _21039_;
  wire _21040_;
  wire _21041_;
  wire _21042_;
  wire _21043_;
  wire _21044_;
  wire _21045_;
  wire _21046_;
  wire _21047_;
  wire _21048_;
  wire _21049_;
  wire _21050_;
  wire _21051_;
  wire _21052_;
  wire _21053_;
  wire _21054_;
  wire _21055_;
  wire _21056_;
  wire _21057_;
  wire _21058_;
  wire _21059_;
  wire _21060_;
  wire _21061_;
  wire _21062_;
  wire _21063_;
  wire _21064_;
  wire _21065_;
  wire _21066_;
  wire _21067_;
  wire _21068_;
  wire _21069_;
  wire _21070_;
  wire _21071_;
  wire _21072_;
  wire _21073_;
  wire _21074_;
  wire _21075_;
  wire _21076_;
  wire _21077_;
  wire _21078_;
  wire _21079_;
  wire _21080_;
  wire _21081_;
  wire _21082_;
  wire _21083_;
  wire _21084_;
  wire _21085_;
  wire _21086_;
  wire _21087_;
  wire _21088_;
  wire _21089_;
  wire _21090_;
  wire _21091_;
  wire _21092_;
  wire _21093_;
  wire _21094_;
  wire _21095_;
  wire _21096_;
  wire _21097_;
  wire _21098_;
  wire _21099_;
  wire _21100_;
  wire _21101_;
  wire _21102_;
  wire _21103_;
  wire _21104_;
  wire _21105_;
  wire _21106_;
  wire _21107_;
  wire _21108_;
  wire _21109_;
  wire _21110_;
  wire _21111_;
  wire _21112_;
  wire _21113_;
  wire _21114_;
  wire _21115_;
  wire _21116_;
  wire _21117_;
  wire _21118_;
  wire _21119_;
  wire _21120_;
  wire _21121_;
  wire _21122_;
  wire _21123_;
  wire _21124_;
  wire _21125_;
  wire _21126_;
  wire _21127_;
  wire _21128_;
  wire _21129_;
  wire _21130_;
  wire _21131_;
  wire _21132_;
  wire _21133_;
  wire _21134_;
  wire _21135_;
  wire _21136_;
  wire _21137_;
  wire _21138_;
  wire _21139_;
  wire _21140_;
  wire _21141_;
  wire _21142_;
  wire _21143_;
  wire _21144_;
  wire _21145_;
  wire _21146_;
  wire _21147_;
  wire _21148_;
  wire _21149_;
  wire _21150_;
  wire _21151_;
  wire _21152_;
  wire _21153_;
  wire _21154_;
  wire _21155_;
  wire _21156_;
  wire _21157_;
  wire _21158_;
  wire _21159_;
  wire _21160_;
  wire _21161_;
  wire _21162_;
  wire _21163_;
  wire _21164_;
  wire _21165_;
  wire _21166_;
  wire _21167_;
  wire _21168_;
  wire _21169_;
  wire _21170_;
  wire _21171_;
  wire _21172_;
  wire _21173_;
  wire _21174_;
  wire _21175_;
  wire _21176_;
  wire _21177_;
  wire _21178_;
  wire _21179_;
  wire _21180_;
  wire _21181_;
  wire _21182_;
  wire _21183_;
  wire _21184_;
  wire _21185_;
  wire _21186_;
  wire _21187_;
  wire _21188_;
  wire _21189_;
  wire _21190_;
  wire _21191_;
  wire _21192_;
  wire _21193_;
  wire _21194_;
  wire _21195_;
  wire _21196_;
  wire _21197_;
  wire _21198_;
  wire _21199_;
  wire _21200_;
  wire _21201_;
  wire _21202_;
  wire _21203_;
  wire _21204_;
  wire _21205_;
  wire _21206_;
  wire _21207_;
  wire _21208_;
  wire _21209_;
  wire _21210_;
  wire _21211_;
  wire _21212_;
  wire _21213_;
  wire _21214_;
  wire _21215_;
  wire _21216_;
  wire _21217_;
  wire _21218_;
  wire _21219_;
  wire _21220_;
  wire _21221_;
  wire _21222_;
  wire _21223_;
  wire _21224_;
  wire _21225_;
  wire _21226_;
  wire _21227_;
  wire _21228_;
  wire _21229_;
  wire _21230_;
  wire _21231_;
  wire _21232_;
  wire _21233_;
  wire _21234_;
  wire _21235_;
  wire _21236_;
  wire _21237_;
  wire _21238_;
  wire _21239_;
  wire _21240_;
  wire _21241_;
  wire _21242_;
  wire _21243_;
  wire _21244_;
  wire _21245_;
  wire _21246_;
  wire _21247_;
  wire _21248_;
  wire _21249_;
  wire _21250_;
  wire _21251_;
  wire _21252_;
  wire _21253_;
  wire _21254_;
  wire _21255_;
  wire _21256_;
  wire _21257_;
  wire _21258_;
  wire _21259_;
  wire _21260_;
  wire _21261_;
  wire _21262_;
  wire _21263_;
  wire _21264_;
  wire _21265_;
  wire _21266_;
  wire _21267_;
  wire _21268_;
  wire _21269_;
  wire _21270_;
  wire _21271_;
  wire _21272_;
  wire _21273_;
  wire _21274_;
  wire _21275_;
  wire _21276_;
  wire _21277_;
  wire _21278_;
  wire _21279_;
  wire _21280_;
  wire _21281_;
  wire _21282_;
  wire _21283_;
  wire _21284_;
  wire _21285_;
  wire _21286_;
  wire _21287_;
  wire _21288_;
  wire _21289_;
  wire _21290_;
  wire _21291_;
  wire _21292_;
  wire _21293_;
  wire _21294_;
  wire _21295_;
  wire _21296_;
  wire _21297_;
  wire _21298_;
  wire _21299_;
  wire _21300_;
  wire _21301_;
  wire _21302_;
  wire _21303_;
  wire _21304_;
  wire _21305_;
  wire _21306_;
  wire _21307_;
  wire _21308_;
  wire _21309_;
  wire _21310_;
  wire _21311_;
  wire _21312_;
  wire _21313_;
  wire _21314_;
  wire _21315_;
  wire _21316_;
  wire _21317_;
  wire _21318_;
  wire _21319_;
  wire _21320_;
  wire _21321_;
  wire _21322_;
  wire _21323_;
  wire _21324_;
  wire _21325_;
  wire _21326_;
  wire _21327_;
  wire _21328_;
  wire _21329_;
  wire _21330_;
  wire _21331_;
  wire _21332_;
  wire _21333_;
  wire _21334_;
  wire _21335_;
  wire _21336_;
  wire _21337_;
  wire _21338_;
  wire _21339_;
  wire _21340_;
  wire _21341_;
  wire _21342_;
  wire _21343_;
  wire _21344_;
  wire _21345_;
  wire _21346_;
  wire _21347_;
  wire _21348_;
  wire _21349_;
  wire _21350_;
  wire _21351_;
  wire _21352_;
  wire _21353_;
  wire _21354_;
  wire _21355_;
  wire _21356_;
  wire _21357_;
  wire _21358_;
  wire _21359_;
  wire _21360_;
  wire _21361_;
  wire _21362_;
  wire _21363_;
  wire _21364_;
  wire _21365_;
  wire _21366_;
  wire _21367_;
  wire _21368_;
  wire _21369_;
  wire _21370_;
  wire _21371_;
  wire _21372_;
  wire _21373_;
  wire _21374_;
  wire _21375_;
  wire _21376_;
  wire _21377_;
  wire _21378_;
  wire _21379_;
  wire _21380_;
  wire _21381_;
  wire _21382_;
  wire _21383_;
  wire _21384_;
  wire _21385_;
  wire _21386_;
  wire _21387_;
  wire _21388_;
  wire _21389_;
  wire _21390_;
  wire _21391_;
  wire _21392_;
  wire _21393_;
  wire _21394_;
  wire _21395_;
  wire _21396_;
  wire _21397_;
  wire _21398_;
  wire _21399_;
  wire _21400_;
  wire _21401_;
  wire _21402_;
  wire _21403_;
  wire _21404_;
  wire _21405_;
  wire _21406_;
  wire _21407_;
  wire _21408_;
  wire _21409_;
  wire _21410_;
  wire _21411_;
  wire _21412_;
  wire _21413_;
  wire _21414_;
  wire _21415_;
  wire _21416_;
  wire _21417_;
  wire _21418_;
  wire _21419_;
  wire _21420_;
  wire _21421_;
  wire _21422_;
  wire _21423_;
  wire _21424_;
  wire _21425_;
  wire _21426_;
  wire _21427_;
  wire _21428_;
  wire _21429_;
  wire _21430_;
  wire _21431_;
  wire _21432_;
  wire _21433_;
  wire _21434_;
  wire _21435_;
  wire _21436_;
  wire _21437_;
  wire _21438_;
  wire _21439_;
  wire _21440_;
  wire _21441_;
  wire _21442_;
  wire _21443_;
  wire _21444_;
  wire _21445_;
  wire _21446_;
  wire _21447_;
  wire _21448_;
  wire _21449_;
  wire _21450_;
  wire _21451_;
  wire _21452_;
  wire _21453_;
  wire _21454_;
  wire _21455_;
  wire _21456_;
  wire _21457_;
  wire _21458_;
  wire _21459_;
  wire _21460_;
  wire _21461_;
  wire _21462_;
  wire _21463_;
  wire _21464_;
  wire _21465_;
  wire _21466_;
  wire _21467_;
  wire _21468_;
  wire _21469_;
  wire _21470_;
  wire _21471_;
  wire _21472_;
  wire _21473_;
  wire _21474_;
  wire _21475_;
  wire _21476_;
  wire _21477_;
  wire _21478_;
  wire _21479_;
  wire _21480_;
  wire _21481_;
  wire _21482_;
  wire _21483_;
  wire _21484_;
  wire _21485_;
  wire _21486_;
  wire _21487_;
  wire _21488_;
  wire _21489_;
  wire _21490_;
  wire _21491_;
  wire _21492_;
  wire _21493_;
  wire _21494_;
  wire _21495_;
  wire _21496_;
  wire _21497_;
  wire _21498_;
  wire _21499_;
  wire _21500_;
  wire _21501_;
  wire _21502_;
  wire _21503_;
  wire _21504_;
  wire _21505_;
  wire _21506_;
  wire _21507_;
  wire _21508_;
  wire _21509_;
  wire _21510_;
  wire _21511_;
  wire _21512_;
  wire _21513_;
  wire _21514_;
  wire _21515_;
  wire _21516_;
  wire _21517_;
  wire _21518_;
  wire _21519_;
  wire _21520_;
  wire _21521_;
  wire _21522_;
  wire _21523_;
  wire _21524_;
  wire _21525_;
  wire _21526_;
  wire _21527_;
  wire _21528_;
  wire _21529_;
  wire _21530_;
  wire _21531_;
  wire _21532_;
  wire _21533_;
  wire _21534_;
  wire _21535_;
  wire _21536_;
  wire _21537_;
  wire _21538_;
  wire _21539_;
  wire _21540_;
  wire _21541_;
  wire _21542_;
  wire _21543_;
  wire _21544_;
  wire _21545_;
  wire _21546_;
  wire _21547_;
  wire _21548_;
  wire _21549_;
  wire _21550_;
  wire _21551_;
  wire _21552_;
  wire _21553_;
  wire _21554_;
  wire _21555_;
  wire _21556_;
  wire _21557_;
  wire _21558_;
  wire _21559_;
  wire _21560_;
  wire _21561_;
  wire _21562_;
  wire _21563_;
  wire _21564_;
  wire _21565_;
  wire _21566_;
  wire _21567_;
  wire _21568_;
  wire _21569_;
  wire _21570_;
  wire _21571_;
  wire _21572_;
  wire _21573_;
  wire _21574_;
  wire _21575_;
  wire _21576_;
  wire _21577_;
  wire _21578_;
  wire _21579_;
  wire _21580_;
  wire _21581_;
  wire _21582_;
  wire _21583_;
  wire _21584_;
  wire _21585_;
  wire _21586_;
  wire _21587_;
  wire _21588_;
  wire _21589_;
  wire _21590_;
  wire _21591_;
  wire _21592_;
  wire _21593_;
  wire _21594_;
  wire _21595_;
  wire _21596_;
  wire _21597_;
  wire _21598_;
  wire _21599_;
  wire _21600_;
  wire _21601_;
  wire _21602_;
  wire _21603_;
  wire _21604_;
  wire _21605_;
  wire _21606_;
  wire _21607_;
  wire _21608_;
  wire _21609_;
  wire _21610_;
  wire _21611_;
  wire _21612_;
  wire _21613_;
  wire _21614_;
  wire _21615_;
  wire _21616_;
  wire _21617_;
  wire _21618_;
  wire _21619_;
  wire _21620_;
  wire _21621_;
  wire _21622_;
  wire _21623_;
  wire _21624_;
  wire _21625_;
  wire _21626_;
  wire _21627_;
  wire _21628_;
  wire _21629_;
  wire _21630_;
  wire _21631_;
  wire _21632_;
  wire _21633_;
  wire _21634_;
  wire _21635_;
  wire _21636_;
  wire _21637_;
  wire _21638_;
  wire _21639_;
  wire _21640_;
  wire _21641_;
  wire _21642_;
  wire _21643_;
  wire _21644_;
  wire _21645_;
  wire _21646_;
  wire _21647_;
  wire _21648_;
  wire _21649_;
  wire _21650_;
  wire _21651_;
  wire _21652_;
  wire _21653_;
  wire _21654_;
  wire _21655_;
  wire _21656_;
  wire _21657_;
  wire _21658_;
  wire _21659_;
  wire _21660_;
  wire _21661_;
  wire _21662_;
  wire _21663_;
  wire _21664_;
  wire _21665_;
  wire _21666_;
  wire _21667_;
  wire _21668_;
  wire _21669_;
  wire _21670_;
  wire _21671_;
  wire _21672_;
  wire _21673_;
  wire _21674_;
  wire _21675_;
  wire _21676_;
  wire _21677_;
  wire _21678_;
  wire _21679_;
  wire _21680_;
  wire _21681_;
  wire _21682_;
  wire _21683_;
  wire _21684_;
  wire _21685_;
  wire _21686_;
  wire _21687_;
  wire _21688_;
  wire _21689_;
  wire _21690_;
  wire _21691_;
  wire _21692_;
  wire _21693_;
  wire _21694_;
  wire _21695_;
  wire _21696_;
  wire _21697_;
  wire _21698_;
  wire _21699_;
  wire _21700_;
  wire _21701_;
  wire _21702_;
  wire _21703_;
  wire _21704_;
  wire _21705_;
  wire _21706_;
  wire _21707_;
  wire _21708_;
  wire _21709_;
  wire _21710_;
  wire _21711_;
  wire _21712_;
  wire _21713_;
  wire _21714_;
  wire _21715_;
  wire _21716_;
  wire _21717_;
  wire _21718_;
  wire _21719_;
  wire _21720_;
  wire _21721_;
  wire _21722_;
  wire _21723_;
  wire _21724_;
  wire _21725_;
  wire _21726_;
  wire _21727_;
  wire _21728_;
  wire _21729_;
  wire _21730_;
  wire _21731_;
  wire _21732_;
  wire _21733_;
  wire _21734_;
  wire _21735_;
  wire _21736_;
  wire _21737_;
  wire _21738_;
  wire _21739_;
  wire _21740_;
  wire _21741_;
  wire _21742_;
  wire _21743_;
  wire _21744_;
  wire _21745_;
  wire _21746_;
  wire _21747_;
  wire _21748_;
  wire _21749_;
  wire _21750_;
  wire _21751_;
  wire _21752_;
  wire _21753_;
  wire _21754_;
  wire _21755_;
  wire _21756_;
  wire _21757_;
  wire _21758_;
  wire _21759_;
  wire _21760_;
  wire _21761_;
  wire _21762_;
  wire _21763_;
  wire _21764_;
  wire _21765_;
  wire _21766_;
  wire _21767_;
  wire _21768_;
  wire _21769_;
  wire _21770_;
  wire _21771_;
  wire _21772_;
  wire _21773_;
  wire _21774_;
  wire _21775_;
  wire _21776_;
  wire _21777_;
  wire _21778_;
  wire _21779_;
  wire _21780_;
  wire _21781_;
  wire _21782_;
  wire _21783_;
  wire _21784_;
  wire _21785_;
  wire _21786_;
  wire _21787_;
  wire _21788_;
  wire _21789_;
  wire _21790_;
  wire _21791_;
  wire _21792_;
  wire _21793_;
  wire _21794_;
  wire _21795_;
  wire _21796_;
  wire _21797_;
  wire _21798_;
  wire _21799_;
  wire _21800_;
  wire _21801_;
  wire _21802_;
  wire _21803_;
  wire _21804_;
  wire _21805_;
  wire _21806_;
  wire _21807_;
  wire _21808_;
  wire _21809_;
  wire _21810_;
  wire _21811_;
  wire _21812_;
  wire _21813_;
  wire _21814_;
  wire _21815_;
  wire _21816_;
  wire _21817_;
  wire _21818_;
  wire _21819_;
  wire _21820_;
  wire _21821_;
  wire _21822_;
  wire _21823_;
  wire _21824_;
  wire _21825_;
  wire _21826_;
  wire _21827_;
  wire _21828_;
  wire _21829_;
  wire _21830_;
  wire _21831_;
  wire _21832_;
  wire _21833_;
  wire _21834_;
  wire _21835_;
  wire _21836_;
  wire _21837_;
  wire _21838_;
  wire _21839_;
  wire _21840_;
  wire _21841_;
  wire _21842_;
  wire _21843_;
  wire _21844_;
  wire _21845_;
  wire _21846_;
  wire _21847_;
  wire _21848_;
  wire _21849_;
  wire _21850_;
  wire _21851_;
  wire _21852_;
  wire _21853_;
  wire _21854_;
  wire _21855_;
  wire _21856_;
  wire _21857_;
  wire _21858_;
  wire _21859_;
  wire _21860_;
  wire _21861_;
  wire _21862_;
  wire _21863_;
  wire _21864_;
  wire _21865_;
  wire _21866_;
  wire _21867_;
  wire _21868_;
  wire _21869_;
  wire _21870_;
  wire _21871_;
  wire _21872_;
  wire _21873_;
  wire _21874_;
  wire _21875_;
  wire _21876_;
  wire _21877_;
  wire _21878_;
  wire _21879_;
  wire _21880_;
  wire _21881_;
  wire _21882_;
  wire _21883_;
  wire _21884_;
  wire _21885_;
  wire _21886_;
  wire _21887_;
  wire _21888_;
  wire _21889_;
  wire _21890_;
  wire _21891_;
  wire _21892_;
  wire _21893_;
  wire _21894_;
  wire _21895_;
  wire _21896_;
  wire _21897_;
  wire _21898_;
  wire _21899_;
  wire _21900_;
  wire _21901_;
  wire _21902_;
  wire _21903_;
  wire _21904_;
  wire _21905_;
  wire _21906_;
  wire _21907_;
  wire _21908_;
  wire _21909_;
  wire _21910_;
  wire _21911_;
  wire _21912_;
  wire _21913_;
  wire _21914_;
  wire _21915_;
  wire _21916_;
  wire _21917_;
  wire _21918_;
  wire _21919_;
  wire _21920_;
  wire _21921_;
  wire _21922_;
  wire _21923_;
  wire _21924_;
  wire _21925_;
  wire _21926_;
  wire _21927_;
  wire _21928_;
  wire _21929_;
  wire _21930_;
  wire _21931_;
  wire _21932_;
  wire _21933_;
  wire _21934_;
  wire _21935_;
  wire _21936_;
  wire _21937_;
  wire _21938_;
  wire _21939_;
  wire _21940_;
  wire _21941_;
  wire _21942_;
  wire _21943_;
  wire _21944_;
  wire _21945_;
  wire _21946_;
  wire _21947_;
  wire _21948_;
  wire _21949_;
  wire _21950_;
  wire _21951_;
  wire _21952_;
  wire _21953_;
  wire _21954_;
  wire _21955_;
  wire _21956_;
  wire _21957_;
  wire _21958_;
  wire _21959_;
  wire _21960_;
  wire _21961_;
  wire _21962_;
  wire _21963_;
  wire _21964_;
  wire _21965_;
  wire _21966_;
  wire _21967_;
  wire _21968_;
  wire _21969_;
  wire _21970_;
  wire _21971_;
  wire _21972_;
  wire _21973_;
  wire _21974_;
  wire _21975_;
  wire _21976_;
  wire _21977_;
  wire _21978_;
  wire _21979_;
  wire _21980_;
  wire _21981_;
  wire _21982_;
  wire _21983_;
  wire _21984_;
  wire _21985_;
  wire _21986_;
  wire _21987_;
  wire _21988_;
  wire _21989_;
  wire _21990_;
  wire _21991_;
  wire _21992_;
  wire _21993_;
  wire _21994_;
  wire _21995_;
  wire _21996_;
  wire _21997_;
  wire _21998_;
  wire _21999_;
  wire _22000_;
  wire _22001_;
  wire _22002_;
  wire _22003_;
  wire _22004_;
  wire _22005_;
  wire _22006_;
  wire _22007_;
  wire _22008_;
  wire _22009_;
  wire _22010_;
  wire _22011_;
  wire _22012_;
  wire _22013_;
  wire _22014_;
  wire _22015_;
  wire _22016_;
  wire _22017_;
  wire _22018_;
  wire _22019_;
  wire _22020_;
  wire _22021_;
  wire _22022_;
  wire _22023_;
  wire _22024_;
  wire _22025_;
  wire _22026_;
  wire _22027_;
  wire _22028_;
  wire _22029_;
  wire _22030_;
  wire _22031_;
  wire _22032_;
  wire _22033_;
  wire _22034_;
  wire _22035_;
  wire _22036_;
  wire _22037_;
  wire _22038_;
  wire _22039_;
  wire _22040_;
  wire _22041_;
  wire _22042_;
  wire _22043_;
  wire _22044_;
  wire _22045_;
  wire _22046_;
  wire _22047_;
  wire _22048_;
  wire _22049_;
  wire _22050_;
  wire _22051_;
  wire _22052_;
  wire _22053_;
  wire _22054_;
  wire _22055_;
  wire _22056_;
  wire _22057_;
  wire _22058_;
  wire _22059_;
  wire _22060_;
  wire _22061_;
  wire _22062_;
  wire _22063_;
  wire _22064_;
  wire _22065_;
  wire _22066_;
  wire _22067_;
  wire _22068_;
  wire _22069_;
  wire _22070_;
  wire _22071_;
  wire _22072_;
  wire _22073_;
  wire _22074_;
  wire _22075_;
  wire _22076_;
  wire _22077_;
  wire _22078_;
  wire _22079_;
  wire _22080_;
  wire _22081_;
  wire _22082_;
  wire _22083_;
  wire _22084_;
  wire _22085_;
  wire _22086_;
  wire _22087_;
  wire _22088_;
  wire _22089_;
  wire _22090_;
  wire _22091_;
  wire _22092_;
  wire _22093_;
  wire _22094_;
  wire _22095_;
  wire _22096_;
  wire _22097_;
  wire _22098_;
  wire _22099_;
  wire _22100_;
  wire _22101_;
  wire _22102_;
  wire _22103_;
  wire _22104_;
  wire _22105_;
  wire _22106_;
  wire _22107_;
  wire _22108_;
  wire _22109_;
  wire _22110_;
  wire _22111_;
  wire _22112_;
  wire _22113_;
  wire _22114_;
  wire _22115_;
  wire _22116_;
  wire _22117_;
  wire _22118_;
  wire _22119_;
  wire _22120_;
  wire _22121_;
  wire _22122_;
  wire _22123_;
  wire _22124_;
  wire _22125_;
  wire _22126_;
  wire _22127_;
  wire _22128_;
  wire _22129_;
  wire _22130_;
  wire _22131_;
  wire _22132_;
  wire _22133_;
  wire _22134_;
  wire _22135_;
  wire _22136_;
  wire _22137_;
  wire _22138_;
  wire _22139_;
  wire _22140_;
  wire _22141_;
  wire _22142_;
  wire _22143_;
  wire _22144_;
  wire _22145_;
  wire _22146_;
  wire _22147_;
  wire _22148_;
  wire _22149_;
  wire _22150_;
  wire _22151_;
  wire _22152_;
  wire _22153_;
  wire _22154_;
  wire _22155_;
  wire _22156_;
  wire _22157_;
  wire _22158_;
  wire _22159_;
  wire _22160_;
  wire _22161_;
  wire _22162_;
  wire _22163_;
  wire _22164_;
  wire _22165_;
  wire _22166_;
  wire _22167_;
  wire _22168_;
  wire _22169_;
  wire _22170_;
  wire _22171_;
  wire _22172_;
  wire _22173_;
  wire _22174_;
  wire _22175_;
  wire _22176_;
  wire _22177_;
  wire _22178_;
  wire _22179_;
  wire _22180_;
  wire _22181_;
  wire _22182_;
  wire _22183_;
  wire _22184_;
  wire _22185_;
  wire _22186_;
  wire _22187_;
  wire _22188_;
  wire _22189_;
  wire _22190_;
  wire _22191_;
  wire _22192_;
  wire _22193_;
  wire _22194_;
  wire _22195_;
  wire _22196_;
  wire _22197_;
  wire _22198_;
  wire _22199_;
  wire _22200_;
  wire _22201_;
  wire _22202_;
  wire _22203_;
  wire _22204_;
  wire _22205_;
  wire _22206_;
  wire _22207_;
  wire _22208_;
  wire _22209_;
  wire _22210_;
  wire _22211_;
  wire _22212_;
  wire _22213_;
  wire _22214_;
  wire _22215_;
  wire _22216_;
  wire _22217_;
  wire _22218_;
  wire _22219_;
  wire _22220_;
  wire _22221_;
  wire _22222_;
  wire _22223_;
  wire _22224_;
  wire _22225_;
  wire _22226_;
  wire _22227_;
  wire _22228_;
  wire _22229_;
  wire _22230_;
  wire _22231_;
  wire _22232_;
  wire _22233_;
  wire _22234_;
  wire _22235_;
  wire _22236_;
  wire _22237_;
  wire _22238_;
  wire _22239_;
  wire _22240_;
  wire _22241_;
  wire _22242_;
  wire _22243_;
  wire _22244_;
  wire _22245_;
  wire _22246_;
  wire _22247_;
  wire _22248_;
  wire _22249_;
  wire _22250_;
  wire _22251_;
  wire _22252_;
  wire _22253_;
  wire _22254_;
  wire _22255_;
  wire _22256_;
  wire _22257_;
  wire _22258_;
  wire _22259_;
  wire _22260_;
  wire _22261_;
  wire _22262_;
  wire _22263_;
  wire _22264_;
  wire _22265_;
  wire _22266_;
  wire _22267_;
  wire _22268_;
  wire _22269_;
  wire _22270_;
  wire _22271_;
  wire _22272_;
  wire _22273_;
  wire _22274_;
  wire _22275_;
  wire _22276_;
  wire _22277_;
  wire _22278_;
  wire _22279_;
  wire _22280_;
  wire _22281_;
  wire _22282_;
  wire _22283_;
  wire _22284_;
  wire _22285_;
  wire _22286_;
  wire _22287_;
  wire _22288_;
  wire _22289_;
  wire _22290_;
  wire _22291_;
  wire _22292_;
  wire _22293_;
  wire _22294_;
  wire _22295_;
  wire _22296_;
  wire _22297_;
  wire _22298_;
  wire _22299_;
  wire _22300_;
  wire _22301_;
  wire _22302_;
  wire _22303_;
  wire _22304_;
  wire _22305_;
  wire _22306_;
  wire _22307_;
  wire _22308_;
  wire _22309_;
  wire _22310_;
  wire _22311_;
  wire _22312_;
  wire _22313_;
  wire _22314_;
  wire _22315_;
  wire _22316_;
  wire _22317_;
  wire _22318_;
  wire _22319_;
  wire _22320_;
  wire _22321_;
  wire _22322_;
  wire _22323_;
  wire _22324_;
  wire _22325_;
  wire _22326_;
  wire _22327_;
  wire _22328_;
  wire _22329_;
  wire _22330_;
  wire _22331_;
  wire _22332_;
  wire _22333_;
  wire _22334_;
  wire _22335_;
  wire _22336_;
  wire _22337_;
  wire _22338_;
  wire _22339_;
  wire _22340_;
  wire _22341_;
  wire _22342_;
  wire _22343_;
  wire _22344_;
  wire _22345_;
  wire _22346_;
  wire _22347_;
  wire _22348_;
  wire _22349_;
  wire _22350_;
  wire _22351_;
  wire _22352_;
  wire _22353_;
  wire _22354_;
  wire _22355_;
  wire _22356_;
  wire _22357_;
  wire _22358_;
  wire _22359_;
  wire _22360_;
  wire _22361_;
  wire _22362_;
  wire _22363_;
  wire _22364_;
  wire _22365_;
  wire _22366_;
  wire _22367_;
  wire _22368_;
  wire _22369_;
  wire _22370_;
  wire _22371_;
  wire _22372_;
  wire _22373_;
  wire _22374_;
  wire _22375_;
  wire _22376_;
  wire _22377_;
  wire _22378_;
  wire _22379_;
  wire _22380_;
  wire _22381_;
  wire _22382_;
  wire _22383_;
  wire _22384_;
  wire _22385_;
  wire _22386_;
  wire _22387_;
  wire _22388_;
  wire _22389_;
  wire _22390_;
  wire _22391_;
  wire _22392_;
  wire _22393_;
  wire _22394_;
  wire _22395_;
  wire _22396_;
  wire _22397_;
  wire _22398_;
  wire _22399_;
  wire _22400_;
  wire _22401_;
  wire _22402_;
  wire _22403_;
  wire _22404_;
  wire _22405_;
  wire _22406_;
  wire _22407_;
  wire _22408_;
  wire _22409_;
  wire _22410_;
  wire _22411_;
  wire _22412_;
  wire _22413_;
  wire _22414_;
  wire _22415_;
  wire _22416_;
  wire _22417_;
  wire _22418_;
  wire _22419_;
  wire _22420_;
  wire _22421_;
  wire _22422_;
  wire _22423_;
  wire _22424_;
  wire _22425_;
  wire _22426_;
  wire _22427_;
  wire _22428_;
  wire _22429_;
  wire _22430_;
  wire _22431_;
  wire _22432_;
  wire _22433_;
  wire _22434_;
  wire _22435_;
  wire _22436_;
  wire _22437_;
  wire _22438_;
  wire _22439_;
  wire _22440_;
  wire _22441_;
  wire _22442_;
  wire _22443_;
  wire _22444_;
  wire _22445_;
  wire _22446_;
  wire _22447_;
  wire _22448_;
  wire _22449_;
  wire _22450_;
  wire _22451_;
  wire _22452_;
  wire _22453_;
  wire _22454_;
  wire _22455_;
  wire _22456_;
  wire _22457_;
  wire _22458_;
  wire _22459_;
  wire _22460_;
  wire _22461_;
  wire _22462_;
  wire _22463_;
  wire _22464_;
  wire _22465_;
  wire _22466_;
  wire _22467_;
  wire _22468_;
  wire _22469_;
  wire _22470_;
  wire _22471_;
  wire _22472_;
  wire _22473_;
  wire _22474_;
  wire _22475_;
  wire _22476_;
  wire _22477_;
  wire _22478_;
  wire _22479_;
  wire _22480_;
  wire _22481_;
  wire _22482_;
  wire _22483_;
  wire _22484_;
  wire _22485_;
  wire _22486_;
  wire _22487_;
  wire _22488_;
  wire _22489_;
  wire _22490_;
  wire _22491_;
  wire _22492_;
  wire _22493_;
  wire _22494_;
  wire _22495_;
  wire _22496_;
  wire _22497_;
  wire _22498_;
  wire _22499_;
  wire _22500_;
  wire _22501_;
  wire _22502_;
  wire _22503_;
  wire _22504_;
  wire _22505_;
  wire _22506_;
  wire _22507_;
  wire _22508_;
  wire _22509_;
  wire _22510_;
  wire _22511_;
  wire _22512_;
  wire _22513_;
  wire _22514_;
  wire _22515_;
  wire _22516_;
  wire _22517_;
  wire _22518_;
  wire _22519_;
  wire _22520_;
  wire _22521_;
  wire _22522_;
  wire _22523_;
  wire _22524_;
  wire _22525_;
  wire _22526_;
  wire _22527_;
  wire _22528_;
  wire _22529_;
  wire _22530_;
  wire _22531_;
  wire _22532_;
  wire _22533_;
  wire _22534_;
  wire _22535_;
  wire _22536_;
  wire _22537_;
  wire _22538_;
  wire _22539_;
  wire _22540_;
  wire _22541_;
  wire _22542_;
  wire _22543_;
  wire _22544_;
  wire _22545_;
  wire _22546_;
  wire _22547_;
  wire _22548_;
  wire _22549_;
  wire _22550_;
  wire _22551_;
  wire _22552_;
  wire _22553_;
  wire _22554_;
  wire _22555_;
  wire _22556_;
  wire _22557_;
  wire _22558_;
  wire _22559_;
  wire _22560_;
  wire _22561_;
  wire _22562_;
  wire _22563_;
  wire _22564_;
  wire _22565_;
  wire _22566_;
  wire _22567_;
  wire _22568_;
  wire _22569_;
  wire _22570_;
  wire _22571_;
  wire _22572_;
  wire _22573_;
  wire _22574_;
  wire _22575_;
  wire _22576_;
  wire _22577_;
  wire _22578_;
  wire _22579_;
  wire _22580_;
  wire _22581_;
  wire _22582_;
  wire _22583_;
  wire _22584_;
  wire _22585_;
  wire _22586_;
  wire _22587_;
  wire _22588_;
  wire _22589_;
  wire _22590_;
  wire _22591_;
  wire _22592_;
  wire _22593_;
  wire _22594_;
  wire _22595_;
  wire _22596_;
  wire _22597_;
  wire _22598_;
  wire _22599_;
  wire _22600_;
  wire _22601_;
  wire _22602_;
  wire _22603_;
  wire _22604_;
  wire _22605_;
  wire _22606_;
  wire _22607_;
  wire _22608_;
  wire _22609_;
  wire _22610_;
  wire _22611_;
  wire _22612_;
  wire _22613_;
  wire _22614_;
  wire _22615_;
  wire _22616_;
  wire _22617_;
  wire _22618_;
  wire _22619_;
  wire _22620_;
  wire _22621_;
  wire _22622_;
  wire _22623_;
  wire _22624_;
  wire _22625_;
  wire _22626_;
  wire _22627_;
  wire _22628_;
  wire _22629_;
  wire _22630_;
  wire _22631_;
  wire _22632_;
  wire _22633_;
  wire _22634_;
  wire _22635_;
  wire _22636_;
  wire _22637_;
  wire _22638_;
  wire _22639_;
  wire _22640_;
  wire _22641_;
  wire _22642_;
  wire _22643_;
  wire _22644_;
  wire _22645_;
  wire _22646_;
  wire _22647_;
  wire _22648_;
  wire _22649_;
  wire _22650_;
  wire _22651_;
  wire _22652_;
  wire _22653_;
  wire _22654_;
  wire _22655_;
  wire _22656_;
  wire _22657_;
  wire _22658_;
  wire _22659_;
  wire _22660_;
  wire _22661_;
  wire _22662_;
  wire _22663_;
  wire _22664_;
  wire _22665_;
  wire _22666_;
  wire _22667_;
  wire _22668_;
  wire _22669_;
  wire _22670_;
  wire _22671_;
  wire _22672_;
  wire _22673_;
  wire _22674_;
  wire _22675_;
  wire _22676_;
  wire _22677_;
  wire _22678_;
  wire _22679_;
  wire _22680_;
  wire _22681_;
  wire _22682_;
  wire _22683_;
  wire _22684_;
  wire _22685_;
  wire _22686_;
  wire _22687_;
  wire _22688_;
  wire _22689_;
  wire _22690_;
  wire _22691_;
  wire _22692_;
  wire _22693_;
  wire _22694_;
  wire _22695_;
  wire _22696_;
  wire _22697_;
  wire _22698_;
  wire _22699_;
  wire _22700_;
  wire _22701_;
  wire _22702_;
  wire _22703_;
  wire _22704_;
  wire _22705_;
  wire _22706_;
  wire _22707_;
  wire _22708_;
  wire _22709_;
  wire _22710_;
  wire _22711_;
  wire _22712_;
  wire _22713_;
  wire _22714_;
  wire _22715_;
  wire _22716_;
  wire _22717_;
  wire _22718_;
  wire _22719_;
  wire _22720_;
  wire _22721_;
  wire _22722_;
  wire _22723_;
  wire _22724_;
  wire _22725_;
  wire _22726_;
  wire _22727_;
  wire _22728_;
  wire _22729_;
  wire _22730_;
  wire _22731_;
  wire _22732_;
  wire _22733_;
  wire _22734_;
  wire _22735_;
  wire _22736_;
  wire _22737_;
  wire _22738_;
  wire _22739_;
  wire _22740_;
  wire _22741_;
  wire _22742_;
  wire _22743_;
  wire _22744_;
  wire _22745_;
  wire _22746_;
  wire _22747_;
  wire _22748_;
  wire _22749_;
  wire _22750_;
  wire _22751_;
  wire _22752_;
  wire _22753_;
  wire _22754_;
  wire _22755_;
  wire _22756_;
  wire _22757_;
  wire _22758_;
  wire _22759_;
  wire _22760_;
  wire _22761_;
  wire _22762_;
  wire _22763_;
  wire _22764_;
  wire _22765_;
  wire _22766_;
  wire _22767_;
  wire _22768_;
  wire _22769_;
  wire _22770_;
  wire _22771_;
  wire _22772_;
  wire _22773_;
  wire _22774_;
  wire _22775_;
  wire _22776_;
  wire _22777_;
  wire _22778_;
  wire _22779_;
  wire _22780_;
  wire _22781_;
  wire _22782_;
  wire _22783_;
  wire _22784_;
  wire _22785_;
  wire _22786_;
  wire _22787_;
  wire _22788_;
  wire _22789_;
  wire _22790_;
  wire _22791_;
  wire _22792_;
  wire _22793_;
  wire _22794_;
  wire _22795_;
  wire _22796_;
  wire _22797_;
  wire _22798_;
  wire _22799_;
  wire _22800_;
  wire _22801_;
  wire _22802_;
  wire _22803_;
  wire _22804_;
  wire _22805_;
  wire _22806_;
  wire _22807_;
  wire _22808_;
  wire _22809_;
  wire _22810_;
  wire _22811_;
  wire _22812_;
  wire _22813_;
  wire _22814_;
  wire _22815_;
  wire _22816_;
  wire _22817_;
  wire _22818_;
  wire _22819_;
  wire _22820_;
  wire _22821_;
  wire _22822_;
  wire _22823_;
  wire _22824_;
  wire _22825_;
  wire _22826_;
  wire _22827_;
  wire _22828_;
  wire _22829_;
  wire _22830_;
  wire _22831_;
  wire _22832_;
  wire _22833_;
  wire _22834_;
  wire _22835_;
  wire _22836_;
  wire _22837_;
  wire _22838_;
  wire _22839_;
  wire _22840_;
  wire _22841_;
  wire _22842_;
  wire _22843_;
  wire _22844_;
  wire _22845_;
  wire _22846_;
  wire _22847_;
  wire _22848_;
  wire _22849_;
  wire _22850_;
  wire _22851_;
  wire _22852_;
  wire _22853_;
  wire _22854_;
  wire _22855_;
  wire _22856_;
  wire _22857_;
  wire _22858_;
  wire _22859_;
  wire _22860_;
  wire _22861_;
  wire _22862_;
  wire _22863_;
  wire _22864_;
  wire _22865_;
  wire _22866_;
  wire _22867_;
  wire _22868_;
  wire _22869_;
  wire _22870_;
  wire _22871_;
  wire _22872_;
  wire _22873_;
  wire _22874_;
  wire _22875_;
  wire _22876_;
  wire _22877_;
  wire _22878_;
  wire _22879_;
  wire _22880_;
  wire _22881_;
  wire _22882_;
  wire _22883_;
  wire _22884_;
  wire _22885_;
  wire _22886_;
  wire _22887_;
  wire _22888_;
  wire _22889_;
  wire _22890_;
  wire _22891_;
  wire _22892_;
  wire _22893_;
  wire _22894_;
  wire _22895_;
  wire _22896_;
  wire _22897_;
  wire _22898_;
  wire _22899_;
  wire _22900_;
  wire _22901_;
  wire _22902_;
  wire _22903_;
  wire _22904_;
  wire _22905_;
  wire _22906_;
  wire _22907_;
  wire _22908_;
  wire _22909_;
  wire _22910_;
  wire _22911_;
  wire _22912_;
  wire _22913_;
  wire _22914_;
  wire _22915_;
  wire _22916_;
  wire _22917_;
  wire _22918_;
  wire _22919_;
  wire _22920_;
  wire _22921_;
  wire _22922_;
  wire _22923_;
  wire _22924_;
  wire _22925_;
  wire _22926_;
  wire _22927_;
  wire _22928_;
  wire _22929_;
  wire _22930_;
  wire _22931_;
  wire _22932_;
  wire _22933_;
  wire _22934_;
  wire _22935_;
  wire _22936_;
  wire _22937_;
  wire _22938_;
  wire _22939_;
  wire _22940_;
  wire _22941_;
  wire _22942_;
  wire _22943_;
  wire _22944_;
  wire _22945_;
  wire _22946_;
  wire _22947_;
  wire _22948_;
  wire _22949_;
  wire _22950_;
  wire _22951_;
  wire _22952_;
  wire _22953_;
  wire _22954_;
  wire _22955_;
  wire _22956_;
  wire _22957_;
  wire _22958_;
  wire _22959_;
  wire _22960_;
  wire _22961_;
  wire _22962_;
  wire _22963_;
  wire _22964_;
  wire _22965_;
  wire _22966_;
  wire _22967_;
  wire _22968_;
  wire _22969_;
  wire _22970_;
  wire _22971_;
  wire _22972_;
  wire _22973_;
  wire _22974_;
  wire _22975_;
  wire _22976_;
  wire _22977_;
  wire _22978_;
  wire _22979_;
  wire _22980_;
  wire _22981_;
  wire _22982_;
  wire _22983_;
  wire _22984_;
  wire _22985_;
  wire _22986_;
  wire _22987_;
  wire _22988_;
  wire _22989_;
  wire _22990_;
  wire _22991_;
  wire _22992_;
  wire _22993_;
  wire _22994_;
  wire _22995_;
  wire _22996_;
  wire _22997_;
  wire _22998_;
  wire _22999_;
  wire _23000_;
  wire _23001_;
  wire _23002_;
  wire _23003_;
  wire _23004_;
  wire _23005_;
  wire _23006_;
  wire _23007_;
  wire _23008_;
  wire _23009_;
  wire _23010_;
  wire _23011_;
  wire _23012_;
  wire _23013_;
  wire _23014_;
  wire _23015_;
  wire _23016_;
  wire _23017_;
  wire _23018_;
  wire _23019_;
  wire _23020_;
  wire _23021_;
  wire _23022_;
  wire _23023_;
  wire _23024_;
  wire _23025_;
  wire _23026_;
  wire _23027_;
  wire _23028_;
  wire _23029_;
  wire _23030_;
  wire _23031_;
  wire _23032_;
  wire _23033_;
  wire _23034_;
  wire _23035_;
  wire _23036_;
  wire _23037_;
  wire _23038_;
  wire _23039_;
  wire _23040_;
  wire _23041_;
  wire _23042_;
  wire _23043_;
  wire _23044_;
  wire _23045_;
  wire _23046_;
  wire _23047_;
  wire _23048_;
  wire _23049_;
  wire _23050_;
  wire _23051_;
  wire _23052_;
  wire _23053_;
  wire _23054_;
  wire _23055_;
  wire _23056_;
  wire _23057_;
  wire _23058_;
  wire _23059_;
  wire _23060_;
  wire _23061_;
  wire _23062_;
  wire _23063_;
  wire _23064_;
  wire _23065_;
  wire _23066_;
  wire _23067_;
  wire _23068_;
  wire _23069_;
  wire _23070_;
  wire _23071_;
  wire _23072_;
  wire _23073_;
  wire _23074_;
  wire _23075_;
  wire _23076_;
  wire _23077_;
  wire _23078_;
  wire _23079_;
  wire _23080_;
  wire _23081_;
  wire _23082_;
  wire _23083_;
  wire _23084_;
  wire _23085_;
  wire _23086_;
  wire _23087_;
  wire _23088_;
  wire _23089_;
  wire _23090_;
  wire _23091_;
  wire _23092_;
  wire _23093_;
  wire _23094_;
  wire _23095_;
  wire _23096_;
  wire _23097_;
  wire _23098_;
  wire _23099_;
  wire _23100_;
  wire _23101_;
  wire _23102_;
  wire _23103_;
  wire _23104_;
  wire _23105_;
  wire _23106_;
  wire _23107_;
  wire _23108_;
  wire _23109_;
  wire _23110_;
  wire _23111_;
  wire _23112_;
  wire _23113_;
  wire _23114_;
  wire _23115_;
  wire _23116_;
  wire _23117_;
  wire _23118_;
  wire _23119_;
  wire _23120_;
  wire _23121_;
  wire _23122_;
  wire _23123_;
  wire _23124_;
  wire _23125_;
  wire _23126_;
  wire _23127_;
  wire _23128_;
  wire _23129_;
  wire _23130_;
  wire _23131_;
  wire _23132_;
  wire _23133_;
  wire _23134_;
  wire _23135_;
  wire _23136_;
  wire _23137_;
  wire _23138_;
  wire _23139_;
  wire _23140_;
  wire _23141_;
  wire _23142_;
  wire _23143_;
  wire _23144_;
  wire _23145_;
  wire _23146_;
  wire _23147_;
  wire _23148_;
  wire _23149_;
  wire _23150_;
  wire _23151_;
  wire _23152_;
  wire _23153_;
  wire _23154_;
  wire _23155_;
  wire _23156_;
  wire _23157_;
  wire _23158_;
  wire _23159_;
  wire _23160_;
  wire _23161_;
  wire _23162_;
  wire _23163_;
  wire _23164_;
  wire _23165_;
  wire _23166_;
  wire _23167_;
  wire _23168_;
  wire _23169_;
  wire _23170_;
  wire _23171_;
  wire _23172_;
  wire _23173_;
  wire _23174_;
  wire _23175_;
  wire _23176_;
  wire _23177_;
  wire _23178_;
  wire _23179_;
  wire _23180_;
  wire _23181_;
  wire _23182_;
  wire _23183_;
  wire _23184_;
  wire _23185_;
  wire _23186_;
  wire _23187_;
  wire _23188_;
  wire _23189_;
  wire _23190_;
  wire _23191_;
  wire _23192_;
  wire _23193_;
  wire _23194_;
  wire _23195_;
  wire _23196_;
  wire _23197_;
  wire _23198_;
  wire _23199_;
  wire _23200_;
  wire _23201_;
  wire _23202_;
  wire _23203_;
  wire _23204_;
  wire _23205_;
  wire _23206_;
  wire _23207_;
  wire _23208_;
  wire _23209_;
  wire _23210_;
  wire _23211_;
  wire _23212_;
  wire _23213_;
  wire _23214_;
  wire _23215_;
  wire _23216_;
  wire _23217_;
  wire _23218_;
  wire _23219_;
  wire _23220_;
  wire _23221_;
  wire _23222_;
  wire _23223_;
  wire _23224_;
  wire _23225_;
  wire _23226_;
  wire _23227_;
  wire _23228_;
  wire _23229_;
  wire _23230_;
  wire _23231_;
  wire _23232_;
  wire _23233_;
  wire _23234_;
  wire _23235_;
  wire _23236_;
  wire _23237_;
  wire _23238_;
  wire _23239_;
  wire _23240_;
  wire _23241_;
  wire _23242_;
  wire _23243_;
  wire _23244_;
  wire _23245_;
  wire _23246_;
  wire _23247_;
  wire _23248_;
  wire _23249_;
  wire _23250_;
  wire _23251_;
  wire _23252_;
  wire _23253_;
  wire _23254_;
  wire _23255_;
  wire _23256_;
  wire _23257_;
  wire _23258_;
  wire _23259_;
  wire _23260_;
  wire _23261_;
  wire _23262_;
  wire _23263_;
  wire _23264_;
  wire _23265_;
  wire _23266_;
  wire _23267_;
  wire _23268_;
  wire _23269_;
  wire _23270_;
  wire _23271_;
  wire _23272_;
  wire _23273_;
  wire _23274_;
  wire _23275_;
  wire _23276_;
  wire _23277_;
  wire _23278_;
  wire _23279_;
  wire _23280_;
  wire _23281_;
  wire _23282_;
  wire _23283_;
  wire _23284_;
  wire _23285_;
  wire _23286_;
  wire _23287_;
  wire _23288_;
  wire _23289_;
  wire _23290_;
  wire _23291_;
  wire _23292_;
  wire _23293_;
  wire _23294_;
  wire _23295_;
  wire _23296_;
  wire _23297_;
  wire _23298_;
  wire _23299_;
  wire _23300_;
  wire _23301_;
  wire _23302_;
  wire _23303_;
  wire _23304_;
  wire _23305_;
  wire _23306_;
  wire _23307_;
  wire _23308_;
  wire _23309_;
  wire _23310_;
  wire _23311_;
  wire _23312_;
  wire _23313_;
  wire _23314_;
  wire _23315_;
  wire _23316_;
  wire _23317_;
  wire _23318_;
  wire _23319_;
  wire _23320_;
  wire _23321_;
  wire _23322_;
  wire _23323_;
  wire _23324_;
  wire _23325_;
  wire _23326_;
  wire _23327_;
  wire _23328_;
  wire _23329_;
  wire _23330_;
  wire _23331_;
  wire _23332_;
  wire _23333_;
  wire _23334_;
  wire _23335_;
  wire _23336_;
  wire _23337_;
  wire _23338_;
  wire _23339_;
  wire _23340_;
  wire _23341_;
  wire _23342_;
  wire _23343_;
  wire _23344_;
  wire _23345_;
  wire _23346_;
  wire _23347_;
  wire _23348_;
  wire _23349_;
  wire _23350_;
  wire _23351_;
  wire _23352_;
  wire _23353_;
  wire _23354_;
  wire _23355_;
  wire _23356_;
  wire _23357_;
  wire _23358_;
  wire _23359_;
  wire _23360_;
  wire _23361_;
  wire _23362_;
  wire _23363_;
  wire _23364_;
  wire _23365_;
  wire _23366_;
  wire _23367_;
  wire _23368_;
  wire _23369_;
  wire _23370_;
  wire _23371_;
  wire _23372_;
  wire _23373_;
  wire _23374_;
  wire _23375_;
  wire _23376_;
  wire _23377_;
  wire _23378_;
  wire _23379_;
  wire _23380_;
  wire _23381_;
  wire _23382_;
  wire _23383_;
  wire _23384_;
  wire _23385_;
  wire _23386_;
  wire _23387_;
  wire _23388_;
  wire _23389_;
  wire _23390_;
  wire _23391_;
  wire _23392_;
  wire _23393_;
  wire _23394_;
  wire _23395_;
  wire _23396_;
  wire _23397_;
  wire _23398_;
  wire _23399_;
  wire _23400_;
  wire _23401_;
  wire _23402_;
  wire _23403_;
  wire _23404_;
  wire _23405_;
  wire _23406_;
  wire _23407_;
  wire _23408_;
  wire _23409_;
  wire _23410_;
  wire _23411_;
  wire _23412_;
  wire _23413_;
  wire _23414_;
  wire _23415_;
  wire _23416_;
  wire _23417_;
  wire _23418_;
  wire _23419_;
  wire _23420_;
  wire _23421_;
  wire _23422_;
  wire _23423_;
  wire _23424_;
  wire _23425_;
  wire _23426_;
  wire _23427_;
  wire _23428_;
  wire _23429_;
  wire _23430_;
  wire _23431_;
  wire _23432_;
  wire _23433_;
  wire _23434_;
  wire _23435_;
  wire _23436_;
  wire _23437_;
  wire _23438_;
  wire _23439_;
  wire _23440_;
  wire _23441_;
  wire _23442_;
  wire _23443_;
  wire _23444_;
  wire _23445_;
  wire _23446_;
  wire _23447_;
  wire _23448_;
  wire _23449_;
  wire _23450_;
  wire _23451_;
  wire _23452_;
  wire _23453_;
  wire _23454_;
  wire _23455_;
  wire _23456_;
  wire _23457_;
  wire _23458_;
  wire _23459_;
  wire _23460_;
  wire _23461_;
  wire _23462_;
  wire _23463_;
  wire _23464_;
  wire _23465_;
  wire _23466_;
  wire _23467_;
  wire _23468_;
  wire _23469_;
  wire _23470_;
  wire _23471_;
  wire _23472_;
  wire _23473_;
  wire _23474_;
  wire _23475_;
  wire _23476_;
  wire _23477_;
  wire _23478_;
  wire _23479_;
  wire _23480_;
  wire _23481_;
  wire _23482_;
  wire _23483_;
  wire _23484_;
  wire _23485_;
  wire _23486_;
  wire _23487_;
  wire _23488_;
  wire _23489_;
  wire _23490_;
  wire _23491_;
  wire _23492_;
  wire _23493_;
  wire _23494_;
  wire _23495_;
  wire _23496_;
  wire _23497_;
  wire _23498_;
  wire _23499_;
  wire _23500_;
  wire _23501_;
  wire _23502_;
  wire _23503_;
  wire _23504_;
  wire _23505_;
  wire _23506_;
  wire _23507_;
  wire _23508_;
  wire _23509_;
  wire _23510_;
  wire _23511_;
  wire _23512_;
  wire _23513_;
  wire _23514_;
  wire _23515_;
  wire _23516_;
  wire _23517_;
  wire _23518_;
  wire _23519_;
  wire _23520_;
  wire _23521_;
  wire _23522_;
  wire _23523_;
  wire _23524_;
  wire _23525_;
  wire _23526_;
  wire _23527_;
  wire _23528_;
  wire _23529_;
  wire _23530_;
  wire _23531_;
  wire _23532_;
  wire _23533_;
  wire _23534_;
  wire _23535_;
  wire _23536_;
  wire _23537_;
  wire _23538_;
  wire _23539_;
  wire _23540_;
  wire _23541_;
  wire _23542_;
  wire _23543_;
  wire _23544_;
  wire _23545_;
  wire _23546_;
  wire _23547_;
  wire _23548_;
  wire _23549_;
  wire _23550_;
  wire _23551_;
  wire _23552_;
  wire _23553_;
  wire _23554_;
  wire _23555_;
  wire _23556_;
  wire _23557_;
  wire _23558_;
  wire _23559_;
  wire _23560_;
  wire _23561_;
  wire _23562_;
  wire _23563_;
  wire _23564_;
  wire _23565_;
  wire _23566_;
  wire _23567_;
  wire _23568_;
  wire _23569_;
  wire _23570_;
  wire _23571_;
  wire _23572_;
  wire _23573_;
  wire _23574_;
  wire _23575_;
  wire _23576_;
  wire _23577_;
  wire _23578_;
  wire _23579_;
  wire _23580_;
  wire _23581_;
  wire _23582_;
  wire _23583_;
  wire _23584_;
  wire _23585_;
  wire _23586_;
  wire _23587_;
  wire _23588_;
  wire _23589_;
  wire _23590_;
  wire _23591_;
  wire _23592_;
  wire _23593_;
  wire _23594_;
  wire _23595_;
  wire _23596_;
  wire _23597_;
  wire _23598_;
  wire _23599_;
  wire _23600_;
  wire _23601_;
  wire _23602_;
  wire _23603_;
  wire _23604_;
  wire _23605_;
  wire _23606_;
  wire _23607_;
  wire _23608_;
  wire _23609_;
  wire _23610_;
  wire _23611_;
  wire _23612_;
  wire _23613_;
  wire _23614_;
  wire _23615_;
  wire _23616_;
  wire _23617_;
  wire _23618_;
  wire _23619_;
  wire _23620_;
  wire _23621_;
  wire _23622_;
  wire _23623_;
  wire _23624_;
  wire _23625_;
  wire _23626_;
  wire _23627_;
  wire _23628_;
  wire _23629_;
  wire _23630_;
  wire _23631_;
  wire _23632_;
  wire _23633_;
  wire _23634_;
  wire _23635_;
  wire _23636_;
  wire _23637_;
  wire _23638_;
  wire _23639_;
  wire _23640_;
  wire _23641_;
  wire _23642_;
  wire _23643_;
  wire _23644_;
  wire _23645_;
  wire _23646_;
  wire _23647_;
  wire _23648_;
  wire _23649_;
  wire _23650_;
  wire _23651_;
  wire _23652_;
  wire _23653_;
  wire _23654_;
  wire _23655_;
  wire _23656_;
  wire _23657_;
  wire _23658_;
  wire _23659_;
  wire _23660_;
  wire _23661_;
  wire _23662_;
  wire _23663_;
  wire _23664_;
  wire _23665_;
  wire _23666_;
  wire _23667_;
  wire _23668_;
  wire _23669_;
  wire _23670_;
  wire _23671_;
  wire _23672_;
  wire _23673_;
  wire _23674_;
  wire _23675_;
  wire _23676_;
  wire _23677_;
  wire _23678_;
  wire _23679_;
  wire _23680_;
  wire _23681_;
  wire _23682_;
  wire _23683_;
  wire _23684_;
  wire _23685_;
  wire _23686_;
  wire _23687_;
  wire _23688_;
  wire _23689_;
  wire _23690_;
  wire _23691_;
  wire _23692_;
  wire _23693_;
  wire _23694_;
  wire _23695_;
  wire _23696_;
  wire _23697_;
  wire _23698_;
  wire _23699_;
  wire _23700_;
  wire _23701_;
  wire _23702_;
  wire _23703_;
  wire _23704_;
  wire _23705_;
  wire _23706_;
  wire _23707_;
  wire _23708_;
  wire _23709_;
  wire _23710_;
  wire _23711_;
  wire _23712_;
  wire _23713_;
  wire _23714_;
  wire _23715_;
  wire _23716_;
  wire _23717_;
  wire _23718_;
  wire _23719_;
  wire _23720_;
  wire _23721_;
  wire _23722_;
  wire _23723_;
  wire _23724_;
  wire _23725_;
  wire _23726_;
  wire _23727_;
  wire _23728_;
  wire _23729_;
  wire _23730_;
  wire _23731_;
  wire _23732_;
  wire _23733_;
  wire _23734_;
  wire _23735_;
  wire _23736_;
  wire _23737_;
  wire _23738_;
  wire _23739_;
  wire _23740_;
  wire _23741_;
  wire _23742_;
  wire _23743_;
  wire _23744_;
  wire _23745_;
  wire _23746_;
  wire _23747_;
  wire _23748_;
  wire _23749_;
  wire _23750_;
  wire _23751_;
  wire _23752_;
  wire _23753_;
  wire _23754_;
  wire _23755_;
  wire _23756_;
  wire _23757_;
  wire _23758_;
  wire _23759_;
  wire _23760_;
  wire _23761_;
  wire _23762_;
  wire _23763_;
  wire _23764_;
  wire _23765_;
  wire _23766_;
  wire _23767_;
  wire _23768_;
  wire _23769_;
  wire _23770_;
  wire _23771_;
  wire _23772_;
  wire _23773_;
  wire _23774_;
  wire _23775_;
  wire _23776_;
  wire _23777_;
  wire _23778_;
  wire _23779_;
  wire _23780_;
  wire _23781_;
  wire _23782_;
  wire _23783_;
  wire _23784_;
  wire _23785_;
  wire _23786_;
  wire _23787_;
  wire _23788_;
  wire _23789_;
  wire _23790_;
  wire _23791_;
  wire _23792_;
  wire _23793_;
  wire _23794_;
  wire _23795_;
  wire _23796_;
  wire _23797_;
  wire _23798_;
  wire _23799_;
  wire _23800_;
  wire _23801_;
  wire _23802_;
  wire _23803_;
  wire _23804_;
  wire _23805_;
  wire _23806_;
  wire _23807_;
  wire _23808_;
  wire _23809_;
  wire _23810_;
  wire _23811_;
  wire _23812_;
  wire _23813_;
  wire _23814_;
  wire _23815_;
  wire _23816_;
  wire _23817_;
  wire _23818_;
  wire _23819_;
  wire _23820_;
  wire _23821_;
  wire _23822_;
  wire _23823_;
  wire _23824_;
  wire _23825_;
  wire _23826_;
  wire _23827_;
  wire _23828_;
  wire _23829_;
  wire _23830_;
  wire _23831_;
  wire _23832_;
  wire _23833_;
  wire _23834_;
  wire _23835_;
  wire _23836_;
  wire _23837_;
  wire _23838_;
  wire _23839_;
  wire _23840_;
  wire _23841_;
  wire _23842_;
  wire _23843_;
  wire _23844_;
  wire _23845_;
  wire _23846_;
  wire _23847_;
  wire _23848_;
  wire _23849_;
  wire _23850_;
  wire _23851_;
  wire _23852_;
  wire _23853_;
  wire _23854_;
  wire _23855_;
  wire _23856_;
  wire _23857_;
  wire _23858_;
  wire _23859_;
  wire _23860_;
  wire _23861_;
  wire _23862_;
  wire _23863_;
  wire _23864_;
  wire _23865_;
  wire _23866_;
  wire _23867_;
  wire _23868_;
  wire _23869_;
  wire _23870_;
  wire _23871_;
  wire _23872_;
  wire _23873_;
  wire _23874_;
  wire _23875_;
  wire _23876_;
  wire _23877_;
  wire _23878_;
  wire _23879_;
  wire _23880_;
  wire _23881_;
  wire _23882_;
  wire _23883_;
  wire _23884_;
  wire _23885_;
  wire _23886_;
  wire _23887_;
  wire _23888_;
  wire _23889_;
  wire _23890_;
  wire _23891_;
  wire _23892_;
  wire _23893_;
  wire _23894_;
  wire _23895_;
  wire _23896_;
  wire _23897_;
  wire _23898_;
  wire _23899_;
  wire _23900_;
  wire _23901_;
  wire _23902_;
  wire _23903_;
  wire _23904_;
  wire _23905_;
  wire _23906_;
  wire _23907_;
  wire _23908_;
  wire _23909_;
  wire _23910_;
  wire _23911_;
  wire _23912_;
  wire _23913_;
  wire _23914_;
  wire _23915_;
  wire _23916_;
  wire _23917_;
  wire _23918_;
  wire _23919_;
  wire _23920_;
  wire _23921_;
  wire _23922_;
  wire _23923_;
  wire _23924_;
  wire _23925_;
  wire _23926_;
  wire _23927_;
  wire _23928_;
  wire _23929_;
  wire _23930_;
  wire _23931_;
  wire _23932_;
  wire _23933_;
  wire _23934_;
  wire _23935_;
  wire _23936_;
  wire _23937_;
  wire _23938_;
  wire _23939_;
  wire _23940_;
  wire _23941_;
  wire _23942_;
  wire _23943_;
  wire _23944_;
  wire _23945_;
  wire _23946_;
  wire _23947_;
  wire _23948_;
  wire _23949_;
  wire _23950_;
  wire _23951_;
  wire _23952_;
  wire _23953_;
  wire _23954_;
  wire _23955_;
  wire _23956_;
  wire _23957_;
  wire _23958_;
  wire _23959_;
  wire _23960_;
  wire _23961_;
  wire _23962_;
  wire _23963_;
  wire _23964_;
  wire _23965_;
  wire _23966_;
  wire _23967_;
  wire _23968_;
  wire _23969_;
  wire _23970_;
  wire _23971_;
  wire _23972_;
  wire _23973_;
  wire _23974_;
  wire _23975_;
  wire _23976_;
  wire _23977_;
  wire _23978_;
  wire _23979_;
  wire _23980_;
  wire _23981_;
  wire _23982_;
  wire _23983_;
  wire _23984_;
  wire _23985_;
  wire _23986_;
  wire _23987_;
  wire _23988_;
  wire _23989_;
  wire _23990_;
  wire _23991_;
  wire _23992_;
  wire _23993_;
  wire _23994_;
  wire _23995_;
  wire _23996_;
  wire _23997_;
  wire _23998_;
  wire _23999_;
  wire _24000_;
  wire _24001_;
  wire _24002_;
  wire _24003_;
  wire _24004_;
  wire _24005_;
  wire _24006_;
  wire _24007_;
  wire _24008_;
  wire _24009_;
  wire _24010_;
  wire _24011_;
  wire _24012_;
  wire _24013_;
  wire _24014_;
  wire _24015_;
  wire _24016_;
  wire _24017_;
  wire _24018_;
  wire _24019_;
  wire _24020_;
  wire _24021_;
  wire _24022_;
  wire _24023_;
  wire _24024_;
  wire _24025_;
  wire _24026_;
  wire _24027_;
  wire _24028_;
  wire _24029_;
  wire _24030_;
  wire _24031_;
  wire _24032_;
  wire _24033_;
  wire _24034_;
  wire _24035_;
  wire _24036_;
  wire _24037_;
  wire _24038_;
  wire _24039_;
  wire _24040_;
  wire _24041_;
  wire _24042_;
  wire _24043_;
  wire _24044_;
  wire _24045_;
  wire _24046_;
  wire _24047_;
  wire _24048_;
  wire _24049_;
  wire _24050_;
  wire _24051_;
  wire _24052_;
  wire _24053_;
  wire _24054_;
  wire _24055_;
  wire _24056_;
  wire _24057_;
  wire _24058_;
  wire _24059_;
  wire _24060_;
  wire _24061_;
  wire _24062_;
  wire _24063_;
  wire _24064_;
  wire _24065_;
  wire _24066_;
  wire _24067_;
  wire _24068_;
  wire _24069_;
  wire _24070_;
  wire _24071_;
  wire _24072_;
  wire _24073_;
  wire _24074_;
  wire _24075_;
  wire _24076_;
  wire _24077_;
  wire _24078_;
  wire _24079_;
  wire _24080_;
  wire _24081_;
  wire _24082_;
  wire _24083_;
  wire _24084_;
  wire _24085_;
  wire _24086_;
  wire _24087_;
  wire _24088_;
  wire _24089_;
  wire _24090_;
  wire _24091_;
  wire _24092_;
  wire _24093_;
  wire _24094_;
  wire _24095_;
  wire _24096_;
  wire _24097_;
  wire _24098_;
  wire _24099_;
  wire _24100_;
  wire _24101_;
  wire _24102_;
  wire _24103_;
  wire _24104_;
  wire _24105_;
  wire _24106_;
  wire _24107_;
  wire _24108_;
  wire _24109_;
  wire _24110_;
  wire _24111_;
  wire _24112_;
  wire _24113_;
  wire _24114_;
  wire _24115_;
  wire _24116_;
  wire _24117_;
  wire _24118_;
  wire _24119_;
  wire _24120_;
  wire _24121_;
  wire _24122_;
  wire _24123_;
  wire _24124_;
  wire _24125_;
  wire _24126_;
  wire _24127_;
  wire _24128_;
  wire _24129_;
  wire _24130_;
  wire _24131_;
  wire _24132_;
  wire _24133_;
  wire _24134_;
  wire _24135_;
  wire _24136_;
  wire _24137_;
  wire _24138_;
  wire _24139_;
  wire _24140_;
  wire _24141_;
  wire _24142_;
  wire _24143_;
  wire _24144_;
  wire _24145_;
  wire _24146_;
  wire _24147_;
  wire _24148_;
  wire _24149_;
  wire _24150_;
  wire _24151_;
  wire _24152_;
  wire _24153_;
  wire _24154_;
  wire _24155_;
  wire _24156_;
  wire _24157_;
  wire _24158_;
  wire _24159_;
  wire _24160_;
  wire _24161_;
  wire _24162_;
  wire _24163_;
  wire _24164_;
  wire _24165_;
  wire _24166_;
  wire _24167_;
  wire _24168_;
  wire _24169_;
  wire _24170_;
  wire _24171_;
  wire _24172_;
  wire _24173_;
  wire _24174_;
  wire _24175_;
  wire _24176_;
  wire _24177_;
  wire _24178_;
  wire _24179_;
  wire _24180_;
  wire _24181_;
  wire _24182_;
  wire _24183_;
  wire _24184_;
  wire _24185_;
  wire _24186_;
  wire _24187_;
  wire _24188_;
  wire _24189_;
  wire _24190_;
  wire _24191_;
  wire _24192_;
  wire _24193_;
  wire _24194_;
  wire _24195_;
  wire _24196_;
  wire _24197_;
  wire _24198_;
  wire _24199_;
  wire _24200_;
  wire _24201_;
  wire _24202_;
  wire _24203_;
  wire _24204_;
  wire _24205_;
  wire _24206_;
  wire _24207_;
  wire _24208_;
  wire _24209_;
  wire _24210_;
  wire _24211_;
  wire _24212_;
  wire _24213_;
  wire _24214_;
  wire _24215_;
  wire _24216_;
  wire _24217_;
  wire _24218_;
  wire _24219_;
  wire _24220_;
  wire _24221_;
  wire _24222_;
  wire _24223_;
  wire _24224_;
  wire _24225_;
  wire _24226_;
  wire _24227_;
  wire _24228_;
  wire _24229_;
  wire _24230_;
  wire _24231_;
  wire _24232_;
  wire _24233_;
  wire _24234_;
  wire _24235_;
  wire _24236_;
  wire _24237_;
  wire _24238_;
  wire _24239_;
  wire _24240_;
  wire _24241_;
  wire _24242_;
  wire _24243_;
  wire _24244_;
  wire _24245_;
  wire _24246_;
  wire _24247_;
  wire _24248_;
  wire _24249_;
  wire _24250_;
  wire _24251_;
  wire _24252_;
  wire _24253_;
  wire _24254_;
  wire _24255_;
  wire _24256_;
  wire _24257_;
  wire _24258_;
  wire _24259_;
  wire _24260_;
  wire _24261_;
  wire _24262_;
  wire _24263_;
  wire _24264_;
  wire _24265_;
  wire _24266_;
  wire _24267_;
  wire _24268_;
  wire _24269_;
  wire _24270_;
  wire _24271_;
  wire _24272_;
  wire _24273_;
  wire _24274_;
  wire _24275_;
  wire _24276_;
  wire _24277_;
  wire _24278_;
  wire _24279_;
  wire _24280_;
  wire _24281_;
  wire _24282_;
  wire _24283_;
  wire _24284_;
  wire _24285_;
  wire _24286_;
  wire _24287_;
  wire _24288_;
  wire _24289_;
  wire _24290_;
  wire _24291_;
  wire _24292_;
  wire _24293_;
  wire _24294_;
  wire _24295_;
  wire _24296_;
  wire _24297_;
  wire _24298_;
  wire _24299_;
  wire _24300_;
  wire _24301_;
  wire _24302_;
  wire _24303_;
  wire _24304_;
  wire _24305_;
  wire _24306_;
  wire _24307_;
  wire _24308_;
  wire _24309_;
  wire _24310_;
  wire _24311_;
  wire _24312_;
  wire _24313_;
  wire _24314_;
  wire _24315_;
  wire _24316_;
  wire _24317_;
  wire _24318_;
  wire _24319_;
  wire _24320_;
  wire _24321_;
  wire _24322_;
  wire _24323_;
  wire _24324_;
  wire _24325_;
  wire _24326_;
  wire _24327_;
  wire _24328_;
  wire _24329_;
  wire _24330_;
  wire _24331_;
  wire _24332_;
  wire _24333_;
  wire _24334_;
  wire _24335_;
  wire _24336_;
  wire _24337_;
  wire _24338_;
  wire _24339_;
  wire _24340_;
  wire _24341_;
  wire _24342_;
  wire _24343_;
  wire _24344_;
  wire _24345_;
  wire _24346_;
  wire _24347_;
  wire _24348_;
  wire _24349_;
  wire _24350_;
  wire _24351_;
  wire _24352_;
  wire _24353_;
  wire _24354_;
  wire _24355_;
  wire _24356_;
  wire _24357_;
  wire _24358_;
  wire _24359_;
  wire _24360_;
  wire _24361_;
  wire _24362_;
  wire _24363_;
  wire _24364_;
  wire _24365_;
  wire _24366_;
  wire _24367_;
  wire _24368_;
  wire _24369_;
  wire _24370_;
  wire _24371_;
  wire _24372_;
  wire _24373_;
  wire _24374_;
  wire _24375_;
  wire _24376_;
  wire _24377_;
  wire _24378_;
  wire _24379_;
  wire _24380_;
  wire _24381_;
  wire _24382_;
  wire _24383_;
  wire _24384_;
  wire _24385_;
  wire _24386_;
  wire _24387_;
  wire _24388_;
  wire _24389_;
  wire _24390_;
  wire _24391_;
  wire _24392_;
  wire _24393_;
  wire _24394_;
  wire _24395_;
  wire _24396_;
  wire _24397_;
  wire _24398_;
  wire _24399_;
  wire _24400_;
  wire _24401_;
  wire _24402_;
  wire _24403_;
  wire _24404_;
  wire _24405_;
  wire _24406_;
  wire _24407_;
  wire _24408_;
  wire _24409_;
  wire _24410_;
  wire _24411_;
  wire _24412_;
  wire _24413_;
  wire _24414_;
  wire _24415_;
  wire _24416_;
  wire _24417_;
  wire _24418_;
  wire _24419_;
  wire _24420_;
  wire _24421_;
  wire _24422_;
  wire _24423_;
  wire _24424_;
  wire _24425_;
  wire _24426_;
  wire _24427_;
  wire _24428_;
  wire _24429_;
  wire _24430_;
  wire _24431_;
  wire _24432_;
  wire _24433_;
  wire _24434_;
  wire _24435_;
  wire _24436_;
  wire _24437_;
  wire _24438_;
  wire _24439_;
  wire _24440_;
  wire _24441_;
  wire _24442_;
  wire _24443_;
  wire _24444_;
  wire _24445_;
  wire _24446_;
  wire _24447_;
  wire _24448_;
  wire _24449_;
  wire _24450_;
  wire _24451_;
  wire _24452_;
  wire _24453_;
  wire _24454_;
  wire _24455_;
  wire _24456_;
  wire _24457_;
  wire _24458_;
  wire _24459_;
  wire _24460_;
  wire _24461_;
  wire _24462_;
  wire _24463_;
  wire _24464_;
  wire _24465_;
  wire _24466_;
  wire _24467_;
  wire _24468_;
  wire _24469_;
  wire _24470_;
  wire _24471_;
  wire _24472_;
  wire _24473_;
  wire _24474_;
  wire _24475_;
  wire _24476_;
  wire _24477_;
  wire _24478_;
  wire _24479_;
  wire _24480_;
  wire _24481_;
  wire _24482_;
  wire _24483_;
  wire _24484_;
  wire _24485_;
  wire _24486_;
  wire _24487_;
  wire _24488_;
  wire _24489_;
  wire _24490_;
  wire _24491_;
  wire _24492_;
  wire _24493_;
  wire _24494_;
  wire _24495_;
  wire _24496_;
  wire _24497_;
  wire _24498_;
  wire _24499_;
  wire _24500_;
  wire _24501_;
  wire _24502_;
  wire _24503_;
  wire _24504_;
  wire _24505_;
  wire _24506_;
  wire _24507_;
  wire _24508_;
  wire _24509_;
  wire _24510_;
  wire _24511_;
  wire _24512_;
  wire _24513_;
  wire _24514_;
  wire _24515_;
  wire _24516_;
  wire _24517_;
  wire _24518_;
  wire _24519_;
  wire _24520_;
  wire _24521_;
  wire _24522_;
  wire _24523_;
  wire _24524_;
  wire _24525_;
  wire _24526_;
  wire _24527_;
  wire _24528_;
  wire _24529_;
  wire _24530_;
  wire _24531_;
  wire _24532_;
  wire _24533_;
  wire _24534_;
  wire _24535_;
  wire _24536_;
  wire _24537_;
  wire _24538_;
  wire _24539_;
  wire _24540_;
  wire _24541_;
  wire _24542_;
  wire _24543_;
  wire _24544_;
  wire _24545_;
  wire _24546_;
  wire _24547_;
  wire _24548_;
  wire _24549_;
  wire _24550_;
  wire _24551_;
  wire _24552_;
  wire _24553_;
  wire _24554_;
  wire _24555_;
  wire _24556_;
  wire _24557_;
  wire _24558_;
  wire _24559_;
  wire _24560_;
  wire _24561_;
  wire _24562_;
  wire _24563_;
  wire _24564_;
  wire _24565_;
  wire _24566_;
  wire _24567_;
  wire _24568_;
  wire _24569_;
  wire _24570_;
  wire _24571_;
  wire _24572_;
  wire _24573_;
  wire _24574_;
  wire _24575_;
  wire _24576_;
  wire _24577_;
  wire _24578_;
  wire _24579_;
  wire _24580_;
  wire _24581_;
  wire _24582_;
  wire _24583_;
  wire _24584_;
  wire _24585_;
  wire _24586_;
  wire _24587_;
  wire _24588_;
  wire _24589_;
  wire _24590_;
  wire _24591_;
  wire _24592_;
  wire _24593_;
  wire _24594_;
  wire _24595_;
  wire _24596_;
  wire _24597_;
  wire _24598_;
  wire _24599_;
  wire _24600_;
  wire _24601_;
  wire _24602_;
  wire _24603_;
  wire _24604_;
  wire _24605_;
  wire _24606_;
  wire _24607_;
  wire _24608_;
  wire _24609_;
  wire _24610_;
  wire _24611_;
  wire _24612_;
  wire _24613_;
  wire _24614_;
  wire _24615_;
  wire _24616_;
  wire _24617_;
  wire _24618_;
  wire _24619_;
  wire _24620_;
  wire _24621_;
  wire _24622_;
  wire _24623_;
  wire _24624_;
  wire _24625_;
  wire _24626_;
  wire _24627_;
  wire _24628_;
  wire _24629_;
  wire _24630_;
  wire _24631_;
  wire _24632_;
  wire _24633_;
  wire _24634_;
  wire _24635_;
  wire _24636_;
  wire _24637_;
  wire _24638_;
  wire _24639_;
  wire _24640_;
  wire _24641_;
  wire _24642_;
  wire _24643_;
  wire _24644_;
  wire _24645_;
  wire _24646_;
  wire _24647_;
  wire _24648_;
  wire _24649_;
  wire _24650_;
  wire _24651_;
  wire _24652_;
  wire _24653_;
  wire _24654_;
  wire _24655_;
  wire _24656_;
  wire _24657_;
  wire _24658_;
  wire _24659_;
  wire _24660_;
  wire _24661_;
  wire _24662_;
  wire _24663_;
  wire _24664_;
  wire _24665_;
  wire _24666_;
  wire _24667_;
  wire _24668_;
  wire _24669_;
  wire _24670_;
  wire _24671_;
  wire _24672_;
  wire _24673_;
  wire _24674_;
  wire _24675_;
  wire _24676_;
  wire _24677_;
  wire _24678_;
  wire _24679_;
  wire _24680_;
  wire _24681_;
  wire _24682_;
  wire _24683_;
  wire _24684_;
  wire _24685_;
  wire _24686_;
  wire _24687_;
  wire _24688_;
  wire _24689_;
  wire _24690_;
  wire _24691_;
  wire _24692_;
  wire _24693_;
  wire _24694_;
  wire _24695_;
  wire _24696_;
  wire _24697_;
  wire _24698_;
  wire _24699_;
  wire _24700_;
  wire _24701_;
  wire _24702_;
  wire _24703_;
  wire _24704_;
  wire _24705_;
  wire _24706_;
  wire _24707_;
  wire _24708_;
  wire _24709_;
  wire _24710_;
  wire _24711_;
  wire _24712_;
  wire _24713_;
  wire _24714_;
  wire _24715_;
  wire _24716_;
  wire _24717_;
  wire _24718_;
  wire _24719_;
  wire _24720_;
  wire _24721_;
  wire _24722_;
  wire _24723_;
  wire _24724_;
  wire _24725_;
  wire _24726_;
  wire _24727_;
  wire _24728_;
  wire _24729_;
  wire _24730_;
  wire _24731_;
  wire _24732_;
  wire _24733_;
  wire _24734_;
  wire _24735_;
  wire _24736_;
  wire _24737_;
  wire _24738_;
  wire _24739_;
  wire _24740_;
  wire _24741_;
  wire _24742_;
  wire _24743_;
  wire _24744_;
  wire _24745_;
  wire _24746_;
  wire _24747_;
  wire _24748_;
  wire _24749_;
  wire _24750_;
  wire _24751_;
  wire _24752_;
  wire _24753_;
  wire _24754_;
  wire _24755_;
  wire _24756_;
  wire _24757_;
  wire _24758_;
  wire _24759_;
  wire _24760_;
  wire _24761_;
  wire _24762_;
  wire _24763_;
  wire _24764_;
  wire _24765_;
  wire _24766_;
  wire _24767_;
  wire _24768_;
  wire _24769_;
  wire _24770_;
  wire _24771_;
  wire _24772_;
  wire _24773_;
  wire _24774_;
  wire _24775_;
  wire _24776_;
  wire _24777_;
  wire _24778_;
  wire _24779_;
  wire _24780_;
  wire _24781_;
  wire _24782_;
  wire _24783_;
  wire _24784_;
  wire _24785_;
  wire _24786_;
  wire _24787_;
  wire _24788_;
  wire _24789_;
  wire _24790_;
  wire _24791_;
  wire _24792_;
  wire _24793_;
  wire _24794_;
  wire _24795_;
  wire _24796_;
  wire _24797_;
  wire _24798_;
  wire _24799_;
  wire _24800_;
  wire _24801_;
  wire _24802_;
  wire _24803_;
  wire _24804_;
  wire _24805_;
  wire _24806_;
  wire _24807_;
  wire _24808_;
  wire _24809_;
  wire _24810_;
  wire _24811_;
  wire _24812_;
  wire _24813_;
  wire _24814_;
  wire _24815_;
  wire _24816_;
  wire _24817_;
  wire _24818_;
  wire _24819_;
  wire _24820_;
  wire _24821_;
  wire _24822_;
  wire _24823_;
  wire _24824_;
  wire _24825_;
  wire _24826_;
  wire _24827_;
  wire _24828_;
  wire _24829_;
  wire _24830_;
  wire _24831_;
  wire _24832_;
  wire _24833_;
  wire _24834_;
  wire _24835_;
  wire _24836_;
  wire _24837_;
  wire _24838_;
  wire _24839_;
  wire _24840_;
  wire _24841_;
  wire _24842_;
  wire _24843_;
  wire _24844_;
  wire _24845_;
  wire _24846_;
  wire _24847_;
  wire _24848_;
  wire _24849_;
  wire _24850_;
  wire _24851_;
  wire _24852_;
  wire _24853_;
  wire _24854_;
  wire _24855_;
  wire _24856_;
  wire _24857_;
  wire _24858_;
  wire _24859_;
  wire _24860_;
  wire _24861_;
  wire _24862_;
  wire _24863_;
  wire _24864_;
  wire _24865_;
  wire _24866_;
  wire _24867_;
  wire _24868_;
  wire _24869_;
  wire _24870_;
  wire _24871_;
  wire _24872_;
  wire _24873_;
  wire _24874_;
  wire _24875_;
  wire _24876_;
  wire _24877_;
  wire _24878_;
  wire _24879_;
  wire _24880_;
  wire _24881_;
  wire _24882_;
  wire _24883_;
  wire _24884_;
  wire _24885_;
  wire _24886_;
  wire _24887_;
  wire _24888_;
  wire _24889_;
  wire _24890_;
  wire _24891_;
  wire _24892_;
  wire _24893_;
  wire _24894_;
  wire _24895_;
  wire _24896_;
  wire _24897_;
  wire _24898_;
  wire _24899_;
  wire _24900_;
  wire _24901_;
  wire _24902_;
  wire _24903_;
  wire _24904_;
  wire _24905_;
  wire _24906_;
  wire _24907_;
  wire _24908_;
  wire _24909_;
  wire _24910_;
  wire _24911_;
  wire _24912_;
  wire _24913_;
  wire _24914_;
  wire _24915_;
  wire _24916_;
  wire _24917_;
  wire _24918_;
  wire _24919_;
  wire _24920_;
  wire _24921_;
  wire _24922_;
  wire _24923_;
  wire _24924_;
  wire _24925_;
  wire _24926_;
  wire _24927_;
  wire _24928_;
  wire _24929_;
  wire _24930_;
  wire _24931_;
  wire _24932_;
  wire _24933_;
  wire _24934_;
  wire _24935_;
  wire _24936_;
  wire _24937_;
  wire _24938_;
  wire _24939_;
  wire _24940_;
  wire _24941_;
  wire _24942_;
  wire _24943_;
  wire _24944_;
  wire _24945_;
  wire _24946_;
  wire _24947_;
  wire _24948_;
  wire _24949_;
  wire _24950_;
  wire _24951_;
  wire _24952_;
  wire _24953_;
  wire _24954_;
  wire _24955_;
  wire _24956_;
  wire _24957_;
  wire _24958_;
  wire _24959_;
  wire _24960_;
  wire _24961_;
  wire _24962_;
  wire _24963_;
  wire [15:0] _24964_;
  wire _24965_;
  wire _24966_;
  wire _24967_;
  wire _24968_;
  wire _24969_;
  wire _24970_;
  wire _24971_;
  wire _24972_;
  wire _24973_;
  wire _24974_;
  wire _24975_;
  wire _24976_;
  wire _24977_;
  wire _24978_;
  wire _24979_;
  wire _24980_;
  wire _24981_;
  wire _24982_;
  wire _24983_;
  wire _24984_;
  wire _24985_;
  wire _24986_;
  wire _24987_;
  wire _24988_;
  wire _24989_;
  wire _24990_;
  wire _24991_;
  wire _24992_;
  wire _24993_;
  wire _24994_;
  wire _24995_;
  wire _24996_;
  wire _24997_;
  wire _24998_;
  wire _24999_;
  wire _25000_;
  wire _25001_;
  wire _25002_;
  wire _25003_;
  wire _25004_;
  wire [7:0] _25005_;
  wire [7:0] _25006_;
  wire [7:0] _25007_;
  wire [7:0] _25008_;
  wire [7:0] _25009_;
  wire [7:0] _25010_;
  wire [7:0] _25011_;
  wire [7:0] _25012_;
  wire [7:0] _25013_;
  wire [7:0] _25014_;
  wire [7:0] _25015_;
  wire [2:0] _25016_;
  wire [2:0] _25017_;
  wire [1:0] _25018_;
  wire [7:0] _25019_;
  wire [1:0] _25020_;
  wire [2:0] _25021_;
  wire [1:0] _25022_;
  wire _25023_;
  wire [7:0] _25024_;
  wire [7:0] _25025_;
  wire [7:0] _25026_;
  wire [7:0] _25027_;
  wire [7:0] _25028_;
  wire [7:0] _25029_;
  wire [7:0] _25030_;
  wire [15:0] _25031_;
  wire [15:0] _25032_;
  wire [7:0] _25033_;
  wire [15:0] _25034_;
  wire _25035_;
  wire [7:0] _25036_;
  wire [2:0] _25037_;
  wire [7:0] _25038_;
  wire [7:0] _25039_;
  wire [7:0] _25040_;
  wire _25041_;
  wire [31:0] _25042_;
  wire [31:0] _25043_;
  wire [7:0] _25044_;
  wire _25045_;
  wire _25046_;
  wire _25047_;
  wire _25048_;
  wire _25049_;
  wire _25050_;
  wire _25051_;
  wire _25052_;
  wire _25053_;
  wire _25054_;
  wire _25055_;
  wire _25056_;
  wire _25057_;
  wire _25058_;
  wire _25059_;
  wire _25060_;
  wire _25061_;
  wire _25062_;
  wire _25063_;
  wire _25064_;
  wire _25065_;
  wire _25066_;
  wire _25067_;
  wire _25068_;
  wire _25069_;
  wire _25070_;
  wire _25071_;
  wire _25072_;
  wire _25073_;
  wire _25074_;
  wire _25075_;
  wire _25076_;
  wire _25077_;
  wire _25078_;
  wire _25079_;
  wire _25080_;
  wire _25081_;
  wire _25082_;
  wire _25083_;
  wire _25084_;
  wire _25085_;
  wire _25086_;
  wire _25087_;
  wire _25088_;
  wire _25089_;
  wire _25090_;
  wire _25091_;
  wire _25092_;
  wire _25093_;
  wire _25094_;
  wire _25095_;
  wire _25096_;
  wire _25097_;
  wire _25098_;
  wire _25099_;
  wire _25100_;
  wire _25101_;
  wire _25102_;
  wire _25103_;
  wire _25104_;
  wire _25105_;
  wire _25106_;
  wire _25107_;
  wire _25108_;
  wire _25109_;
  wire _25110_;
  wire _25111_;
  wire _25112_;
  wire _25113_;
  wire _25114_;
  wire _25115_;
  wire _25116_;
  wire _25117_;
  wire _25118_;
  wire _25119_;
  wire _25120_;
  wire _25121_;
  wire _25122_;
  wire _25123_;
  wire _25124_;
  wire _25125_;
  wire _25126_;
  wire _25127_;
  wire _25128_;
  wire _25129_;
  wire _25130_;
  wire _25131_;
  wire _25132_;
  wire _25133_;
  wire _25134_;
  wire _25135_;
  wire _25136_;
  wire _25137_;
  wire _25138_;
  wire _25139_;
  wire _25140_;
  wire _25141_;
  wire _25142_;
  wire _25143_;
  wire _25144_;
  wire _25145_;
  wire _25146_;
  wire _25147_;
  wire _25148_;
  wire _25149_;
  wire _25150_;
  wire _25151_;
  wire _25152_;
  wire _25153_;
  wire _25154_;
  wire _25155_;
  wire _25156_;
  wire _25157_;
  wire _25158_;
  wire _25159_;
  wire _25160_;
  wire _25161_;
  wire _25162_;
  wire _25163_;
  wire _25164_;
  wire _25165_;
  wire _25166_;
  wire _25167_;
  wire _25168_;
  wire _25169_;
  wire _25170_;
  wire _25171_;
  wire _25172_;
  wire _25173_;
  wire _25174_;
  wire _25175_;
  wire _25176_;
  wire _25177_;
  wire _25178_;
  wire _25179_;
  wire _25180_;
  wire _25181_;
  wire _25182_;
  wire _25183_;
  wire _25184_;
  wire _25185_;
  wire _25186_;
  wire _25187_;
  wire _25188_;
  wire _25189_;
  wire _25190_;
  wire _25191_;
  wire _25192_;
  wire _25193_;
  wire _25194_;
  wire _25195_;
  wire _25196_;
  wire _25197_;
  wire _25198_;
  wire _25199_;
  wire _25200_;
  wire _25201_;
  wire _25202_;
  wire _25203_;
  wire _25204_;
  wire _25205_;
  wire _25206_;
  wire _25207_;
  wire _25208_;
  wire _25209_;
  wire _25210_;
  wire _25211_;
  wire _25212_;
  wire _25213_;
  wire _25214_;
  wire _25215_;
  wire _25216_;
  wire _25217_;
  wire _25218_;
  wire _25219_;
  wire _25220_;
  wire _25221_;
  wire _25222_;
  wire _25223_;
  wire _25224_;
  wire _25225_;
  wire _25226_;
  wire _25227_;
  wire _25228_;
  wire _25229_;
  wire _25230_;
  wire _25231_;
  wire _25232_;
  wire _25233_;
  wire _25234_;
  wire _25235_;
  wire _25236_;
  wire _25237_;
  wire _25238_;
  wire _25239_;
  wire _25240_;
  wire _25241_;
  wire _25242_;
  wire _25243_;
  wire _25244_;
  wire _25245_;
  wire _25246_;
  wire _25247_;
  wire _25248_;
  wire _25249_;
  wire _25250_;
  wire _25251_;
  wire _25252_;
  wire _25253_;
  wire _25254_;
  wire _25255_;
  wire _25256_;
  wire _25257_;
  wire _25258_;
  wire _25259_;
  wire _25260_;
  wire _25261_;
  wire _25262_;
  wire _25263_;
  wire _25264_;
  wire _25265_;
  wire _25266_;
  wire _25267_;
  wire _25268_;
  wire _25269_;
  wire _25270_;
  wire _25271_;
  wire _25272_;
  wire _25273_;
  wire _25274_;
  wire _25275_;
  wire _25276_;
  wire _25277_;
  wire _25278_;
  wire _25279_;
  wire _25280_;
  wire _25281_;
  wire _25282_;
  wire _25283_;
  wire _25284_;
  wire _25285_;
  wire _25286_;
  wire _25287_;
  wire _25288_;
  wire _25289_;
  wire _25290_;
  wire _25291_;
  wire _25292_;
  wire _25293_;
  wire _25294_;
  wire _25295_;
  wire _25296_;
  wire _25297_;
  wire _25298_;
  wire _25299_;
  wire _25300_;
  wire _25301_;
  wire _25302_;
  wire _25303_;
  wire _25304_;
  wire _25305_;
  wire _25306_;
  wire _25307_;
  wire _25308_;
  wire _25309_;
  wire _25310_;
  wire _25311_;
  wire _25312_;
  wire _25313_;
  wire _25314_;
  wire _25315_;
  wire _25316_;
  wire _25317_;
  wire _25318_;
  wire _25319_;
  wire _25320_;
  wire _25321_;
  wire _25322_;
  wire _25323_;
  wire _25324_;
  wire _25325_;
  wire _25326_;
  wire _25327_;
  wire _25328_;
  wire _25329_;
  wire _25330_;
  wire _25331_;
  wire _25332_;
  wire _25333_;
  wire _25334_;
  wire _25335_;
  wire _25336_;
  wire _25337_;
  wire _25338_;
  wire _25339_;
  wire _25340_;
  wire _25341_;
  wire _25342_;
  wire _25343_;
  wire _25344_;
  wire _25345_;
  wire _25346_;
  wire _25347_;
  wire _25348_;
  wire _25349_;
  wire _25350_;
  wire _25351_;
  wire _25352_;
  wire _25353_;
  wire _25354_;
  wire _25355_;
  wire _25356_;
  wire _25357_;
  wire _25358_;
  wire _25359_;
  wire _25360_;
  wire _25361_;
  wire _25362_;
  wire _25363_;
  wire _25364_;
  wire _25365_;
  wire _25366_;
  wire _25367_;
  wire _25368_;
  wire _25369_;
  wire _25370_;
  wire _25371_;
  wire _25372_;
  wire _25373_;
  wire _25374_;
  wire _25375_;
  wire _25376_;
  wire _25377_;
  wire _25378_;
  wire _25379_;
  wire _25380_;
  wire _25381_;
  wire _25382_;
  wire _25383_;
  wire _25384_;
  wire _25385_;
  wire _25386_;
  wire _25387_;
  wire _25388_;
  wire _25389_;
  wire _25390_;
  wire _25391_;
  wire _25392_;
  wire _25393_;
  wire _25394_;
  wire _25395_;
  wire _25396_;
  wire _25397_;
  wire _25398_;
  wire _25399_;
  wire _25400_;
  wire _25401_;
  wire _25402_;
  wire _25403_;
  wire _25404_;
  wire _25405_;
  wire _25406_;
  wire _25407_;
  wire _25408_;
  wire _25409_;
  wire _25410_;
  wire _25411_;
  wire _25412_;
  wire _25413_;
  wire _25414_;
  wire _25415_;
  wire _25416_;
  wire _25417_;
  wire _25418_;
  wire _25419_;
  wire _25420_;
  wire _25421_;
  wire _25422_;
  wire _25423_;
  wire _25424_;
  wire _25425_;
  wire _25426_;
  wire _25427_;
  wire _25428_;
  wire _25429_;
  wire _25430_;
  wire _25431_;
  wire _25432_;
  wire _25433_;
  wire _25434_;
  wire _25435_;
  wire _25436_;
  wire _25437_;
  wire _25438_;
  wire _25439_;
  wire _25440_;
  wire _25441_;
  wire _25442_;
  wire _25443_;
  wire _25444_;
  wire _25445_;
  wire _25446_;
  wire _25447_;
  wire _25448_;
  wire _25449_;
  wire _25450_;
  wire _25451_;
  wire _25452_;
  wire _25453_;
  wire [7:0] _25454_;
  wire [3:0] _25455_;
  input [34:0] ABINPUT;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [34:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [7:0] \oc8051_top_1.des1 ;
  wire [7:0] \oc8051_top_1.des2 ;
  wire \oc8051_top_1.desAc ;
  wire \oc8051_top_1.desCy ;
  wire \oc8051_top_1.desOv ;
  wire [7:0] \oc8051_top_1.des_acc ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.des ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.data_in ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.alu ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des1 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des2 ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.des_acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.wr_dat ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_addr_r ;
  wire \oc8051_top_1.oc8051_ram_top1.bit_data_in ;
  wire [2:0] \oc8051_top_1.oc8051_ram_top1.bit_select ;
  wire \oc8051_top_1.oc8051_ram_top1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data ;
  wire \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.rd_data_m ;
  wire \oc8051_top_1.oc8051_ram_top1.rd_en_r ;
  wire \oc8051_top_1.oc8051_ram_top1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data ;
  wire [7:0] \oc8051_top_1.oc8051_ram_top1.wr_data_r ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat2 ;
  wire \oc8051_top_1.oc8051_sfr1.desAc ;
  wire \oc8051_top_1.oc8051_sfr1.desOv ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.des_acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.bit_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.p ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire \oc8051_top_1.srcAc ;
  wire [7:0] \oc8051_top_1.sub_result ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  wire [7:0] \oc8051_top_1.wr_dat ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc2;
  output property_invalid;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not (_21183_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_21184_, \oc8051_top_1.oc8051_decoder1.wr , _21183_);
  nand (_21185_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _21183_);
  nor (_21186_, _21185_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_21187_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  not (_21188_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nand (_21189_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nand (_21190_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_21191_, _21190_, _21189_);
  nand (_21192_, _21191_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_21193_, _21192_, _21188_);
  nand (_21194_, _21193_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_21195_, _21194_, _21187_);
  not (_21196_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  not (_21197_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_21198_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  nor (_21199_, _21198_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_21200_, _21199_, _21197_);
  nor (_21202_, _21200_, _21196_);
  nand (_21203_, _21194_, _21187_);
  nand (_21205_, _21203_, _21202_);
  nor (_21206_, _21205_, _21195_);
  nor (_21207_, _21197_, _21196_);
  nand (_21208_, _21207_, _21199_);
  not (_21209_, _21208_);
  not (_21210_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  nand (_21212_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _21183_);
  nor (_21213_, _21212_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  nand (_21214_, _21213_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nor (_21215_, _21214_, _21210_);
  nor (_21216_, _21215_, _21209_);
  nor (_21217_, _21196_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_21218_, _21217_, _21198_);
  nor (_21219_, _21218_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nand (_21220_, _21219_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_21221_, _21200_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  nand (_21222_, _21221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nand (_21223_, _21222_, _21220_);
  not (_21224_, _21223_);
  nand (_21226_, _21224_, _21216_);
  nor (_21227_, _21226_, _21206_);
  nor (_21229_, _21227_, _21186_);
  nor (_21230_, _21229_, _21184_);
  not (_21231_, _21230_);
  not (_21232_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  not (_21233_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_21234_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_21235_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_21236_, _21189_, _21235_);
  nand (_21237_, _21236_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_21238_, _21237_, _21234_);
  nand (_21239_, _21238_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_21240_, _21239_, _21233_);
  nor (_21241_, _21240_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_21242_, _21241_, _21195_);
  nand (_21243_, _21242_, _21202_);
  not (_21244_, _21216_);
  nor (_21245_, _21223_, _21244_);
  nand (_21246_, _21245_, _21243_);
  nor (_21247_, _21246_, _21232_);
  not (_21248_, _21247_);
  nand (_21249_, _21237_, _21234_);
  nand (_21250_, _21249_, _21202_);
  nor (_21251_, _21250_, _21238_);
  not (_21252_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_21253_, _21197_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_21254_, _21253_, _21199_);
  nand (_21255_, _21254_, _21212_);
  nor (_21256_, _21255_, _21252_);
  nor (_21257_, _21256_, _21209_);
  not (_21258_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nand (_21259_, _21186_, _21196_);
  nor (_21260_, _21259_, _21258_);
  nor (_21261_, _21218_, _21197_);
  nand (_21262_, _21261_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nand (_21263_, _21219_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nand (_21264_, _21263_, _21262_);
  nor (_21266_, _21264_, _21260_);
  nand (_21267_, _21266_, _21257_);
  nor (_21268_, _21267_, _21251_);
  nor (_21269_, _21268_, _21248_);
  nand (_21270_, _21219_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  nand (_21271_, _21221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nand (_21272_, _21271_, _21270_);
  not (_21273_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  not (_21274_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_21275_, _21274_, _21273_);
  nor (_21276_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_21277_, _21276_, _21275_);
  nand (_21278_, _21277_, _21202_);
  not (_21279_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nor (_21280_, _21214_, _21279_);
  not (_21281_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  nor (_21282_, _21255_, _21281_);
  nor (_21283_, _21282_, _21280_);
  nand (_21284_, _21283_, _21278_);
  nor (_21285_, _21284_, _21272_);
  nor (_21286_, _21285_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_21287_, _21286_, _21269_);
  nor (_21288_, _21287_, _21231_);
  not (_21289_, _21288_);
  nand (_21290_, _21186_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  not (_21291_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nand (_21292_, _21275_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nand (_21293_, _21292_, _21291_);
  nand (_21294_, _21293_, _21237_);
  nor (_21295_, _21294_, _21290_);
  nand (_21296_, _21219_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  not (_21297_, _21296_);
  not (_21298_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor (_21300_, _21255_, _21298_);
  nor (_21301_, _21300_, _21297_);
  not (_21302_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  nor (_21303_, _21214_, _21302_);
  not (_21304_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_21305_, _21259_, _21304_);
  nor (_21306_, _21305_, _21303_);
  nand (_21307_, _21306_, _21301_);
  nor (_21308_, _21307_, _21295_);
  nor (_21309_, _21308_, _21248_);
  nand (_21310_, _21261_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  nand (_21311_, _21219_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nand (_21312_, _21311_, _21310_);
  nand (_21313_, _21221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_21314_, _21290_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  not (_21315_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_21316_, _21255_, _21315_);
  nor (_21318_, _21316_, _21314_);
  nand (_21319_, _21318_, _21313_);
  nor (_21320_, _21319_, _21312_);
  nor (_21321_, _21320_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_21322_, _21321_, _21309_);
  nor (_21323_, _21322_, _21231_);
  nor (_21324_, _21323_, _21289_);
  not (_21325_, _21324_);
  nor (_21327_, _21238_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_21328_, _21327_, _21193_);
  nand (_21329_, _21328_, _21202_);
  nand (_21330_, _21219_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nand (_21331_, _21330_, _21208_);
  nand (_21332_, _21221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  nand (_21333_, _21261_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nand (_21334_, _21333_, _21332_);
  nor (_21335_, _21334_, _21331_);
  nand (_21336_, _21335_, _21329_);
  not (_21337_, _21336_);
  nor (_21338_, _21337_, _21248_);
  nand (_21339_, _21219_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  nand (_21340_, _21221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nand (_21341_, _21340_, _21339_);
  nor (_21342_, _21275_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_21343_, _21342_, _21236_);
  nand (_21344_, _21343_, _21202_);
  not (_21345_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  nor (_21346_, _21214_, _21345_);
  not (_21347_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  nor (_21348_, _21255_, _21347_);
  nor (_21349_, _21348_, _21346_);
  nand (_21350_, _21349_, _21344_);
  nor (_21351_, _21350_, _21341_);
  nor (_21352_, _21351_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_21353_, _21352_, _21338_);
  nor (_21354_, _21353_, _21231_);
  nand (_21355_, _21239_, _21233_);
  nand (_21356_, _21355_, _21202_);
  nor (_21357_, _21356_, _21240_);
  nand (_21358_, _21219_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  nand (_21359_, _21358_, _21208_);
  nand (_21360_, _21221_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  nand (_21361_, _21261_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  nand (_21362_, _21361_, _21360_);
  nor (_21363_, _21362_, _21359_);
  not (_21364_, _21363_);
  nor (_21365_, _21364_, _21357_);
  nor (_21366_, _21365_, _21248_);
  nor (_21367_, _21308_, _21247_);
  nor (_21368_, _21367_, _21366_);
  nor (_21370_, _21368_, _21231_);
  nor (_21371_, _21370_, _21354_);
  not (_21372_, _21371_);
  nor (_21373_, _21372_, _21325_);
  not (_21374_, _21373_);
  nor (_21375_, _21290_, _21240_);
  nand (_21376_, _21375_, _21355_);
  nand (_21377_, _21363_, _21376_);
  nor (_21378_, _21377_, _21227_);
  not (_21379_, _21378_);
  nor (_21380_, _21268_, _21247_);
  not (_21381_, _21380_);
  nor (_21382_, _21381_, _21231_);
  not (_21383_, _21382_);
  nor (_21384_, _21383_, _21336_);
  not (_21385_, _21384_);
  nor (_21386_, _21385_, _21379_);
  not (_21388_, _21386_);
  nor (_21389_, _21388_, _21374_);
  nor (_21390_, _21389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  not (_21391_, _21389_);
  nor (_21392_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  not (_21393_, \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_21394_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _21393_);
  nor (_21395_, _21394_, _21392_);
  not (_21396_, _21395_);
  not (_21397_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_21398_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  not (_21400_, _21398_);
  nor (_21401_, _21400_, _21397_);
  not (_21403_, _21401_);
  nand (_21404_, _21403_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_21406_, _21404_, _21396_);
  nand (_21407_, \oc8051_top_1.oc8051_ram_top1.bit_select [2], \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_21409_, _21407_, _21400_);
  nand (_21410_, _21409_, ABINPUT[0]);
  nand (_21411_, _21232_, ABINPUT[7]);
  nand (_21412_, _21411_, _21410_);
  nor (_21413_, _21412_, _21406_);
  nor (_21414_, _21413_, _21231_);
  nor (_21417_, _21414_, _21391_);
  nor (_19577_, _21417_, _21390_);
  nor (_21418_, _21323_, _21288_);
  not (_21419_, _21418_);
  not (_21420_, _21354_);
  not (_21421_, _21370_);
  nor (_21422_, _21421_, _21420_);
  not (_21423_, _21422_);
  nor (_21424_, _21423_, _21419_);
  not (_21425_, _21424_);
  nor (_21426_, _21365_, _21227_);
  not (_21427_, _21426_);
  nor (_21428_, _21427_, _21385_);
  not (_21429_, _21428_);
  nor (_21430_, _21429_, _21425_);
  nor (_21431_, _21430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  not (_21432_, _21430_);
  nor (_21433_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_21434_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _21393_);
  nor (_21435_, _21434_, _21433_);
  not (_21437_, _21435_);
  not (_21438_, \oc8051_top_1.oc8051_ram_top1.bit_select [0]);
  nor (_21439_, _21438_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  not (_21440_, _21439_);
  nor (_21441_, _21440_, _21397_);
  not (_21442_, _21441_);
  nand (_21443_, _21442_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_21444_, _21443_, _21437_);
  nor (_21445_, _21440_, _21407_);
  nand (_21446_, _21445_, ABINPUT[0]);
  nand (_21448_, _21232_, ABINPUT[8]);
  nand (_21449_, _21448_, _21446_);
  nor (_21450_, _21449_, _21444_);
  nor (_21451_, _21450_, _21231_);
  nor (_21452_, _21451_, _21432_);
  nor (_22384_, _21452_, _21431_);
  nor (_21453_, _21430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  nor (_21454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_21455_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _21393_);
  nor (_21456_, _21455_, _21454_);
  not (_21458_, _21456_);
  nor (_21459_, _21440_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_21461_, _21459_);
  nand (_21462_, _21461_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_21464_, _21462_, _21458_);
  nor (_21465_, \oc8051_top_1.oc8051_ram_top1.bit_select [2], _21232_);
  not (_21466_, _21465_);
  nor (_21467_, _21466_, _21440_);
  nand (_21468_, _21467_, ABINPUT[0]);
  nand (_21469_, _21232_, ABINPUT[4]);
  nand (_21472_, _21469_, _21468_);
  nor (_21473_, _21472_, _21464_);
  nor (_21474_, _21473_, _21231_);
  nor (_21475_, _21474_, _21432_);
  nor (_03003_, _21475_, _21453_);
  not (_21476_, _21323_);
  nor (_21477_, _21476_, _21289_);
  not (_21478_, _21477_);
  nor (_21479_, _21421_, _21354_);
  not (_21480_, _21479_);
  nor (_21481_, _21480_, _21478_);
  not (_21482_, _21481_);
  nor (_21483_, _21482_, _21429_);
  nor (_21484_, _21483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  not (_21485_, _21483_);
  nor (_21486_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_21487_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _21393_);
  nor (_21488_, _21487_, _21486_);
  not (_21490_, _21488_);
  not (_21491_, \oc8051_top_1.oc8051_ram_top1.bit_select [1]);
  nor (_21493_, \oc8051_top_1.oc8051_ram_top1.bit_select [0], _21491_);
  not (_21494_, _21493_);
  nor (_21495_, _21494_, _21397_);
  not (_21496_, _21495_);
  nand (_21497_, _21496_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_21498_, _21497_, _21490_);
  nor (_21499_, _21494_, _21407_);
  nand (_21500_, _21499_, ABINPUT[0]);
  nand (_21501_, _21232_, ABINPUT[9]);
  nand (_21502_, _21501_, _21500_);
  nor (_21503_, _21502_, _21498_);
  nor (_21504_, _21503_, _21231_);
  nor (_21505_, _21504_, _21485_);
  nor (_10367_, _21505_, _21484_);
  nor (_21506_, _21389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  not (_21507_, ABINPUT[0]);
  nor (_21508_, _21438_, _21491_);
  nand (_21510_, _21465_, _21508_);
  nor (_21511_, _21510_, _21507_);
  nor (_21512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_21514_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _21393_);
  nor (_21515_, _21514_, _21512_);
  not (_21517_, _21515_);
  not (_21518_, _21508_);
  nor (_21519_, _21518_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  nor (_21520_, _21519_, _21517_);
  nor (_21521_, _21520_, _21232_);
  nor (_21523_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r , ABINPUT[6]);
  nor (_21524_, _21523_, _21521_);
  nor (_21525_, _21524_, _21511_);
  nor (_21526_, _21525_, _21231_);
  nor (_21528_, _21526_, _21391_);
  nor (_20896_, _21528_, _21506_);
  nor (_21529_, _21480_, _21325_);
  not (_21530_, _21529_);
  nor (_21531_, _21530_, _21429_);
  nor (_21532_, _21531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  not (_21533_, _21531_);
  nor (_21534_, _21533_, _21451_);
  nor (_21018_, _21534_, _21532_);
  nor (_21536_, _21531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  nor (_21537_, _21533_, _21526_);
  nor (_25256_, _21537_, _21536_);
  nor (_21538_, _21389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  nor (_21540_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_21541_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _21393_);
  nor (_21542_, _21541_, _21540_);
  not (_21544_, _21542_);
  nor (_21545_, _21494_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_21546_, _21545_);
  nand (_21547_, _21546_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_21548_, _21547_, _21544_);
  nor (_21549_, _21466_, _21494_);
  nand (_21550_, _21549_, ABINPUT[0]);
  nand (_21551_, _21232_, ABINPUT[5]);
  nand (_21552_, _21551_, _21550_);
  nor (_21553_, _21552_, _21548_);
  nor (_21554_, _21553_, _21231_);
  nor (_21555_, _21554_, _21391_);
  nor (_21061_, _21555_, _21538_);
  nor (_21557_, _21480_, _21419_);
  not (_21558_, _21557_);
  nor (_21559_, _21558_, _21429_);
  nor (_21560_, _21559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  not (_21561_, _21559_);
  nor (_21562_, _21561_, _21414_);
  nor (_21091_, _21562_, _21560_);
  nor (_21563_, _21370_, _21420_);
  not (_21564_, _21563_);
  nor (_21565_, _21564_, _21478_);
  not (_21566_, _21565_);
  nor (_21567_, _21566_, _21429_);
  nor (_21568_, _21567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  not (_21569_, _21567_);
  nor (_21570_, _21569_, _21451_);
  nor (_21415_, _21570_, _21568_);
  nor (_21571_, _21567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  nand (_21572_, _21232_, ABINPUT[3]);
  nor (_21573_, _21466_, _21400_);
  nand (_21574_, _21573_, ABINPUT[0]);
  nand (_21576_, _21574_, _21572_);
  nor (_21577_, _21400_, \oc8051_top_1.oc8051_ram_top1.bit_select [2]);
  not (_21578_, _21577_);
  nand (_21579_, _21578_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_21580_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], \oc8051_top_1.oc8051_ram_top1.rd_en_r );
  nor (_21581_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _21393_);
  nor (_21582_, _21581_, _21580_);
  not (_21583_, _21582_);
  nor (_21584_, _21583_, _21579_);
  nor (_21585_, _21584_, _21576_);
  nor (_21586_, _21585_, _21231_);
  nor (_21587_, _21586_, _21569_);
  nor (_22154_, _21587_, _21571_);
  nor (_21588_, _21564_, _21325_);
  not (_21589_, _21588_);
  nor (_21590_, _21589_, _21429_);
  nor (_21591_, _21590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  not (_21592_, _21590_);
  nor (_21593_, _21592_, _21414_);
  nor (_22554_, _21593_, _21591_);
  nor (_21596_, _21476_, _21288_);
  not (_21597_, _21596_);
  nor (_21598_, _21597_, _21564_);
  not (_21599_, _21598_);
  nor (_21600_, _21599_, _21429_);
  nor (_21601_, _21600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  not (_21602_, _21600_);
  nor (_21603_, _21602_, _21504_);
  nor (_23451_, _21603_, _21601_);
  nor (_21604_, _21600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  nor (_21605_, _21602_, _21414_);
  nor (_23633_, _21605_, _21604_);
  nor (_21606_, _21597_, _21480_);
  not (_21607_, _21606_);
  nor (_21608_, _21607_, _21429_);
  nor (_21609_, _21608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  not (_21610_, _21608_);
  nor (_21611_, \oc8051_top_1.oc8051_ram_top1.rd_en_r , \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nor (_21612_, _21393_, \oc8051_top_1.oc8051_ram_top1.wr_data_r [7]);
  nor (_21613_, _21612_, _21611_);
  not (_21614_, _21613_);
  nor (_21615_, _21518_, _21397_);
  not (_21616_, _21615_);
  nand (_21617_, _21616_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  nor (_21618_, _21617_, _21614_);
  nor (_21619_, _21518_, _21407_);
  nand (_21620_, _21619_, ABINPUT[0]);
  nand (_21621_, ABINPUT[10], _21232_);
  nand (_21622_, _21621_, _21620_);
  nor (_21623_, _21622_, _21618_);
  nor (_21626_, _21623_, _21231_);
  nor (_21627_, _21626_, _21610_);
  nor (_24106_, _21627_, _21609_);
  nor (_21629_, _21597_, _21423_);
  not (_21631_, _21629_);
  nor (_21632_, _21631_, _21429_);
  nor (_21634_, _21632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  not (_21635_, _21632_);
  nor (_21636_, _21635_, _21586_);
  nor (_24338_, _21636_, _21634_);
  nor (_21637_, _21419_, _21372_);
  not (_21638_, _21637_);
  nor (_21639_, _21336_, _21247_);
  nor (_21640_, _21639_, _21231_);
  not (_21641_, _21640_);
  nor (_21642_, _21641_, _21382_);
  not (_21643_, _21642_);
  nor (_21644_, _21643_, _21427_);
  not (_21645_, _21644_);
  nor (_21646_, _21645_, _21638_);
  nor (_21647_, _21646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  not (_21648_, _21646_);
  nor (_21649_, _21648_, _21626_);
  nor (_00635_, _21649_, _21647_);
  nor (_21651_, _21478_, _21423_);
  not (_21652_, _21651_);
  nor (_21653_, _21652_, _21429_);
  nor (_21654_, _21653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  not (_21655_, _21653_);
  nor (_21656_, _21655_, _21451_);
  nor (_25270_, _21656_, _21654_);
  nor (_21657_, _21597_, _21372_);
  not (_21658_, _21657_);
  nor (_21659_, _21658_, _21388_);
  nor (_21660_, _21659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  not (_21661_, _21659_);
  nor (_21662_, _21661_, _21554_);
  nor (_01751_, _21662_, _21660_);
  nor (_21663_, _21632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  nor (_21664_, _21635_, _21554_);
  nor (_02301_, _21664_, _21663_);
  nor (_21666_, _21430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  nor (_21667_, _21626_, _21432_);
  nor (_02483_, _21667_, _21666_);
  nor (_21668_, _21430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  nor (_21669_, _21526_, _21432_);
  nor (_02651_, _21669_, _21668_);
  nor (_21670_, _21483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  nor (_21671_, _21554_, _21485_);
  nor (_03577_, _21671_, _21670_);
  nor (_21672_, _21531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  nor (_21673_, _21626_, _21533_);
  nor (_25258_, _21673_, _21672_);
  nor (_21674_, _21559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  nor (_21675_, _21561_, _21474_);
  nor (_04410_, _21675_, _21674_);
  nor (_21677_, _21567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  nor (_21678_, _21569_, _21554_);
  nor (_04956_, _21678_, _21677_);
  nor (_21679_, _21590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  nor (_21681_, _21592_, _21504_);
  nor (_25253_, _21681_, _21679_);
  nor (_21682_, _21608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  nor (_21683_, _21610_, _21474_);
  nor (_06469_, _21683_, _21682_);
  nor (_21684_, _21646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  nor (_21685_, _21648_, _21586_);
  nor (_06997_, _21685_, _21684_);
  nor (_21686_, _21653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  nor (_21687_, _21655_, _21474_);
  nor (_07190_, _21687_, _21686_);
  nor (_21688_, _21423_, _21325_);
  not (_21689_, _21688_);
  nor (_21690_, _21689_, _21429_);
  nor (_21691_, _21690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  not (_21692_, _21690_);
  nor (_21693_, _21692_, _21554_);
  nor (_07486_, _21693_, _21691_);
  nor (_21694_, _21643_, _21379_);
  not (_21695_, _21694_);
  nor (_21697_, _21695_, _21425_);
  nor (_21698_, _21697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  not (_21699_, _21697_);
  nor (_21700_, _21699_, _21526_);
  nor (_08454_, _21700_, _21698_);
  nor (_21701_, _21559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  nor (_21702_, _21561_, _21451_);
  nor (_08929_, _21702_, _21701_);
  nor (_21703_, _21567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  nor (_21704_, _21569_, _21504_);
  nor (_09148_, _21704_, _21703_);
  nor (_21706_, _21659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  nor (_21707_, _21661_, _21451_);
  nor (_25121_, _21707_, _21706_);
  nor (_21708_, _21590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  nor (_21709_, _21592_, _21586_);
  nor (_09528_, _21709_, _21708_);
  nor (_21711_, _21608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  nor (_21712_, _21610_, _21554_);
  nor (_09726_, _21712_, _21711_);
  nor (_21714_, _21659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  nor (_21716_, _21661_, _21414_);
  nor (_09923_, _21716_, _21714_);
  nor (_21717_, _21632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  nor (_21718_, _21635_, _21526_);
  nor (_10116_, _21718_, _21717_);
  nor (_21719_, _21590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  nor (_21720_, _21626_, _21592_);
  nor (_10441_, _21720_, _21719_);
  nor (_21722_, _21531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  nor (_21723_, _21586_, _21533_);
  nor (_10576_, _21723_, _21722_);
  nor (_21724_, _21559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  nor (_21725_, _21561_, _21504_);
  nor (_11258_, _21725_, _21724_);
  nor (_21726_, _21697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  nor (_21727_, _21699_, _21451_);
  nor (_11410_, _21727_, _21726_);
  nor (_21728_, _21658_, _21429_);
  nor (_21729_, _21728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  not (_21731_, _21728_);
  nor (_21732_, _21731_, _21414_);
  nor (_13311_, _21732_, _21729_);
  nor (_21733_, _21638_, _21429_);
  nor (_21734_, _21733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  not (_21735_, _21733_);
  nor (_21736_, _21735_, _21586_);
  nor (_13642_, _21736_, _21734_);
  nor (_21737_, _21427_, _21231_);
  nor (_21738_, _21640_, _21382_);
  nand (_21739_, _21738_, _21737_);
  nor (_21741_, _21739_, _21652_);
  nor (_21742_, _21741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  not (_21744_, _21741_);
  nor (_21745_, _21744_, _21526_);
  nor (_13930_, _21745_, _21742_);
  nor (_21747_, _21739_, _21631_);
  nor (_21748_, _21747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  not (_21749_, _21747_);
  nor (_21750_, _21749_, _21451_);
  nor (_14445_, _21750_, _21748_);
  nor (_21752_, _21739_, _21425_);
  nor (_21753_, _21752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  not (_21754_, _21752_);
  nor (_21756_, _21754_, _21626_);
  nor (_14712_, _21756_, _21753_);
  nor (_21757_, _21739_, _21530_);
  nor (_21758_, _21757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  not (_21759_, _21757_);
  nor (_21760_, _21759_, _21414_);
  nor (_15202_, _21760_, _21758_);
  nor (_21761_, _21739_, _21566_);
  nor (_21762_, _21761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  not (_21763_, _21761_);
  nor (_21764_, _21763_, _21554_);
  nor (_15777_, _21764_, _21762_);
  nor (_21766_, _21739_, _21638_);
  nor (_21767_, _21766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  not (_21768_, _21766_);
  nor (_21769_, _21768_, _21526_);
  nor (_17169_, _21769_, _21767_);
  nor (_21771_, _21377_, _21337_);
  not (_21772_, _21771_);
  nor (_21773_, _21772_, _21227_);
  not (_21774_, _21773_);
  nor (_21775_, _21774_, _21383_);
  not (_21776_, _21775_);
  nor (_21777_, _21776_, _21652_);
  nor (_21778_, _21777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  not (_21779_, _21777_);
  nor (_21780_, _21779_, _21504_);
  nor (_17464_, _21780_, _21778_);
  nor (_21782_, _21776_, _21689_);
  nor (_21783_, _21782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  not (_21784_, _21782_);
  nor (_21785_, _21784_, _21474_);
  nor (_18078_, _21785_, _21783_);
  nor (_21786_, _21776_, _21631_);
  nor (_21787_, _21786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  not (_21788_, _21786_);
  nor (_21789_, _21788_, _21451_);
  nor (_25214_, _21789_, _21787_);
  nor (_21790_, _21776_, _21425_);
  nor (_21791_, _21790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  not (_21792_, _21790_);
  nor (_21794_, _21792_, _21554_);
  nor (_18979_, _21794_, _21791_);
  nor (_21796_, _21776_, _21558_);
  nor (_21798_, _21796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  not (_21799_, _21796_);
  nor (_21801_, _21799_, _21414_);
  nor (_19290_, _21801_, _21798_);
  nor (_21804_, _21776_, _21566_);
  nor (_21805_, _21804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  not (_21806_, _21804_);
  nor (_21808_, _21806_, _21504_);
  nor (_19578_, _21808_, _21805_);
  nor (_21810_, _21776_, _21589_);
  nor (_21811_, _21810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  not (_21812_, _21810_);
  nor (_21814_, _21812_, _21554_);
  nor (_20168_, _21814_, _21811_);
  nor (_21816_, _21776_, _21599_);
  nor (_21817_, _21816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  not (_21818_, _21816_);
  nor (_21819_, _21818_, _21414_);
  nor (_20470_, _21819_, _21817_);
  nor (_21820_, _21564_, _21419_);
  not (_21821_, _21820_);
  nor (_21822_, _21821_, _21776_);
  nor (_21823_, _21822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  not (_21824_, _21822_);
  nor (_21825_, _21824_, _21526_);
  nor (_20866_, _21825_, _21823_);
  nor (_21826_, _21389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  nor (_21827_, _21626_, _21391_);
  nor (_25122_, _21827_, _21826_);
  nor (_21829_, _21776_, _21374_);
  nor (_21830_, _21829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  not (_21831_, _21829_);
  nor (_21832_, _21831_, _21504_);
  nor (_20879_, _21832_, _21830_);
  nor (_21834_, _21776_, _21658_);
  nor (_21835_, _21834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  not (_21836_, _21834_);
  nor (_21837_, _21836_, _21451_);
  nor (_20894_, _21837_, _21835_);
  nor (_21838_, _21834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  nor (_21839_, _21836_, _21586_);
  nor (_20898_, _21839_, _21838_);
  nor (_21842_, _21776_, _21638_);
  nor (_21843_, _21842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  not (_21844_, _21842_);
  nor (_21846_, _21844_, _21414_);
  nor (_20909_, _21846_, _21843_);
  nor (_21847_, _21389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  nor (_21849_, _21504_, _21391_);
  nor (_20914_, _21849_, _21847_);
  nor (_21850_, _21695_, _21652_);
  nor (_21852_, _21850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  not (_21853_, _21850_);
  nor (_21855_, _21853_, _21451_);
  nor (_20923_, _21855_, _21852_);
  nor (_21856_, _21776_, _21607_);
  nor (_21857_, _21856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  not (_21858_, _21856_);
  nor (_21859_, _21858_, _21526_);
  nor (_20947_, _21859_, _21857_);
  nor (_21860_, _21810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  nor (_21861_, _21812_, _21526_);
  nor (_20953_, _21861_, _21860_);
  nor (_21863_, _21478_, _21372_);
  not (_21864_, _21863_);
  nor (_21865_, _21864_, _21429_);
  nor (_21866_, _21865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  not (_21867_, _21865_);
  nor (_21868_, _21867_, _21554_);
  nor (_20962_, _21868_, _21866_);
  nor (_21869_, _21739_, _21689_);
  nor (_21870_, _21869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  not (_21871_, _21869_);
  nor (_21872_, _21871_, _21414_);
  nor (_20964_, _21872_, _21870_);
  nor (_21873_, _21739_, _21482_);
  nor (_21874_, _21873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  not (_21875_, _21873_);
  nor (_21876_, _21875_, _21554_);
  nor (_20979_, _21876_, _21874_);
  nor (_21877_, _21739_, _21607_);
  nor (_21878_, _21877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  not (_21880_, _21877_);
  nor (_21881_, _21880_, _21504_);
  nor (_20987_, _21881_, _21878_);
  nor (_21882_, _21739_, _21589_);
  nor (_21883_, _21882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  not (_21884_, _21882_);
  nor (_21885_, _21884_, _21504_);
  nor (_25226_, _21885_, _21883_);
  nor (_21887_, _21864_, _21739_);
  nor (_21889_, _21887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  not (_21891_, _21887_);
  nor (_21892_, _21891_, _21526_);
  nor (_20992_, _21892_, _21889_);
  nor (_21893_, _21739_, _21658_);
  nor (_21894_, _21893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  not (_21895_, _21893_);
  nor (_21897_, _21895_, _21526_);
  nor (_21001_, _21897_, _21894_);
  nor (_21899_, _21864_, _21388_);
  nor (_21900_, _21899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  not (_21902_, _21899_);
  nor (_21903_, _21902_, _21474_);
  nor (_21019_, _21903_, _21900_);
  nor (_21904_, _21864_, _21776_);
  nor (_21905_, _21904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  not (_21906_, _21904_);
  nor (_21907_, _21906_, _21554_);
  nor (_21021_, _21907_, _21905_);
  nor (_21910_, _21829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  nor (_21911_, _21831_, _21554_);
  nor (_21022_, _21911_, _21910_);
  nor (_21913_, _21776_, _21482_);
  nor (_21914_, _21913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  not (_21915_, _21913_);
  nor (_21917_, _21915_, _21414_);
  nor (_21027_, _21917_, _21914_);
  nor (_21919_, _21776_, _21530_);
  nor (_21920_, _21919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  not (_21922_, _21919_);
  nor (_21923_, _21922_, _21626_);
  nor (_21029_, _21923_, _21920_);
  nor (_21926_, _21856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  nor (_21928_, _21858_, _21626_);
  nor (_21030_, _21928_, _21926_);
  nor (_21929_, _21728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  nor (_21930_, _21731_, _21451_);
  nor (_21031_, _21930_, _21929_);
  nor (_21931_, _21810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  nor (_21932_, _21812_, _21414_);
  nor (_21032_, _21932_, _21931_);
  nor (_21933_, _21739_, _21558_);
  nor (_21934_, _21933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  not (_21935_, _21933_);
  nor (_21937_, _21935_, _21586_);
  nor (_21033_, _21937_, _21934_);
  nor (_21938_, _21739_, _21599_);
  nor (_21939_, _21938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  not (_21940_, _21938_);
  nor (_21942_, _21940_, _21586_);
  nor (_21036_, _21942_, _21939_);
  nor (_21943_, _21899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  nor (_21944_, _21902_, _21586_);
  nor (_21038_, _21944_, _21943_);
  nor (_21945_, _21782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  nor (_21946_, _21784_, _21554_);
  nor (_21040_, _21946_, _21945_);
  nor (_21947_, _21697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  nor (_21948_, _21699_, _21626_);
  nor (_25188_, _21948_, _21947_);
  nor (_21949_, _21821_, _21429_);
  nor (_21951_, _21949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  not (_21952_, _21949_);
  nor (_21954_, _21952_, _21451_);
  nor (_21053_, _21954_, _21951_);
  nor (_21955_, _21893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  nor (_21956_, _21895_, _21414_);
  nor (_21064_, _21956_, _21955_);
  nor (_21957_, _21913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  nor (_21958_, _21915_, _21451_);
  nor (_21066_, _21958_, _21957_);
  nor (_21959_, _21933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  nor (_21960_, _21935_, _21474_);
  nor (_21068_, _21960_, _21959_);
  nor (_21961_, _21856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  nor (_21962_, _21858_, _21586_);
  nor (_21088_, _21962_, _21961_);
  nor (_21963_, _21856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  nor (_21964_, _21858_, _21504_);
  nor (_21090_, _21964_, _21963_);
  nor (_21965_, _21919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  nor (_21966_, _21922_, _21554_);
  nor (_25210_, _21966_, _21965_);
  nor (_21967_, _21919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  nor (_21968_, _21922_, _21474_);
  nor (_21092_, _21968_, _21967_);
  nor (_21969_, _21919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  nor (_21970_, _21922_, _21504_);
  nor (_21094_, _21970_, _21969_);
  nor (_21971_, _21919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  nor (_21972_, _21922_, _21451_);
  nor (_21095_, _21972_, _21971_);
  nor (_21973_, _21913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  nor (_21974_, _21915_, _21586_);
  nor (_21097_, _21974_, _21973_);
  nor (_21975_, _21913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  nor (_21976_, _21915_, _21526_);
  nor (_21098_, _21976_, _21975_);
  nor (_21977_, _21822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  nor (_21978_, _21824_, _21504_);
  nor (_21110_, _21978_, _21977_);
  nor (_21979_, _21842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  nor (_21980_, _21844_, _21554_);
  nor (_25198_, _21980_, _21979_);
  nor (_21981_, _21842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  nor (_21982_, _21844_, _21504_);
  nor (_21117_, _21982_, _21981_);
  nor (_21983_, _21834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  nor (_21984_, _21836_, _21526_);
  nor (_21118_, _21984_, _21983_);
  nor (_21985_, _21829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  nor (_21986_, _21831_, _21474_);
  nor (_21119_, _21986_, _21985_);
  nor (_21987_, _21829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  nor (_21988_, _21831_, _21526_);
  nor (_21128_, _21988_, _21987_);
  nor (_21989_, _21904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  nor (_21990_, _21906_, _21474_);
  nor (_25201_, _21990_, _21989_);
  nor (_21991_, _21904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  nor (_21992_, _21906_, _21504_);
  nor (_21132_, _21992_, _21991_);
  nor (_21993_, _21904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  nor (_21994_, _21906_, _21414_);
  nor (_21133_, _21994_, _21993_);
  not (_21995_, _21738_);
  nand (_21996_, _21377_, _21248_);
  nor (_21997_, _21996_, _21231_);
  not (_21998_, _21997_);
  nor (_21999_, _21998_, _21246_);
  not (_22000_, _21999_);
  nor (_22002_, _22000_, _21995_);
  not (_22003_, _22002_);
  nor (_22004_, _22003_, _21530_);
  nor (_22005_, _22004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  not (_22006_, _22004_);
  nor (_22007_, _22006_, _21414_);
  nor (_25411_, _22007_, _22005_);
  nor (_22008_, _21822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  nor (_22009_, _21824_, _21586_);
  nor (_21137_, _22009_, _22008_);
  nor (_22010_, _21822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  nor (_22011_, _21824_, _21626_);
  nor (_21138_, _22011_, _22010_);
  nor (_22012_, _21822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  nor (_22013_, _21824_, _21451_);
  nor (_21139_, _22013_, _22012_);
  nor (_22014_, _22004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  nor (_22015_, _22006_, _21526_);
  nor (_21146_, _22015_, _22014_);
  nor (_22016_, _21383_, _21337_);
  not (_22018_, _22016_);
  nor (_22019_, _22000_, _22018_);
  not (_22020_, _22019_);
  nor (_22021_, _22020_, _21658_);
  nor (_22022_, _22021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  not (_22023_, _22021_);
  nor (_22024_, _22023_, _21451_);
  nor (_21172_, _22024_, _22022_);
  nor (_22025_, _21796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  nor (_22026_, _21799_, _21474_);
  nor (_21173_, _22026_, _22025_);
  nor (_22027_, _21913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  nor (_22028_, _21915_, _21626_);
  nor (_21177_, _22028_, _22027_);
  nor (_22029_, _21790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  nor (_22030_, _21792_, _21626_);
  nor (_25213_, _22030_, _22029_);
  nor (_22031_, _21786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  nor (_22032_, _21788_, _21554_);
  nor (_21180_, _22032_, _22031_);
  nor (_22034_, _21786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  nor (_22035_, _21788_, _21626_);
  nor (_21181_, _22035_, _22034_);
  nor (_22036_, _21782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  nor (_22037_, _21784_, _21626_);
  nor (_21182_, _22037_, _22036_);
  nor (_22038_, _21777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  nor (_22039_, _21779_, _21554_);
  nor (_21265_, _22039_, _22038_);
  nor (_22040_, _21893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  nor (_22041_, _21895_, _21554_);
  nor (_21317_, _22041_, _22040_);
  nor (_22042_, _21739_, _21374_);
  nor (_22043_, _22042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  not (_22044_, _22042_);
  nor (_22045_, _22044_, _21554_);
  nor (_21369_, _22045_, _22043_);
  nor (_22046_, _21887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  nor (_22047_, _21891_, _21554_);
  nor (_21416_, _22047_, _22046_);
  nor (_22048_, _22000_, _21643_);
  not (_22049_, _22048_);
  nor (_22050_, _22049_, _21658_);
  nor (_22051_, _22050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  not (_22052_, _22050_);
  nor (_22053_, _22052_, _21414_);
  nor (_21436_, _22053_, _22051_);
  nor (_22054_, _21821_, _21739_);
  nor (_22055_, _22054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  not (_22056_, _22054_);
  nor (_22058_, _22056_, _21586_);
  nor (_21470_, _22058_, _22055_);
  nor (_22059_, _22050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  nor (_22060_, _22052_, _21504_);
  nor (_25447_, _22060_, _22059_);
  nor (_22061_, _22054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  nor (_22062_, _22056_, _21626_);
  nor (_21513_, _22062_, _22061_);
  nor (_22063_, _21938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  nor (_22064_, _21940_, _21626_);
  nor (_21535_, _22064_, _22063_);
  nor (_22065_, _21882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  nor (_22066_, _21884_, _21451_);
  nor (_21556_, _22066_, _22065_);
  nor (_22067_, _21882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  nor (_22068_, _21884_, _21474_);
  nor (_21575_, _22068_, _22067_);
  nor (_22069_, _22049_, _21374_);
  nor (_22070_, _22069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  not (_22071_, _22069_);
  nor (_22072_, _22071_, _21474_);
  nor (_21595_, _22072_, _22070_);
  nor (_22073_, _21761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  nor (_22074_, _21763_, _21626_);
  nor (_21624_, _22074_, _22073_);
  nor (_22075_, _21761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  nor (_22076_, _21763_, _21414_);
  nor (_25227_, _22076_, _22075_);
  nor (_22077_, _21933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  nor (_22078_, _21935_, _21626_);
  nor (_21665_, _22078_, _22077_);
  nor (_22080_, _21933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  nor (_22081_, _21935_, _21414_);
  nor (_21680_, _22081_, _22080_);
  nor (_22082_, _21877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  nor (_22083_, _21880_, _21451_);
  nor (_21696_, _22083_, _22082_);
  nor (_22084_, _22069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  nor (_22085_, _22071_, _21526_);
  nor (_21713_, _22085_, _22084_);
  nor (_22086_, _22069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  nor (_22087_, _22071_, _21451_);
  nor (_21730_, _22087_, _22086_);
  nor (_22088_, _21873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  nor (_22090_, _21875_, _21474_);
  nor (_21751_, _22090_, _22088_);
  nor (_22091_, _21757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  nor (_22092_, _21759_, _21626_);
  nor (_25234_, _22092_, _22091_);
  nor (_22094_, _21752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  nor (_22096_, _21754_, _21586_);
  nor (_25235_, _22096_, _22094_);
  nor (_22098_, _21752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  nor (_22099_, _21754_, _21526_);
  nor (_21840_, _22099_, _22098_);
  nor (_22100_, _22069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  nor (_22101_, _22071_, _21504_);
  nor (_21862_, _22101_, _22100_);
  nor (_22102_, _21747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  nor (_22103_, _21749_, _21554_);
  nor (_21879_, _22103_, _22102_);
  nor (_22105_, _21869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  nor (_22106_, _21871_, _21526_);
  nor (_21901_, _22106_, _22105_);
  nor (_22108_, _21869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  nor (_22109_, _21871_, _21586_);
  nor (_21924_, _22109_, _22108_);
  nor (_22111_, _22000_, _21385_);
  not (_22113_, _22111_);
  nor (_22114_, _22113_, _21631_);
  nor (_22115_, _22114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  not (_22116_, _22114_);
  nor (_22117_, _22116_, _21626_);
  nor (_25438_, _22117_, _22115_);
  nor (_22118_, _21733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  nor (_22119_, _21735_, _21626_);
  nor (_22001_, _22119_, _22118_);
  nor (_22121_, _22113_, _21689_);
  nor (_22122_, _22121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  not (_22123_, _22121_);
  nor (_22124_, _22123_, _21586_);
  nor (_22017_, _22124_, _22122_);
  nor (_22125_, _22121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  nor (_22126_, _22123_, _21554_);
  nor (_22033_, _22126_, _22125_);
  nor (_22127_, _21429_, _21374_);
  nor (_22128_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  not (_22130_, _22127_);
  nor (_22131_, _22130_, _21526_);
  nor (_22057_, _22131_, _22128_);
  nor (_22132_, _21865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  nor (_22133_, _21867_, _21474_);
  nor (_22079_, _22133_, _22132_);
  nor (_22134_, _22121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  nor (_22135_, _22123_, _21414_);
  nor (_22095_, _22135_, _22134_);
  nor (_22136_, _21865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  nor (_22137_, _21867_, _21626_);
  nor (_25248_, _22137_, _22136_);
  nor (_22138_, _22121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  nor (_22139_, _22123_, _21504_);
  nor (_25439_, _22139_, _22138_);
  nor (_22140_, _21695_, _21631_);
  nor (_22141_, _22140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  not (_22142_, _22140_);
  nor (_22143_, _22142_, _21474_);
  nor (_22171_, _22143_, _22141_);
  nor (_22144_, _22140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  nor (_22145_, _22142_, _21526_);
  nor (_25190_, _22145_, _22144_);
  nor (_22146_, _21804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  nor (_22147_, _21806_, _21414_);
  nor (_22445_, _22147_, _22146_);
  nor (_22148_, _21804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  nor (_22149_, _21806_, _21451_);
  nor (_25207_, _22149_, _22148_);
  nor (_22150_, _22113_, _21652_);
  nor (_22151_, _22150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  not (_22152_, _22150_);
  nor (_22153_, _22152_, _21474_);
  nor (_22662_, _22153_, _22151_);
  nor (_22155_, _22150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  nor (_22156_, _22152_, _21526_);
  nor (_22704_, _22156_, _22155_);
  nor (_22158_, _21804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  nor (_22159_, _21806_, _21526_);
  nor (_22746_, _22159_, _22158_);
  nor (_22160_, _22150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  nor (_22161_, _22152_, _21504_);
  nor (_22913_, _22161_, _22160_);
  nor (_22162_, _22020_, _21589_);
  nor (_22164_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  not (_22165_, _22162_);
  nor (_22166_, _22165_, _21474_);
  nor (_25070_, _22166_, _22164_);
  nor (_22167_, _22150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  nor (_22168_, _22152_, _21626_);
  nor (_23254_, _22168_, _22167_);
  nor (_22169_, _21804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  nor (_22170_, _21806_, _21474_);
  nor (_23463_, _22170_, _22169_);
  nor (_22172_, _21804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  nor (_22173_, _21806_, _21554_);
  nor (_23559_, _22173_, _22172_);
  nor (_22174_, _21804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  nor (_22175_, _21806_, _21586_);
  nor (_23576_, _22175_, _22174_);
  nor (_22176_, _22049_, _21638_);
  nor (_22178_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  not (_22179_, _22176_);
  nor (_22180_, _22179_, _21586_);
  nor (_23665_, _22180_, _22178_);
  nor (_22181_, _21796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  nor (_22182_, _21799_, _21554_);
  nor (_23778_, _22182_, _22181_);
  nor (_22183_, _21796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  nor (_22184_, _21799_, _21526_);
  nor (_23814_, _22184_, _22183_);
  nor (_22186_, _22049_, _21530_);
  nor (_22187_, _22186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  not (_22188_, _22186_);
  nor (_22189_, _22188_, _21626_);
  nor (_23962_, _22189_, _22187_);
  nor (_22190_, _21600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  nor (_22191_, _21602_, _21474_);
  nor (_25251_, _22191_, _22190_);
  nor (_22192_, _21949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  nor (_22193_, _21952_, _21504_);
  nor (_25249_, _22193_, _22192_);
  nor (_22194_, _21949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  nor (_22195_, _21952_, _21626_);
  nor (_25250_, _22195_, _22194_);
  nor (_22196_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  nor (_22197_, _22179_, _21554_);
  nor (_25443_, _22197_, _22196_);
  nor (_22198_, _21695_, _21689_);
  nor (_22199_, _22198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  not (_22200_, _22198_);
  nor (_22201_, _22200_, _21504_);
  nor (_25195_, _22201_, _22199_);
  nor (_22202_, _22198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  nor (_22203_, _22200_, _21474_);
  nor (_25192_, _22203_, _22202_);
  nor (_22204_, _22140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  nor (_22205_, _22142_, _21626_);
  nor (_25191_, _22205_, _22204_);
  nor (_22206_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  nor (_22207_, _22179_, _21414_);
  nor (_25444_, _22207_, _22206_);
  nor (_22208_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  nor (_22209_, _22179_, _21504_);
  nor (_25445_, _22209_, _22208_);
  nor (_22210_, _22140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  nor (_22211_, _22142_, _21554_);
  nor (_25189_, _22211_, _22210_);
  nor (_22212_, _21697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  nor (_22213_, _21699_, _21504_);
  nor (_25187_, _22213_, _22212_);
  nor (_22214_, _21697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  nor (_22215_, _21699_, _21414_);
  nor (_25186_, _22215_, _22214_);
  nor (_22216_, _21697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  nor (_22217_, _21699_, _21586_);
  nor (_25184_, _22217_, _22216_);
  nor (_22219_, _21695_, _21482_);
  nor (_22220_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  not (_22221_, _22219_);
  nor (_22222_, _22221_, _21626_);
  nor (_25183_, _22222_, _22220_);
  nor (_22223_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  nor (_22224_, _22221_, _21451_);
  nor (_25182_, _22224_, _22223_);
  nor (_22225_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  nor (_22226_, _22221_, _21586_);
  nor (_25181_, _22226_, _22225_);
  nor (_22227_, _21695_, _21530_);
  nor (_22228_, _22227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  not (_22229_, _22227_);
  nor (_22230_, _22229_, _21626_);
  nor (_25180_, _22230_, _22228_);
  nor (_22231_, _22227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  nor (_22232_, _22229_, _21451_);
  nor (_25178_, _22232_, _22231_);
  nor (_22233_, _22227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  nor (_22234_, _22229_, _21474_);
  nor (_25176_, _22234_, _22233_);
  nor (_22235_, _22050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  nor (_22236_, _22052_, _21474_);
  nor (_25446_, _22236_, _22235_);
  nor (_22238_, _21695_, _21607_);
  nor (_22239_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  not (_22240_, _22238_);
  nor (_22241_, _22240_, _21504_);
  nor (_25175_, _22241_, _22239_);
  nor (_22242_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  nor (_22243_, _22240_, _21586_);
  nor (_25172_, _22243_, _22242_);
  nor (_22245_, _22049_, _21864_);
  nor (_22246_, _22245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  not (_22248_, _22245_);
  nor (_22249_, _22248_, _21474_);
  nor (_25448_, _22249_, _22246_);
  nor (_22250_, _21695_, _21558_);
  nor (_22251_, _22250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  not (_22252_, _22250_);
  nor (_22253_, _22252_, _21451_);
  nor (_25171_, _22253_, _22251_);
  nor (_22255_, _22245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  nor (_22256_, _22248_, _21526_);
  nor (_25449_, _22256_, _22255_);
  nor (_22257_, _22250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  nor (_22258_, _22252_, _21474_);
  nor (_25170_, _22258_, _22257_);
  nor (_22259_, _21695_, _21566_);
  nor (_22260_, _22259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  not (_22261_, _22259_);
  nor (_22262_, _22261_, _21504_);
  nor (_25169_, _22262_, _22260_);
  nor (_22263_, _21695_, _21599_);
  nor (_22264_, _22263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  not (_22265_, _22263_);
  nor (_22266_, _22265_, _21414_);
  nor (_25161_, _22266_, _22264_);
  nor (_22268_, _22263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  nor (_22269_, _22265_, _21554_);
  nor (_25160_, _22269_, _22268_);
  nor (_22270_, _22245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  nor (_22271_, _22248_, _21451_);
  nor (_25450_, _22271_, _22270_);
  nor (_22272_, _21821_, _21695_);
  nor (_22273_, _22272_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  not (_22274_, _22272_);
  nor (_22275_, _22274_, _21451_);
  nor (_25158_, _22275_, _22273_);
  nor (_22276_, _22272_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  nor (_22277_, _22274_, _21526_);
  nor (_25157_, _22277_, _22276_);
  nor (_22278_, _21864_, _21695_);
  nor (_22279_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  not (_22280_, _22278_);
  nor (_22281_, _22280_, _21626_);
  nor (_25156_, _22281_, _22279_);
  nor (_22282_, _22245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  nor (_22283_, _22248_, _21504_);
  nor (_25451_, _22283_, _22282_);
  nor (_22284_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  nor (_22285_, _22280_, _21554_);
  nor (_25155_, _22285_, _22284_);
  nor (_22286_, _22049_, _21821_);
  nor (_22287_, _22286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  not (_22288_, _22286_);
  nor (_22289_, _22288_, _21586_);
  nor (_25045_, _22289_, _22287_);
  nor (_22290_, _22286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  nor (_22291_, _22288_, _21554_);
  nor (_25046_, _22291_, _22290_);
  nor (_22292_, _21695_, _21374_);
  nor (_22293_, _22292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  not (_22294_, _22292_);
  nor (_22295_, _22294_, _21526_);
  nor (_25153_, _22295_, _22293_);
  nor (_22296_, _22286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  nor (_22297_, _22288_, _21414_);
  nor (_25047_, _22297_, _22296_);
  nor (_22298_, _22259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  nor (_22299_, _22261_, _21474_);
  nor (_25168_, _22299_, _22298_);
  nor (_22300_, _21695_, _21589_);
  nor (_22301_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  not (_22302_, _22300_);
  nor (_22303_, _22302_, _21504_);
  nor (_25166_, _22303_, _22301_);
  nor (_22305_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  nor (_22306_, _22302_, _21554_);
  nor (_25164_, _22306_, _22305_);
  nor (_22307_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  nor (_22308_, _22302_, _21414_);
  nor (_00001_, _22308_, _22307_);
  nor (_22310_, _22198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  nor (_22311_, _22200_, _21526_);
  nor (_25194_, _22311_, _22310_);
  nor (_22312_, _22140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  nor (_22313_, _22142_, _21414_);
  nor (_00087_, _22313_, _22312_);
  nor (_22314_, _22286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  nor (_22315_, _22288_, _21451_);
  nor (_00109_, _22315_, _22314_);
  nor (_22316_, _22049_, _21599_);
  nor (_22317_, _22316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  not (_22318_, _22316_);
  nor (_22319_, _22318_, _21586_);
  nor (_00140_, _22319_, _22317_);
  nor (_22320_, _22316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  nor (_22321_, _22318_, _21474_);
  nor (_00172_, _22321_, _22320_);
  nor (_22322_, _22316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  nor (_22323_, _22318_, _21526_);
  nor (_00193_, _22323_, _22322_);
  nor (_22324_, _22316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  nor (_22325_, _22318_, _21451_);
  nor (_00214_, _22325_, _22324_);
  nor (_22326_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  nor (_22327_, _22240_, _21554_);
  nor (_00236_, _22327_, _22326_);
  nor (_22328_, _22250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  nor (_22329_, _22252_, _21626_);
  nor (_00257_, _22329_, _22328_);
  nor (_22330_, _22250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  nor (_22331_, _22252_, _21526_);
  nor (_00278_, _22331_, _22330_);
  nor (_22332_, _22263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  nor (_22333_, _22265_, _21504_);
  nor (_25163_, _22333_, _22332_);
  nor (_22334_, _22272_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  nor (_22335_, _22274_, _21626_);
  nor (_00330_, _22335_, _22334_);
  nor (_22336_, _22316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  nor (_22337_, _22318_, _21626_);
  nor (_00351_, _22337_, _22336_);
  nor (_22338_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  nor (_22339_, _22280_, _21414_);
  nor (_00392_, _22339_, _22338_);
  nor (_22341_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  nor (_22342_, _22280_, _21586_);
  nor (_00414_, _22342_, _22341_);
  nor (_22343_, _22292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  nor (_22344_, _22294_, _21451_);
  nor (_00436_, _22344_, _22343_);
  nor (_22346_, _22259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  nor (_22347_, _22261_, _21526_);
  nor (_00457_, _22347_, _22346_);
  nor (_22348_, _22049_, _21589_);
  nor (_22349_, _22348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  not (_22351_, _22348_);
  nor (_22352_, _22351_, _21586_);
  nor (_00488_, _22352_, _22349_);
  nor (_22353_, _22198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  nor (_22354_, _22200_, _21626_);
  nor (_00509_, _22354_, _22353_);
  nor (_22355_, _22140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  nor (_22356_, _22142_, _21586_);
  nor (_00530_, _22356_, _22355_);
  nor (_22357_, _21697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  nor (_22358_, _21699_, _21474_);
  nor (_25185_, _22358_, _22357_);
  nor (_22359_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  nor (_22360_, _22221_, _21474_);
  nor (_00571_, _22360_, _22359_);
  nor (_22361_, _22227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  nor (_22362_, _22229_, _21554_);
  nor (_25177_, _22362_, _22361_);
  nor (_22363_, _22348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  nor (_22364_, _22351_, _21554_);
  nor (_00612_, _22364_, _22363_);
  nor (_22365_, _22348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  nor (_22366_, _22351_, _21414_);
  nor (_00636_, _22366_, _22365_);
  nor (_22367_, _22348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  nor (_22368_, _22351_, _21626_);
  nor (_00700_, _22368_, _22367_);
  nor (_22369_, _22049_, _21566_);
  nor (_22370_, _22369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  not (_22371_, _22369_);
  nor (_22372_, _22371_, _21586_);
  nor (_00729_, _22372_, _22370_);
  nor (_22373_, _22369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  nor (_22374_, _22371_, _21554_);
  nor (_00761_, _22374_, _22373_);
  nor (_22376_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  nor (_22377_, _22240_, _21526_);
  nor (_00776_, _22377_, _22376_);
  nor (_22378_, _22263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  nor (_22379_, _22265_, _21626_);
  nor (_00792_, _22379_, _22378_);
  nor (_22380_, _22272_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  nor (_22381_, _22274_, _21586_);
  nor (_00807_, _22381_, _22380_);
  nor (_22382_, _22259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  nor (_22383_, _22261_, _21414_);
  nor (_00823_, _22383_, _22382_);
  nor (_22385_, _22369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  nor (_22386_, _22371_, _21414_);
  nor (_00838_, _22386_, _22385_);
  nor (_22387_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  nor (_22388_, _22221_, _21554_);
  nor (_00854_, _22388_, _22387_);
  nor (_22389_, _21850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  nor (_22390_, _21853_, _21586_);
  nor (_25196_, _22390_, _22389_);
  nor (_22392_, _21231_, _21227_);
  not (_22393_, _22392_);
  nor (_22394_, _22393_, _21377_);
  nand (_22395_, _21738_, _22394_);
  nor (_22396_, _22395_, _21652_);
  nor (_22397_, _22396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  not (_22398_, _22396_);
  nor (_22399_, _22398_, _21414_);
  nor (_00951_, _22399_, _22397_);
  nor (_22401_, _22369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  nor (_22402_, _22371_, _21504_);
  nor (_00972_, _22402_, _22401_);
  nor (_22403_, _22395_, _21631_);
  nor (_22404_, _22403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  not (_22406_, _22403_);
  nor (_22407_, _22406_, _21474_);
  nor (_01024_, _22407_, _22404_);
  nor (_22408_, _22395_, _21530_);
  nor (_22409_, _22408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  not (_22410_, _22408_);
  nor (_22411_, _22410_, _21504_);
  nor (_01082_, _22411_, _22409_);
  nor (_22412_, _22395_, _21607_);
  nor (_22413_, _22412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  not (_22414_, _22412_);
  nor (_22415_, _22414_, _21626_);
  nor (_01109_, _22415_, _22413_);
  nor (_22416_, _22049_, _21558_);
  nor (_22417_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  not (_22418_, _22416_);
  nor (_22420_, _22418_, _21474_);
  nor (_01126_, _22420_, _22417_);
  nor (_22421_, _22395_, _21558_);
  nor (_22422_, _22421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  not (_22423_, _22421_);
  nor (_22424_, _22423_, _21554_);
  nor (_01155_, _22424_, _22422_);
  nor (_22425_, _22395_, _21566_);
  nor (_22426_, _22425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  not (_22427_, _22425_);
  nor (_22428_, _22427_, _21554_);
  nor (_01180_, _22428_, _22426_);
  nor (_22429_, _22395_, _21589_);
  nor (_22430_, _22429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  not (_22431_, _22429_);
  nor (_22432_, _22431_, _21414_);
  nor (_25104_, _22432_, _22430_);
  nor (_22434_, _22395_, _21599_);
  nor (_22435_, _22434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  not (_22437_, _22434_);
  nor (_22438_, _22437_, _21504_);
  nor (_01232_, _22438_, _22435_);
  nor (_22439_, _22434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  nor (_22440_, _22437_, _21586_);
  nor (_25101_, _22440_, _22439_);
  nor (_22441_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  nor (_22442_, _22418_, _21526_);
  nor (_01270_, _22442_, _22441_);
  nor (_22443_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  nor (_22444_, _22418_, _21504_);
  nor (_01313_, _22444_, _22443_);
  nor (_22446_, _22395_, _21658_);
  nor (_22447_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  not (_22448_, _22446_);
  nor (_22449_, _22448_, _21586_);
  nor (_01368_, _22449_, _22447_);
  nor (_22450_, _22020_, _21652_);
  nor (_22451_, _22450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  not (_22452_, _22450_);
  nor (_22453_, _22452_, _21414_);
  nor (_01399_, _22453_, _22451_);
  nor (_22454_, _22020_, _21689_);
  nor (_22455_, _22454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  not (_22456_, _22454_);
  nor (_22457_, _22456_, _21504_);
  nor (_01421_, _22457_, _22455_);
  nor (_22458_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  nor (_22459_, _22418_, _21626_);
  nor (_01443_, _22459_, _22458_);
  nor (_22461_, _22049_, _21607_);
  nor (_22462_, _22461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  not (_22463_, _22461_);
  nor (_22464_, _22463_, _21474_);
  nor (_01478_, _22464_, _22462_);
  nor (_22465_, _22020_, _21482_);
  nor (_22466_, _22465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  not (_22467_, _22465_);
  nor (_22468_, _22467_, _21474_);
  nor (_01511_, _22468_, _22466_);
  nor (_22470_, _22020_, _21530_);
  nor (_22471_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  not (_22473_, _22470_);
  nor (_22474_, _22473_, _21554_);
  nor (_01544_, _22474_, _22471_);
  nor (_22475_, _22461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  nor (_22476_, _22463_, _21554_);
  nor (_01600_, _22476_, _22475_);
  nor (_22477_, _22461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  nor (_22478_, _22463_, _21451_);
  nor (_25054_, _22478_, _22477_);
  nor (_22479_, _22020_, _21864_);
  nor (_22481_, _22479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  not (_22482_, _22479_);
  nor (_22483_, _22482_, _21526_);
  nor (_01684_, _22483_, _22481_);
  nor (_22484_, _22020_, _21374_);
  nor (_22485_, _22484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  not (_22486_, _22484_);
  nor (_22487_, _22486_, _21451_);
  nor (_01717_, _22487_, _22485_);
  nor (_22488_, _22021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  nor (_22489_, _22023_, _21474_);
  nor (_01763_, _22489_, _22488_);
  nor (_22490_, _22049_, _21652_);
  nor (_22491_, _22490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  not (_22492_, _22490_);
  nor (_22493_, _22492_, _21626_);
  nor (_01827_, _22493_, _22491_);
  nor (_22494_, _22461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  nor (_22495_, _22463_, _21504_);
  nor (_01849_, _22495_, _22494_);
  nor (_22496_, _22049_, _21689_);
  nor (_22497_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  not (_22498_, _22496_);
  nor (_22499_, _22498_, _21504_);
  nor (_01870_, _22499_, _22497_);
  nor (_22500_, _22049_, _21631_);
  nor (_22501_, _22500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  not (_22502_, _22500_);
  nor (_22503_, _22502_, _21626_);
  nor (_01935_, _22503_, _22501_);
  nor (_22504_, _22186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  nor (_22505_, _22188_, _21586_);
  nor (_01968_, _22505_, _22504_);
  nor (_22506_, _22049_, _21482_);
  nor (_22507_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  not (_22508_, _22506_);
  nor (_22509_, _22508_, _21586_);
  nor (_25056_, _22509_, _22507_);
  nor (_22510_, _22186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  nor (_22511_, _22188_, _21474_);
  nor (_02089_, _22511_, _22510_);
  nor (_22512_, _22020_, _21566_);
  nor (_22513_, _22512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  not (_22514_, _22512_);
  nor (_22515_, _22514_, _21474_);
  nor (_02123_, _22515_, _22513_);
  nor (_22516_, _22004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  nor (_22517_, _22006_, _21451_);
  nor (_25412_, _22517_, _22516_);
  nor (_22519_, _22004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  nor (_22520_, _22006_, _21626_);
  nor (_02200_, _22520_, _22519_);
  nor (_22521_, _22020_, _21821_);
  nor (_22523_, _22521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  not (_22524_, _22521_);
  nor (_22525_, _22524_, _21626_);
  nor (_02233_, _22525_, _22523_);
  nor (_22526_, _22020_, _21599_);
  nor (_22527_, _22526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  not (_22528_, _22526_);
  nor (_22529_, _22528_, _21626_);
  nor (_02266_, _22529_, _22527_);
  nor (_22531_, _22395_, _21689_);
  nor (_22532_, _22531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  not (_22533_, _22531_);
  nor (_22534_, _22533_, _21586_);
  nor (_02355_, _22534_, _22532_);
  nor (_22535_, _22395_, _21425_);
  nor (_22536_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  not (_22537_, _22535_);
  nor (_22538_, _22537_, _21414_);
  nor (_02378_, _22538_, _22536_);
  nor (_22539_, _22004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  nor (_22540_, _22006_, _21504_);
  nor (_02396_, _22540_, _22539_);
  nor (_22541_, _22412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  nor (_22542_, _22414_, _21586_);
  nor (_02417_, _22542_, _22541_);
  nor (_22543_, _22395_, _21821_);
  nor (_22544_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  not (_22545_, _22543_);
  nor (_22546_, _22545_, _21586_);
  nor (_25099_, _22546_, _22544_);
  nor (_22547_, _22395_, _21374_);
  nor (_22548_, _22547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  not (_22549_, _22547_);
  nor (_22550_, _22549_, _21504_);
  nor (_25095_, _22550_, _22548_);
  nor (_22551_, _22020_, _21631_);
  nor (_22553_, _22551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  not (_22555_, _22551_);
  nor (_22556_, _22555_, _21451_);
  nor (_25083_, _22556_, _22553_);
  nor (_22557_, _22020_, _21425_);
  nor (_22558_, _22557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  not (_22559_, _22557_);
  nor (_22560_, _22559_, _21586_);
  nor (_02571_, _22560_, _22558_);
  nor (_22561_, _22020_, _21607_);
  nor (_22562_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  not (_22563_, _22561_);
  nor (_22564_, _22563_, _21586_);
  nor (_02592_, _22564_, _22562_);
  nor (_22565_, _22521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  nor (_22566_, _22524_, _21554_);
  nor (_02608_, _22566_, _22565_);
  nor (_22567_, _22049_, _21425_);
  nor (_22568_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  not (_22569_, _22567_);
  nor (_22570_, _22569_, _21451_);
  nor (_02695_, _22570_, _22568_);
  nor (_22571_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  nor (_22572_, _22508_, _21414_);
  nor (_02721_, _22572_, _22571_);
  nor (_22573_, _22512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  nor (_22574_, _22514_, _21451_);
  nor (_02742_, _22574_, _22573_);
  nor (_22576_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  nor (_22577_, _22165_, _21626_);
  nor (_02764_, _22577_, _22576_);
  nor (_22578_, _22526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  nor (_22579_, _22528_, _21554_);
  nor (_02791_, _22579_, _22578_);
  nor (_22581_, _21659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  nor (_22582_, _21661_, _21586_);
  nor (_25120_, _22582_, _22581_);
  nor (_22583_, _22408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  nor (_22584_, _22410_, _21626_);
  nor (_02842_, _22584_, _22583_);
  nor (_22585_, _22425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  nor (_22586_, _22427_, _21526_);
  nor (_25107_, _22586_, _22585_);
  nor (_22587_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  nor (_22588_, _22448_, _21474_);
  nor (_02894_, _22588_, _22587_);
  nor (_22590_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  nor (_22591_, _22473_, _21526_);
  nor (_02916_, _22591_, _22590_);
  nor (_22592_, _22003_, _21607_);
  nor (_22593_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  not (_22594_, _22592_);
  nor (_22595_, _22594_, _21451_);
  nor (_02949_, _22595_, _22593_);
  nor (_22596_, _22484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  nor (_22598_, _22486_, _21526_);
  nor (_02970_, _22598_, _22596_);
  nor (_22599_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  nor (_22600_, _22594_, _21626_);
  nor (_03016_, _22600_, _22599_);
  nor (_22601_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  nor (_22602_, _22545_, _21474_);
  nor (_03091_, _22602_, _22601_);
  nor (_22603_, _22551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  nor (_22604_, _22555_, _21504_);
  nor (_03113_, _22604_, _22603_);
  nor (_22605_, _22521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  nor (_22606_, _22524_, _21526_);
  nor (_03140_, _22606_, _22605_);
  nor (_22607_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  nor (_22608_, _22594_, _21504_);
  nor (_03163_, _22608_, _22607_);
  nor (_22609_, _22512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  nor (_22611_, _22514_, _21504_);
  nor (_03187_, _22611_, _22609_);
  nor (_22612_, _21659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  nor (_22613_, _21661_, _21474_);
  nor (_03210_, _22613_, _22612_);
  nor (_22614_, _21652_, _21388_);
  nor (_22615_, _22614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  not (_22616_, _22614_);
  nor (_22617_, _22616_, _21504_);
  nor (_25149_, _22617_, _22615_);
  nor (_22619_, _22614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  nor (_22620_, _22616_, _21554_);
  nor (_03422_, _22620_, _22619_);
  nor (_22621_, _22614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  nor (_22622_, _22616_, _21586_);
  nor (_03448_, _22622_, _22621_);
  nor (_22623_, _21689_, _21388_);
  nor (_22624_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  not (_22625_, _22623_);
  nor (_22626_, _22625_, _21626_);
  nor (_03487_, _22626_, _22624_);
  nor (_22627_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  nor (_22628_, _22625_, _21414_);
  nor (_03520_, _22628_, _22627_);
  nor (_22629_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  nor (_22630_, _22625_, _21474_);
  nor (_03578_, _22630_, _22629_);
  nor (_22631_, _21631_, _21388_);
  nor (_22632_, _22631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  not (_22633_, _22631_);
  nor (_22634_, _22633_, _21626_);
  nor (_03612_, _22634_, _22632_);
  nor (_22635_, _22631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  nor (_22636_, _22633_, _21554_);
  nor (_03645_, _22636_, _22635_);
  nor (_22637_, _22631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  nor (_22638_, _22633_, _21586_);
  nor (_03671_, _22638_, _22637_);
  nor (_22639_, _21425_, _21388_);
  nor (_22640_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  not (_22641_, _22639_);
  nor (_22642_, _22641_, _21414_);
  nor (_03725_, _22642_, _22640_);
  nor (_22644_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  nor (_22645_, _22641_, _21586_);
  nor (_25143_, _22645_, _22644_);
  nor (_22646_, _21482_, _21388_);
  nor (_22647_, _22646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  not (_22648_, _22646_);
  nor (_22649_, _22648_, _21451_);
  nor (_03815_, _22649_, _22647_);
  nor (_22650_, _22646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  nor (_22651_, _22648_, _21554_);
  nor (_25141_, _22651_, _22650_);
  nor (_22652_, _22646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  nor (_22653_, _22648_, _21586_);
  nor (_03877_, _22653_, _22652_);
  nor (_22654_, _21530_, _21388_);
  nor (_22655_, _22654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  not (_22656_, _22654_);
  nor (_22657_, _22656_, _21626_);
  nor (_03920_, _22657_, _22655_);
  nor (_22658_, _22654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  nor (_22659_, _22656_, _21451_);
  nor (_03949_, _22659_, _22658_);
  nor (_22660_, _22654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  nor (_22661_, _22656_, _21586_);
  nor (_03987_, _22661_, _22660_);
  nor (_22663_, _21558_, _21388_);
  nor (_22664_, _22663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  not (_22665_, _22663_);
  nor (_22666_, _22665_, _21474_);
  nor (_04024_, _22666_, _22664_);
  nor (_22667_, _21566_, _21388_);
  nor (_22668_, _22667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  not (_22669_, _22667_);
  nor (_22670_, _22669_, _21451_);
  nor (_04083_, _22670_, _22668_);
  nor (_22671_, _22667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  nor (_22672_, _22669_, _21474_);
  nor (_04130_, _22672_, _22671_);
  nor (_22673_, _21589_, _21388_);
  nor (_22674_, _22673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  not (_22675_, _22673_);
  nor (_22676_, _22675_, _21504_);
  nor (_04164_, _22676_, _22674_);
  nor (_22677_, _22673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  nor (_22678_, _22675_, _21526_);
  nor (_25134_, _22678_, _22677_);
  nor (_22679_, _21599_, _21388_);
  nor (_22680_, _22679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  not (_22681_, _22679_);
  nor (_22682_, _22681_, _21414_);
  nor (_04244_, _22682_, _22680_);
  nor (_22683_, _21607_, _21388_);
  nor (_22684_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  not (_22685_, _22683_);
  nor (_22686_, _22685_, _21504_);
  nor (_04298_, _22686_, _22684_);
  nor (_22688_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  nor (_22689_, _22685_, _21474_);
  nor (_04341_, _22689_, _22688_);
  nor (_22690_, _22663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  nor (_22692_, _22665_, _21414_);
  nor (_04376_, _22692_, _22690_);
  nor (_22693_, _21695_, _21638_);
  nor (_22695_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  not (_22696_, _22693_);
  nor (_22697_, _22696_, _21554_);
  nor (_04397_, _22697_, _22695_);
  nor (_22698_, _22614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  nor (_22699_, _22616_, _21414_);
  nor (_04422_, _22699_, _22698_);
  nor (_22700_, _22631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  nor (_22701_, _22633_, _21414_);
  nor (_25146_, _22701_, _22700_);
  nor (_22702_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  nor (_22703_, _22641_, _21504_);
  nor (_04548_, _22703_, _22702_);
  nor (_22705_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  nor (_22706_, _22641_, _21554_);
  nor (_04569_, _22706_, _22705_);
  nor (_22707_, _22646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  nor (_22708_, _22648_, _21626_);
  nor (_25142_, _22708_, _22707_);
  nor (_22709_, _22004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  nor (_22710_, _22006_, _21474_);
  nor (_04635_, _22710_, _22709_);
  nor (_22712_, _22654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  nor (_22713_, _22656_, _21554_);
  nor (_04689_, _22713_, _22712_);
  nor (_22714_, _22667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  nor (_22716_, _22669_, _21626_);
  nor (_04725_, _22716_, _22714_);
  nor (_22717_, _22667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  nor (_22718_, _22669_, _21526_);
  nor (_04747_, _22718_, _22717_);
  nor (_22719_, _22021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  nor (_22721_, _22023_, _21504_);
  nor (_04771_, _22721_, _22719_);
  nor (_22723_, _22004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  nor (_22724_, _22006_, _21586_);
  nor (_04792_, _22724_, _22723_);
  nor (_22725_, _22673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  nor (_22726_, _22675_, _21586_);
  nor (_04816_, _22726_, _22725_);
  nor (_22728_, _22679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  nor (_22730_, _22681_, _21474_);
  nor (_04837_, _22730_, _22728_);
  nor (_22731_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  nor (_22732_, _22685_, _21526_);
  nor (_04871_, _22732_, _22731_);
  nor (_22733_, _22663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  nor (_22734_, _22665_, _21504_);
  nor (_04890_, _22734_, _22733_);
  nor (_22735_, _22663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  nor (_22736_, _22665_, _21554_);
  nor (_25137_, _22736_, _22735_);
  nor (_22738_, _22673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  nor (_22739_, _22675_, _21414_);
  nor (_25135_, _22739_, _22738_);
  nor (_22740_, _22679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  nor (_22741_, _22681_, _21451_);
  nor (_05039_, _22741_, _22740_);
  nor (_22743_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  nor (_22744_, _22685_, _21626_);
  nor (_25140_, _22744_, _22743_);
  nor (_22745_, _22663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  nor (_22747_, _22665_, _21626_);
  nor (_05200_, _22747_, _22745_);
  nor (_22749_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  nor (_22750_, _22594_, _21586_);
  nor (_05218_, _22750_, _22749_);
  nor (_22751_, _22663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  nor (_22752_, _22665_, _21526_);
  nor (_05249_, _22752_, _22751_);
  nor (_22754_, _22663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  nor (_22756_, _22665_, _21451_);
  nor (_05271_, _22756_, _22754_);
  nor (_22757_, _22526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  nor (_22758_, _22528_, _21474_);
  nor (_05292_, _22758_, _22757_);
  nor (_22759_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  nor (_22760_, _22165_, _21554_);
  nor (_05327_, _22760_, _22759_);
  nor (_22761_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  nor (_22762_, _22685_, _21586_);
  nor (_25138_, _22762_, _22761_);
  nor (_22763_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  nor (_22764_, _22165_, _21586_);
  nor (_05359_, _22764_, _22763_);
  nor (_22765_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  nor (_22766_, _22685_, _21554_);
  nor (_25139_, _22766_, _22765_);
  nor (_22767_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  nor (_22768_, _22165_, _21504_);
  nor (_05392_, _22768_, _22767_);
  nor (_22769_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  nor (_22770_, _22685_, _21414_);
  nor (_05410_, _22770_, _22769_);
  nor (_22771_, _22512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  nor (_22772_, _22514_, _21586_);
  nor (_25072_, _22772_, _22771_);
  nor (_22773_, _22512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  nor (_22775_, _22514_, _21414_);
  nor (_05451_, _22775_, _22773_);
  nor (_22776_, _22683_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  nor (_22778_, _22685_, _21451_);
  nor (_05466_, _22778_, _22776_);
  nor (_22779_, _22512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  nor (_22780_, _22514_, _21526_);
  nor (_05480_, _22780_, _22779_);
  nor (_22781_, _21821_, _21388_);
  nor (_22782_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  not (_22783_, _22781_);
  nor (_22784_, _22783_, _21626_);
  nor (_05504_, _22784_, _22782_);
  nor (_22785_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  nor (_22786_, _22594_, _21526_);
  nor (_05524_, _22786_, _22785_);
  nor (_22787_, _22186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  nor (_22789_, _22188_, _21504_);
  nor (_05542_, _22789_, _22787_);
  nor (_22790_, _22679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  nor (_22791_, _22681_, _21586_);
  nor (_25129_, _22791_, _22790_);
  nor (_22792_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  nor (_22793_, _22508_, _21526_);
  nor (_05578_, _22793_, _22792_);
  nor (_22794_, _22679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  nor (_22795_, _22681_, _21554_);
  nor (_25130_, _22795_, _22794_);
  nor (_22796_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  nor (_22797_, _22569_, _21586_);
  nor (_05618_, _22797_, _22796_);
  nor (_22798_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  nor (_22799_, _22594_, _21554_);
  nor (_05640_, _22799_, _22798_);
  nor (_22800_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  nor (_22801_, _22508_, _21504_);
  nor (_05662_, _22801_, _22800_);
  nor (_22802_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  nor (_22803_, _22569_, _21414_);
  nor (_05683_, _22803_, _22802_);
  nor (_22804_, _22679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  nor (_22805_, _22681_, _21526_);
  nor (_05705_, _22805_, _22804_);
  nor (_22806_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  nor (_22807_, _22569_, _21554_);
  nor (_05720_, _22807_, _22806_);
  nor (_22808_, _22679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  nor (_22810_, _22681_, _21504_);
  nor (_05739_, _22810_, _22808_);
  nor (_22811_, _22500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  nor (_22812_, _22502_, _21586_);
  nor (_05792_, _22812_, _22811_);
  nor (_22813_, _22679_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  nor (_22815_, _22681_, _21626_);
  nor (_25131_, _22815_, _22813_);
  nor (_22816_, _22500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  nor (_22817_, _22502_, _21451_);
  nor (_25060_, _22817_, _22816_);
  nor (_22818_, _22673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  nor (_22819_, _22675_, _21474_);
  nor (_25133_, _22819_, _22818_);
  nor (_22820_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  nor (_22821_, _22498_, _21554_);
  nor (_05875_, _22821_, _22820_);
  nor (_22822_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  nor (_22823_, _22498_, _21474_);
  nor (_05896_, _22823_, _22822_);
  nor (_22824_, _22673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  nor (_22825_, _22675_, _21554_);
  nor (_05916_, _22825_, _22824_);
  nor (_22826_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  nor (_22827_, _22498_, _21414_);
  nor (_05936_, _22827_, _22826_);
  nor (_22828_, _22490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  nor (_22829_, _22492_, _21554_);
  nor (_05959_, _22829_, _22828_);
  nor (_22830_, _22673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  nor (_22831_, _22675_, _21451_);
  nor (_05980_, _22831_, _22830_);
  nor (_22832_, _22673_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  nor (_22833_, _22675_, _21626_);
  nor (_05999_, _22833_, _22832_);
  nor (_22834_, _22003_, _21558_);
  nor (_22835_, _22834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  not (_22836_, _22834_);
  nor (_22837_, _22836_, _21414_);
  nor (_06035_, _22837_, _22835_);
  nor (_22838_, _22020_, _21638_);
  nor (_22839_, _22838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  not (_22840_, _22838_);
  nor (_22841_, _22840_, _21554_);
  nor (_25066_, _22841_, _22839_);
  nor (_22842_, _22667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  nor (_22843_, _22669_, _21586_);
  nor (_06105_, _22843_, _22842_);
  nor (_22844_, _22834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  nor (_22845_, _22836_, _21526_);
  nor (_25408_, _22845_, _22844_);
  nor (_22846_, _22667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  nor (_22847_, _22669_, _21554_);
  nor (_06157_, _22847_, _22846_);
  nor (_22848_, _22838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  nor (_22849_, _22840_, _21504_);
  nor (_06182_, _22849_, _22848_);
  nor (_22851_, _22834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  nor (_22852_, _22836_, _21554_);
  nor (_06204_, _22852_, _22851_);
  nor (_22853_, _22021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  nor (_22854_, _22023_, _21626_);
  nor (_06232_, _22854_, _22853_);
  nor (_22855_, _22667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  nor (_22856_, _22669_, _21414_);
  nor (_06259_, _22856_, _22855_);
  nor (_22857_, _22667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  nor (_22858_, _22669_, _21504_);
  nor (_06301_, _22858_, _22857_);
  nor (_22860_, _22484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  nor (_22861_, _22486_, _21554_);
  nor (_06324_, _22861_, _22860_);
  nor (_22862_, _22521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  nor (_22863_, _22524_, _21474_);
  nor (_06383_, _22863_, _22862_);
  nor (_22864_, _22663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  nor (_22865_, _22665_, _21586_);
  nor (_25136_, _22865_, _22864_);
  nor (_22866_, _22479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  nor (_22867_, _22482_, _21504_);
  nor (_25068_, _22867_, _22866_);
  nor (_22869_, _22020_, _21558_);
  nor (_22870_, _22869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  not (_22872_, _22869_);
  nor (_22873_, _22872_, _21554_);
  nor (_06511_, _22873_, _22870_);
  nor (_22874_, _22869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  nor (_22876_, _22872_, _21586_);
  nor (_25074_, _22876_, _22874_);
  nor (_22877_, _22654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  nor (_22878_, _22656_, _21474_);
  nor (_06565_, _22878_, _22877_);
  nor (_22879_, _22869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  nor (_22881_, _22872_, _21451_);
  nor (_06632_, _22881_, _22879_);
  nor (_22882_, _22654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  nor (_22883_, _22656_, _21526_);
  nor (_06649_, _22883_, _22882_);
  nor (_22884_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  nor (_22885_, _22563_, _21451_);
  nor (_06672_, _22885_, _22884_);
  nor (_22886_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  nor (_22887_, _22563_, _21554_);
  nor (_06726_, _22887_, _22886_);
  nor (_22889_, _22834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  nor (_22890_, _22836_, _21504_);
  nor (_06776_, _22890_, _22889_);
  nor (_22891_, _22654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  nor (_22892_, _22656_, _21414_);
  nor (_06801_, _22892_, _22891_);
  nor (_22893_, _22834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  nor (_22894_, _22836_, _21451_);
  nor (_25409_, _22894_, _22893_);
  nor (_22895_, _22654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  nor (_22896_, _22656_, _21504_);
  nor (_06899_, _22896_, _22895_);
  nor (_22897_, _22557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  nor (_22898_, _22559_, _21504_);
  nor (_06998_, _22898_, _22897_);
  nor (_22899_, _22646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  nor (_22900_, _22648_, _21474_);
  nor (_07017_, _22900_, _22899_);
  nor (_22901_, _22557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  nor (_22902_, _22559_, _21414_);
  nor (_07036_, _22902_, _22901_);
  nor (_22903_, _22646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  nor (_22904_, _22648_, _21526_);
  nor (_07055_, _22904_, _22903_);
  nor (_22905_, _22551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  nor (_22907_, _22555_, _21414_);
  nor (_07070_, _22907_, _22905_);
  nor (_22908_, _22646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  nor (_22909_, _22648_, _21414_);
  nor (_07150_, _22909_, _22908_);
  nor (_22910_, _22003_, _21566_);
  nor (_22911_, _22910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  not (_22912_, _22910_);
  nor (_22914_, _22912_, _21504_);
  nor (_07181_, _22914_, _22911_);
  nor (_22915_, _22646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  nor (_22917_, _22648_, _21504_);
  nor (_07199_, _22917_, _22915_);
  nor (_22918_, _22910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  nor (_22919_, _22912_, _21451_);
  nor (_07223_, _22919_, _22918_);
  nor (_22920_, _22910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  nor (_22921_, _22912_, _21414_);
  nor (_07237_, _22921_, _22920_);
  nor (_22922_, _22395_, _21638_);
  nor (_22923_, _22922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  not (_22924_, _22922_);
  nor (_22925_, _22924_, _21474_);
  nor (_25089_, _22925_, _22923_);
  nor (_22927_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  nor (_22928_, _22641_, _21474_);
  nor (_25144_, _22928_, _22927_);
  nor (_22929_, _22910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  nor (_22930_, _22912_, _21526_);
  nor (_07371_, _22930_, _22929_);
  nor (_22931_, _22922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  nor (_22932_, _22924_, _21451_);
  nor (_07391_, _22932_, _22931_);
  nor (_22933_, _22547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  nor (_22934_, _22549_, _21586_);
  nor (_07423_, _22934_, _22933_);
  nor (_22936_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  nor (_22937_, _22641_, _21526_);
  nor (_07444_, _22937_, _22936_);
  nor (_22938_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  nor (_22939_, _22448_, _21451_);
  nor (_07466_, _22939_, _22938_);
  nor (_22940_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  nor (_22941_, _22641_, _21451_);
  nor (_07487_, _22941_, _22940_);
  nor (_22942_, _22547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  nor (_22943_, _22549_, _21451_);
  nor (_07506_, _22943_, _22942_);
  nor (_22945_, _22547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  nor (_22946_, _22549_, _21526_);
  nor (_07557_, _22946_, _22945_);
  nor (_22947_, _22639_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  nor (_22948_, _22641_, _21626_);
  nor (_25145_, _22948_, _22947_);
  nor (_22949_, _22395_, _21864_);
  nor (_22950_, _22949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  not (_22951_, _22949_);
  nor (_22952_, _22951_, _21554_);
  nor (_25096_, _22952_, _22950_);
  nor (_22953_, _22227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  nor (_22954_, _22229_, _21526_);
  nor (_07695_, _22954_, _22953_);
  nor (_22955_, _22631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  nor (_22956_, _22633_, _21474_);
  nor (_07717_, _22956_, _22955_);
  nor (_22957_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  nor (_22958_, _22545_, _21451_);
  nor (_07739_, _22958_, _22957_);
  nor (_22960_, _22631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  nor (_22961_, _22633_, _21526_);
  nor (_07760_, _22961_, _22960_);
  nor (_22962_, _22834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  nor (_22963_, _22836_, _21586_);
  nor (_07780_, _22963_, _22962_);
  nor (_22965_, _22434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  nor (_22966_, _22437_, _21526_);
  nor (_07822_, _22966_, _22965_);
  nor (_22967_, _22631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  nor (_22968_, _22633_, _21451_);
  nor (_07848_, _22968_, _22967_);
  nor (_22969_, _21822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  nor (_22970_, _21824_, _21414_);
  nor (_25204_, _22970_, _22969_);
  nor (_22971_, _22910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  nor (_22972_, _22912_, _21626_);
  nor (_07913_, _22972_, _22971_);
  nor (_22973_, _22631_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  nor (_22974_, _22633_, _21504_);
  nor (_25147_, _22974_, _22973_);
  nor (_22975_, _22429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  nor (_22976_, _22431_, _21626_);
  nor (_07956_, _22976_, _22975_);
  nor (_22977_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  nor (_22978_, _22625_, _21586_);
  nor (_07999_, _22978_, _22977_);
  nor (_22980_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  nor (_22981_, _22625_, _21554_);
  nor (_08057_, _22981_, _22980_);
  nor (_22982_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  nor (_22983_, _22625_, _21526_);
  nor (_08144_, _22983_, _22982_);
  nor (_22984_, _22412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  nor (_22986_, _22414_, _21526_);
  nor (_08168_, _22986_, _22984_);
  nor (_22987_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  nor (_22988_, _22625_, _21451_);
  nor (_08188_, _22988_, _22987_);
  nor (_22989_, _22408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  nor (_22990_, _22410_, _21554_);
  nor (_08212_, _22990_, _22989_);
  nor (_22991_, _22395_, _21482_);
  nor (_22992_, _22991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  not (_22993_, _22991_);
  nor (_22994_, _22993_, _21451_);
  nor (_08247_, _22994_, _22992_);
  nor (_22995_, _22623_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  nor (_22996_, _22625_, _21504_);
  nor (_25148_, _22996_, _22995_);
  nor (_22997_, _22991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  nor (_22998_, _22993_, _21554_);
  nor (_08292_, _22998_, _22997_);
  nor (_22999_, _22003_, _21589_);
  nor (_23000_, _22999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  not (_23001_, _22999_);
  nor (_23002_, _23001_, _21626_);
  nor (_25407_, _23002_, _23000_);
  nor (_23003_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  nor (_23004_, _22537_, _21526_);
  nor (_08344_, _23004_, _23003_);
  nor (_23005_, _22999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  nor (_23006_, _23001_, _21504_);
  nor (_08383_, _23006_, _23005_);
  nor (_23007_, _22614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  nor (_23008_, _22616_, _21474_);
  nor (_08407_, _23008_, _23007_);
  nor (_23009_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  nor (_23010_, _22537_, _21504_);
  nor (_08427_, _23010_, _23009_);
  nor (_23011_, _22614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  nor (_23012_, _22616_, _21526_);
  nor (_08455_, _23012_, _23011_);
  nor (_23013_, _22403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  nor (_23014_, _22406_, _21451_);
  nor (_08490_, _23014_, _23013_);
  nor (_23015_, _22531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  nor (_23016_, _22533_, _21504_);
  nor (_08527_, _23016_, _23015_);
  nor (_23017_, _22614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  nor (_23018_, _22616_, _21451_);
  nor (_08549_, _23018_, _23017_);
  nor (_23020_, _22614_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  nor (_23021_, _22616_, _21626_);
  nor (_25150_, _23021_, _23020_);
  nor (_23022_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  nor (_23023_, _22696_, _21586_);
  nor (_08656_, _23023_, _23022_);
  nor (_23025_, _21638_, _21388_);
  nor (_23026_, _23025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  not (_23027_, _23025_);
  nor (_23028_, _23027_, _21474_);
  nor (_25118_, _23028_, _23026_);
  nor (_23029_, _23025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  nor (_23030_, _23027_, _21626_);
  nor (_08758_, _23030_, _23029_);
  nor (_23031_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  nor (_23032_, _22696_, _21474_);
  nor (_08790_, _23032_, _23031_);
  nor (_23034_, _23025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  nor (_23035_, _23027_, _21414_);
  nor (_08820_, _23035_, _23034_);
  nor (_23036_, _22910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  nor (_23037_, _22912_, _21586_);
  nor (_08905_, _23037_, _23036_);
  not (_23038_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_23039_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nand (_23040_, _23039_, _23038_);
  not (_23041_, _23040_);
  nor (_23042_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  not (_23043_, _23042_);
  nor (_23044_, _23043_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_23045_, _23044_, _23041_);
  not (_23046_, _23045_);
  not (_23047_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_23048_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_23049_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_23050_, _23049_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_23051_, _23050_, _23048_);
  not (_23052_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  not (_23054_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not (_23055_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  not (_23056_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_23057_, _23056_, _23055_);
  nand (_23058_, _23057_, _23054_);
  nor (_23059_, _23058_, _23052_);
  nor (_23060_, _23059_, _23051_);
  nand (_23061_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _23055_);
  nor (_23062_, _23061_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_23063_, _23062_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nand (_23064_, _23063_, _23060_);
  not (_23065_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_23066_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _23055_);
  nand (_23067_, _23066_, _23054_);
  nor (_23068_, _23067_, _23065_);
  nor (_23069_, _23068_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_23070_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nand (_23072_, _23056_, _23055_);
  nand (_23073_, _23072_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_23074_, _23073_, _23070_);
  not (_23075_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nand (_23076_, _23049_, _23054_);
  nor (_23077_, _23076_, _23075_);
  nor (_23078_, _23077_, _23074_);
  nand (_23079_, _23078_, _23069_);
  nor (_23080_, _23079_, _23064_);
  nand (_23081_, _23080_, _23047_);
  nor (_23082_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _23047_);
  not (_23083_, _23082_);
  nand (_23084_, _23083_, _23081_);
  nand (_23085_, _23084_, _23046_);
  nor (_23086_, _23044_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_23087_, _23086_, _23040_);
  nand (_23088_, _23087_, _23085_);
  not (_23090_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nor (_23091_, _23076_, _23090_);
  not (_23092_, _23091_);
  nand (_23094_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_23095_, _23094_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_23096_, _23095_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nand (_23097_, _23096_, _23092_);
  not (_23098_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_23099_, _23073_, _23098_);
  not (_23100_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_23101_, _23067_, _23100_);
  nor (_23102_, _23101_, _23099_);
  not (_23103_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_23104_, _23050_, _23103_);
  not (_23105_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_23106_, _23056_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_23107_, _23106_, _23054_);
  nor (_23108_, _23107_, _23105_);
  nor (_23109_, _23108_, _23104_);
  nand (_23110_, _23109_, _23102_);
  nor (_23111_, _23110_, _23097_);
  nor (_23112_, _23111_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_23113_, _23112_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_23114_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _23047_);
  nor (_23115_, _23114_, _23113_);
  nor (_23116_, _23115_, _23045_);
  nor (_23117_, _23044_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_23118_, _23117_, _23040_);
  not (_23119_, _23118_);
  nor (_23120_, _23119_, _23116_);
  nor (_23121_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_23122_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_23123_, _23076_, _23122_);
  not (_23124_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_23125_, _23067_, _23124_);
  nor (_23126_, _23125_, _23123_);
  nor (_23127_, _23049_, _23054_);
  nand (_23128_, _23127_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_23129_, _23095_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nand (_23130_, _23129_, _23128_);
  nor (_23131_, _23072_, _23054_);
  nand (_23132_, _23131_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand (_23133_, _23062_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nand (_23134_, _23133_, _23132_);
  nor (_23135_, _23134_, _23130_);
  nand (_23137_, _23135_, _23126_);
  nand (_23138_, _23137_, _23121_);
  not (_23139_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  nor (_23140_, _23139_, _23047_);
  not (_23141_, _23140_);
  nand (_23143_, _23141_, _23138_);
  nor (_23144_, _23143_, _23045_);
  nor (_23145_, _23044_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_23146_, _23145_, _23040_);
  not (_23147_, _23146_);
  nor (_23148_, _23147_, _23144_);
  nand (_23149_, _23148_, _23120_);
  nor (_23150_, _23149_, _23088_);
  not (_23151_, \oc8051_top_1.oc8051_memory_interface1.cdata [0]);
  nor (_23152_, _23151_, _23047_);
  not (_23153_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_23154_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_23155_, _23076_, _23154_);
  not (_23156_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_23157_, _23067_, _23156_);
  nor (_23159_, _23157_, _23155_);
  nand (_23160_, _23127_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_23161_, _23131_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nand (_23162_, _23161_, _23160_);
  nand (_23163_, _23095_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nand (_23164_, _23062_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nand (_23165_, _23164_, _23163_);
  nor (_23166_, _23165_, _23162_);
  nand (_23167_, _23166_, _23159_);
  nand (_23168_, _23167_, _23153_);
  nor (_23169_, _23168_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_23170_, _23169_, _23152_);
  nand (_23172_, _23170_, _23046_);
  nor (_23173_, _23044_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_23174_, _23173_, _23040_);
  nand (_23175_, _23174_, _23172_);
  not (_23176_, _23121_);
  nor (_23177_, _23072_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_23178_, _23177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_23179_, _23056_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_23180_, _23179_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_23181_, _23180_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nand (_23182_, _23181_, _23178_);
  not (_23183_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_23184_, _23073_, _23183_);
  not (_23185_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_23186_, _23058_, _23185_);
  nor (_23187_, _23186_, _23184_);
  not (_23188_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_23189_, _23050_, _23188_);
  not (_23190_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_23191_, _23107_, _23190_);
  nor (_23192_, _23191_, _23189_);
  nand (_23193_, _23192_, _23187_);
  nor (_23194_, _23193_, _23182_);
  nor (_23195_, _23194_, _23176_);
  not (_23197_, \oc8051_top_1.oc8051_memory_interface1.cdata [3]);
  nor (_23198_, _23197_, _23047_);
  nor (_23199_, _23198_, _23195_);
  nand (_23200_, _23199_, _23046_);
  nor (_23201_, _23044_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_23202_, _23201_, _23040_);
  nand (_23203_, _23202_, _23200_);
  not (_23204_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_23206_, _23076_, _23204_);
  not (_23207_, _23206_);
  nand (_23208_, _23180_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nand (_23209_, _23208_, _23207_);
  not (_23210_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_23211_, _23073_, _23210_);
  not (_23212_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_23213_, _23058_, _23212_);
  nor (_23214_, _23213_, _23211_);
  not (_23215_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_23216_, _23050_, _23215_);
  not (_23217_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_23218_, _23107_, _23217_);
  nor (_23219_, _23218_, _23216_);
  nand (_23220_, _23219_, _23214_);
  nor (_23221_, _23220_, _23209_);
  nor (_23222_, _23221_, _23176_);
  not (_23223_, \oc8051_top_1.oc8051_memory_interface1.cdata [2]);
  nor (_23224_, _23223_, _23047_);
  nor (_23225_, _23224_, _23222_);
  nand (_23226_, _23225_, _23046_);
  nor (_23227_, _23044_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_23228_, _23227_, _23040_);
  nand (_23229_, _23228_, _23226_);
  nand (_23230_, _23131_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand (_23231_, _23095_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nand (_23232_, _23231_, _23230_);
  not (_23233_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_23234_, _23073_, _23233_);
  nor (_23235_, _23234_, _23232_);
  nand (_23236_, _23180_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nand (_23237_, _23177_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nand (_23238_, _23237_, _23236_);
  nand (_23239_, _23062_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nand (_23240_, _23239_, _23153_);
  nor (_23241_, _23240_, _23238_);
  nand (_23242_, _23241_, _23235_);
  nor (_23243_, _23242_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_23244_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _23047_);
  nor (_23245_, _23244_, _23243_);
  nor (_23246_, _23245_, _23045_);
  nor (_23247_, _23044_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_23248_, _23247_, _23040_);
  not (_23249_, _23248_);
  nor (_23250_, _23249_, _23246_);
  nor (_23251_, _23250_, _23229_);
  nand (_23253_, _23251_, _23203_);
  nor (_23255_, _23253_, _23175_);
  nand (_23256_, _23255_, _23150_);
  not (_23257_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_23258_, _23050_, _23257_);
  not (_23259_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_23261_, _23058_, _23259_);
  nor (_23262_, _23261_, _23258_);
  nand (_23263_, _23239_, _23262_);
  not (_23264_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_23265_, _23067_, _23264_);
  nor (_23266_, _23265_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_23268_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_23269_, _23076_, _23268_);
  nor (_23271_, _23269_, _23234_);
  nand (_23272_, _23271_, _23266_);
  nor (_23273_, _23272_, _23263_);
  nand (_23275_, _23273_, _23047_);
  not (_23276_, _23244_);
  nand (_23277_, _23276_, _23275_);
  nand (_23278_, _23277_, _23046_);
  nand (_23279_, _23248_, _23278_);
  nand (_23280_, _23229_, _23203_);
  nor (_23282_, _23280_, _23279_);
  not (_23283_, _23088_);
  not (_23284_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_23285_, _23076_, _23284_);
  not (_23286_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_23287_, _23067_, _23286_);
  nor (_23288_, _23287_, _23285_);
  nand (_23289_, _23127_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_23290_, _23131_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nand (_23292_, _23290_, _23289_);
  nand (_23293_, _23095_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nand (_23294_, _23062_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nand (_23295_, _23294_, _23293_);
  nor (_23296_, _23295_, _23292_);
  nand (_23297_, _23296_, _23288_);
  nand (_23298_, _23297_, _23153_);
  nand (_23299_, _23298_, _23047_);
  nor (_23300_, _23047_, \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  not (_23301_, _23300_);
  nand (_23302_, _23301_, _23299_);
  nand (_23303_, _23302_, _23046_);
  nor (_23304_, _23044_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_23305_, _23304_, _23040_);
  nand (_23306_, _23305_, _23303_);
  nor (_23307_, _23101_, _23091_);
  nand (_23308_, _23127_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_23309_, _23131_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand (_23310_, _23309_, _23308_);
  nand (_23312_, _23062_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nand (_23313_, _23312_, _23096_);
  nor (_23315_, _23313_, _23310_);
  nand (_23316_, _23315_, _23307_);
  nand (_23317_, _23316_, _23153_);
  nand (_23318_, _23317_, _23047_);
  not (_23319_, _23114_);
  nand (_23320_, _23319_, _23318_);
  nand (_23321_, _23320_, _23046_);
  nand (_23323_, _23118_, _23321_);
  nor (_23324_, _23148_, _23323_);
  nand (_23326_, _23324_, _23306_);
  nor (_23327_, _23326_, _23283_);
  nand (_23328_, _23327_, _23282_);
  nand (_23329_, _23328_, _23256_);
  nand (_23330_, _23282_, _23175_);
  nand (_23331_, _23306_, _23323_);
  nor (_23332_, _23331_, _23148_);
  nand (_23333_, _23332_, _23283_);
  nor (_23334_, _23333_, _23330_);
  not (_23335_, _23334_);
  not (_23337_, _23148_);
  nor (_23338_, _23306_, _23120_);
  nand (_23339_, _23338_, _23337_);
  nor (_23341_, _23339_, _23283_);
  nand (_23342_, _23341_, _23255_);
  nand (_23343_, _23342_, _23335_);
  nor (_23345_, _23343_, _23329_);
  not (_23346_, _23152_);
  nand (_23347_, _23167_, _23121_);
  nand (_23348_, _23347_, _23346_);
  nor (_23349_, _23348_, _23045_);
  not (_23350_, _23174_);
  nor (_23351_, _23350_, _23349_);
  nor (_23352_, _23194_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_23353_, _23352_, _23047_);
  not (_23354_, _23198_);
  nand (_23355_, _23354_, _23353_);
  nor (_23356_, _23355_, _23045_);
  not (_23358_, _23202_);
  nor (_23359_, _23358_, _23356_);
  not (_23360_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_23362_, _23067_, _23360_);
  nor (_23364_, _23362_, _23206_);
  nand (_23365_, _23127_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand (_23366_, _23095_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nand (_23367_, _23366_, _23365_);
  nand (_23368_, _23131_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand (_23369_, _23062_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nand (_23370_, _23369_, _23368_);
  nor (_23371_, _23370_, _23367_);
  nand (_23372_, _23371_, _23364_);
  nand (_23373_, _23372_, _23121_);
  not (_23374_, _23224_);
  nand (_23375_, _23374_, _23373_);
  nor (_23376_, _23375_, _23045_);
  not (_23377_, _23228_);
  nor (_23378_, _23377_, _23376_);
  nand (_23379_, _23279_, _23378_);
  nor (_23381_, _23379_, _23359_);
  nand (_23382_, _23381_, _23351_);
  not (_23383_, _23285_);
  nand (_23384_, _23293_, _23383_);
  not (_23385_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_23386_, _23073_, _23385_);
  nor (_23387_, _23287_, _23386_);
  not (_23388_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_23389_, _23050_, _23388_);
  not (_23391_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_23392_, _23107_, _23391_);
  nor (_23393_, _23392_, _23389_);
  nand (_23394_, _23393_, _23387_);
  nor (_23396_, _23394_, _23384_);
  nor (_23397_, _23396_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_23398_, _23397_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_23400_, _23300_, _23398_);
  nor (_23402_, _23400_, _23045_);
  not (_23403_, _23305_);
  nor (_23404_, _23403_, _23402_);
  nor (_23405_, _23404_, _23120_);
  nand (_23407_, _23405_, _23337_);
  nor (_23408_, _23407_, _23088_);
  nand (_23409_, _23324_, _23404_);
  nor (_23410_, _23409_, _23088_);
  nor (_23411_, _23410_, _23408_);
  nor (_23412_, _23411_, _23382_);
  nor (_23413_, _23409_, _23283_);
  nor (_23414_, _23337_, _23088_);
  nand (_23415_, _23338_, _23414_);
  not (_23416_, _23415_);
  nor (_23418_, _23416_, _23413_);
  nor (_23419_, _23418_, _23330_);
  nor (_23420_, _23419_, _23412_);
  nand (_23421_, _23420_, _23345_);
  not (_23422_, _23282_);
  nor (_23423_, _23404_, _23149_);
  nand (_23424_, _23423_, _23088_);
  nor (_23425_, _23424_, _23422_);
  nand (_23426_, _23413_, _23255_);
  nand (_23427_, _23337_, _23120_);
  nor (_23428_, _23427_, _23306_);
  nor (_23429_, _23250_, _23351_);
  not (_23430_, _23429_);
  nor (_23431_, _23430_, _23280_);
  nand (_23432_, _23431_, _23428_);
  nand (_23433_, _23432_, _23426_);
  nor (_23434_, _23433_, _23425_);
  nand (_23435_, _23332_, _23088_);
  nor (_23436_, _23435_, _23382_);
  nand (_23438_, _23250_, _23175_);
  nor (_23440_, _23438_, _23280_);
  nand (_23441_, _23410_, _23440_);
  nor (_23442_, _23339_, _23088_);
  nand (_23443_, _23442_, _23440_);
  nand (_23444_, _23443_, _23441_);
  nor (_23445_, _23444_, _23436_);
  nand (_23447_, _23445_, _23434_);
  nor (_23448_, _23447_, _23421_);
  nor (_23449_, _23326_, _23088_);
  nand (_23450_, _23449_, _23282_);
  nor (_23452_, _23279_, _23229_);
  nand (_23454_, _23452_, _23203_);
  nor (_23455_, _23454_, _23409_);
  nor (_23456_, _23203_, _23283_);
  not (_23457_, _23456_);
  nor (_23458_, _23457_, _23409_);
  nor (_23459_, _23458_, _23455_);
  not (_23460_, _23459_);
  nand (_23461_, _23404_, _23323_);
  nor (_23462_, _23461_, _23148_);
  nand (_23464_, _23462_, _23088_);
  nor (_23465_, _23454_, _23464_);
  nor (_23466_, _23465_, _23460_);
  nand (_23467_, _23466_, _23450_);
  nor (_23468_, _23410_, _23332_);
  nor (_23469_, _23468_, _23203_);
  nor (_23470_, _23250_, _23175_);
  not (_23471_, _23280_);
  nand (_23472_, _23471_, _23470_);
  nor (_23473_, _23472_, _23088_);
  nor (_23474_, _23457_, _23461_);
  nor (_23475_, _23474_, _23473_);
  nand (_23476_, _23359_, _23150_);
  nand (_23477_, _23476_, _23475_);
  nor (_23478_, _23477_, _23469_);
  nand (_23479_, _23250_, _23378_);
  nor (_23480_, _23479_, _23359_);
  nor (_23481_, _23461_, _23337_);
  nand (_23482_, _23481_, _23088_);
  nor (_23484_, _23332_, _23150_);
  nand (_23485_, _23484_, _23482_);
  nand (_23486_, _23485_, _23480_);
  nand (_23487_, _23486_, _23478_);
  nor (_23488_, _23487_, _23467_);
  nand (_23489_, _23488_, _23448_);
  not (_23490_, _23044_);
  nor (_23491_, _23490_, rst);
  nand (_23492_, _23491_, _23489_);
  not (_23493_, rst);
  nand (_23495_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_23496_, \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_23497_, _23496_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_23498_, _23497_);
  nor (_23499_, _23498_, \oc8051_top_1.oc8051_decoder1.state [0]);
  not (_23500_, _23499_);
  nand (_23501_, _23431_, _23408_);
  nor (_23502_, _23501_, _23500_);
  not (_23504_, _23473_);
  nand (_23505_, _23504_, _23335_);
  not (_23507_, _23505_);
  nor (_23508_, _23507_, _23500_);
  not (_23509_, \oc8051_top_1.oc8051_decoder1.state [0]);
  nor (_23510_, \oc8051_top_1.oc8051_sfr1.wait_data , _23509_);
  not (_23512_, _23510_);
  nor (_23513_, _23512_, \oc8051_top_1.oc8051_decoder1.state [1]);
  nor (_23514_, _23253_, _23351_);
  nand (_23515_, _23514_, _23338_);
  nor (_23516_, _23515_, _23283_);
  nand (_23517_, _23516_, _23513_);
  not (_23518_, _23517_);
  nor (_23519_, _23518_, _23508_);
  not (_23520_, _23519_);
  nor (_23521_, _23520_, _23502_);
  nand (_23522_, _23521_, _23495_);
  nand (_23523_, _23522_, _23493_);
  nand (_25023_, _23523_, _23492_);
  nor (_23524_, _22910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  nor (_23525_, _22912_, _21474_);
  nor (_09578_, _23525_, _23524_);
  nor (_23527_, _23422_, _23175_);
  not (_23528_, _23527_);
  nor (_23529_, _23482_, _23528_);
  not (_23531_, _23529_);
  nand (_23532_, _23442_, _23431_);
  nand (_23534_, _23532_, _23531_);
  nand (_23535_, _23413_, _23381_);
  nand (_23536_, _23535_, _23459_);
  nor (_23537_, _23536_, _23534_);
  nor (_23539_, _23537_, _23490_);
  nand (_23540_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_23541_, _23540_, _23517_);
  nor (_23542_, _23541_, _23539_);
  nor (_25020_[1], _23542_, rst);
  nor (_23543_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  nor (_23544_, _22508_, _21626_);
  nor (_10241_, _23544_, _23543_);
  nor (_23545_, _21645_, _21425_);
  nor (_23546_, _23545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  not (_23547_, _23545_);
  nor (_23549_, _23547_, _21414_);
  nor (_25294_, _23549_, _23546_);
  nor (_23551_, _23057_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_23552_, _23551_, _23490_);
  nor (_23553_, _23552_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_23554_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand (_23555_, _23553_, _23210_);
  nand (_23556_, _23555_, _23493_);
  nor (_10326_, _23556_, _23554_);
  nor (_23557_, _21695_, _21658_);
  nor (_23558_, _23557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  not (_23560_, _23557_);
  nor (_23561_, _23560_, _21526_);
  nor (_10590_, _23561_, _23558_);
  nor (_23562_, _21899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  nor (_23563_, _21902_, _21504_);
  nor (_10631_, _23563_, _23562_);
  nor (_23564_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  nor (_23565_, _22783_, _21451_);
  nor (_10652_, _23565_, _23564_);
  nor (_23567_, _23557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  nor (_23568_, _23560_, _21586_);
  nor (_10666_, _23568_, _23567_);
  nor (_23569_, _23557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  nor (_23570_, _23560_, _21626_);
  nor (_10757_, _23570_, _23569_);
  nor (_23571_, _22292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  nor (_23572_, _22294_, _21586_);
  nor (_10779_, _23572_, _23571_);
  nor (_23574_, _21389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  nor (_23575_, _21451_, _21391_);
  nor (_10849_, _23575_, _23574_);
  nor (_23577_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  nor (_23578_, _22696_, _21451_);
  nor (_10894_, _23578_, _23577_);
  nor (_23579_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  nor (_23580_, _22696_, _21504_);
  nor (_10912_, _23580_, _23579_);
  nor (_23581_, _21899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  nor (_23582_, _21902_, _21554_);
  nor (_25123_, _23582_, _23581_);
  nor (_23583_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  nor (_23584_, _22696_, _21526_);
  nor (_25152_, _23584_, _23583_);
  nor (_23585_, _21659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  nor (_23586_, _21661_, _21504_);
  nor (_10974_, _23586_, _23585_);
  nor (_23587_, _22999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  nor (_23588_, _23001_, _21554_);
  nor (_10995_, _23588_, _23587_);
  nor (_23589_, _21659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  nor (_23590_, _21661_, _21526_);
  nor (_11010_, _23590_, _23589_);
  nor (_23591_, _22999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  nor (_23592_, _23001_, _21474_);
  nor (_11025_, _23592_, _23591_);
  nor (_23593_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  nor (_23594_, _22696_, _21414_);
  nor (_11041_, _23594_, _23593_);
  nor (_23595_, _21389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  nor (_23596_, _21474_, _21391_);
  nor (_11057_, _23596_, _23595_);
  nor (_23597_, _22999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  nor (_23598_, _23001_, _21586_);
  nor (_11073_, _23598_, _23597_);
  nor (_23599_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  nor (_23600_, _22783_, _21504_);
  nor (_11142_, _23600_, _23599_);
  nor (_23601_, _23557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  nor (_23602_, _23560_, _21474_);
  nor (_11157_, _23602_, _23601_);
  nor (_23603_, _21899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  nor (_23604_, _21902_, _21414_);
  nor (_11228_, _23604_, _23603_);
  nor (_23606_, _22186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  nor (_23607_, _22188_, _21554_);
  nor (_11290_, _23607_, _23606_);
  nor (_23608_, _22461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  nor (_23609_, _22463_, _21626_);
  nor (_25055_, _23609_, _23608_);
  nor (_23610_, _22461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  nor (_23611_, _22463_, _21526_);
  nor (_25053_, _23611_, _23610_);
  nor (_23612_, _22999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  nor (_23613_, _23001_, _21414_);
  nor (_11366_, _23613_, _23612_);
  nor (_23614_, _22999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  nor (_23615_, _23001_, _21451_);
  nor (_11417_, _23615_, _23614_);
  nor (_23616_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  nor (_23617_, _22418_, _21554_);
  nor (_11432_, _23617_, _23616_);
  nor (_23619_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  nor (_23620_, _22418_, _21586_);
  nor (_11446_, _23620_, _23619_);
  nor (_23622_, _22369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  nor (_23623_, _22371_, _21626_);
  nor (_11460_, _23623_, _23622_);
  nor (_23624_, _22369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  nor (_23625_, _22371_, _21526_);
  nor (_11497_, _23625_, _23624_);
  nor (_23626_, _22369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  nor (_23627_, _22371_, _21474_);
  nor (_11515_, _23627_, _23626_);
  nor (_23628_, _22348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  nor (_23629_, _22351_, _21526_);
  nor (_11583_, _23629_, _23628_);
  nor (_23630_, _22348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  nor (_23631_, _22351_, _21474_);
  nor (_11602_, _23631_, _23630_);
  nor (_23632_, _22316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  nor (_23634_, _22318_, _21414_);
  nor (_25049_, _23634_, _23632_);
  nor (_23636_, _22316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  nor (_23637_, _22318_, _21554_);
  nor (_11665_, _23637_, _23636_);
  nor (_23638_, _22286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  nor (_23639_, _22288_, _21504_);
  nor (_25048_, _23639_, _23638_);
  nor (_23640_, _22286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  nor (_23641_, _22288_, _21474_);
  nor (_11740_, _23641_, _23640_);
  nor (_23642_, _22245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  nor (_23643_, _22248_, _21626_);
  nor (_11757_, _23643_, _23642_);
  nor (_23644_, _22245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  nor (_23646_, _22248_, _21554_);
  nor (_11797_, _23646_, _23644_);
  nor (_23647_, _22050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  nor (_23648_, _22052_, _21586_);
  nor (_11828_, _23648_, _23647_);
  nor (_23650_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  nor (_23651_, _22179_, _21451_);
  nor (_11869_, _23651_, _23650_);
  nor (_23652_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  nor (_23653_, _22179_, _21474_);
  nor (_11909_, _23653_, _23652_);
  nor (_23654_, _22003_, _21599_);
  nor (_23655_, _23654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  not (_23657_, _23654_);
  nor (_23658_, _23657_, _21414_);
  nor (_11930_, _23658_, _23655_);
  nor (_23659_, _22150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  nor (_23660_, _22152_, _21554_);
  nor (_25441_, _23660_, _23659_);
  nor (_23661_, _22150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  nor (_23662_, _22152_, _21586_);
  nor (_11971_, _23662_, _23661_);
  nor (_23663_, _22121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  nor (_23664_, _22123_, _21626_);
  nor (_25440_, _23664_, _23663_);
  nor (_23666_, _22121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  nor (_23667_, _22123_, _21526_);
  nor (_12012_, _23667_, _23666_);
  nor (_23668_, _22121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  nor (_23669_, _22123_, _21474_);
  nor (_12033_, _23669_, _23668_);
  nor (_23670_, _23654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  nor (_23671_, _23657_, _21526_);
  nor (_12054_, _23671_, _23670_);
  nor (_23672_, _22069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  nor (_23673_, _22071_, _21626_);
  nor (_12075_, _23673_, _23672_);
  nor (_23675_, _23654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  nor (_23676_, _23657_, _21554_);
  nor (_12096_, _23676_, _23675_);
  nor (_23677_, _22069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  nor (_23678_, _22071_, _21554_);
  nor (_12117_, _23678_, _23677_);
  nor (_23679_, _22050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  nor (_23680_, _22052_, _21451_);
  nor (_12147_, _23680_, _23679_);
  nor (_23681_, _22069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  nor (_23682_, _22071_, _21586_);
  nor (_12168_, _23682_, _23681_);
  nor (_23683_, _22461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  nor (_23684_, _22463_, _21586_);
  nor (_25052_, _23684_, _23683_);
  nor (_23685_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  nor (_23686_, _22418_, _21414_);
  nor (_12269_, _23686_, _23685_);
  nor (_23687_, _22369_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  nor (_23689_, _22371_, _21451_);
  nor (_25051_, _23689_, _23687_);
  nor (_23690_, _22348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  nor (_23691_, _22351_, _21451_);
  nor (_12340_, _23691_, _23690_);
  nor (_23692_, _22316_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  nor (_23693_, _22318_, _21504_);
  nor (_12378_, _23693_, _23692_);
  nor (_23694_, _22286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  nor (_23695_, _22288_, _21526_);
  nor (_12450_, _23695_, _23694_);
  nor (_23696_, _22245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  nor (_23697_, _22248_, _21414_);
  nor (_12470_, _23697_, _23696_);
  nor (_23698_, _22050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  nor (_23700_, _22052_, _21554_);
  nor (_12485_, _23700_, _23698_);
  nor (_23701_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  nor (_23702_, _22179_, _21626_);
  nor (_12499_, _23702_, _23701_);
  nor (_23704_, _22176_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  nor (_23705_, _22179_, _21526_);
  nor (_12513_, _23705_, _23704_);
  nor (_23707_, _23654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  nor (_23708_, _23657_, _21626_);
  nor (_12529_, _23708_, _23707_);
  nor (_23709_, _22150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  nor (_23710_, _22152_, _21414_);
  nor (_25442_, _23710_, _23709_);
  nor (_23711_, _22121_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  nor (_23713_, _22123_, _21451_);
  nor (_12557_, _23713_, _23711_);
  nor (_23714_, _22069_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  nor (_23716_, _22071_, _21414_);
  nor (_12581_, _23716_, _23714_);
  nor (_23717_, _22050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  nor (_23718_, _22052_, _21626_);
  nor (_12602_, _23718_, _23717_);
  nor (_23719_, _22186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  nor (_23721_, _22188_, _21526_);
  nor (_12623_, _23721_, _23719_);
  nor (_23722_, _22461_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  nor (_23723_, _22463_, _21414_);
  nor (_12644_, _23723_, _23722_);
  nor (_23725_, _23654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  nor (_23726_, _23657_, _21504_);
  nor (_12665_, _23726_, _23725_);
  nor (_23727_, _23654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  nor (_23728_, _23657_, _21451_);
  nor (_12696_, _23728_, _23727_);
  nor (_23729_, _22286_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  nor (_23730_, _22288_, _21626_);
  nor (_12717_, _23730_, _23729_);
  nor (_23732_, _22416_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  nor (_23733_, _22418_, _21451_);
  nor (_12828_, _23733_, _23732_);
  nor (_23735_, _22348_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  nor (_23736_, _22351_, _21504_);
  nor (_25050_, _23736_, _23735_);
  nor (_23737_, _22050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  nor (_23738_, _22052_, _21526_);
  nor (_12869_, _23738_, _23737_);
  nor (_23739_, _22150_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  nor (_23740_, _22152_, _21451_);
  nor (_12890_, _23740_, _23739_);
  nor (_23741_, _22245_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  nor (_23742_, _22248_, _21586_);
  nor (_12911_, _23742_, _23741_);
  nor (_23743_, _22186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  nor (_23744_, _22188_, _21414_);
  nor (_12932_, _23744_, _23743_);
  nor (_23745_, _22021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  nor (_23746_, _22023_, _21526_);
  nor (_12953_, _23746_, _23745_);
  nor (_23747_, _22003_, _21821_);
  nor (_23748_, _23747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  not (_23749_, _23747_);
  nor (_23750_, _23749_, _21414_);
  nor (_12974_, _23750_, _23748_);
  nor (_23751_, _22004_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  nor (_23752_, _22006_, _21554_);
  nor (_13005_, _23752_, _23751_);
  nor (_23753_, _23747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  nor (_23754_, _23749_, _21526_);
  nor (_13026_, _23754_, _23753_);
  nor (_23755_, _22834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  nor (_23756_, _22836_, _21474_);
  nor (_13057_, _23756_, _23755_);
  nor (_23757_, _23747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  nor (_23758_, _23749_, _21554_);
  nor (_13108_, _23758_, _23757_);
  nor (_23759_, _22003_, _21374_);
  nor (_23760_, _23759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  not (_23761_, _23759_);
  nor (_23763_, _23761_, _21451_);
  nor (_13189_, _23763_, _23760_);
  nor (_23764_, _21997_, _22392_);
  not (_23766_, _23764_);
  nor (_23767_, _23766_, _22018_);
  not (_23768_, _23767_);
  nor (_23769_, _23768_, _21689_);
  nor (_23770_, _23769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  not (_23771_, _23769_);
  nor (_23772_, _23771_, _21474_);
  nor (_13250_, _23772_, _23770_);
  nor (_23774_, _23768_, _21631_);
  nor (_23775_, _23774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  not (_23776_, _23774_);
  nor (_23777_, _23776_, _21414_);
  nor (_25392_, _23777_, _23775_);
  nor (_23779_, _23768_, _21482_);
  nor (_23781_, _23779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  not (_23782_, _23779_);
  nor (_23783_, _23782_, _21626_);
  nor (_13332_, _23783_, _23781_);
  nor (_23784_, _23779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  nor (_23785_, _23782_, _21586_);
  nor (_13353_, _23785_, _23784_);
  nor (_23786_, _23768_, _21558_);
  nor (_23788_, _23786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  not (_23789_, _23786_);
  nor (_23790_, _23789_, _21554_);
  nor (_13391_, _23790_, _23788_);
  nor (_23791_, _23768_, _21566_);
  nor (_23792_, _23791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  not (_23793_, _23791_);
  nor (_23794_, _23793_, _21414_);
  nor (_13414_, _23794_, _23792_);
  nor (_23795_, _23768_, _21589_);
  nor (_23796_, _23795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  not (_23797_, _23795_);
  nor (_23798_, _23797_, _21504_);
  nor (_13437_, _23798_, _23796_);
  nor (_23799_, _23768_, _21599_);
  nor (_23800_, _23799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  not (_23801_, _23799_);
  nor (_23802_, _23801_, _21474_);
  nor (_13467_, _23802_, _23800_);
  nor (_23803_, _23766_, _21643_);
  not (_23805_, _23803_);
  nor (_23806_, _23805_, _21652_);
  nor (_23807_, _23806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  not (_23808_, _23806_);
  nor (_23809_, _23808_, _21451_);
  nor (_13516_, _23809_, _23807_);
  nor (_23810_, _23805_, _21689_);
  nor (_23811_, _23810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  not (_23812_, _23810_);
  nor (_23813_, _23812_, _21474_);
  nor (_13555_, _23813_, _23811_);
  nor (_23815_, _23747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  nor (_23816_, _23749_, _21626_);
  nor (_25404_, _23816_, _23815_);
  nor (_23817_, _23805_, _21482_);
  nor (_23818_, _23817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  not (_23819_, _23817_);
  nor (_23821_, _23819_, _21626_);
  nor (_13602_, _23821_, _23818_);
  nor (_23822_, _23747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  nor (_23824_, _23749_, _21504_);
  nor (_13622_, _23824_, _23822_);
  nor (_23825_, _23805_, _21530_);
  nor (_23826_, _23825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  not (_23827_, _23825_);
  nor (_23828_, _23827_, _21474_);
  nor (_13653_, _23828_, _23826_);
  nor (_23829_, _23805_, _21589_);
  nor (_23830_, _23829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  not (_23831_, _23829_);
  nor (_23832_, _23831_, _21414_);
  nor (_13730_, _23832_, _23830_);
  nor (_23833_, _23768_, _21374_);
  nor (_23834_, _23833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  not (_23835_, _23833_);
  nor (_23836_, _23835_, _21451_);
  nor (_13760_, _23836_, _23834_);
  nor (_23837_, _23768_, _21658_);
  nor (_23838_, _23837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  not (_23839_, _23837_);
  nor (_23840_, _23839_, _21626_);
  nor (_13790_, _23840_, _23838_);
  nor (_23841_, _23837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  nor (_23842_, _23839_, _21526_);
  nor (_13810_, _23842_, _23841_);
  nor (_23843_, _22003_, _21482_);
  nor (_23844_, _23843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  not (_23845_, _23843_);
  nor (_23846_, _23845_, _21586_);
  nor (_13878_, _23846_, _23844_);
  nor (_23847_, _23654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  nor (_23848_, _23657_, _21474_);
  nor (_13949_, _23848_, _23847_);
  nor (_23849_, _22003_, _21864_);
  nor (_23850_, _23849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  not (_23851_, _23849_);
  nor (_23852_, _23851_, _21526_);
  nor (_13976_, _23852_, _23850_);
  nor (_23853_, _22003_, _21658_);
  nor (_23854_, _23853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  not (_23855_, _23853_);
  nor (_23856_, _23855_, _21504_);
  nor (_25400_, _23856_, _23854_);
  nor (_23857_, _23768_, _21530_);
  nor (_23858_, _23857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  not (_23859_, _23857_);
  nor (_23860_, _23859_, _21474_);
  nor (_14074_, _23860_, _23858_);
  nor (_23861_, _21804_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  nor (_23862_, _21806_, _21626_);
  nor (_25208_, _23862_, _23861_);
  nor (_23863_, _23849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  nor (_23864_, _23851_, _21451_);
  nor (_14124_, _23864_, _23863_);
  nor (_23865_, _23805_, _21425_);
  nor (_23867_, _23865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  not (_23868_, _23865_);
  nor (_23870_, _23868_, _21504_);
  nor (_14171_, _23870_, _23867_);
  nor (_23871_, _23817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  nor (_23872_, _23819_, _21526_);
  nor (_14190_, _23872_, _23871_);
  nor (_23873_, _23805_, _21607_);
  nor (_23874_, _23873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  not (_23875_, _23873_);
  nor (_23876_, _23875_, _21554_);
  nor (_14225_, _23876_, _23874_);
  nor (_23877_, _23849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  nor (_23878_, _23851_, _21414_);
  nor (_14252_, _23878_, _23877_);
  nor (_23879_, _21796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  nor (_23880_, _21799_, _21586_);
  nor (_14320_, _23880_, _23879_);
  nor (_23881_, _23769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  nor (_23882_, _23771_, _21626_);
  nor (_14341_, _23882_, _23881_);
  nor (_23883_, _23825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  nor (_23884_, _23827_, _21554_);
  nor (_14386_, _23884_, _23883_);
  nor (_23885_, _23833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  nor (_23887_, _23835_, _21504_);
  nor (_14428_, _23887_, _23885_);
  nor (_23888_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  nor (_23889_, _22165_, _21451_);
  nor (_14465_, _23889_, _23888_);
  nor (_23890_, _22113_, _21482_);
  nor (_23891_, _23890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  not (_23892_, _23890_);
  nor (_23893_, _23892_, _21586_);
  nor (_14546_, _23893_, _23891_);
  nor (_23894_, _22113_, _21530_);
  nor (_23895_, _23894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  not (_23896_, _23894_);
  nor (_23897_, _23896_, _21626_);
  nor (_25431_, _23897_, _23895_);
  nor (_23898_, _23894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  nor (_23899_, _23896_, _21474_);
  nor (_14627_, _23899_, _23898_);
  nor (_23900_, _22113_, _21607_);
  nor (_23901_, _23900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  not (_23902_, _23900_);
  nor (_23903_, _23902_, _21626_);
  nor (_25429_, _23903_, _23901_);
  nor (_23904_, _23900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  nor (_23905_, _23902_, _21526_);
  nor (_14704_, _23905_, _23904_);
  nor (_23906_, _23900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  nor (_23907_, _23902_, _21474_);
  nor (_14720_, _23907_, _23906_);
  nor (_23908_, _22113_, _21558_);
  nor (_23909_, _23908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  not (_23910_, _23908_);
  nor (_23911_, _23910_, _21504_);
  nor (_14739_, _23911_, _23909_);
  nor (_23912_, _22113_, _21566_);
  nor (_23913_, _23912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  not (_23914_, _23912_);
  nor (_23915_, _23914_, _21451_);
  nor (_14800_, _23915_, _23913_);
  nor (_23917_, _23912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  nor (_23918_, _23914_, _21474_);
  nor (_14819_, _23918_, _23917_);
  nor (_23919_, _22113_, _21589_);
  nor (_23920_, _23919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  not (_23921_, _23919_);
  nor (_23922_, _23921_, _21504_);
  nor (_14844_, _23922_, _23920_);
  nor (_23923_, _23747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  nor (_23924_, _23749_, _21586_);
  nor (_14868_, _23924_, _23923_);
  nor (_23925_, _23919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  nor (_23926_, _23921_, _21474_);
  nor (_14883_, _23926_, _23925_);
  nor (_23927_, _22113_, _21599_);
  nor (_23928_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  not (_23929_, _23927_);
  nor (_23930_, _23929_, _21451_);
  nor (_14909_, _23930_, _23928_);
  nor (_23931_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  nor (_23932_, _23929_, _21554_);
  nor (_25424_, _23932_, _23931_);
  nor (_23933_, _23849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  nor (_23934_, _23851_, _21626_);
  nor (_25403_, _23934_, _23933_);
  nor (_23935_, _22113_, _21864_);
  nor (_23936_, _23935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  not (_23937_, _23935_);
  nor (_23938_, _23937_, _21451_);
  nor (_25422_, _23938_, _23936_);
  nor (_23939_, _22113_, _21374_);
  nor (_23940_, _23939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  not (_23941_, _23939_);
  nor (_23942_, _23941_, _21626_);
  nor (_15003_, _23942_, _23940_);
  nor (_23943_, _23939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  nor (_23944_, _23941_, _21451_);
  nor (_15020_, _23944_, _23943_);
  nor (_23945_, _23939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  nor (_23946_, _23941_, _21586_);
  nor (_15042_, _23946_, _23945_);
  nor (_23947_, _22113_, _21658_);
  nor (_23948_, _23947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  not (_23949_, _23947_);
  nor (_23950_, _23949_, _21451_);
  nor (_15074_, _23950_, _23948_);
  nor (_23951_, _22113_, _21821_);
  nor (_23952_, _23951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  not (_23953_, _23951_);
  nor (_23954_, _23953_, _21504_);
  nor (_15144_, _23954_, _23952_);
  nor (_23955_, _23951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  nor (_23956_, _23953_, _21414_);
  nor (_15165_, _23956_, _23955_);
  nor (_23957_, _23951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  nor (_23958_, _23953_, _21474_);
  nor (_25423_, _23958_, _23957_);
  nor (_23959_, _23894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  nor (_23960_, _23896_, _21526_);
  nor (_15292_, _23960_, _23959_);
  nor (_23961_, _23900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  nor (_23963_, _23902_, _21451_);
  nor (_15337_, _23963_, _23961_);
  nor (_23964_, _23759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  nor (_23965_, _23761_, _21626_);
  nor (_25402_, _23965_, _23964_);
  nor (_23966_, _23908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  nor (_23967_, _23910_, _21526_);
  nor (_25427_, _23967_, _23966_);
  nor (_23968_, _23908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  nor (_23969_, _23910_, _21586_);
  nor (_15400_, _23969_, _23968_);
  nor (_23970_, _23919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  nor (_23971_, _23921_, _21526_);
  nor (_15481_, _23971_, _23970_);
  nor (_23972_, _23759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  nor (_23973_, _23761_, _21504_);
  nor (_15502_, _23973_, _23972_);
  nor (_23974_, _23935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  nor (_23975_, _23937_, _21586_);
  nor (_15573_, _23975_, _23974_);
  nor (_23976_, _21790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  nor (_23977_, _21792_, _21586_);
  nor (_15614_, _23977_, _23976_);
  nor (_23978_, _23947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  nor (_23979_, _23949_, _21626_);
  nor (_15635_, _23979_, _23978_);
  nor (_23980_, _23947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  nor (_23981_, _23949_, _21474_);
  nor (_25420_, _23981_, _23980_);
  nor (_23982_, _21790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  nor (_23983_, _21792_, _21474_);
  nor (_25212_, _23983_, _23982_);
  nor (_23984_, _23912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  nor (_23985_, _23914_, _21554_);
  nor (_15736_, _23985_, _23984_);
  nor (_23987_, _23939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  nor (_23989_, _23941_, _21554_);
  nor (_15788_, _23989_, _23987_);
  nor (_23990_, _23849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  nor (_23991_, _23851_, _21474_);
  nor (_15959_, _23991_, _23990_);
  nor (_23992_, _23768_, _21638_);
  nor (_23993_, _23992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  not (_23994_, _23992_);
  nor (_23996_, _23994_, _21626_);
  nor (_15990_, _23996_, _23993_);
  nor (_23997_, _23951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  nor (_23998_, _23953_, _21586_);
  nor (_16011_, _23998_, _23997_);
  nor (_23999_, _23992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  nor (_24000_, _23994_, _21451_);
  nor (_16032_, _24000_, _23999_);
  nor (_24002_, _23849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  nor (_24003_, _23851_, _21586_);
  nor (_16053_, _24003_, _24002_);
  nor (_24004_, _23935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  nor (_24005_, _23937_, _21504_);
  nor (_16074_, _24005_, _24004_);
  nor (_24006_, _23806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  nor (_24008_, _23808_, _21626_);
  nor (_25372_, _24008_, _24006_);
  nor (_24010_, _23992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  nor (_24011_, _23994_, _21554_);
  nor (_25373_, _24011_, _24010_);
  nor (_24012_, _23935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  nor (_24013_, _23937_, _21626_);
  nor (_16135_, _24013_, _24012_);
  nor (_24014_, _23951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  nor (_24015_, _23953_, _21554_);
  nor (_16154_, _24015_, _24014_);
  nor (_24016_, _23951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  nor (_24017_, _23953_, _21526_);
  nor (_16224_, _24017_, _24016_);
  nor (_24018_, _23837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  nor (_24019_, _23839_, _21414_);
  nor (_16244_, _24019_, _24018_);
  nor (_24020_, _23833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  nor (_24021_, _23835_, _21474_);
  nor (_16271_, _24021_, _24020_);
  nor (_24022_, _23951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  nor (_24023_, _23953_, _21451_);
  nor (_16291_, _24023_, _24022_);
  nor (_24025_, _23951_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  nor (_24026_, _23953_, _21626_);
  nor (_16318_, _24026_, _24025_);
  nor (_24027_, _22113_, _21638_);
  nor (_24028_, _24027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  not (_24029_, _24027_);
  nor (_24030_, _24029_, _21626_);
  nor (_16384_, _24030_, _24028_);
  nor (_24031_, _23759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  nor (_24032_, _23761_, _21586_);
  nor (_16404_, _24032_, _24031_);
  nor (_24033_, _23947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  nor (_24034_, _23949_, _21586_);
  nor (_16443_, _24034_, _24033_);
  nor (_24035_, _23829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  nor (_24036_, _23831_, _21626_);
  nor (_25358_, _24036_, _24035_);
  nor (_24038_, _23853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  nor (_24039_, _23855_, _21626_);
  nor (_16478_, _24039_, _24038_);
  nor (_24041_, _23947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  nor (_24042_, _23949_, _21554_);
  nor (_16519_, _24042_, _24041_);
  nor (_24043_, _23805_, _21566_);
  nor (_24044_, _24043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  not (_24045_, _24043_);
  nor (_24046_, _24045_, _21414_);
  nor (_16550_, _24046_, _24044_);
  nor (_24048_, _23947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  nor (_24049_, _23949_, _21526_);
  nor (_16601_, _24049_, _24048_);
  nor (_24050_, _23805_, _21558_);
  nor (_24051_, _24050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  not (_24052_, _24050_);
  nor (_24053_, _24052_, _21451_);
  nor (_16672_, _24053_, _24051_);
  nor (_24054_, _23947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  nor (_24055_, _23949_, _21414_);
  nor (_16693_, _24055_, _24054_);
  nor (_24057_, _23947_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  nor (_24058_, _23949_, _21504_);
  nor (_16724_, _24058_, _24057_);
  nor (_24059_, _23873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  nor (_24060_, _23875_, _21474_);
  nor (_25366_, _24060_, _24059_);
  nor (_24061_, _23759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  nor (_24062_, _23761_, _21414_);
  nor (_25401_, _24062_, _24061_);
  nor (_24063_, _23873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  nor (_24064_, _23875_, _21451_);
  nor (_16825_, _24064_, _24063_);
  nor (_24065_, _23873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  nor (_24066_, _23875_, _21414_);
  nor (_16846_, _24066_, _24065_);
  nor (_24067_, _23939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  nor (_24068_, _23941_, _21474_);
  nor (_16867_, _24068_, _24067_);
  nor (_24069_, _23939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  nor (_24070_, _23941_, _21526_);
  nor (_16908_, _24070_, _24069_);
  nor (_24071_, _23825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  nor (_24072_, _23827_, _21504_);
  nor (_16929_, _24072_, _24071_);
  nor (_24073_, _23759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  nor (_24074_, _23761_, _21526_);
  nor (_16950_, _24074_, _24073_);
  nor (_24075_, _23759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  nor (_24076_, _23761_, _21554_);
  nor (_16971_, _24076_, _24075_);
  nor (_24077_, _23817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  nor (_24078_, _23819_, _21554_);
  nor (_16992_, _24078_, _24077_);
  nor (_24079_, _23939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  nor (_24080_, _23941_, _21414_);
  nor (_17013_, _24080_, _24079_);
  nor (_24081_, _23817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  nor (_24082_, _23819_, _21586_);
  nor (_17034_, _24082_, _24081_);
  nor (_24083_, _23939_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  nor (_24084_, _23941_, _21504_);
  nor (_17085_, _24084_, _24083_);
  nor (_24085_, _23817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  nor (_24086_, _23819_, _21451_);
  nor (_17106_, _24086_, _24085_);
  nor (_24087_, _23865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  nor (_24088_, _23868_, _21451_);
  nor (_17137_, _24088_, _24087_);
  nor (_24089_, _23865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  nor (_24090_, _23868_, _21554_);
  nor (_17158_, _24090_, _24089_);
  nor (_24091_, _23935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  nor (_24092_, _23937_, _21474_);
  nor (_17180_, _24092_, _24091_);
  nor (_24094_, _23805_, _21631_);
  nor (_24095_, _24094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  not (_24096_, _24094_);
  nor (_24097_, _24096_, _21526_);
  nor (_17211_, _24097_, _24095_);
  nor (_24098_, _23935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  nor (_24100_, _23937_, _21554_);
  nor (_17232_, _24100_, _24098_);
  nor (_24101_, _23935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  nor (_24102_, _23937_, _21526_);
  nor (_17258_, _24102_, _24101_);
  nor (_24103_, _23853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  nor (_24104_, _23855_, _21474_);
  nor (_17393_, _24104_, _24103_);
  nor (_24105_, _23935_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  nor (_24107_, _23937_, _21414_);
  nor (_25421_, _24107_, _24105_);
  nor (_24108_, _23806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  nor (_24109_, _23808_, _21474_);
  nor (_25371_, _24109_, _24108_);
  nor (_24110_, _23768_, _21864_);
  nor (_24111_, _24110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  not (_24112_, _24110_);
  nor (_24113_, _24112_, _21554_);
  nor (_25379_, _24113_, _24111_);
  nor (_24115_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  nor (_24117_, _23929_, _21586_);
  nor (_17515_, _24117_, _24115_);
  nor (_24118_, _24110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  nor (_24119_, _24112_, _21586_);
  nor (_17536_, _24119_, _24118_);
  nor (_24120_, _23853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  nor (_24121_, _23855_, _21586_);
  nor (_17557_, _24121_, _24120_);
  nor (_24122_, _24110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  nor (_24123_, _24112_, _21626_);
  nor (_17578_, _24123_, _24122_);
  nor (_24125_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  nor (_24126_, _23929_, _21474_);
  nor (_17599_, _24126_, _24125_);
  nor (_24127_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  nor (_24128_, _23929_, _21526_);
  nor (_17650_, _24128_, _24127_);
  nor (_24129_, _23768_, _21821_);
  nor (_24130_, _24129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  not (_24131_, _24129_);
  nor (_24132_, _24131_, _21414_);
  nor (_17681_, _24132_, _24130_);
  nor (_24133_, _24129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  nor (_24134_, _24131_, _21474_);
  nor (_25380_, _24134_, _24133_);
  nor (_24135_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  nor (_24136_, _23929_, _21414_);
  nor (_25425_, _24136_, _24135_);
  nor (_24137_, _24129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  nor (_24138_, _24131_, _21626_);
  nor (_17752_, _24138_, _24137_);
  nor (_24140_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  nor (_24142_, _23929_, _21504_);
  nor (_17777_, _24142_, _24140_);
  nor (_24143_, _23799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  nor (_24144_, _23801_, _21451_);
  nor (_17798_, _24144_, _24143_);
  nor (_24145_, _23927_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  nor (_24146_, _23929_, _21626_);
  nor (_17819_, _24146_, _24145_);
  nor (_24147_, _23919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  nor (_24148_, _23921_, _21586_);
  nor (_17840_, _24148_, _24147_);
  nor (_24149_, _23919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  nor (_24150_, _23921_, _21554_);
  nor (_17871_, _24150_, _24149_);
  nor (_24151_, _23853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  nor (_24152_, _23855_, _21414_);
  nor (_17892_, _24152_, _24151_);
  nor (_24153_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  not (_24154_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_24155_, _23553_, _24154_);
  nand (_24156_, _24155_, _23493_);
  nor (_25042_[13], _24156_, _24153_);
  nor (_24157_, _23919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  nor (_24158_, _23921_, _21414_);
  nor (_25426_, _24158_, _24157_);
  nor (_24159_, _23768_, _21607_);
  nor (_24160_, _24159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  not (_24161_, _24159_);
  nor (_24162_, _24161_, _21554_);
  nor (_25386_, _24162_, _24160_);
  nor (_24163_, _23853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  nor (_24164_, _23855_, _21526_);
  nor (_17983_, _24164_, _24163_);
  nor (_24165_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand (_24166_, _23553_, _23098_);
  nand (_24167_, _24166_, _23493_);
  nor (_18004_, _24167_, _24165_);
  nand (_24168_, _23490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_24169_, _24168_);
  not (_24170_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  nor (_24171_, _23153_, _24170_);
  nor (_24172_, _23058_, _23070_);
  nor (_24173_, _23067_, _23052_);
  nor (_24174_, _24173_, _24172_);
  not (_24175_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nor (_24176_, _23050_, _24175_);
  nor (_24177_, _23107_, _23048_);
  nor (_24178_, _24177_, _24176_);
  nand (_24179_, _24178_, _24174_);
  not (_24180_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor (_24181_, _23073_, _24180_);
  not (_24183_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_24184_, _23076_, _24183_);
  nor (_24185_, _24184_, _24181_);
  not (_24186_, _24185_);
  nor (_24187_, _24186_, _24179_);
  nor (_24188_, _24187_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_24189_, _24188_, _24171_);
  nor (_24190_, _24189_, _23490_);
  nor (_24191_, _24190_, _24169_);
  nor (_18025_, _24191_, rst);
  nor (_24192_, _23857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  nor (_24193_, _23859_, _21586_);
  nor (_18046_, _24193_, _24192_);
  nor (_24194_, _23919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  nor (_24195_, _23921_, _21451_);
  nor (_18067_, _24195_, _24194_);
  nor (_24196_, _21757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  nor (_24197_, _21759_, _21504_);
  nor (_18089_, _24197_, _24196_);
  nor (_24198_, _23919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  nor (_24199_, _23921_, _21626_);
  nor (_18110_, _24199_, _24198_);
  nor (_24200_, _22227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  nor (_24201_, _22229_, _21586_);
  nor (_18131_, _24201_, _24200_);
  nor (_24202_, _23912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  nor (_24203_, _23914_, _21586_);
  nor (_18152_, _24203_, _24202_);
  nor (_24204_, _23912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  nor (_24205_, _23914_, _21526_);
  nor (_18183_, _24205_, _24204_);
  nor (_24206_, _23768_, _21425_);
  nor (_24207_, _24206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  not (_24208_, _24206_);
  nor (_24209_, _24208_, _21626_);
  nor (_25389_, _24209_, _24207_);
  nor (_24210_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  nor (_24211_, _22240_, _21626_);
  nor (_18264_, _24211_, _24210_);
  nor (_24212_, _22003_, _21638_);
  nor (_24213_, _24212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  not (_24214_, _24212_);
  nor (_24215_, _24214_, _21526_);
  nor (_18305_, _24215_, _24213_);
  nor (_24216_, _23912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  nor (_24217_, _23914_, _21414_);
  nor (_18326_, _24217_, _24216_);
  nor (_24218_, _23912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  nor (_24219_, _23914_, _21504_);
  nor (_18347_, _24219_, _24218_);
  nor (_24220_, _24212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  nor (_24221_, _24214_, _21554_);
  nor (_18368_, _24221_, _24220_);
  nor (_24222_, _23769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  nor (_24223_, _23771_, _21504_);
  nor (_18409_, _24223_, _24222_);
  nor (_24224_, _23912_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  nor (_24225_, _23914_, _21626_);
  nor (_18430_, _24225_, _24224_);
  nor (_24226_, _23769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  nor (_24227_, _23771_, _21414_);
  nor (_25394_, _24227_, _24226_);
  nor (_24229_, _23908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  nor (_24230_, _23910_, _21474_);
  nor (_18471_, _24230_, _24229_);
  nor (_24231_, _23768_, _21652_);
  nor (_24232_, _24231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  not (_24233_, _24231_);
  nor (_24234_, _24233_, _21451_);
  nor (_25397_, _24234_, _24232_);
  nor (_24235_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  nor (_24236_, _22240_, _21451_);
  nor (_18522_, _24236_, _24235_);
  nor (_24238_, _24231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  nor (_24239_, _24233_, _21554_);
  nor (_25396_, _24239_, _24238_);
  nor (_24240_, _24212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  nor (_24241_, _24214_, _21474_);
  nor (_18587_, _24241_, _24240_);
  nor (_24242_, _23908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  nor (_24243_, _23910_, _21554_);
  nor (_18605_, _24243_, _24242_);
  nor (_24244_, _23908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  nor (_24245_, _23910_, _21414_);
  nor (_18629_, _24245_, _24244_);
  nor (_24246_, _24212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  nor (_24247_, _24214_, _21626_);
  nor (_18645_, _24247_, _24246_);
  nor (_24248_, _24212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  nor (_24249_, _24214_, _21414_);
  nor (_18659_, _24249_, _24248_);
  nor (_24250_, _23853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  nor (_24251_, _23855_, _21451_);
  nor (_18690_, _24251_, _24250_);
  nor (_24252_, _23908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  nor (_24253_, _23910_, _21451_);
  nor (_18711_, _24253_, _24252_);
  nor (_24254_, _23853_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  nor (_24255_, _23855_, _21554_);
  nor (_25399_, _24255_, _24254_);
  nor (_24256_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  nor (_24257_, _22240_, _21414_);
  nor (_25174_, _24257_, _24256_);
  nor (_24258_, _23908_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  nor (_24260_, _23910_, _21626_);
  nor (_25428_, _24260_, _24258_);
  nor (_24261_, _23759_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  nor (_24263_, _23761_, _21474_);
  nor (_18792_, _24263_, _24261_);
  nor (_24264_, _23849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  nor (_24265_, _23851_, _21554_);
  nor (_18833_, _24265_, _24264_);
  nor (_24266_, _23900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  nor (_24267_, _23902_, _21586_);
  nor (_18854_, _24267_, _24266_);
  nor (_24268_, _23747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  nor (_24269_, _23749_, _21474_);
  nor (_18895_, _24269_, _24268_);
  nor (_24271_, _23900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  nor (_24272_, _23902_, _21554_);
  nor (_18916_, _24272_, _24271_);
  nor (_24273_, _23849_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  nor (_24274_, _23851_, _21504_);
  nor (_18937_, _24274_, _24273_);
  nor (_24275_, _23900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  nor (_24276_, _23902_, _21414_);
  nor (_18958_, _24276_, _24275_);
  nor (_24277_, _23654_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  nor (_24278_, _23657_, _21586_);
  nor (_18980_, _24278_, _24277_);
  nor (_24279_, _22238_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  nor (_24280_, _22240_, _21474_);
  nor (_25173_, _24280_, _24279_);
  nor (_24282_, _23747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  nor (_24283_, _23749_, _21451_);
  nor (_19021_, _24283_, _24282_);
  nor (_24284_, _23900_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  nor (_24286_, _23902_, _21504_);
  nor (_19072_, _24286_, _24284_);
  nor (_24287_, _24212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  nor (_24288_, _24214_, _21504_);
  nor (_25398_, _24288_, _24287_);
  nor (_24289_, _22999_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  nor (_24290_, _23001_, _21526_);
  nor (_19153_, _24290_, _24289_);
  nor (_24291_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand (_24292_, _23553_, _23385_);
  nand (_24293_, _24292_, _23493_);
  nor (_19174_, _24293_, _24291_);
  nor (_24294_, _22910_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  nor (_24295_, _22912_, _21554_);
  nor (_19195_, _24295_, _24294_);
  nor (_24296_, _23894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  nor (_24297_, _23896_, _21586_);
  nor (_19216_, _24297_, _24296_);
  nor (_24298_, _23894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  nor (_24299_, _23896_, _21554_);
  nor (_19237_, _24299_, _24298_);
  nor (_24300_, _24212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  nor (_24301_, _24214_, _21451_);
  nor (_19258_, _24301_, _24300_);
  nor (_24302_, _21757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  nor (_24303_, _21759_, _21451_);
  nor (_19279_, _24303_, _24302_);
  nor (_24304_, _23894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  nor (_24305_, _23896_, _21414_);
  nor (_19301_, _24305_, _24304_);
  nor (_24306_, _22834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  nor (_24307_, _22836_, _21626_);
  nor (_19322_, _24307_, _24306_);
  nor (_24308_, _23894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  nor (_24309_, _23896_, _21451_);
  nor (_25430_, _24309_, _24308_);
  nor (_24310_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  nor (_24312_, _22594_, _21414_);
  nor (_25410_, _24312_, _24310_);
  nor (_24313_, _22592_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  nor (_24314_, _22594_, _21474_);
  nor (_19393_, _24314_, _24313_);
  nor (_24315_, _23894_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  nor (_24316_, _23896_, _21504_);
  nor (_19452_, _24316_, _24315_);
  nor (_24317_, _24231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  nor (_24318_, _24233_, _21626_);
  nor (_19806_, _24318_, _24317_);
  nor (_24319_, _24231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  nor (_24320_, _24233_, _21504_);
  nor (_19837_, _24320_, _24319_);
  nor (_24322_, _22186_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  nor (_24324_, _22188_, _21451_);
  nor (_20369_, _24324_, _24322_);
  nor (_24325_, _22113_, _21425_);
  nor (_24326_, _24325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  not (_24327_, _24325_);
  nor (_24328_, _24327_, _21451_);
  nor (_20867_, _24328_, _24326_);
  nor (_24329_, _23890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  nor (_24330_, _23892_, _21451_);
  nor (_25432_, _24330_, _24329_);
  nor (_24331_, _22003_, _21631_);
  nor (_24332_, _24331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  not (_24333_, _24331_);
  nor (_24335_, _24333_, _21626_);
  nor (_20868_, _24335_, _24332_);
  nor (_24336_, _23890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  nor (_24337_, _23892_, _21414_);
  nor (_20869_, _24337_, _24336_);
  nor (_24340_, _23890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  nor (_24342_, _23892_, _21504_);
  nor (_25433_, _24342_, _24340_);
  nor (_24343_, _22003_, _21689_);
  nor (_24344_, _24343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  not (_24345_, _24343_);
  nor (_24346_, _24345_, _21554_);
  nor (_20870_, _24346_, _24344_);
  nor (_24348_, _22250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  nor (_24349_, _22252_, _21504_);
  nor (_20871_, _24349_, _24348_);
  nor (_24350_, _22250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  nor (_24351_, _22252_, _21414_);
  nor (_20872_, _24351_, _24350_);
  nor (_24352_, _22114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  nor (_24353_, _22116_, _21474_);
  nor (_20873_, _24353_, _24352_);
  nor (_24355_, _24212_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  nor (_24357_, _24214_, _21586_);
  nor (_20874_, _24357_, _24355_);
  nor (_24359_, _24325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  nor (_24360_, _24327_, _21586_);
  nor (_20875_, _24360_, _24359_);
  nor (_24361_, _23890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  nor (_24362_, _23892_, _21626_);
  nor (_20876_, _24362_, _24361_);
  nor (_24363_, _21741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  nor (_24364_, _21744_, _21626_);
  nor (_20877_, _24364_, _24363_);
  nor (_24365_, _22003_, _21652_);
  nor (_24366_, _24365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  not (_24367_, _24365_);
  nor (_24368_, _24367_, _21626_);
  nor (_20878_, _24368_, _24366_);
  nor (_24369_, _24325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  nor (_24370_, _24327_, _21474_);
  nor (_25434_, _24370_, _24369_);
  nor (_24372_, _24027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  nor (_24373_, _24029_, _21451_);
  nor (_25418_, _24373_, _24372_);
  nor (_24375_, _22114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  nor (_24376_, _22116_, _21451_);
  nor (_20880_, _24376_, _24375_);
  nor (_24378_, _24231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  nor (_24379_, _24233_, _21474_);
  nor (_20881_, _24379_, _24378_);
  nor (_24380_, _21645_, _21482_);
  nor (_24381_, _24380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  not (_24382_, _24380_);
  nor (_24383_, _24382_, _21626_);
  nor (_20882_, _24383_, _24381_);
  nor (_24384_, _24231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  nor (_24385_, _24233_, _21586_);
  nor (_20883_, _24385_, _24384_);
  nand (_24386_, _23043_, _21183_);
  nand (_24387_, _23405_, _23148_);
  nor (_24389_, _24387_, _23330_);
  nor (_24390_, _24389_, _23455_);
  nor (_24391_, _23454_, _23407_);
  nor (_24393_, _24387_, _23454_);
  nor (_24394_, _24393_, _24391_);
  nand (_24395_, _24394_, _24390_);
  not (_24396_, _23465_);
  nand (_24397_, _23429_, _23471_);
  nor (_24398_, _24397_, _23409_);
  nand (_24399_, _24398_, _23283_);
  nand (_24400_, _24399_, _24396_);
  nor (_24401_, _24400_, _24395_);
  nand (_24402_, _23480_, _23449_);
  nor (_24403_, _23306_, _23149_);
  nor (_24404_, _23454_, _23283_);
  nand (_24405_, _24404_, _24403_);
  nand (_24406_, _24405_, _24402_);
  nor (_24407_, _23454_, _23415_);
  nor (_24408_, _23454_, _23424_);
  nor (_24409_, _24408_, _24407_);
  nand (_24410_, _23462_, _23283_);
  nor (_24411_, _23454_, _24410_);
  nand (_24412_, _23480_, _23088_);
  nor (_24413_, _24412_, _23326_);
  nor (_24414_, _24413_, _24411_);
  nand (_24416_, _24414_, _24409_);
  nor (_24417_, _24416_, _24406_);
  nand (_24419_, _24417_, _24401_);
  nand (_24420_, _24419_, _24386_);
  nor (_24421_, _23528_, _24410_);
  nand (_24422_, _23423_, _23283_);
  nor (_24423_, _24422_, _23528_);
  nor (_24424_, _24423_, _24421_);
  nand (_24425_, _24424_, _23531_);
  nand (_24426_, _24425_, _24386_);
  nand (_24427_, _24426_, _24420_);
  nand (_24428_, _23431_, _23423_);
  nor (_24429_, _24428_, _23500_);
  nor (_24430_, _23498_, _23509_);
  nand (_24431_, _24430_, _24389_);
  not (_24432_, _24431_);
  nor (_24433_, _24432_, _24429_);
  not (_24434_, _24433_);
  nor (_24435_, _24434_, _24427_);
  nor (_25016_[0], _24435_, rst);
  nor (_24436_, _24331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  nor (_24437_, _24333_, _21586_);
  nor (_20884_, _24437_, _24436_);
  nor (_24438_, _23890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  nor (_24439_, _23892_, _21526_);
  nor (_20885_, _24439_, _24438_);
  nor (_24440_, _22003_, _21425_);
  nor (_24441_, _24440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  not (_24442_, _24440_);
  nor (_24443_, _24442_, _21504_);
  nor (_25414_, _24443_, _24441_);
  nor (_24444_, _23843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  nor (_24445_, _23845_, _21451_);
  nor (_20886_, _24445_, _24444_);
  nor (_24446_, _23890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  nor (_24447_, _23892_, _21474_);
  nor (_20887_, _24447_, _24446_);
  nor (_24448_, _23843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  nor (_24449_, _23845_, _21554_);
  nor (_20888_, _24449_, _24448_);
  nor (_24450_, _22250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  nor (_24451_, _22252_, _21554_);
  nor (_20889_, _24451_, _24450_);
  nor (_24452_, _24440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  nor (_24453_, _24442_, _21526_);
  nor (_20890_, _24453_, _24452_);
  nor (_24454_, _23890_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  nor (_24455_, _23892_, _21554_);
  nor (_20891_, _24455_, _24454_);
  nor (_24456_, _21913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  nor (_24457_, _21915_, _21504_);
  nor (_20892_, _24457_, _24456_);
  nor (_24458_, _22250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  nor (_24459_, _22252_, _21586_);
  nor (_20893_, _24459_, _24458_);
  not (_24460_, _24386_);
  nor (_24461_, _23482_, _24397_);
  not (_24462_, _24461_);
  nand (_24463_, _23306_, _23150_);
  nand (_24464_, _24463_, _23464_);
  nand (_24465_, _24464_, _23440_);
  nand (_24466_, _24465_, _24462_);
  not (_24467_, _24466_);
  nand (_24468_, _23428_, _23283_);
  nand (_24469_, _24468_, _23333_);
  nand (_24470_, _24469_, _23255_);
  nand (_24471_, _23428_, _23088_);
  nand (_24472_, _23415_, _24471_);
  nand (_24473_, _24472_, _23440_);
  nand (_24474_, _24473_, _24470_);
  nand (_24475_, _23327_, _23255_);
  nor (_24476_, _24397_, _23415_);
  nor (_24477_, _23326_, _23422_);
  nor (_24478_, _24477_, _24476_);
  nand (_24479_, _24478_, _24475_);
  nor (_24480_, _24479_, _24474_);
  nand (_24481_, _24480_, _24467_);
  nor (_24482_, _23337_, _23323_);
  nand (_24483_, _23306_, _24482_);
  nor (_24484_, _24483_, _23283_);
  nor (_24485_, _23331_, _23337_);
  nor (_24486_, _24485_, _24484_);
  nand (_24487_, _24410_, _23415_);
  nor (_24488_, _23427_, _23404_);
  nand (_24489_, _24488_, _23283_);
  nand (_24490_, _24403_, _23088_);
  nand (_24491_, _24490_, _24489_);
  nor (_24492_, _24491_, _24487_);
  nand (_24493_, _24492_, _24486_);
  nand (_24494_, _24493_, _23255_);
  nor (_24495_, _24397_, _23333_);
  nor (_24496_, _24387_, _24397_);
  nor (_24497_, _24496_, _24495_);
  nor (_24498_, _23440_, _23359_);
  nor (_24499_, _24498_, _23482_);
  nand (_24500_, _23338_, _23148_);
  nor (_24501_, _24412_, _24500_);
  nor (_24502_, _24501_, _24389_);
  nand (_24503_, _24502_, _23342_);
  nor (_24504_, _24503_, _24499_);
  nand (_24505_, _24504_, _24497_);
  nor (_24506_, _24505_, _23447_);
  nand (_24507_, _24506_, _24494_);
  nor (_24508_, _24507_, _24481_);
  nor (_24509_, _24508_, _24460_);
  nand (_24510_, _24485_, _23440_);
  nor (_24511_, _24510_, _23498_);
  nand (_24512_, _24511_, \oc8051_top_1.oc8051_decoder1.state [0]);
  nor (_24513_, _24397_, _23326_);
  nand (_24514_, _24513_, _23499_);
  not (_24515_, _24514_);
  nor (_24516_, _24515_, _24429_);
  nand (_24517_, _24516_, _24512_);
  nor (_24518_, _24517_, _24509_);
  nor (_25016_[1], _24518_, rst);
  nor (_24519_, _24231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  nor (_24520_, _24233_, _21414_);
  nor (_20895_, _24520_, _24519_);
  nor (_24521_, _23805_, _21599_);
  nor (_24522_, _24521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  not (_24523_, _24521_);
  nor (_24524_, _24523_, _21626_);
  nor (_20897_, _24524_, _24522_);
  nor (_24525_, _24521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  nor (_24526_, _24523_, _21414_);
  nor (_20899_, _24526_, _24525_);
  nor (_24527_, _24521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  nor (_24528_, _24523_, _21586_);
  nor (_20900_, _24528_, _24527_);
  nor (_24529_, _23805_, _21821_);
  nor (_24530_, _24529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  not (_24531_, _24529_);
  nor (_24532_, _24531_, _21626_);
  nor (_20901_, _24532_, _24530_);
  nor (_24533_, _24529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  nor (_24534_, _24531_, _21451_);
  nor (_20902_, _24534_, _24533_);
  nor (_24535_, _24231_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  nor (_24536_, _24233_, _21526_);
  nor (_20903_, _24536_, _24535_);
  nor (_24537_, _23805_, _21864_);
  nor (_24538_, _24537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  not (_24539_, _24537_);
  nor (_24540_, _24539_, _21414_);
  nor (_20904_, _24540_, _24538_);
  nor (_24541_, _24537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  nor (_24542_, _24539_, _21586_);
  nor (_20905_, _24542_, _24541_);
  nor (_24543_, _22259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  nor (_24544_, _22261_, _21626_);
  nor (_20906_, _24544_, _24543_);
  nor (_24545_, _23805_, _21374_);
  nor (_24546_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  not (_24547_, _24545_);
  nor (_24548_, _24547_, _21451_);
  nor (_20907_, _24548_, _24546_);
  nor (_24549_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  nor (_24550_, _24547_, _21554_);
  nor (_20908_, _24550_, _24549_);
  nor (_24551_, _23805_, _21658_);
  nor (_24552_, _24551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  not (_24553_, _24551_);
  nor (_24554_, _24553_, _21626_);
  nor (_20910_, _24554_, _24552_);
  nor (_24555_, _24551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  nor (_24556_, _24553_, _21526_);
  nor (_25353_, _24556_, _24555_);
  nor (_24557_, _24551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  nor (_24558_, _24553_, _21586_);
  nor (_20911_, _24558_, _24557_);
  nor (_24559_, _23805_, _21638_);
  nor (_24560_, _24559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  not (_24561_, _24559_);
  nor (_24562_, _24561_, _21626_);
  nor (_20912_, _24562_, _24560_);
  nor (_24563_, _24559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  nor (_24564_, _24561_, _21451_);
  nor (_20913_, _24564_, _24563_);
  nor (_24565_, _24559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  nor (_24566_, _24561_, _21586_);
  nor (_20915_, _24566_, _24565_);
  nor (_24567_, _23766_, _21385_);
  not (_24568_, _24567_);
  nor (_24569_, _24568_, _21652_);
  nor (_24570_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  not (_24571_, _24569_);
  nor (_24572_, _24571_, _21504_);
  nor (_20916_, _24572_, _24570_);
  nor (_24573_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  nor (_24574_, _24571_, _21414_);
  nor (_20917_, _24574_, _24573_);
  nor (_24575_, _24568_, _21631_);
  nor (_24576_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  not (_24577_, _24575_);
  nor (_24578_, _24577_, _21504_);
  nor (_20918_, _24578_, _24576_);
  nor (_24579_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  nor (_24580_, _24577_, _21414_);
  nor (_20919_, _24580_, _24579_);
  nor (_24581_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  nor (_24582_, _24577_, _21586_);
  nor (_20920_, _24582_, _24581_);
  nor (_24583_, _24568_, _21425_);
  nor (_24584_, _24583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  not (_24585_, _24583_);
  nor (_24586_, _24585_, _21626_);
  nor (_25345_, _24586_, _24584_);
  nor (_24587_, _24583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  nor (_24588_, _24585_, _21451_);
  nor (_20921_, _24588_, _24587_);
  nor (_24589_, _23769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  nor (_24590_, _23771_, _21526_);
  nor (_25393_, _24590_, _24589_);
  nor (_24591_, _24583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  nor (_24592_, _24585_, _21474_);
  nor (_20922_, _24592_, _24591_);
  nor (_24593_, _24568_, _21482_);
  nor (_24594_, _24593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  not (_24595_, _24593_);
  nor (_24596_, _24595_, _21504_);
  nor (_20924_, _24596_, _24594_);
  nor (_24597_, _23769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  nor (_24598_, _23771_, _21554_);
  nor (_20925_, _24598_, _24597_);
  nor (_24599_, _24593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  nor (_24600_, _24595_, _21554_);
  nor (_20926_, _24600_, _24599_);
  nor (_24601_, _24568_, _21530_);
  nor (_24602_, _24601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  not (_24603_, _24601_);
  nor (_24604_, _24603_, _21626_);
  nor (_20927_, _24604_, _24602_);
  nor (_24605_, _22259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  nor (_24606_, _22261_, _21451_);
  nor (_20928_, _24606_, _24605_);
  nor (_24607_, _24568_, _21689_);
  nor (_24608_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  not (_24609_, _24607_);
  nor (_24610_, _24609_, _21554_);
  nor (_20929_, _24610_, _24608_);
  nor (_24611_, _23528_, _23339_);
  nor (_24612_, _24490_, _23422_);
  nor (_24613_, _24612_, _24611_);
  nand (_24614_, _23404_, _24482_);
  nor (_24615_, _24614_, _24397_);
  nand (_24616_, _24615_, _23088_);
  nand (_24617_, _24616_, _24613_);
  nand (_25017_[0], _24617_, _23491_);
  nor (_24618_, _24529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  nor (_24619_, _24531_, _21474_);
  nor (_20930_, _24619_, _24618_);
  nor (_24620_, _24537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  nor (_24621_, _24539_, _21504_);
  nor (_20931_, _24621_, _24620_);
  nor (_24622_, _24537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  nor (_24623_, _24539_, _21554_);
  nor (_25356_, _24623_, _24622_);
  nor (_24624_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  nor (_24625_, _24547_, _21626_);
  nor (_20932_, _24625_, _24624_);
  nor (_24626_, _24559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  nor (_24627_, _24561_, _21554_);
  nor (_25350_, _24627_, _24626_);
  nor (_24628_, _23769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  nor (_24629_, _23771_, _21451_);
  nor (_25395_, _24629_, _24628_);
  nor (_24630_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  nor (_24631_, _24609_, _21626_);
  nor (_20933_, _24631_, _24630_);
  nor (_24632_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  nor (_24633_, _24609_, _21414_);
  nor (_20934_, _24633_, _24632_);
  nor (_24634_, _24521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  nor (_24635_, _24523_, _21474_);
  nor (_20935_, _24635_, _24634_);
  not (_24636_, _24611_);
  not (_24637_, _24615_);
  nand (_24638_, _24637_, _24636_);
  nand (_25017_[1], _24638_, _23491_);
  nor (_24640_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  nor (_24641_, _24547_, _21526_);
  nor (_20936_, _24641_, _24640_);
  nor (_24642_, _24551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  nor (_24643_, _24553_, _21414_);
  nor (_20937_, _24643_, _24642_);
  nor (_24644_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  nor (_24645_, _24609_, _21586_);
  nor (_20938_, _24645_, _24644_);
  nor (_24646_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  nor (_24647_, _24577_, _21474_);
  nor (_20939_, _24647_, _24646_);
  nor (_24648_, _24583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  nor (_24649_, _24585_, _21554_);
  nor (_20940_, _24649_, _24648_);
  nor (_24650_, _24593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  nor (_24651_, _24595_, _21526_);
  nor (_20941_, _24651_, _24650_);
  nor (_24652_, _24529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  nor (_24653_, _24531_, _21554_);
  nor (_25357_, _24653_, _24652_);
  nor (_24654_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  nor (_24655_, _24571_, _21474_);
  nor (_20942_, _24655_, _24654_);
  nor (_24657_, _22869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  nor (_24659_, _22872_, _21526_);
  nor (_20943_, _24659_, _24657_);
  nor (_24661_, _24568_, _21558_);
  nor (_24662_, _24661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  not (_24663_, _24661_);
  nor (_24665_, _24663_, _21451_);
  nor (_20944_, _24665_, _24662_);
  nor (_24666_, _24568_, _21566_);
  nor (_24667_, _24666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  not (_24668_, _24666_);
  nor (_24669_, _24668_, _21474_);
  nor (_20945_, _24669_, _24667_);
  nor (_24670_, _24568_, _21589_);
  nor (_24671_, _24670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  not (_24672_, _24670_);
  nor (_24673_, _24672_, _21526_);
  nor (_20946_, _24673_, _24671_);
  nor (_24674_, _24568_, _21864_);
  nor (_24675_, _24674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  not (_24676_, _24674_);
  nor (_24677_, _24676_, _21504_);
  nor (_20948_, _24677_, _24675_);
  nor (_24678_, _24674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  nor (_24679_, _24676_, _21586_);
  nor (_20949_, _24679_, _24678_);
  nor (_24680_, _23774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  nor (_24681_, _23776_, _21626_);
  nor (_20950_, _24681_, _24680_);
  nor (_24682_, _22263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  nor (_24683_, _22265_, _21451_);
  nor (_25162_, _24683_, _24682_);
  nor (_24684_, _24568_, _21638_);
  nor (_24685_, _24684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  not (_24686_, _24684_);
  nor (_24687_, _24686_, _21414_);
  nor (_20951_, _24687_, _24685_);
  nor (_24688_, _23766_, _21995_);
  not (_24689_, _24688_);
  nor (_24690_, _24689_, _21689_);
  nor (_24691_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  not (_24692_, _24690_);
  nor (_24693_, _24692_, _21414_);
  nor (_25132_, _24693_, _24691_);
  nor (_24694_, _23774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  nor (_24695_, _23776_, _21504_);
  nor (_20952_, _24695_, _24694_);
  nor (_24696_, _24689_, _21425_);
  nor (_24697_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  not (_24698_, _24696_);
  nor (_24699_, _24698_, _21554_);
  nor (_20954_, _24699_, _24697_);
  nor (_24700_, _23774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  nor (_24701_, _23776_, _21451_);
  nor (_20955_, _24701_, _24700_);
  nor (_24702_, _24689_, _21530_);
  nor (_24703_, _24702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  not (_24704_, _24702_);
  nor (_24705_, _24704_, _21451_);
  nor (_20956_, _24705_, _24703_);
  nor (_24706_, _24689_, _21566_);
  nor (_24707_, _24706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  not (_24708_, _24706_);
  nor (_24709_, _24708_, _21451_);
  nor (_20957_, _24709_, _24707_);
  nor (_24710_, _24689_, _21821_);
  nor (_24711_, _24710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  not (_24712_, _24710_);
  nor (_24713_, _24712_, _21626_);
  nor (_20958_, _24713_, _24711_);
  nor (_24714_, _24387_, _23088_);
  not (_24715_, _24714_);
  nor (_24716_, _24715_, _24397_);
  nor (_24717_, _24716_, _24495_);
  nor (_24718_, _24717_, _23500_);
  nor (_24719_, _23464_, _23330_);
  nor (_24720_, _24719_, _24476_);
  not (_24721_, _24720_);
  nor (_24722_, _24410_, _23330_);
  nor (_24723_, _23404_, _23323_);
  nand (_24724_, _24723_, _23414_);
  nor (_24725_, _24724_, _23330_);
  nor (_24726_, _24725_, _24461_);
  nand (_24727_, _24726_, _23441_);
  nor (_24728_, _24727_, _24722_);
  nor (_24729_, _23482_, _23330_);
  not (_24730_, _24717_);
  nor (_24731_, _24730_, _24729_);
  not (_24732_, _24731_);
  nor (_24733_, _23415_, _23330_);
  nor (_24734_, _24471_, _23330_);
  nor (_24735_, _24734_, _24733_);
  nor (_24736_, _24387_, _23283_);
  nand (_24737_, _24736_, _23431_);
  nand (_24738_, _24737_, _24735_);
  nor (_24739_, _24738_, _24732_);
  nand (_24740_, _24739_, _24728_);
  nor (_24741_, _24740_, _24721_);
  nor (_24742_, _24741_, _24460_);
  nor (_24743_, _24742_, _24718_);
  nand (_24744_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_24745_, _24479_);
  nand (_24746_, _24745_, _23420_);
  nor (_24747_, _24746_, _24466_);
  not (_24748_, _24486_);
  nor (_24749_, _23442_, _23416_);
  nor (_24750_, _24614_, _23283_);
  nor (_24751_, _24750_, _23449_);
  nand (_24752_, _24751_, _24749_);
  nor (_24753_, _24752_, _24748_);
  nor (_24754_, _24753_, _23382_);
  nand (_24755_, _24484_, _23282_);
  nor (_24756_, _24471_, _23382_);
  nor (_24757_, _24398_, _24756_);
  nand (_24758_, _24757_, _24755_);
  nor (_24759_, _23407_, _23283_);
  nand (_24760_, _24759_, _23255_);
  nor (_24761_, _24468_, _23330_);
  nor (_24762_, _24722_, _24761_);
  nand (_24763_, _24762_, _24760_);
  nor (_24764_, _24763_, _24758_);
  not (_24765_, _24496_);
  nand (_24766_, _24765_, _23501_);
  nor (_24767_, _23482_, _23203_);
  nor (_24768_, _24729_, _24767_);
  nor (_24769_, _23464_, _23382_);
  nand (_24770_, _24404_, _23481_);
  nand (_24771_, _24770_, _24510_);
  nor (_24773_, _24771_, _24769_);
  nand (_24774_, _24773_, _24768_);
  nor (_24775_, _24774_, _24766_);
  nand (_24776_, _24775_, _24764_);
  nor (_24777_, _24776_, _24754_);
  nand (_24778_, _24777_, _24747_);
  nand (_24779_, _24778_, _24386_);
  not (_24780_, _24517_);
  nand (_24781_, _24780_, _24779_);
  nand (_24782_, _24781_, _21183_);
  nand (_24783_, _24782_, _24744_);
  nand (_24784_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_24785_, _24784_);
  not (_24786_, _24429_);
  nor (_24788_, _24463_, _23528_);
  not (_24789_, _24788_);
  nor (_24790_, _24421_, _23529_);
  nand (_24791_, _24790_, _24789_);
  nand (_24792_, _24791_, _24386_);
  nand (_24793_, _24792_, _24786_);
  nor (_24794_, _23461_, _23283_);
  nand (_24795_, _24794_, _23514_);
  not (_24796_, _24795_);
  nor (_24797_, _24515_, _24796_);
  not (_24798_, _24797_);
  nor (_24799_, _24798_, _24793_);
  nor (_24800_, _24799_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_24801_, _24800_, _24785_);
  nand (_24802_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_24803_, _24802_);
  nor (_24804_, _24435_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_24805_, _24804_, _24803_);
  nand (_24807_, _24805_, _24801_);
  nor (_24808_, _24807_, _24783_);
  not (_24809_, _24808_);
  nor (_24810_, _24809_, _23279_);
  not (_24811_, _24512_);
  nor (_24812_, _24793_, _24811_);
  nand (_24813_, _24812_, _24420_);
  nand (_24814_, _24813_, _21183_);
  nand (_24815_, _24814_, _24802_);
  not (_24816_, _24744_);
  nor (_24817_, _24518_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_24818_, _24817_, _24816_);
  nor (_24819_, _24818_, _24815_);
  nand (_24820_, _24819_, _24801_);
  nand (_24821_, _23490_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  not (_24822_, _24821_);
  nor (_24823_, _23490_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_24824_, _24823_);
  nor (_24826_, _23058_, _23257_);
  nor (_24827_, _23107_, _23259_);
  nor (_24828_, _24827_, _24826_);
  not (_24829_, _24828_);
  not (_24830_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nor (_24831_, _23073_, _24830_);
  nor (_24832_, _23076_, _23264_);
  nor (_24833_, _24832_, _24831_);
  nor (_24834_, _23050_, _23233_);
  not (_24835_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_24836_, _23067_, _24835_);
  nor (_24837_, _24836_, _24834_);
  nand (_24838_, _24837_, _24833_);
  nor (_24839_, _24838_, _24829_);
  nor (_24840_, _24839_, _24824_);
  nor (_24841_, _24840_, _24822_);
  nor (_24842_, _24841_, _24820_);
  nor (_24843_, _24842_, _24810_);
  nor (_24844_, _24783_, _24805_);
  nand (_24845_, _24844_, _24801_);
  not (_24847_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_24848_, _21336_, _21268_);
  not (_24849_, _24848_);
  nand (_24850_, _21278_, _21270_);
  nor (_24851_, _24850_, _21280_);
  not (_24852_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_24853_, _21259_, _24852_);
  nor (_24854_, _21282_, _24853_);
  nand (_24855_, _24854_, _24851_);
  not (_24856_, _21320_);
  nor (_24857_, _24856_, _24855_);
  nand (_24858_, _24857_, _21351_);
  nor (_24859_, _21184_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  not (_24860_, _24859_);
  nor (_24861_, _24860_, _21186_);
  nand (_24862_, _24861_, _21308_);
  nor (_24863_, _24862_, _24858_);
  nand (_24864_, _24863_, _21426_);
  nor (_24865_, _24864_, _24849_);
  nor (_24866_, _24865_, _24847_);
  not (_24867_, ABINPUT[6]);
  not (_24868_, _24865_);
  nor (_24869_, _24868_, _24867_);
  nor (_24870_, _24869_, _24866_);
  not (_24871_, _24870_);
  nor (_24872_, _24871_, _21308_);
  not (_24873_, _21295_);
  nand (_24874_, _21296_, _24873_);
  nor (_24875_, _24874_, _21303_);
  nor (_24876_, _21305_, _21300_);
  nand (_24877_, _24876_, _24875_);
  nor (_24878_, _24870_, _24877_);
  nor (_24879_, _24878_, _24872_);
  nor (_24880_, _23175_, _24856_);
  nor (_24881_, _23351_, _21320_);
  nor (_24882_, _24860_, _21336_);
  nand (_24883_, _21351_, _21285_);
  nor (_24884_, _24883_, _21377_);
  nand (_24885_, _24884_, _24882_);
  nor (_24886_, _24885_, _21246_);
  not (_24887_, _24886_);
  nor (_24888_, _24887_, _24881_);
  not (_24889_, _24888_);
  nor (_24890_, _24889_, _24880_);
  not (_24891_, _24890_);
  nand (_24892_, _21262_, _21208_);
  not (_24893_, _21251_);
  nand (_24894_, _21263_, _24893_);
  nor (_24895_, _24894_, _24892_);
  nor (_24896_, _21260_, _21256_);
  nand (_24897_, _24896_, _24895_);
  not (_24898_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_24899_, _24865_, _24898_);
  not (_24900_, ABINPUT[7]);
  nor (_24901_, _21268_, _21227_);
  nor (_24902_, _24858_, _24877_);
  not (_24903_, _24902_);
  nor (_24904_, _21365_, _21336_);
  nand (_24905_, _24904_, _24861_);
  nor (_24906_, _24905_, _24903_);
  nand (_24907_, _24906_, _24901_);
  nor (_24908_, _24907_, _24900_);
  nor (_24909_, _24908_, _24899_);
  nor (_24910_, _24909_, _24897_);
  not (_24911_, _24910_);
  nand (_24912_, _24909_, _24897_);
  nand (_24913_, _24912_, _24911_);
  nor (_24914_, _24913_, _24891_);
  nand (_24915_, _24914_, _24879_);
  nor (_24916_, _24915_, ABINPUT[4]);
  not (_24917_, _24916_);
  not (_24918_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nand (_24919_, _24870_, _23175_);
  nor (_24920_, _24919_, _24909_);
  not (_24921_, _24920_);
  nor (_24922_, _24921_, _24918_);
  not (_24923_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_24924_, _24870_, _23351_);
  nand (_24925_, _24924_, _24909_);
  nor (_24926_, _24925_, _24923_);
  nor (_24927_, _24926_, _24922_);
  not (_24928_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  not (_24929_, _24909_);
  nor (_24930_, _24871_, _23175_);
  nand (_24931_, _24930_, _24929_);
  nor (_24932_, _24931_, _24928_);
  not (_24933_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nand (_24934_, _24930_, _24909_);
  nor (_24935_, _24934_, _24933_);
  nor (_24936_, _24935_, _24932_);
  nand (_24937_, _24936_, _24927_);
  not (_24938_, _24937_);
  not (_24939_, _24915_);
  not (_24940_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_24941_, _24870_, _23175_);
  not (_24942_, _24941_);
  nor (_24943_, _24942_, _24909_);
  not (_24944_, _24943_);
  nor (_24945_, _24944_, _24940_);
  not (_24946_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_24947_, _24942_, _24929_);
  not (_24948_, _24947_);
  nor (_24949_, _24948_, _24946_);
  nor (_24950_, _24949_, _24945_);
  not (_24951_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nand (_24952_, _24924_, _24929_);
  nor (_24953_, _24952_, _24951_);
  not (_24954_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_24955_, _24919_, _24929_);
  not (_24956_, _24955_);
  nor (_24957_, _24956_, _24954_);
  nor (_24958_, _24957_, _24953_);
  nand (_24959_, _24958_, _24950_);
  nor (_24960_, _24959_, _24939_);
  nand (_24961_, _24960_, _24938_);
  nand (_24962_, _24961_, _24917_);
  nor (_24963_, _24962_, _24845_);
  not (_00002_, _24801_);
  nand (_00003_, _24844_, _00002_);
  nand (_00004_, _24783_, _24815_);
  nor (_00005_, _00004_, _00002_);
  not (_00006_, ABINPUT[4]);
  nand (_00007_, _21365_, _21337_);
  nand (_00008_, _21268_, _21246_);
  nor (_00009_, _00008_, _00007_);
  not (_00010_, _24861_);
  nor (_00011_, _24883_, _21320_);
  nand (_00013_, _00011_, _21308_);
  nor (_00014_, _00013_, _00010_);
  nand (_00015_, _00014_, _00009_);
  nor (_00016_, _00015_, _00006_);
  nor (_00017_, _21336_, _24897_);
  nand (_00018_, _00017_, _21378_);
  nor (_00019_, _21320_, _24855_);
  nand (_00020_, _00019_, _21351_);
  nor (_00021_, _00020_, _24877_);
  nand (_00022_, _00021_, _24861_);
  nor (_00023_, _00022_, _00018_);
  not (_00024_, _21278_);
  nand (_00025_, _00015_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nand (_00026_, _00023_, ABINPUT[4]);
  nand (_00027_, _00026_, _00025_);
  nor (_00028_, _00023_, _21274_);
  not (_00029_, ABINPUT[3]);
  nor (_00030_, _00015_, _00029_);
  nor (_00031_, _00030_, _00028_);
  nand (_00032_, _00031_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_00033_, _00032_, _00027_);
  nor (_00034_, _00023_, _21273_);
  nor (_00035_, _00016_, _00034_);
  not (_00036_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nand (_00037_, _00015_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nand (_00038_, _00023_, ABINPUT[3]);
  nand (_00039_, _00038_, _00037_);
  nor (_00040_, _00039_, _00036_);
  nor (_00041_, _00040_, _00035_);
  nor (_00042_, _00041_, _00033_);
  nor (_00043_, _00042_, _21202_);
  nor (_00045_, _00043_, _00024_);
  nor (_00046_, _00045_, _00023_);
  nor (_00047_, _00046_, _00016_);
  not (_00048_, _00047_);
  nand (_00049_, _00048_, _00005_);
  nand (_00050_, _00049_, _00003_);
  nor (_00051_, _00050_, _24963_);
  nand (_00052_, _00051_, _24843_);
  nand (_00053_, _00052_, _24743_);
  not (_00054_, \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  nor (_00055_, _23044_, _00054_);
  nor (_00056_, _23058_, _23388_);
  not (_00057_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_00058_, _23107_, _00057_);
  nor (_00059_, _00058_, _00056_);
  not (_00060_, _00059_);
  not (_00062_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nor (_00063_, _23073_, _00062_);
  nor (_00064_, _23067_, _23391_);
  nor (_00066_, _00064_, _00063_);
  nor (_00067_, _23076_, _23286_);
  nor (_00068_, _23050_, _23385_);
  nor (_00069_, _00068_, _00067_);
  nand (_00070_, _00069_, _00066_);
  nor (_00071_, _00070_, _00060_);
  nor (_00072_, _00071_, _24824_);
  nor (_00073_, _00072_, _00055_);
  not (_00074_, _00073_);
  nand (_00075_, _00074_, _24819_);
  nor (_00076_, _24915_, ABINPUT[10]);
  not (_00077_, _00076_);
  nand (_00078_, _24955_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  not (_00079_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_00080_, _24925_, _00079_);
  nand (_00081_, _24947_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  not (_00083_, _00081_);
  nor (_00084_, _00083_, _00080_);
  nand (_00085_, _00084_, _00078_);
  nand (_00086_, _24943_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  not (_00088_, _00086_);
  not (_00089_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor (_00090_, _24952_, _00089_);
  nor (_00091_, _00090_, _00088_);
  nand (_00092_, _24920_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nand (_00093_, _00092_, _00091_);
  nor (_00094_, _00093_, _00085_);
  not (_00095_, _24931_);
  nand (_00096_, _00095_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  not (_00097_, _24934_);
  nand (_00098_, _00097_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nand (_00099_, _00098_, _00096_);
  nor (_00100_, _00099_, _24939_);
  nand (_00101_, _00100_, _00094_);
  nand (_00103_, _00101_, _00077_);
  nor (_00104_, _00103_, _24845_);
  nor (_00105_, _24818_, _24805_);
  not (_00106_, ABINPUT[10]);
  nor (_00107_, _00015_, _00106_);
  not (_00108_, _00107_);
  nor (_00110_, _00023_, _21187_);
  nor (_00111_, _00110_, _00107_);
  not (_00112_, _00111_);
  nor (_00113_, _00023_, _21233_);
  not (_00114_, ABINPUT[9]);
  nor (_00115_, _00015_, _00114_);
  nor (_00116_, _00115_, _00113_);
  nor (_00117_, _00015_, _24867_);
  nor (_00118_, _00023_, _21291_);
  nor (_00119_, _00118_, _00117_);
  nor (_00120_, _00023_, _21235_);
  not (_00121_, ABINPUT[5]);
  nor (_00122_, _00015_, _00121_);
  nor (_00123_, _00122_, _00120_);
  not (_00124_, _00123_);
  nand (_00125_, _00040_, _00035_);
  nor (_00126_, _00125_, _00124_);
  nand (_00127_, _00126_, _00119_);
  nor (_00128_, _00023_, _21188_);
  not (_00129_, ABINPUT[8]);
  nor (_00130_, _00015_, _00129_);
  nor (_00131_, _00130_, _00128_);
  nor (_00132_, _00023_, _21234_);
  nor (_00133_, _00015_, _24900_);
  nor (_00134_, _00133_, _00132_);
  nand (_00135_, _00134_, _00131_);
  nor (_00136_, _00135_, _00127_);
  nand (_00137_, _00136_, _00116_);
  nand (_00138_, _00137_, _00112_);
  not (_00139_, _00116_);
  not (_00141_, _00119_);
  nand (_00142_, _00033_, _00123_);
  nor (_00143_, _00142_, _00141_);
  not (_00144_, _00135_);
  nand (_00145_, _00144_, _00143_);
  nor (_00146_, _00145_, _00139_);
  nand (_00147_, _00146_, _00111_);
  nand (_00148_, _00147_, _00138_);
  nand (_00149_, _00148_, _21290_);
  nand (_00150_, _00149_, _21243_);
  nand (_00151_, _00150_, _00015_);
  nand (_00152_, _00151_, _00108_);
  nand (_00153_, _00152_, _00105_);
  nand (_00154_, _00153_, _24801_);
  nor (_00155_, _00154_, _00104_);
  nand (_00156_, _00155_, _00075_);
  nor (_00157_, _24743_, _00156_);
  nand (_00158_, _23490_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  not (_00159_, _00158_);
  nor (_00160_, _23058_, _23048_);
  nor (_00161_, _23107_, _23052_);
  nor (_00162_, _00161_, _00160_);
  not (_00163_, _00162_);
  nor (_00164_, _23073_, _24175_);
  nor (_00165_, _23067_, _24183_);
  nor (_00167_, _00165_, _00164_);
  nor (_00168_, _23076_, _23065_);
  nor (_00169_, _23050_, _23070_);
  nor (_00170_, _00169_, _00168_);
  nand (_00171_, _00170_, _00167_);
  nor (_00173_, _00171_, _00163_);
  nor (_00174_, _00173_, _24824_);
  nor (_00175_, _00174_, _00159_);
  nor (_00176_, _00175_, _24820_);
  nor (_00177_, _24809_, _24909_);
  nor (_00178_, _00177_, _00176_);
  nor (_00179_, _24915_, ABINPUT[7]);
  not (_00180_, _00179_);
  not (_00181_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor (_00182_, _24944_, _00181_);
  not (_00183_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_00184_, _24956_, _00183_);
  nor (_00185_, _00184_, _00182_);
  not (_00186_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor (_00187_, _24952_, _00186_);
  not (_00188_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_00189_, _24934_, _00188_);
  nor (_00190_, _00189_, _00187_);
  nand (_00191_, _00190_, _00185_);
  not (_00192_, _00191_);
  not (_00194_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_00195_, _24948_, _00194_);
  not (_00196_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_00197_, _24925_, _00196_);
  nor (_00198_, _00197_, _00195_);
  not (_00199_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_00200_, _24931_, _00199_);
  not (_00201_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  nor (_00202_, _24921_, _00201_);
  nor (_00203_, _00202_, _00200_);
  nand (_00204_, _00203_, _00198_);
  nor (_00205_, _00204_, _24939_);
  nand (_00206_, _00205_, _00192_);
  nand (_00207_, _00206_, _00180_);
  nor (_00208_, _00207_, _24845_);
  not (_00209_, _00134_);
  nor (_00210_, _00209_, _00127_);
  nor (_00211_, _00134_, _00143_);
  nor (_00212_, _00211_, _00210_);
  nor (_00213_, _00212_, _21202_);
  nor (_00216_, _00213_, _21251_);
  nor (_00217_, _00216_, _00023_);
  nor (_00218_, _00217_, _00133_);
  not (_00219_, _00218_);
  nand (_00220_, _00219_, _00005_);
  nor (_00221_, _24815_, _24801_);
  not (_00222_, _00221_);
  nand (_00223_, _00222_, _00220_);
  nor (_00224_, _00223_, _00208_);
  nand (_00225_, _00224_, _00178_);
  nand (_00226_, _00225_, _00157_);
  nand (_00227_, _00226_, _00053_);
  nor (_00228_, _00227_, _21287_);
  not (_00229_, _00228_);
  nand (_00230_, _00227_, _21287_);
  nand (_00231_, _00230_, _00229_);
  nor (_00232_, _23331_, _23088_);
  nor (_00233_, _23510_, _24397_);
  nand (_00234_, _00233_, _00232_);
  nor (_00235_, _24476_, _24466_);
  nor (_00237_, _24765_, _23283_);
  nor (_00238_, _00237_, _24729_);
  nand (_00239_, _00238_, _24473_);
  nor (_00240_, _00239_, _23444_);
  nand (_00241_, _00240_, _00235_);
  nand (_00242_, _00241_, _24386_);
  nand (_00243_, _00242_, _00234_);
  not (_00244_, _00243_);
  nor (_00245_, _00244_, _00156_);
  not (_00246_, _00225_);
  nor (_00247_, _00246_, _00245_);
  not (_00248_, _00247_);
  nor (_00249_, _00248_, _21380_);
  nor (_00250_, _24915_, ABINPUT[8]);
  not (_00251_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_00252_, _24931_, _00251_);
  not (_00253_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  nor (_00254_, _24925_, _00253_);
  nor (_00255_, _00254_, _00252_);
  not (_00256_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_00258_, _24944_, _00256_);
  not (_00259_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_00260_, _24934_, _00259_);
  nor (_00261_, _00260_, _00258_);
  nand (_00262_, _00261_, _00255_);
  not (_00263_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor (_00264_, _24921_, _00263_);
  not (_00265_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nor (_00266_, _24956_, _00265_);
  nor (_00267_, _00266_, _00264_);
  not (_00268_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor (_00269_, _24952_, _00268_);
  not (_00270_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_00271_, _24948_, _00270_);
  nor (_00272_, _00271_, _00269_);
  nand (_00273_, _00272_, _00267_);
  nor (_00274_, _00273_, _24939_);
  not (_00275_, _00274_);
  nor (_00276_, _00275_, _00262_);
  nor (_00277_, _00276_, _00250_);
  not (_00279_, _00277_);
  nor (_00280_, _00279_, _24845_);
  nand (_00281_, _23490_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  not (_00282_, _00281_);
  not (_00283_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_00284_, _23058_, _00283_);
  not (_00285_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_00286_, _23107_, _00285_);
  nor (_00287_, _00286_, _00284_);
  not (_00288_, _00287_);
  not (_00290_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nor (_00291_, _23073_, _00290_);
  not (_00292_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_00293_, _23067_, _00292_);
  nor (_00294_, _00293_, _00291_);
  nor (_00295_, _23076_, _23124_);
  nor (_00296_, _23050_, _24154_);
  nor (_00297_, _00296_, _00295_);
  nand (_00298_, _00297_, _00294_);
  nor (_00299_, _00298_, _00288_);
  nor (_00300_, _00299_, _24824_);
  nor (_00301_, _00300_, _00282_);
  nor (_00302_, _00301_, _24820_);
  nor (_00303_, _00302_, _00280_);
  not (_00304_, _00303_);
  not (_00305_, _21329_);
  nor (_00306_, _00210_, _00131_);
  nor (_00307_, _00306_, _00136_);
  nor (_00308_, _00307_, _21202_);
  nor (_00309_, _00308_, _00305_);
  nor (_00310_, _00309_, _00023_);
  nor (_00311_, _00310_, _00130_);
  nor (_00312_, _00311_, _24805_);
  nor (_00313_, _00312_, _00002_);
  nor (_00314_, _24819_, _24844_);
  not (_00315_, _00314_);
  nor (_00316_, _00315_, _00313_);
  nor (_00317_, _00316_, _00304_);
  not (_00318_, _00317_);
  nor (_00319_, _00318_, _00245_);
  not (_00320_, _00319_);
  nor (_00321_, _00320_, _21639_);
  nor (_00322_, _00321_, _00249_);
  nor (_00323_, _24915_, ABINPUT[9]);
  not (_00324_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_00325_, _24944_, _00324_);
  not (_00326_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_00327_, _24934_, _00326_);
  nor (_00328_, _00327_, _00325_);
  not (_00329_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nor (_00331_, _24952_, _00329_);
  not (_00332_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_00333_, _24948_, _00332_);
  nor (_00334_, _00333_, _00331_);
  nand (_00335_, _00334_, _00328_);
  not (_00336_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor (_00337_, _24931_, _00336_);
  not (_00338_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_00339_, _24956_, _00338_);
  nor (_00340_, _00339_, _00337_);
  not (_00341_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor (_00342_, _24921_, _00341_);
  not (_00343_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  nor (_00344_, _24925_, _00343_);
  nor (_00345_, _00344_, _00342_);
  nand (_00346_, _00345_, _00340_);
  nor (_00347_, _00346_, _24939_);
  not (_00348_, _00347_);
  nor (_00349_, _00348_, _00335_);
  nor (_00350_, _00349_, _00323_);
  not (_00352_, _00350_);
  nor (_00353_, _00352_, _24845_);
  nand (_00354_, _00105_, _24801_);
  nor (_00355_, _00136_, _00116_);
  nor (_00356_, _00355_, _00146_);
  nor (_00357_, _00356_, _21202_);
  nor (_00358_, _00357_, _21357_);
  nor (_00359_, _00358_, _00023_);
  nor (_00360_, _00359_, _00115_);
  nor (_00361_, _00360_, _00354_);
  nor (_00362_, _00361_, _00353_);
  nand (_00363_, _23490_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  not (_00364_, _00363_);
  nor (_00365_, _23058_, _23103_);
  not (_00366_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_00367_, _23107_, _00366_);
  nor (_00368_, _00367_, _00365_);
  not (_00369_, _00368_);
  not (_00370_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nor (_00371_, _23073_, _00370_);
  nor (_00372_, _23067_, _23105_);
  nor (_00373_, _00372_, _00371_);
  nor (_00374_, _23076_, _23100_);
  nor (_00375_, _23050_, _23098_);
  nor (_00376_, _00375_, _00374_);
  nand (_00377_, _00376_, _00373_);
  nor (_00378_, _00377_, _00369_);
  nor (_00379_, _00378_, _24824_);
  nor (_00380_, _00379_, _00364_);
  nor (_00381_, _00380_, _24820_);
  nor (_00382_, _24844_, _24801_);
  nor (_00383_, _00382_, _00381_);
  nand (_00384_, _00383_, _00362_);
  not (_00385_, _00384_);
  nor (_00386_, _00385_, _00245_);
  nor (_00387_, _00386_, _21996_);
  nand (_00388_, _00386_, _21996_);
  not (_00389_, _00388_);
  nor (_00390_, _00389_, _00387_);
  nand (_00391_, _00390_, _00322_);
  nor (_00393_, _00391_, _00231_);
  not (_00394_, _21368_);
  nor (_00395_, _24915_, ABINPUT[6]);
  not (_00397_, _00395_);
  not (_00398_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_00399_, _24921_, _00398_);
  not (_00400_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_00401_, _24925_, _00400_);
  nor (_00402_, _00401_, _00399_);
  not (_00403_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_00404_, _24944_, _00403_);
  not (_00405_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_00406_, _24934_, _00405_);
  nor (_00407_, _00406_, _00404_);
  nand (_00408_, _00407_, _00402_);
  not (_00409_, _00408_);
  not (_00410_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor (_00411_, _24931_, _00410_);
  not (_00412_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_00413_, _24956_, _00412_);
  nor (_00415_, _00413_, _00411_);
  not (_00416_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor (_00417_, _24952_, _00416_);
  not (_00418_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_00420_, _24948_, _00418_);
  nor (_00421_, _00420_, _00417_);
  nand (_00422_, _00421_, _00415_);
  nor (_00423_, _00422_, _24939_);
  nand (_00424_, _00423_, _00409_);
  nand (_00425_, _00424_, _00397_);
  nor (_00426_, _00425_, _24845_);
  not (_00427_, _00426_);
  nor (_00428_, _00126_, _00119_);
  nor (_00429_, _00428_, _00143_);
  nor (_00430_, _00429_, _21202_);
  nor (_00431_, _00430_, _21295_);
  nor (_00432_, _00431_, _00023_);
  nor (_00433_, _00432_, _00117_);
  nor (_00434_, _00433_, _00354_);
  nand (_00435_, _24808_, _24871_);
  nor (_00437_, _24807_, _24818_);
  not (_00438_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_00439_, _23044_, _00438_);
  nor (_00440_, _23058_, _23188_);
  nor (_00441_, _23107_, _23185_);
  nor (_00442_, _00441_, _00440_);
  not (_00443_, _00442_);
  not (_00444_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_00445_, _23073_, _00444_);
  nor (_00446_, _23067_, _23190_);
  nor (_00447_, _00446_, _00445_);
  not (_00448_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_00449_, _23076_, _00448_);
  nor (_00450_, _23050_, _23183_);
  nor (_00451_, _00450_, _00449_);
  nand (_00452_, _00451_, _00447_);
  nor (_00453_, _00452_, _00443_);
  nor (_00454_, _24824_, _00453_);
  nor (_00455_, _00454_, _00439_);
  not (_00456_, _00455_);
  nand (_00458_, _00456_, _00437_);
  nand (_00459_, _00458_, _00435_);
  nor (_00460_, _00459_, _00434_);
  nand (_00461_, _00460_, _00427_);
  nor (_00462_, _00245_, _00461_);
  nand (_00463_, _00385_, _00245_);
  not (_00464_, _00463_);
  nor (_00465_, _00464_, _00462_);
  not (_00466_, _00465_);
  nor (_00467_, _00466_, _00394_);
  nor (_00468_, _00465_, _21368_);
  nor (_00469_, _00468_, _00467_);
  nor (_00470_, _24915_, ABINPUT[5]);
  not (_00471_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_00472_, _24944_, _00471_);
  not (_00473_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_00474_, _24934_, _00473_);
  nor (_00475_, _00474_, _00472_);
  not (_00476_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor (_00477_, _24952_, _00476_);
  not (_00478_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_00479_, _24948_, _00478_);
  nor (_00480_, _00479_, _00477_);
  nand (_00481_, _00480_, _00475_);
  not (_00482_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor (_00483_, _24931_, _00482_);
  not (_00484_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  nor (_00485_, _24956_, _00484_);
  nor (_00486_, _00485_, _00483_);
  not (_00487_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_00489_, _24921_, _00487_);
  not (_00490_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_00491_, _24925_, _00490_);
  nor (_00492_, _00491_, _00489_);
  nand (_00493_, _00492_, _00486_);
  nor (_00494_, _00493_, _24939_);
  not (_00495_, _00494_);
  nor (_00496_, _00495_, _00481_);
  nor (_00497_, _00496_, _00470_);
  not (_00498_, _00497_);
  nor (_00499_, _00498_, _24845_);
  nand (_00500_, _23490_, \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  not (_00501_, _00500_);
  nor (_00502_, _23058_, _23215_);
  nor (_00503_, _23107_, _23212_);
  nor (_00504_, _00503_, _00502_);
  not (_00505_, _00504_);
  not (_00506_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor (_00507_, _23073_, _00506_);
  nor (_00508_, _23076_, _23360_);
  nor (_00510_, _00508_, _00507_);
  nor (_00511_, _23050_, _23210_);
  nor (_00512_, _23067_, _23217_);
  nor (_00513_, _00512_, _00511_);
  nand (_00514_, _00513_, _00510_);
  nor (_00515_, _00514_, _00505_);
  nor (_00516_, _00515_, _24824_);
  nor (_00517_, _00516_, _00501_);
  nor (_00518_, _00517_, _24820_);
  nor (_00519_, _00518_, _00499_);
  not (_00520_, _21344_);
  nor (_00521_, _00033_, _00123_);
  nor (_00522_, _00521_, _00126_);
  nor (_00523_, _00522_, _21202_);
  nor (_00524_, _00523_, _00520_);
  nor (_00525_, _00524_, _00023_);
  nor (_00526_, _00525_, _00122_);
  nor (_00527_, _00526_, _00354_);
  nor (_00528_, _24809_, _23229_);
  nor (_00529_, _00528_, _00527_);
  nand (_00531_, _00529_, _00519_);
  nand (_00532_, _00531_, _24743_);
  not (_00533_, _00532_);
  not (_00534_, _00075_);
  nand (_00535_, _24818_, _24815_);
  nor (_00536_, _00535_, _00002_);
  not (_00537_, _00078_);
  nor (_00538_, _00080_, _00537_);
  nand (_00539_, _00538_, _00091_);
  nand (_00540_, _00092_, _00081_);
  nor (_00541_, _00099_, _00540_);
  nand (_00542_, _00541_, _24915_);
  nor (_00543_, _00542_, _00539_);
  nor (_00544_, _00543_, _00076_);
  nand (_00545_, _00544_, _00536_);
  nor (_00546_, _00146_, _00111_);
  nor (_00547_, _00137_, _00112_);
  nor (_00548_, _00547_, _00546_);
  nor (_00549_, _00548_, _21202_);
  nor (_00550_, _00549_, _21206_);
  nor (_00551_, _00550_, _00023_);
  nor (_00552_, _00551_, _00107_);
  nor (_00553_, _00552_, _00004_);
  nor (_00554_, _00553_, _00002_);
  nand (_00555_, _00554_, _00545_);
  nor (_00556_, _00555_, _00534_);
  not (_00557_, _24743_);
  nand (_00558_, _00557_, _00556_);
  nor (_00559_, _00317_, _00558_);
  nor (_00560_, _00559_, _00533_);
  not (_00561_, _00560_);
  nor (_00562_, _00561_, _21353_);
  nand (_00563_, _00561_, _21353_);
  not (_00564_, _00563_);
  nor (_00565_, _00564_, _00562_);
  nand (_00566_, _00565_, _00469_);
  not (_00567_, _21322_);
  nor (_00568_, _24915_, ABINPUT[3]);
  not (_00569_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_00570_, _24948_, _00569_);
  not (_00572_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_00573_, _24925_, _00572_);
  nor (_00574_, _00573_, _00570_);
  not (_00575_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_00576_, _24931_, _00575_);
  not (_00577_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_00578_, _24934_, _00577_);
  nor (_00579_, _00578_, _00576_);
  nand (_00580_, _00579_, _00574_);
  nand (_00581_, _24943_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  not (_00582_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_00583_, _24921_, _00582_);
  not (_00584_, _00583_);
  nand (_00585_, _00584_, _00581_);
  not (_00586_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  nor (_00587_, _24952_, _00586_);
  nand (_00588_, _24955_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  not (_00589_, _00588_);
  nor (_00590_, _00589_, _00587_);
  not (_00591_, _00590_);
  nor (_00592_, _00591_, _00585_);
  nand (_00593_, _00592_, _24915_);
  nor (_00594_, _00593_, _00580_);
  nor (_00595_, _00594_, _00568_);
  nand (_00596_, _00595_, _00536_);
  not (_00597_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_00598_, _23044_, _00597_);
  not (_00599_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_00600_, _23058_, _00599_);
  not (_00601_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_00602_, _23107_, _00601_);
  nor (_00603_, _00602_, _00600_);
  not (_00604_, _00603_);
  not (_00605_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nor (_00606_, _23073_, _00605_);
  not (_00607_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_00608_, _23067_, _00607_);
  nor (_00609_, _00608_, _00606_);
  nor (_00610_, _23076_, _23156_);
  not (_00611_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_00613_, _23050_, _00611_);
  nor (_00615_, _00613_, _00610_);
  nand (_00616_, _00615_, _00609_);
  nor (_00617_, _00616_, _00604_);
  nor (_00618_, _00617_, _24824_);
  nor (_00619_, _00618_, _00598_);
  not (_00620_, _00619_);
  nand (_00621_, _00620_, _00437_);
  nand (_00622_, _00621_, _00596_);
  nor (_00623_, _00031_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_00624_, _00623_, _00040_);
  nor (_00625_, _00624_, _21202_);
  nor (_00626_, _00625_, _21314_);
  nor (_00627_, _00626_, _00023_);
  nor (_00628_, _00627_, _00030_);
  not (_00629_, _00628_);
  nand (_00631_, _00629_, _00005_);
  nand (_00632_, _24808_, _23351_);
  nand (_00633_, _00632_, _00631_);
  nor (_00634_, _00633_, _00622_);
  nor (_00637_, _00634_, _00557_);
  nor (_00638_, _00455_, _24820_);
  nor (_00639_, _00638_, _00434_);
  nand (_00640_, _00639_, _00435_);
  nor (_00641_, _00640_, _00426_);
  nor (_00642_, _00558_, _00641_);
  nor (_00643_, _00642_, _00637_);
  nor (_00644_, _00643_, _00567_);
  not (_00645_, _00632_);
  nor (_00646_, _00622_, _00645_);
  nand (_00647_, _00646_, _00631_);
  nand (_00648_, _00647_, _24743_);
  nand (_00649_, _00157_, _00461_);
  nand (_00650_, _00649_, _00648_);
  nor (_00651_, _00650_, _21322_);
  nor (_00652_, _00651_, _00644_);
  not (_00653_, _21639_);
  nor (_00654_, _00319_, _00653_);
  nor (_00655_, _00556_, _21227_);
  nor (_00656_, _00156_, _21246_);
  nor (_00657_, _00656_, _00655_);
  nor (_00658_, _00657_, _21231_);
  not (_00659_, _00658_);
  nor (_00660_, _00247_, _21381_);
  nor (_00661_, _00660_, _00659_);
  not (_00662_, _00661_);
  nor (_00663_, _00662_, _00654_);
  nand (_00664_, _00663_, _00652_);
  nor (_00665_, _00664_, _00566_);
  nand (_00666_, _00665_, _00393_);
  nor (_20959_, _00666_, rst);
  nor (_20960_, _21623_, rst);
  nor (_20961_, _00244_, rst);
  nor (_00667_, _24689_, _21658_);
  nor (_00668_, _00667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  not (_00669_, _00667_);
  nor (_00670_, _00669_, _21626_);
  nor (_25231_, _00670_, _00668_);
  not (_00671_, _00531_);
  nor (_20963_, _00671_, rst);
  nor (_00672_, _23769_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  nor (_00673_, _23771_, _21586_);
  nor (_20965_, _00673_, _00672_);
  nor (_00674_, _24568_, _21599_);
  nor (_00675_, _00674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  not (_00676_, _00674_);
  nor (_00677_, _00676_, _21451_);
  nor (_20966_, _00677_, _00675_);
  nor (_00678_, _24568_, _21374_);
  nor (_00680_, _00678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  not (_00681_, _00678_);
  nor (_00682_, _00681_, _21474_);
  nor (_20967_, _00682_, _00680_);
  nor (_00683_, _23040_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_00684_, _00683_);
  nor (_00685_, _00684_, \oc8051_top_1.oc8051_decoder1.state [0]);
  nor (_00686_, _23302_, _23115_);
  not (_00687_, _00686_);
  nor (_00688_, _00687_, _23143_);
  nor (_00689_, _23375_, _23355_);
  not (_00690_, _00689_);
  nor (_00691_, _00690_, _23277_);
  not (_00692_, _00691_);
  nor (_00693_, _00692_, _23170_);
  nand (_00694_, _00693_, _00688_);
  nor (_00695_, _00692_, _23348_);
  not (_00696_, _00695_);
  not (_00697_, _23143_);
  nor (_00698_, _00697_, _23084_);
  not (_00699_, _00698_);
  nor (_00701_, _23400_, _23115_);
  not (_00702_, _00701_);
  nor (_00703_, _00702_, _00699_);
  not (_00704_, _23084_);
  nor (_00705_, _00697_, _00704_);
  not (_00706_, _00705_);
  nor (_00707_, _00706_, _00702_);
  nor (_00708_, _00707_, _00703_);
  nor (_00709_, _00708_, _00696_);
  nor (_00710_, _23225_, _23355_);
  not (_00711_, _00710_);
  nor (_00712_, _23245_, _23348_);
  not (_00713_, _00712_);
  nor (_00714_, _00713_, _00711_);
  nor (_00715_, _00687_, _00704_);
  nand (_00716_, _00715_, _00714_);
  nand (_00717_, _00716_, _23496_);
  nor (_00718_, _00717_, _00709_);
  nand (_00719_, _00718_, _00694_);
  nand (_00720_, _00719_, _00685_);
  nor (_00721_, _00683_, _23509_);
  nor (_00722_, _00721_, rst);
  nand (_25018_[0], _00722_, _00720_);
  nor (_00723_, _24689_, _21652_);
  nor (_00724_, _00723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  not (_00725_, _00723_);
  nor (_00726_, _00725_, _21474_);
  nor (_20968_, _00726_, _00724_);
  nor (_00727_, _24689_, _21631_);
  nor (_00728_, _00727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  not (_00730_, _00727_);
  nor (_00731_, _00730_, _21626_);
  nor (_20969_, _00731_, _00728_);
  nor (_00732_, _24689_, _21589_);
  nor (_00733_, _00732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  not (_00734_, _00732_);
  nor (_00736_, _00734_, _21474_);
  nor (_20970_, _00736_, _00733_);
  nor (_00737_, _21377_, _21246_);
  nand (_00738_, _00017_, _00737_);
  nor (_00739_, _00738_, _24903_);
  nand (_00740_, _00739_, _24859_);
  nor (_00741_, _00740_, ABINPUT[5]);
  not (_00742_, _00740_);
  nor (_00743_, _00742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nor (_20971_, _00743_, _00741_);
  nor (_00744_, _21697_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  nor (_00745_, _21699_, _21554_);
  nor (_20972_, _00745_, _00744_);
  nor (_00746_, _21810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  nor (_00747_, _21812_, _21504_);
  nor (_20973_, _00747_, _00746_);
  nor (_00748_, _00667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nor (_00749_, _00669_, _21586_);
  nor (_25229_, _00749_, _00748_);
  nor (_00750_, _21790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  nor (_00751_, _21792_, _21451_);
  nor (_20974_, _00751_, _00750_);
  nor (_00752_, _24674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  nor (_00753_, _24676_, _21626_);
  nor (_20975_, _00753_, _00752_);
  nor (_00754_, _24684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  nor (_00755_, _24686_, _21451_);
  nor (_20976_, _00755_, _00754_);
  nor (_00756_, _24702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_00757_, _24704_, _21504_);
  nor (_25063_, _00757_, _00756_);
  nor (_00759_, _22484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  nor (_00760_, _22486_, _21414_);
  nor (_20977_, _00760_, _00759_);
  nor (_00762_, _21790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  nor (_00763_, _21792_, _21504_);
  nor (_20978_, _00763_, _00762_);
  nor (_00764_, _24689_, _21374_);
  nor (_00765_, _00764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  not (_00766_, _00764_);
  nor (_00767_, _00766_, _21526_);
  nor (_20980_, _00767_, _00765_);
  nor (_00768_, _00764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nor (_00769_, _00766_, _21554_);
  nor (_20981_, _00769_, _00768_);
  nor (_00770_, _00764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nor (_00771_, _00766_, _21586_);
  nor (_20982_, _00771_, _00770_);
  nor (_00772_, _00740_, ABINPUT[9]);
  nor (_00773_, _00742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nor (_20983_, _00773_, _00772_);
  nor (_00774_, _00740_, ABINPUT[7]);
  nor (_00775_, _00742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nor (_20984_, _00775_, _00774_);
  nor (_00777_, _00667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nor (_00778_, _00669_, _21526_);
  nor (_25230_, _00778_, _00777_);
  nor (_00779_, _00667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nor (_00780_, _00669_, _21474_);
  nor (_20985_, _00780_, _00779_);
  nor (_00781_, _00667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nor (_00782_, _00669_, _21414_);
  nor (_20986_, _00782_, _00781_);
  nor (_00783_, _21810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  nor (_00784_, _21812_, _21626_);
  nor (_25206_, _00784_, _00783_);
  nor (_00785_, _00742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nor (_00786_, _00740_, ABINPUT[4]);
  nor (_20988_, _00786_, _00785_);
  nor (_00788_, _24689_, _21864_);
  nor (_00789_, _00788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  not (_00790_, _00788_);
  nor (_00791_, _00790_, _21504_);
  nor (_20989_, _00791_, _00789_);
  nor (_00793_, _24710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nor (_00794_, _24712_, _21474_);
  nor (_20990_, _00794_, _00793_);
  nor (_00795_, _24710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nor (_00796_, _24712_, _21414_);
  nor (_20991_, _00796_, _00795_);
  nor (_00797_, _24689_, _21599_);
  nor (_00798_, _00797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  not (_00799_, _00797_);
  nor (_00800_, _00799_, _21414_);
  nor (_20993_, _00800_, _00798_);
  nor (_00801_, _00797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nor (_00802_, _00799_, _21474_);
  nor (_20994_, _00802_, _00801_);
  nor (_00803_, _00732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nor (_00804_, _00734_, _21586_);
  nor (_20995_, _00804_, _00803_);
  nor (_00805_, _00797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nor (_00806_, _00799_, _21626_);
  nor (_20996_, _00806_, _00805_);
  nor (_00808_, _00732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nor (_00809_, _00734_, _21626_);
  nor (_25406_, _00809_, _00808_);
  nor (_00810_, _23774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  nor (_00811_, _23776_, _21474_);
  nor (_25390_, _00811_, _00810_);
  nor (_00812_, _24689_, _21558_);
  nor (_00813_, _00812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  not (_00814_, _00812_);
  nor (_00815_, _00814_, _21474_);
  nor (_20997_, _00815_, _00813_);
  nor (_00816_, _00812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nor (_00817_, _00814_, _21414_);
  nor (_20998_, _00817_, _00816_);
  nor (_00818_, _24689_, _21607_);
  nor (_00819_, _00818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  not (_00820_, _00818_);
  nor (_00821_, _00820_, _21626_);
  nor (_20999_, _00821_, _00819_);
  nor (_00822_, _00818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nor (_00824_, _00820_, _21526_);
  nor (_21000_, _00824_, _00822_);
  nor (_00825_, _23774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  nor (_00826_, _23776_, _21586_);
  nor (_21002_, _00826_, _00825_);
  nor (_00827_, _24689_, _21482_);
  nor (_00828_, _00827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  not (_00829_, _00827_);
  nor (_00830_, _00829_, _21414_);
  nor (_21003_, _00830_, _00828_);
  nor (_00831_, _00727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nor (_00832_, _00730_, _21474_);
  nor (_21004_, _00832_, _00831_);
  nor (_00833_, _00727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_00834_, _00730_, _21504_);
  nor (_21005_, _00834_, _00833_);
  nor (_00835_, _00727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nor (_00836_, _00730_, _21414_);
  nor (_21006_, _00836_, _00835_);
  nor (_00837_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_00839_, _24692_, _21554_);
  nor (_21007_, _00839_, _00837_);
  nor (_00840_, _00723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_00841_, _00725_, _21586_);
  nor (_21008_, _00841_, _00840_);
  nor (_00842_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nor (_00843_, _24692_, _21626_);
  nor (_21009_, _00843_, _00842_);
  nor (_00844_, _24684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  nor (_00845_, _24686_, _21474_);
  nor (_21010_, _00845_, _00844_);
  nor (_00847_, _24568_, _21658_);
  not (_00848_, _00847_);
  nand (_00849_, _00848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  nor (_00850_, _00848_, _00121_);
  not (_00851_, _00850_);
  nand (_21011_, _00851_, _00849_);
  nor (_00852_, _00678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  nor (_00853_, _00681_, _21586_);
  nor (_21012_, _00853_, _00852_);
  nor (_00855_, _24568_, _21821_);
  nor (_00856_, _00855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  not (_00857_, _00855_);
  nor (_00858_, _00857_, _21451_);
  nor (_21013_, _00858_, _00856_);
  nor (_00859_, _00674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  nor (_00860_, _00676_, _21414_);
  nor (_21014_, _00860_, _00859_);
  nor (_00861_, _23774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  nor (_00862_, _23776_, _21526_);
  nor (_25391_, _00862_, _00861_);
  nor (_00863_, _23774_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  nor (_00864_, _23776_, _21554_);
  nor (_21015_, _00864_, _00863_);
  nand (_00865_, _24663_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  nor (_00866_, _24663_, _00121_);
  not (_00867_, _00866_);
  nand (_25327_, _00867_, _00865_);
  nor (_00868_, _24568_, _21607_);
  nor (_00869_, _00868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  not (_00870_, _00868_);
  nor (_00871_, _00870_, _21554_);
  nor (_21016_, _00871_, _00869_);
  nor (_00872_, _22454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  nor (_00873_, _22456_, _21474_);
  nor (_21017_, _00873_, _00872_);
  nor (_00874_, _24206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  nor (_00875_, _24208_, _21526_);
  nor (_21020_, _00875_, _00874_);
  nor (_00876_, _24380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  nor (_00877_, _24382_, _21504_);
  nor (_21023_, _00877_, _00876_);
  nor (_00878_, _21790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  nor (_00879_, _21792_, _21526_);
  nor (_21024_, _00879_, _00878_);
  nor (_00880_, _21645_, _21530_);
  nor (_00881_, _00880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  not (_00882_, _00880_);
  nor (_00883_, _00882_, _21414_);
  nor (_21025_, _00883_, _00881_);
  nor (_00884_, _21790_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  nor (_00885_, _21792_, _21414_);
  nor (_21026_, _00885_, _00884_);
  nor (_00886_, _24601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  nor (_00887_, _24603_, _21414_);
  nor (_25341_, _00887_, _00886_);
  nor (_00888_, _24601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  nor (_00889_, _24603_, _21554_);
  nor (_25339_, _00889_, _00888_);
  nor (_00890_, _24206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  nor (_00891_, _24208_, _21554_);
  nor (_21028_, _00891_, _00890_);
  nor (_00892_, _24601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  nor (_00893_, _24603_, _21474_);
  nor (_25338_, _00893_, _00892_);
  nor (_00894_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  nor (_00895_, _22165_, _21526_);
  nor (_21034_, _00895_, _00894_);
  nor (_00896_, _21786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  nor (_00897_, _21788_, _21526_);
  nor (_21035_, _00897_, _00896_);
  nor (_00898_, _21786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  nor (_00899_, _21788_, _21414_);
  nor (_21037_, _00899_, _00898_);
  nor (_00900_, _24206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  nor (_00901_, _24208_, _21474_);
  nor (_21039_, _00901_, _00900_);
  nor (_00902_, _24206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  nor (_00903_, _24208_, _21586_);
  nor (_21041_, _00903_, _00902_);
  not (_00904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  not (_00905_, _21351_);
  nor (_00906_, _21320_, _21285_);
  not (_00907_, _00906_);
  nor (_00908_, _00907_, _00905_);
  not (_00909_, _00908_);
  nor (_00910_, _21308_, _24897_);
  not (_00911_, _24904_);
  nor (_00912_, _21186_, _21184_);
  not (_00913_, _00912_);
  nor (_00914_, _00913_, _21232_);
  not (_00915_, _00914_);
  nor (_00916_, _00915_, _21227_);
  not (_00917_, _00916_);
  nor (_00918_, _00917_, _00911_);
  nand (_00919_, _00918_, _00910_);
  nor (_00920_, _00919_, _00909_);
  nor (_00921_, _00920_, _00904_);
  nor (_00922_, _00008_, _00911_);
  not (_00923_, _00922_);
  nor (_00924_, _00010_, _21308_);
  not (_00925_, _00924_);
  nor (_00926_, _00925_, _24858_);
  not (_00927_, _00926_);
  nor (_00928_, _00927_, _00923_);
  not (_00929_, _00928_);
  not (_00930_, _00919_);
  nor (_00931_, _00909_, _21507_);
  nand (_00932_, _00931_, _00930_);
  nand (_00933_, _00932_, _00929_);
  nor (_00934_, _00933_, _00921_);
  nand (_00935_, _00928_, _24867_);
  nand (_00936_, _00935_, _23493_);
  nor (_21042_, _00936_, _00934_);
  nor (_00937_, _23545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  nor (_00938_, _23547_, _21586_);
  nor (_21043_, _00938_, _00937_);
  nor (_00939_, _24206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  nor (_00940_, _24208_, _21504_);
  nor (_21044_, _00940_, _00939_);
  not (_00941_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nor (_00942_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  not (_00943_, _00942_);
  nor (_00944_, _00943_, _00941_);
  not (_00945_, _00944_);
  nand (_00946_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  not (_00947_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  nand (_00948_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not (_00949_, _00948_);
  not (_00950_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  nor (_00952_, _00950_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  nor (_00953_, _00952_, _00949_);
  nor (_00954_, _00953_, _00947_);
  not (_00955_, _00954_);
  not (_00956_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  not (_00957_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  not (_00958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  not (_00959_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  not (_00960_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  not (_00961_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  not (_00962_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  not (_00963_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  not (_00964_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor (_00965_, _00964_, _00963_);
  nand (_00966_, _00965_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_00967_, _00966_, _00962_);
  not (_00968_, _00967_);
  nor (_00969_, _00968_, _00961_);
  not (_00970_, _00969_);
  nor (_00971_, _00970_, _00960_);
  nand (_00973_, _00971_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_00974_, _00973_, _00959_);
  nand (_00975_, _00974_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor (_00976_, _00975_, _00958_);
  nand (_00977_, _00976_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_00978_, _00977_, _00957_);
  nand (_00979_, _00978_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_00980_, _00979_, _00956_);
  nand (_00981_, _00980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  not (_00982_, _00981_);
  nand (_00983_, _00982_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor (_00984_, _00983_, _00955_);
  not (_00985_, _00984_);
  nor (_00986_, _00985_, _00946_);
  nor (_00987_, _00968_, _00955_);
  nand (_00988_, _00987_, _00961_);
  nand (_00989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nand (_00990_, _00942_, _00941_);
  nor (_00991_, _00990_, _00989_);
  nor (_00992_, _00987_, _00961_);
  nor (_00993_, _00992_, _00991_);
  nand (_00994_, _00993_, _00988_);
  nor (_00995_, _00994_, _00986_);
  not (_00996_, _00991_);
  nor (_00997_, _00996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nor (_00998_, _00997_, _00995_);
  not (_00999_, _24857_);
  nor (_01000_, _00999_, _21351_);
  not (_01001_, _01000_);
  nor (_01002_, _01001_, _00925_);
  not (_01003_, _01002_);
  nor (_01004_, _01003_, _00923_);
  nor (_01005_, _01004_, _00998_);
  not (_01006_, _01004_);
  nor (_01007_, _01006_, ABINPUT[7]);
  nor (_01009_, _01007_, _01005_);
  nand (_01010_, _00019_, _00905_);
  nor (_01011_, _01010_, _00925_);
  not (_01012_, _01011_);
  nor (_01013_, _01012_, _00923_);
  nor (_01014_, _01013_, _01009_);
  nand (_01015_, _01013_, _00961_);
  nand (_01016_, _01015_, _23493_);
  nor (_21045_, _01016_, _01014_);
  nor (_01017_, _00989_, _00945_);
  nand (_01018_, _01017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  not (_01020_, _01017_);
  nand (_01021_, _01020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand (_01022_, _01021_, _01018_);
  nor (_01023_, _24856_, _21285_);
  not (_01025_, _01023_);
  nor (_01026_, _01025_, _00905_);
  not (_01027_, _01026_);
  nor (_01028_, _01027_, _00925_);
  not (_01029_, _01028_);
  nor (_01030_, _01029_, _00923_);
  nor (_01031_, _01030_, _01022_);
  not (_01032_, _01030_);
  nor (_01033_, _01032_, ABINPUT[7]);
  nor (_01034_, _01033_, _01031_);
  nor (_01035_, _00909_, _00925_);
  not (_01036_, _01035_);
  nor (_01037_, _01036_, _00923_);
  nor (_01038_, _01037_, _01034_);
  not (_01039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  nand (_01040_, _01037_, _01039_);
  nand (_01041_, _01040_, _23493_);
  nor (_21046_, _01041_, _01038_);
  nor (_01042_, _01030_, _01020_);
  nor (_01043_, _01042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not (_01044_, _01042_);
  nor (_01045_, _01044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor (_01046_, _01045_, _01043_);
  nor (_01047_, _01046_, _01037_);
  nand (_01048_, _01037_, _00029_);
  nand (_01049_, _01048_, _23493_);
  nor (_21047_, _01049_, _01047_);
  nor (_01050_, _24206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  nor (_01051_, _24208_, _21451_);
  nor (_25388_, _01051_, _01050_);
  not (_01052_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  not (_01053_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_01054_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor (_01055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_01056_, _01055_, _01054_);
  not (_01057_, _01056_);
  nor (_01058_, _01057_, _01053_);
  not (_01059_, _01055_);
  not (_01060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_01061_, _01060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_01062_, _01061_, _01054_);
  nor (_01063_, _01062_, _01059_);
  nor (_01064_, _01053_, _01060_);
  nand (_01065_, _01064_, _01059_);
  not (_01066_, _01065_);
  nor (_01067_, _01066_, _01063_);
  nor (_01068_, _01067_, _01058_);
  nor (_01069_, _01059_, _01054_);
  not (_01070_, _01069_);
  nor (_01071_, _01070_, _00950_);
  not (_01072_, _01058_);
  not (_01073_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_01074_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01073_);
  not (_01075_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_01076_, _01075_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nand (_01077_, _01076_, _01074_);
  nor (_01078_, _01077_, _01072_);
  nor (_01079_, _01078_, _01071_);
  not (_01080_, _01079_);
  nor (_01081_, _01080_, _01068_);
  nor (_01083_, _01081_, _01052_);
  nor (_01084_, _01083_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  nor (_01085_, _01052_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nand (_01086_, _01085_, _01080_);
  nand (_01087_, _01086_, _23493_);
  nor (_21048_, _01087_, _01084_);
  nor (_01088_, _24206_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  nor (_01089_, _24208_, _21414_);
  nor (_21049_, _01089_, _01088_);
  not (_01090_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor (_01091_, _01001_, _00919_);
  nor (_01092_, _01091_, _01090_);
  nor (_01093_, _01001_, _21507_);
  nand (_01094_, _01093_, _00930_);
  nand (_01095_, _01094_, _00929_);
  nor (_01096_, _01095_, _01092_);
  nand (_01097_, _00928_, _24900_);
  nand (_01098_, _01097_, _23493_);
  nor (_21050_, _01098_, _01096_);
  nor (_01099_, _23348_, _23043_);
  not (_01100_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nand (_01101_, _23043_, _01100_);
  nand (_01102_, _01101_, _23493_);
  nor (_25019_[0], _01102_, _01099_);
  nand (_01103_, _01017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand (_01104_, _01020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nand (_01105_, _01104_, _01103_);
  nor (_01106_, _01105_, _01030_);
  nor (_01107_, _01032_, ABINPUT[8]);
  nor (_01108_, _01107_, _01106_);
  nor (_01110_, _01108_, _01037_);
  not (_01111_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nand (_01112_, _01037_, _01111_);
  nand (_01113_, _01112_, _23493_);
  nor (_21051_, _01113_, _01110_);
  nor (_01114_, _01042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_01115_, _01044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_01116_, _01115_, _01114_);
  nor (_01117_, _01116_, _01037_);
  nand (_01118_, _01037_, _00006_);
  nand (_01119_, _01118_, _23493_);
  nor (_21052_, _01119_, _01117_);
  nor (_01120_, _21786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  nor (_01121_, _21788_, _21586_);
  nor (_21054_, _01121_, _01120_);
  nor (_01122_, _22263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  nor (_01123_, _22265_, _21526_);
  nor (_21055_, _01123_, _01122_);
  not (_01124_, _24901_);
  nor (_01125_, _01124_, _00007_);
  not (_01127_, _01125_);
  nor (_01128_, _00925_, _00020_);
  not (_01129_, _01128_);
  nor (_01130_, _01129_, _01127_);
  not (_01131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_01132_, _01131_, _00950_);
  nand (_01133_, _01132_, _01055_);
  not (_01134_, _01133_);
  nand (_01135_, _01059_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  nor (_01136_, _01135_, _01131_);
  not (_01137_, _01136_);
  nor (_01138_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_01139_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nand (_01140_, _01139_, _01138_);
  nor (_01141_, _01140_, _01137_);
  nor (_01142_, _01141_, _01134_);
  not (_01143_, _01142_);
  nand (_01144_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nand (_01145_, _01142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nand (_01146_, _01145_, _01144_);
  nor (_01147_, _01146_, _01130_);
  nor (_01148_, _01059_, _00106_);
  nor (_01149_, _01055_, _00114_);
  nor (_01150_, _01149_, _01148_);
  nand (_01151_, _01150_, _01130_);
  nand (_01152_, _01151_, _23493_);
  nor (_21056_, _01152_, _01147_);
  nor (_01153_, _23779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  nor (_01154_, _23782_, _21526_);
  nor (_21057_, _01154_, _01153_);
  nor (_01156_, _23779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  nor (_01157_, _23782_, _21554_);
  nor (_21058_, _01157_, _01156_);
  nor (_01158_, _23779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  nor (_01159_, _23782_, _21474_);
  nor (_21059_, _01159_, _01158_);
  nor (_01160_, _23245_, _23043_);
  not (_01161_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nand (_01162_, _23043_, _01161_);
  nand (_01163_, _01162_, _23493_);
  nor (_25019_[1], _01163_, _01160_);
  nor (_01164_, _21786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  nor (_01165_, _21788_, _21474_);
  nor (_21060_, _01165_, _01164_);
  nor (_01166_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand (_01167_, _23553_, _23103_);
  nand (_01168_, _01167_, _23493_);
  nor (_21062_, _01168_, _01166_);
  nor (_01169_, _22512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  nor (_01170_, _22514_, _21554_);
  nor (_21063_, _01170_, _01169_);
  not (_01171_, _23486_);
  not (_01172_, _23455_);
  nand (_01173_, _24398_, _23088_);
  nand (_01174_, _01173_, _01172_);
  nor (_01175_, _01174_, _01171_);
  nand (_01176_, _01175_, _23507_);
  nand (_01177_, _01176_, _23491_);
  nand (_01178_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_01179_, _01178_, _23519_);
  nand (_01181_, _01179_, _23493_);
  nand (_25021_[1], _01181_, _01177_);
  nor (_01182_, _22018_, _21427_);
  not (_01183_, _01182_);
  nor (_01184_, _01183_, _21689_);
  nor (_01185_, _01184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  not (_01186_, _01184_);
  nor (_01187_, _01186_, _21414_);
  nor (_21065_, _01187_, _01185_);
  nor (_01188_, _23779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  nor (_01189_, _23782_, _21414_);
  nor (_25387_, _01189_, _01188_);
  nor (_01190_, _23779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  nor (_01191_, _23782_, _21504_);
  nor (_21067_, _01191_, _01190_);
  nor (_01192_, _21782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  nor (_01193_, _21784_, _21586_);
  nor (_25217_, _01193_, _01192_);
  nor (_01194_, _01183_, _21425_);
  nor (_01195_, _01194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  not (_01196_, _01194_);
  nor (_01197_, _01196_, _21586_);
  nor (_21069_, _01197_, _01195_);
  nor (_01198_, _01183_, _21589_);
  nor (_01199_, _01198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  not (_01200_, _01198_);
  nor (_01201_, _01200_, _21626_);
  nor (_21070_, _01201_, _01199_);
  nand (_01202_, _01017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nand (_01203_, _01020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nand (_01204_, _01203_, _01202_);
  nor (_01205_, _01204_, _01030_);
  nor (_01206_, _01032_, ABINPUT[6]);
  nor (_01207_, _01206_, _01205_);
  nor (_01208_, _01207_, _01037_);
  not (_01209_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  nand (_01210_, _01037_, _01209_);
  nand (_01211_, _01210_, _23493_);
  nor (_21071_, _01211_, _01208_);
  nand (_01212_, _01017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_01213_, _01020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_01214_, _01213_, _01212_);
  nor (_01215_, _01214_, _01030_);
  nor (_01216_, _01032_, ABINPUT[3]);
  nor (_01217_, _01216_, _01215_);
  nor (_01218_, _01217_, _01037_);
  not (_01219_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_01220_, _01037_, _01219_);
  nand (_01222_, _01220_, _23493_);
  nor (_21072_, _01222_, _01218_);
  nor (_01223_, _23779_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  nor (_01224_, _23782_, _21451_);
  nor (_21073_, _01224_, _01223_);
  nor (_01226_, _01042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_01227_, _01044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nor (_01228_, _01227_, _01226_);
  nor (_01229_, _01228_, _01037_);
  nand (_01230_, _01037_, _24867_);
  nand (_01231_, _01230_, _23493_);
  nor (_21074_, _01231_, _01229_);
  nor (_01233_, _01183_, _21607_);
  nor (_01234_, _01233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  not (_01235_, _01233_);
  nor (_01236_, _01235_, _21504_);
  nor (_21075_, _01236_, _01234_);
  nor (_01237_, _22526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  nor (_01238_, _22528_, _21504_);
  nor (_21076_, _01238_, _01237_);
  nor (_01239_, _01013_, _01004_);
  not (_01240_, _01239_);
  nor (_01241_, _00944_, _01209_);
  nand (_01242_, _01241_, _00984_);
  nor (_01243_, _00966_, _00955_);
  nor (_01244_, _01243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_01245_, _01244_, _00987_);
  nor (_01246_, _01245_, _00991_);
  nand (_01247_, _01246_, _01242_);
  nand (_01248_, _00991_, _01209_);
  nand (_01249_, _01248_, _01247_);
  nor (_01250_, _01249_, _01240_);
  nand (_01251_, _01013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nand (_01252_, _01004_, ABINPUT[6]);
  nand (_01253_, _01252_, _01251_);
  nor (_01254_, _01253_, _01250_);
  nor (_21077_, _01254_, rst);
  nand (_01255_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nor (_01256_, _01255_, _00985_);
  not (_01257_, _01243_);
  not (_01258_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand (_01259_, _00965_, _00954_);
  nand (_01260_, _01259_, _01258_);
  nand (_01261_, _01260_, _01257_);
  nand (_01262_, _01261_, _00996_);
  nor (_01263_, _01262_, _01256_);
  not (_01264_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand (_01265_, _00991_, _01264_);
  nand (_01266_, _01265_, _01006_);
  nor (_01267_, _01266_, _01263_);
  nor (_01268_, _01013_, ABINPUT[5]);
  nor (_01269_, _01268_, _01239_);
  nor (_01271_, _01269_, _01267_);
  nand (_01272_, _01013_, _01258_);
  nand (_01273_, _01272_, _23493_);
  nor (_21078_, _01273_, _01271_);
  nor (_01274_, _22263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  nor (_01275_, _22265_, _21474_);
  nor (_21079_, _01275_, _01274_);
  nand (_01276_, _23504_, _23450_);
  nor (_01277_, _23452_, _23359_);
  nor (_01278_, _01277_, _23464_);
  nor (_01279_, _01278_, _01276_);
  nand (_01280_, _01279_, _23448_);
  nand (_01281_, _01280_, _23491_);
  nand (_01282_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_01283_, _01282_, _23521_);
  nand (_01284_, _01283_, _23493_);
  nand (_25021_[0], _01284_, _01281_);
  nor (_01285_, _23375_, _23043_);
  not (_01286_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nand (_01287_, _23043_, _01286_);
  nand (_01288_, _01287_, _23493_);
  nor (_25019_[2], _01288_, _01285_);
  nor (_01289_, _23857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  nor (_01290_, _23859_, _21414_);
  nor (_21080_, _01290_, _01289_);
  nor (_01291_, _23857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  nor (_01292_, _23859_, _21526_);
  nor (_21081_, _01292_, _01291_);
  nor (_01293_, _22263_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  nor (_01294_, _22265_, _21586_);
  nor (_21082_, _01294_, _01293_);
  nor (_01295_, _23857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  nor (_01296_, _23859_, _21554_);
  nor (_21083_, _01296_, _01295_);
  not (_01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_01298_, _00944_, _01297_);
  nand (_01299_, _01298_, _00954_);
  nor (_01300_, _01299_, _00983_);
  nor (_01301_, _00977_, _00955_);
  not (_01302_, _01301_);
  nand (_01303_, _01302_, _00957_);
  nand (_01304_, _01301_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand (_01305_, _01304_, _01303_);
  nand (_01306_, _01305_, _00996_);
  nor (_01307_, _01306_, _01300_);
  nand (_01308_, _00991_, _01297_);
  nand (_01309_, _01308_, _01239_);
  nor (_01310_, _01309_, _01307_);
  nand (_01311_, _01013_, ABINPUT[6]);
  nand (_01312_, _01004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand (_01314_, _01312_, _01311_);
  nor (_01315_, _01314_, _01310_);
  nor (_21084_, _01315_, rst);
  nor (_01316_, _01027_, _00919_);
  nor (_01317_, _01316_, _00947_);
  nor (_01318_, _01027_, _21507_);
  nand (_01319_, _01318_, _00930_);
  nand (_01320_, _01319_, _00929_);
  nor (_01321_, _01320_, _01317_);
  nand (_01322_, _00928_, _00121_);
  nand (_01323_, _01322_, _23493_);
  nor (_21085_, _01323_, _01321_);
  nor (_01324_, _01083_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nor (_01325_, _01052_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  nand (_01326_, _01325_, _01080_);
  nand (_01327_, _01326_, _23493_);
  nor (_21086_, _01327_, _01324_);
  nand (_01328_, _23490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  not (_01329_, _01328_);
  not (_01330_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  nor (_01331_, _23153_, _01330_);
  nor (_01333_, _23050_, _00290_);
  nor (_01334_, _23067_, _00285_);
  nor (_01335_, _01334_, _01333_);
  not (_01336_, _01335_);
  not (_01337_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor (_01338_, _23073_, _01337_);
  nor (_01340_, _23107_, _00283_);
  nor (_01341_, _01340_, _01338_);
  nor (_01342_, _23076_, _00292_);
  nor (_01344_, _23058_, _24154_);
  nor (_01345_, _01344_, _01342_);
  nand (_01346_, _01345_, _01341_);
  nor (_01347_, _01346_, _01336_);
  nor (_01348_, _01347_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_01350_, _01348_, _01331_);
  nor (_01351_, _01350_, _23490_);
  nor (_01352_, _01351_, _01329_);
  nor (_21087_, _01352_, rst);
  nor (_01353_, _23355_, _23043_);
  not (_01354_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nand (_01355_, _23043_, _01354_);
  nand (_01356_, _01355_, _23493_);
  nor (_25019_[3], _01356_, _01353_);
  nor (_01357_, _22838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  nor (_01358_, _22840_, _21526_);
  nor (_21089_, _01358_, _01357_);
  nor (_01359_, _22272_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  nor (_01360_, _22274_, _21504_);
  nor (_25159_, _01360_, _01359_);
  nor (_01361_, _22272_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  nor (_01362_, _22274_, _21414_);
  nor (_21093_, _01362_, _01361_);
  nor (_01363_, _21816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  nor (_01364_, _21818_, _21504_);
  nor (_21096_, _01364_, _01363_);
  nor (_01365_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  nand (_01366_, _23553_, _00605_);
  nand (_01367_, _01366_, _23493_);
  nor (_21099_, _01367_, _01365_);
  nor (_01369_, _23857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  nor (_01370_, _23859_, _21626_);
  nor (_21100_, _01370_, _01369_);
  nor (_01371_, _23857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  nor (_01372_, _23859_, _21504_);
  nor (_21101_, _01372_, _01371_);
  nor (_01373_, _23857_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  nor (_01374_, _23859_, _21451_);
  nor (_21102_, _01374_, _01373_);
  nor (_01375_, _21645_, _21599_);
  nor (_01376_, _01375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  not (_01377_, _01375_);
  nor (_01378_, _01377_, _21586_);
  nor (_21103_, _01378_, _01376_);
  nor (_01379_, _00704_, _23043_);
  not (_01380_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nand (_01381_, _23043_, _01380_);
  nand (_01382_, _01381_, _23493_);
  nor (_25019_[4], _01382_, _01379_);
  nor (_01383_, _21658_, _21645_);
  nor (_01384_, _01383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  not (_01385_, _01383_);
  nor (_01386_, _01385_, _21586_);
  nor (_25271_, _01386_, _01384_);
  nor (_01387_, _24159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  nor (_01388_, _24161_, _21526_);
  nor (_21104_, _01388_, _01387_);
  nor (_01389_, _22272_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  nor (_01390_, _22274_, _21554_);
  nor (_21105_, _01390_, _01389_);
  nor (_01391_, _24159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  nor (_01392_, _24161_, _21414_);
  nor (_21106_, _01392_, _01391_);
  nor (_01393_, _21904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  nor (_01394_, _21906_, _21626_);
  nor (_21107_, _01394_, _01393_);
  nor (_01395_, _23143_, _23043_);
  not (_01396_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nand (_01397_, _23043_, _01396_);
  nand (_01398_, _01397_, _23493_);
  nor (_25019_[5], _01398_, _01395_);
  nor (_01400_, _22557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  nor (_01401_, _22559_, _21554_);
  nor (_21108_, _01401_, _01400_);
  nor (_01402_, _24159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  nor (_01403_, _24161_, _21451_);
  nor (_21109_, _01403_, _01402_);
  nor (_01404_, _24159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  nor (_01405_, _24161_, _21626_);
  nor (_21111_, _01405_, _01404_);
  nor (_01406_, _24159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  nor (_01407_, _24161_, _21504_);
  nor (_21112_, _01407_, _01406_);
  nor (_01408_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  nor (_01409_, _22221_, _21414_);
  nor (_21113_, _01409_, _01408_);
  nor (_01410_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  nor (_01411_, _22563_, _21626_);
  nor (_25078_, _01411_, _01410_);
  nor (_01412_, _21842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  nor (_01413_, _21844_, _21451_);
  nor (_21114_, _01413_, _01412_);
  nor (_01414_, _21822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  nor (_01415_, _21824_, _21474_);
  nor (_21115_, _01415_, _01414_);
  not (_01416_, _00666_);
  not (_01417_, _00227_);
  nand (_01418_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7]);
  nand (_01419_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7]);
  nand (_01420_, _01419_, _01418_);
  nand (_01422_, _01420_, _01417_);
  nand (_01423_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7]);
  nand (_01424_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  nand (_01425_, _01424_, _01423_);
  nand (_01426_, _01425_, _00227_);
  nand (_01427_, _01426_, _01422_);
  nand (_01428_, _01427_, _00560_);
  nand (_01429_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7]);
  nand (_01430_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  nand (_01431_, _01430_, _01429_);
  nand (_01432_, _01431_, _01417_);
  nand (_01433_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  nand (_01434_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  nand (_01435_, _01434_, _01433_);
  nand (_01436_, _01435_, _00227_);
  nand (_01437_, _01436_, _01432_);
  nand (_01438_, _01437_, _00561_);
  nand (_01439_, _01438_, _01428_);
  nand (_01441_, _01439_, _00466_);
  nor (_01442_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  nor (_01444_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7]);
  nor (_01445_, _01444_, _01442_);
  nand (_01446_, _01445_, _01417_);
  nor (_01447_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7]);
  nor (_01448_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7]);
  nor (_01449_, _01448_, _01447_);
  nand (_01450_, _01449_, _00227_);
  nand (_01451_, _01450_, _01446_);
  nand (_01452_, _01451_, _00560_);
  nor (_01453_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7]);
  nor (_01455_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7]);
  nor (_01456_, _01455_, _01453_);
  nand (_01457_, _01456_, _01417_);
  nor (_01459_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7]);
  nor (_01460_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7]);
  nor (_01461_, _01460_, _01459_);
  nand (_01462_, _01461_, _00227_);
  nand (_01463_, _01462_, _01457_);
  nand (_01464_, _01463_, _00561_);
  nand (_01465_, _01464_, _01452_);
  nand (_01466_, _01465_, _00465_);
  nand (_01467_, _01466_, _01441_);
  nand (_01468_, _01467_, _00247_);
  nand (_01469_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7]);
  nand (_01470_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7]);
  nand (_01471_, _01470_, _01469_);
  nand (_01473_, _01471_, _01417_);
  nand (_01475_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7]);
  nand (_01476_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  nand (_01477_, _01476_, _01475_);
  nand (_01479_, _01477_, _00227_);
  nand (_01480_, _01479_, _01473_);
  nand (_01481_, _01480_, _00560_);
  nand (_01482_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7]);
  nand (_01483_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7]);
  nand (_01484_, _01483_, _01482_);
  nand (_01485_, _01484_, _01417_);
  nand (_01486_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7]);
  nand (_01487_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  nand (_01488_, _01487_, _01486_);
  nand (_01489_, _01488_, _00227_);
  nand (_01490_, _01489_, _01485_);
  nand (_01491_, _01490_, _00561_);
  nand (_01492_, _01491_, _01481_);
  nand (_01493_, _01492_, _00466_);
  nor (_01494_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  nor (_01495_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7]);
  nor (_01496_, _01495_, _01494_);
  nand (_01498_, _01496_, _00227_);
  nand (_01499_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  nand (_01500_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  nand (_01501_, _01500_, _01499_);
  nand (_01502_, _01501_, _01417_);
  nand (_01503_, _01502_, _01498_);
  nand (_01504_, _01503_, _00560_);
  nor (_01505_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  nor (_01506_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7]);
  nor (_01508_, _01506_, _01505_);
  nand (_01509_, _01508_, _00227_);
  nand (_01510_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  nand (_01513_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  nand (_01514_, _01513_, _01510_);
  nand (_01515_, _01514_, _01417_);
  nand (_01516_, _01515_, _01509_);
  nand (_01517_, _01516_, _00561_);
  nand (_01518_, _01517_, _01504_);
  nand (_01519_, _01518_, _00465_);
  nand (_01520_, _01519_, _01493_);
  nand (_01521_, _01520_, _00248_);
  nand (_01522_, _01521_, _01468_);
  nand (_01523_, _01522_, _00320_);
  nand (_01524_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7]);
  nand (_01525_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nand (_01526_, _01525_, _01524_);
  nand (_01527_, _01526_, _01417_);
  nand (_01528_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nand (_01529_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nand (_01530_, _01529_, _01528_);
  nand (_01531_, _01530_, _00227_);
  nand (_01532_, _01531_, _01527_);
  nand (_01533_, _01532_, _00560_);
  nand (_01534_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7]);
  nand (_01535_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7]);
  nand (_01536_, _01535_, _01534_);
  nand (_01537_, _01536_, _01417_);
  nand (_01538_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7]);
  nand (_01539_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nand (_01540_, _01539_, _01538_);
  nand (_01541_, _01540_, _00227_);
  nand (_01543_, _01541_, _01537_);
  nand (_01545_, _01543_, _00561_);
  nand (_01546_, _01545_, _01533_);
  nand (_01547_, _01546_, _00466_);
  nor (_01548_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nor (_01549_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_01550_, _01549_, _01548_);
  nand (_01551_, _01550_, _00227_);
  nand (_01552_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nand (_01553_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7]);
  nand (_01554_, _01553_, _01552_);
  nand (_01555_, _01554_, _01417_);
  nand (_01556_, _01555_, _01551_);
  nand (_01557_, _01556_, _00560_);
  nor (_01558_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7]);
  nor (_01559_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_01560_, _01559_, _01558_);
  nand (_01561_, _01560_, _00227_);
  nand (_01562_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nand (_01563_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7]);
  nand (_01564_, _01563_, _01562_);
  nand (_01565_, _01564_, _01417_);
  nand (_01566_, _01565_, _01561_);
  nand (_01568_, _01566_, _00561_);
  nand (_01570_, _01568_, _01557_);
  nand (_01571_, _01570_, _00465_);
  nand (_01573_, _01571_, _01547_);
  nand (_01574_, _01573_, _00248_);
  nand (_01575_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  nand (_01576_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  nand (_01577_, _01576_, _01575_);
  nand (_01578_, _01577_, _01417_);
  nand (_01580_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7]);
  nand (_01581_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  nand (_01582_, _01581_, _01580_);
  nand (_01583_, _01582_, _00227_);
  nand (_01584_, _01583_, _01578_);
  nand (_01585_, _01584_, _00560_);
  nand (_01586_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  nand (_01587_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  nand (_01588_, _01587_, _01586_);
  nand (_01589_, _01588_, _01417_);
  nand (_01590_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  nand (_01591_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  nand (_01592_, _01591_, _01590_);
  nand (_01593_, _01592_, _00227_);
  nand (_01594_, _01593_, _01589_);
  nand (_01596_, _01594_, _00561_);
  nand (_01597_, _01596_, _01585_);
  nand (_01598_, _01597_, _00466_);
  nor (_01599_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  nor (_01601_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  nor (_01602_, _01601_, _01599_);
  nand (_01603_, _01602_, _01417_);
  nor (_01604_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  nor (_01605_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7]);
  nor (_01606_, _01605_, _01604_);
  nand (_01607_, _01606_, _00227_);
  nand (_01608_, _01607_, _01603_);
  nand (_01609_, _01608_, _00560_);
  nor (_01610_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7]);
  nor (_01611_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  nor (_01612_, _01611_, _01610_);
  nand (_01613_, _01612_, _01417_);
  nor (_01614_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  nor (_01615_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7]);
  nor (_01616_, _01615_, _01614_);
  nand (_01617_, _01616_, _00227_);
  nand (_01618_, _01617_, _01613_);
  nand (_01619_, _01618_, _00561_);
  nand (_01620_, _01619_, _01609_);
  nand (_01622_, _01620_, _00465_);
  nand (_01623_, _01622_, _01598_);
  nand (_01624_, _01623_, _00247_);
  nand (_01625_, _01624_, _01574_);
  nand (_01626_, _01625_, _00319_);
  nand (_01627_, _01626_, _01523_);
  nor (_01628_, _01627_, _00386_);
  not (_01629_, _00386_);
  nand (_01630_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7]);
  nand (_01631_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7]);
  nand (_01632_, _01631_, _01630_);
  nand (_01633_, _01632_, _01417_);
  nand (_01634_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7]);
  nand (_01635_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7]);
  nand (_01636_, _01635_, _01634_);
  nand (_01637_, _01636_, _00227_);
  nand (_01638_, _01637_, _01633_);
  nand (_01639_, _01638_, _00560_);
  nand (_01640_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7]);
  nand (_01641_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7]);
  nand (_01642_, _01641_, _01640_);
  nand (_01643_, _01642_, _01417_);
  nand (_01644_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7]);
  nand (_01645_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7]);
  nand (_01646_, _01645_, _01644_);
  nand (_01647_, _01646_, _00227_);
  nand (_01649_, _01647_, _01643_);
  nand (_01650_, _01649_, _00561_);
  nand (_01651_, _01650_, _01639_);
  nand (_01652_, _01651_, _00466_);
  nor (_01653_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7]);
  nor (_01654_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7]);
  nor (_01655_, _01654_, _01653_);
  nand (_01656_, _01655_, _00227_);
  nand (_01657_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7]);
  nand (_01658_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7]);
  nand (_01659_, _01658_, _01657_);
  nand (_01660_, _01659_, _01417_);
  nand (_01661_, _01660_, _01656_);
  nand (_01662_, _01661_, _00560_);
  nor (_01663_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  nor (_01664_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7]);
  nor (_01665_, _01664_, _01663_);
  nand (_01666_, _01665_, _00227_);
  nand (_01667_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  nand (_01668_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7]);
  nand (_01669_, _01668_, _01667_);
  nand (_01670_, _01669_, _01417_);
  nand (_01671_, _01670_, _01666_);
  nand (_01672_, _01671_, _00561_);
  nand (_01674_, _01672_, _01662_);
  nand (_01675_, _01674_, _00465_);
  nand (_01676_, _01675_, _01652_);
  nand (_01677_, _01676_, _00248_);
  nand (_01678_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  nand (_01679_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7]);
  nand (_01680_, _01679_, _01678_);
  nand (_01681_, _01680_, _01417_);
  nand (_01682_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  nand (_01683_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  nand (_01685_, _01683_, _01682_);
  nand (_01686_, _01685_, _00227_);
  nand (_01687_, _01686_, _01681_);
  nand (_01688_, _01687_, _00560_);
  nand (_01689_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7]);
  nand (_01690_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7]);
  nand (_01691_, _01690_, _01689_);
  nand (_01692_, _01691_, _01417_);
  nand (_01693_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  nand (_01694_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7]);
  nand (_01696_, _01694_, _01693_);
  nand (_01697_, _01696_, _00227_);
  nand (_01698_, _01697_, _01692_);
  nand (_01699_, _01698_, _00561_);
  nand (_01700_, _01699_, _01688_);
  nand (_01702_, _01700_, _00466_);
  nor (_01703_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  nor (_01704_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7]);
  nor (_01705_, _01704_, _01703_);
  nand (_01706_, _01705_, _01417_);
  nor (_01707_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  nor (_01708_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  nor (_01709_, _01708_, _01707_);
  nand (_01710_, _01709_, _00227_);
  nand (_01711_, _01710_, _01706_);
  nand (_01712_, _01711_, _00560_);
  nor (_01713_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  nor (_01714_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  nor (_01715_, _01714_, _01713_);
  nand (_01716_, _01715_, _01417_);
  nor (_01718_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  nor (_01719_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  nor (_01720_, _01719_, _01718_);
  nand (_01721_, _01720_, _00227_);
  nand (_01722_, _01721_, _01716_);
  nand (_01723_, _01722_, _00561_);
  nand (_01724_, _01723_, _01712_);
  nand (_01725_, _01724_, _00465_);
  nand (_01726_, _01725_, _01702_);
  nand (_01727_, _01726_, _00247_);
  nand (_01728_, _01727_, _01677_);
  nand (_01729_, _01728_, _00320_);
  nor (_01731_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  nor (_01732_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7]);
  nor (_01733_, _01732_, _01731_);
  nand (_01734_, _01733_, _01417_);
  nor (_01736_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7]);
  nor (_01737_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7]);
  nor (_01738_, _01737_, _01736_);
  nand (_01739_, _01738_, _00227_);
  nand (_01740_, _01739_, _01734_);
  nand (_01741_, _01740_, _00561_);
  nor (_01742_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7]);
  nor (_01743_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7]);
  nor (_01745_, _01743_, _01742_);
  nand (_01746_, _01745_, _01417_);
  nor (_01747_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7]);
  nor (_01748_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7]);
  nor (_01749_, _01748_, _01747_);
  nand (_01750_, _01749_, _00227_);
  nand (_01752_, _01750_, _01746_);
  nand (_01753_, _01752_, _00560_);
  nand (_01754_, _01753_, _01741_);
  nand (_01755_, _01754_, _00465_);
  nand (_01756_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7]);
  nand (_01757_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7]);
  nand (_01758_, _01757_, _01756_);
  nand (_01759_, _01758_, _01417_);
  nand (_01760_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7]);
  nand (_01762_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7]);
  nand (_01764_, _01762_, _01760_);
  nand (_01765_, _01764_, _00227_);
  nand (_01766_, _01765_, _01759_);
  nand (_01767_, _01766_, _00561_);
  nand (_01768_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7]);
  nand (_01769_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7]);
  nand (_01770_, _01769_, _01768_);
  nand (_01771_, _01770_, _01417_);
  nand (_01773_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7]);
  nand (_01774_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7]);
  nand (_01775_, _01774_, _01773_);
  nand (_01776_, _01775_, _00227_);
  nand (_01777_, _01776_, _01771_);
  nand (_01778_, _01777_, _00560_);
  nand (_01779_, _01778_, _01767_);
  nand (_01780_, _01779_, _00466_);
  nand (_01781_, _01780_, _01755_);
  nand (_01782_, _01781_, _00247_);
  nor (_01783_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  nor (_01784_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7]);
  nor (_01786_, _01784_, _01783_);
  nand (_01787_, _01786_, _00227_);
  nand (_01789_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  nand (_01790_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7]);
  nand (_01791_, _01790_, _01789_);
  nand (_01792_, _01791_, _01417_);
  nand (_01793_, _01792_, _01787_);
  nand (_01794_, _01793_, _00561_);
  nor (_01795_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7]);
  nor (_01796_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  nor (_01797_, _01796_, _01795_);
  nand (_01798_, _01797_, _00227_);
  nand (_01799_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7]);
  nand (_01800_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7]);
  nand (_01801_, _01800_, _01799_);
  nand (_01802_, _01801_, _01417_);
  nand (_01803_, _01802_, _01798_);
  nand (_01804_, _01803_, _00560_);
  nand (_01805_, _01804_, _01794_);
  nand (_01806_, _01805_, _00465_);
  nand (_01807_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7]);
  nand (_01808_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7]);
  nand (_01809_, _01808_, _01807_);
  nand (_01810_, _01809_, _01417_);
  nand (_01811_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7]);
  nand (_01812_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7]);
  nand (_01813_, _01812_, _01811_);
  nand (_01814_, _01813_, _00227_);
  nand (_01815_, _01814_, _01810_);
  nand (_01816_, _01815_, _00561_);
  nand (_01817_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7]);
  nand (_01818_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7]);
  nand (_01819_, _01818_, _01817_);
  nand (_01820_, _01819_, _01417_);
  nand (_01821_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7]);
  nand (_01822_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7]);
  nand (_01823_, _01822_, _01821_);
  nand (_01824_, _01823_, _00227_);
  nand (_01825_, _01824_, _01820_);
  nand (_01826_, _01825_, _00560_);
  nand (_01828_, _01826_, _01816_);
  nand (_01829_, _01828_, _00466_);
  nand (_01830_, _01829_, _01806_);
  nand (_01831_, _01830_, _00248_);
  nand (_01832_, _01831_, _01782_);
  nand (_01833_, _01832_, _00319_);
  nand (_01834_, _01833_, _01729_);
  nor (_01836_, _01834_, _01629_);
  nor (_01837_, _01836_, _01628_);
  nor (_01838_, _01837_, _00156_);
  nand (_01839_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  nand (_01840_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  nand (_01841_, _01840_, _01839_);
  nand (_01842_, _01841_, _01417_);
  nand (_01843_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  nand (_01844_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  nand (_01845_, _01844_, _01843_);
  nand (_01846_, _01845_, _00227_);
  nand (_01847_, _01846_, _01842_);
  nand (_01848_, _01847_, _00560_);
  nand (_01850_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  nand (_01851_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  nand (_01852_, _01851_, _01850_);
  nand (_01853_, _01852_, _01417_);
  nand (_01854_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7]);
  nand (_01855_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  nand (_01856_, _01855_, _01854_);
  nand (_01857_, _01856_, _00227_);
  nand (_01858_, _01857_, _01853_);
  nand (_01859_, _01858_, _00561_);
  nand (_01860_, _01859_, _01848_);
  nand (_01861_, _01860_, _00466_);
  nor (_01862_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7]);
  nor (_01863_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  nor (_01864_, _01863_, _01862_);
  nand (_01865_, _01864_, _00227_);
  nand (_01866_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  nand (_01867_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7]);
  nand (_01868_, _01867_, _01866_);
  nand (_01869_, _01868_, _01417_);
  nand (_01871_, _01869_, _01865_);
  nand (_01872_, _01871_, _00560_);
  nor (_01873_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  nor (_01874_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  nor (_01875_, _01874_, _01873_);
  nand (_01876_, _01875_, _00227_);
  nand (_01878_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  nand (_01879_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  nand (_01880_, _01879_, _01878_);
  nand (_01881_, _01880_, _01417_);
  nand (_01882_, _01881_, _01876_);
  nand (_01883_, _01882_, _00561_);
  nand (_01884_, _01883_, _01872_);
  nand (_01885_, _01884_, _00465_);
  nand (_01887_, _01885_, _01861_);
  nand (_01888_, _01887_, _00248_);
  nand (_01889_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7]);
  nand (_01890_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  nand (_01891_, _01890_, _01889_);
  nand (_01892_, _01891_, _01417_);
  nand (_01893_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  nand (_01894_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7]);
  nand (_01895_, _01894_, _01893_);
  nand (_01896_, _01895_, _00227_);
  nand (_01897_, _01896_, _01892_);
  nand (_01898_, _01897_, _00560_);
  nand (_01899_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7]);
  nand (_01900_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7]);
  nand (_01901_, _01900_, _01899_);
  nand (_01902_, _01901_, _01417_);
  nand (_01904_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7]);
  nand (_01905_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7]);
  nand (_01906_, _01905_, _01904_);
  nand (_01907_, _01906_, _00227_);
  nand (_01909_, _01907_, _01902_);
  nand (_01910_, _01909_, _00561_);
  nand (_01911_, _01910_, _01898_);
  nand (_01912_, _01911_, _00466_);
  nor (_01913_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7]);
  nor (_01914_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7]);
  nor (_01915_, _01914_, _01913_);
  nand (_01916_, _01915_, _01417_);
  nor (_01917_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7]);
  nor (_01918_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7]);
  nor (_01919_, _01918_, _01917_);
  nand (_01920_, _01919_, _00227_);
  nand (_01921_, _01920_, _01916_);
  nand (_01922_, _01921_, _00560_);
  nor (_01923_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7]);
  nor (_01924_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7]);
  nor (_01925_, _01924_, _01923_);
  nand (_01926_, _01925_, _01417_);
  nor (_01927_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7]);
  nor (_01928_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7]);
  nor (_01929_, _01928_, _01927_);
  nand (_01930_, _01929_, _00227_);
  nand (_01931_, _01930_, _01926_);
  nand (_01932_, _01931_, _00561_);
  nand (_01933_, _01932_, _01922_);
  nand (_01934_, _01933_, _00465_);
  nand (_01936_, _01934_, _01912_);
  nand (_01937_, _01936_, _00247_);
  nand (_01939_, _01937_, _01888_);
  nand (_01940_, _01939_, _00319_);
  nand (_01941_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  nand (_01942_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  nand (_01943_, _01942_, _01941_);
  nand (_01944_, _01943_, _01417_);
  nand (_01945_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7]);
  nand (_01946_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  nand (_01947_, _01946_, _01945_);
  nand (_01948_, _01947_, _00227_);
  nand (_01949_, _01948_, _01944_);
  nand (_01950_, _01949_, _00560_);
  nand (_01951_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7]);
  nand (_01952_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  nand (_01953_, _01952_, _01951_);
  nand (_01954_, _01953_, _01417_);
  nand (_01956_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7]);
  nand (_01957_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7]);
  nand (_01958_, _01957_, _01956_);
  nand (_01959_, _01958_, _00227_);
  nand (_01960_, _01959_, _01954_);
  nand (_01961_, _01960_, _00561_);
  nand (_01962_, _01961_, _01950_);
  nand (_01963_, _01962_, _00466_);
  nor (_01964_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  nor (_01965_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7]);
  nor (_01966_, _01965_, _01964_);
  nand (_01967_, _01966_, _01417_);
  nor (_01969_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7]);
  nor (_01970_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7]);
  nor (_01971_, _01970_, _01969_);
  nand (_01972_, _01971_, _00227_);
  nand (_01973_, _01972_, _01967_);
  nand (_01974_, _01973_, _00560_);
  nor (_01975_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7]);
  nor (_01976_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7]);
  nor (_01978_, _01976_, _01975_);
  nand (_01979_, _01978_, _01417_);
  nor (_01980_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  nor (_01981_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7]);
  nor (_01982_, _01981_, _01980_);
  nand (_01983_, _01982_, _00227_);
  nand (_01984_, _01983_, _01979_);
  nand (_01985_, _01984_, _00561_);
  nand (_01986_, _01985_, _01974_);
  nand (_01987_, _01986_, _00465_);
  nand (_01988_, _01987_, _01963_);
  nand (_01989_, _01988_, _00247_);
  nand (_01990_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7]);
  nand (_01991_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  nand (_01992_, _01991_, _01990_);
  nand (_01993_, _01992_, _01417_);
  nand (_01994_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  nand (_01995_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7]);
  nand (_01996_, _01995_, _01994_);
  nand (_01997_, _01996_, _00227_);
  nand (_01998_, _01997_, _01993_);
  nand (_01999_, _01998_, _00560_);
  nand (_02000_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7]);
  nand (_02001_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7]);
  nand (_02002_, _02001_, _02000_);
  nand (_02003_, _02002_, _01417_);
  nand (_02004_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  nand (_02005_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7]);
  nand (_02006_, _02005_, _02004_);
  nand (_02007_, _02006_, _00227_);
  nand (_02008_, _02007_, _02003_);
  nand (_02009_, _02008_, _00561_);
  nand (_02010_, _02009_, _01999_);
  nand (_02011_, _02010_, _00466_);
  nor (_02013_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7]);
  nor (_02014_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7]);
  nor (_02015_, _02014_, _02013_);
  nand (_02016_, _02015_, _00227_);
  nand (_02017_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7]);
  nand (_02019_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7]);
  nand (_02020_, _02019_, _02017_);
  nand (_02021_, _02020_, _01417_);
  nand (_02022_, _02021_, _02016_);
  nand (_02023_, _02022_, _00560_);
  nor (_02024_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7]);
  nor (_02026_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  nor (_02027_, _02026_, _02024_);
  nand (_02028_, _02027_, _00227_);
  nand (_02029_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7]);
  nand (_02030_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7]);
  nand (_02031_, _02030_, _02029_);
  nand (_02032_, _02031_, _01417_);
  nand (_02033_, _02032_, _02028_);
  nand (_02034_, _02033_, _00561_);
  nand (_02035_, _02034_, _02023_);
  nand (_02036_, _02035_, _00465_);
  nand (_02037_, _02036_, _02011_);
  nand (_02038_, _02037_, _00248_);
  nand (_02039_, _02038_, _01989_);
  nand (_02040_, _02039_, _00320_);
  nand (_02041_, _02040_, _01940_);
  nor (_02042_, _02041_, _00386_);
  nand (_02043_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  nand (_02045_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  nand (_02046_, _02045_, _02043_);
  nand (_02047_, _02046_, _00227_);
  nand (_02048_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  nand (_02049_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7]);
  nand (_02051_, _02049_, _02048_);
  nand (_02053_, _02051_, _01417_);
  nand (_02054_, _02053_, _02047_);
  nand (_02055_, _02054_, _00560_);
  nand (_02056_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  nand (_02057_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  nand (_02058_, _02057_, _02056_);
  nand (_02059_, _02058_, _00227_);
  nand (_02060_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  nand (_02061_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  nand (_02062_, _02061_, _02060_);
  nand (_02063_, _02062_, _01417_);
  nand (_02064_, _02063_, _02059_);
  nand (_02065_, _02064_, _00561_);
  nand (_02066_, _02065_, _02055_);
  nand (_02067_, _02066_, _00466_);
  nand (_02068_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  nand (_02069_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  nand (_02070_, _02069_, _02068_);
  nand (_02071_, _02070_, _01417_);
  nor (_02072_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  nor (_02073_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7]);
  nor (_02075_, _02073_, _02072_);
  nand (_02076_, _02075_, _00227_);
  nand (_02078_, _02076_, _02071_);
  nand (_02079_, _02078_, _00560_);
  nand (_02080_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  nand (_02081_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  nand (_02082_, _02081_, _02080_);
  nand (_02084_, _02082_, _01417_);
  nor (_02085_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  nor (_02086_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  nor (_02087_, _02086_, _02085_);
  nand (_02088_, _02087_, _00227_);
  nand (_02091_, _02088_, _02084_);
  nand (_02092_, _02091_, _00561_);
  nand (_02093_, _02092_, _02079_);
  nand (_02094_, _02093_, _00465_);
  nand (_02095_, _02094_, _02067_);
  nand (_02096_, _02095_, _00248_);
  nand (_02097_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  nand (_02098_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  nand (_02099_, _02098_, _02097_);
  nand (_02100_, _02099_, _01417_);
  nand (_02101_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  nand (_02102_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  nand (_02104_, _02102_, _02101_);
  nand (_02105_, _02104_, _00227_);
  nand (_02106_, _02105_, _02100_);
  nand (_02107_, _02106_, _00560_);
  nand (_02108_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  nand (_02110_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  nand (_02111_, _02110_, _02108_);
  nand (_02112_, _02111_, _01417_);
  nand (_02113_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  nand (_02114_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7]);
  nand (_02115_, _02114_, _02113_);
  nand (_02116_, _02115_, _00227_);
  nand (_02117_, _02116_, _02112_);
  nand (_02118_, _02117_, _00561_);
  nand (_02119_, _02118_, _02107_);
  nand (_02120_, _02119_, _00466_);
  nor (_02121_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  nor (_02122_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  nor (_02124_, _02122_, _02121_);
  nand (_02125_, _02124_, _01417_);
  nor (_02126_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  nor (_02127_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  nor (_02128_, _02127_, _02126_);
  nand (_02129_, _02128_, _00227_);
  nand (_02130_, _02129_, _02125_);
  nand (_02131_, _02130_, _00560_);
  nor (_02132_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  nor (_02133_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  nor (_02134_, _02133_, _02132_);
  nor (_02135_, _02134_, _00227_);
  nor (_02136_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  nor (_02137_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  nor (_02138_, _02137_, _02136_);
  nor (_02140_, _02138_, _01417_);
  nor (_02141_, _02140_, _02135_);
  nand (_02142_, _02141_, _00561_);
  nand (_02143_, _02142_, _02131_);
  nand (_02144_, _02143_, _00465_);
  nand (_02146_, _02144_, _02120_);
  nand (_02148_, _02146_, _00247_);
  nand (_02149_, _02148_, _02096_);
  nand (_02150_, _02149_, _00320_);
  nand (_02151_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7]);
  nand (_02152_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  nand (_02153_, _02152_, _02151_);
  nand (_02154_, _02153_, _01417_);
  nand (_02155_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7]);
  nand (_02156_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  nand (_02157_, _02156_, _02155_);
  nand (_02158_, _02157_, _00227_);
  nand (_02159_, _02158_, _02154_);
  nand (_02160_, _02159_, _00560_);
  nand (_02161_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7]);
  nand (_02162_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  nand (_02163_, _02162_, _02161_);
  nand (_02164_, _02163_, _01417_);
  nand (_02165_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  nand (_02167_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7]);
  nand (_02168_, _02167_, _02165_);
  nand (_02169_, _02168_, _00227_);
  nand (_02171_, _02169_, _02164_);
  nand (_02172_, _02171_, _00561_);
  nand (_02173_, _02172_, _02160_);
  nand (_02174_, _02173_, _00466_);
  nor (_02175_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  nor (_02176_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7]);
  nor (_02177_, _02176_, _02175_);
  nand (_02178_, _02177_, _01417_);
  nor (_02180_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  nor (_02181_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7]);
  nor (_02182_, _02181_, _02180_);
  nand (_02183_, _02182_, _00227_);
  nand (_02184_, _02183_, _02178_);
  nand (_02185_, _02184_, _00560_);
  nor (_02186_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7]);
  nor (_02187_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  nor (_02188_, _02187_, _02186_);
  nand (_02189_, _02188_, _01417_);
  nor (_02190_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  nor (_02191_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  nor (_02192_, _02191_, _02190_);
  nand (_02193_, _02192_, _00227_);
  nand (_02194_, _02193_, _02189_);
  nand (_02195_, _02194_, _00561_);
  nand (_02196_, _02195_, _02185_);
  nand (_02197_, _02196_, _00465_);
  nand (_02198_, _02197_, _02174_);
  nand (_02199_, _02198_, _00247_);
  nand (_02201_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  nand (_02202_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  nand (_02203_, _02202_, _02201_);
  nand (_02204_, _02203_, _01417_);
  nand (_02205_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  nand (_02206_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  nand (_02207_, _02206_, _02205_);
  nand (_02208_, _02207_, _00227_);
  nand (_02209_, _02208_, _02204_);
  nand (_02210_, _02209_, _00560_);
  nand (_02211_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7]);
  nand (_02212_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7]);
  nand (_02213_, _02212_, _02211_);
  nand (_02214_, _02213_, _01417_);
  nand (_02215_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7]);
  nand (_02216_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  nand (_02217_, _02216_, _02215_);
  nand (_02218_, _02217_, _00227_);
  nand (_02219_, _02218_, _02214_);
  nand (_02221_, _02219_, _00561_);
  nand (_02222_, _02221_, _02210_);
  nand (_02223_, _02222_, _00466_);
  nor (_02224_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7]);
  nor (_02225_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  nor (_02226_, _02225_, _02224_);
  nand (_02228_, _02226_, _01417_);
  nor (_02229_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  nor (_02230_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7]);
  nor (_02231_, _02230_, _02229_);
  nand (_02232_, _02231_, _00227_);
  nand (_02234_, _02232_, _02228_);
  nand (_02235_, _02234_, _00560_);
  nor (_02236_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7]);
  nor (_02237_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  nor (_02238_, _02237_, _02236_);
  nand (_02239_, _02238_, _01417_);
  nor (_02240_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7]);
  nor (_02241_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  nor (_02242_, _02241_, _02240_);
  nand (_02244_, _02242_, _00227_);
  nand (_02245_, _02244_, _02239_);
  nand (_02246_, _02245_, _00561_);
  nand (_02247_, _02246_, _02235_);
  nand (_02248_, _02247_, _00465_);
  nand (_02249_, _02248_, _02223_);
  nand (_02250_, _02249_, _00248_);
  nand (_02251_, _02250_, _02199_);
  nand (_02252_, _02251_, _00319_);
  nand (_02253_, _02252_, _02150_);
  nor (_02254_, _02253_, _01629_);
  nor (_02256_, _02254_, _02042_);
  nor (_02257_, _02256_, _00556_);
  nor (_02258_, _02257_, _01838_);
  nor (_02259_, _02258_, _01416_);
  not (_02261_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  nand (_02262_, _01416_, _02261_);
  nand (_02263_, _02262_, _23493_);
  nor (_21116_, _02263_, _02259_);
  nor (_02264_, _23115_, _23043_);
  not (_02265_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nand (_02268_, _23043_, _02265_);
  nand (_02269_, _02268_, _23493_);
  nor (_25019_[6], _02269_, _02264_);
  nor (_02271_, _21786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  nor (_02272_, _21788_, _21504_);
  nor (_21120_, _02272_, _02271_);
  nor (_02274_, _22454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  nor (_02275_, _22456_, _21451_);
  nor (_21121_, _02275_, _02274_);
  nor (_02276_, _22838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  nor (_02278_, _22840_, _21474_);
  nor (_21122_, _02278_, _02276_);
  nor (_02280_, _23786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  nor (_02281_, _23789_, _21504_);
  nor (_21123_, _02281_, _02280_);
  nand (_02283_, _23490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  not (_02284_, _02283_);
  not (_02286_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  nor (_02287_, _23153_, _02286_);
  not (_02288_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor (_02289_, _23073_, _02288_);
  nor (_02290_, _23067_, _00366_);
  nor (_02291_, _02290_, _02289_);
  not (_02292_, _02291_);
  nor (_02293_, _23058_, _23098_);
  nor (_02295_, _23076_, _23105_);
  nor (_02296_, _02295_, _02293_);
  nor (_02298_, _23050_, _00370_);
  nor (_02299_, _23107_, _23103_);
  nor (_02300_, _02299_, _02298_);
  nand (_02302_, _02300_, _02296_);
  nor (_02303_, _02302_, _02292_);
  nor (_02304_, _02303_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_02305_, _02304_, _02287_);
  nor (_02306_, _02305_, _23490_);
  nor (_02307_, _02306_, _02284_);
  nor (_21124_, _02307_, rst);
  nor (_02308_, _23786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  nor (_02309_, _23789_, _21451_);
  nor (_21125_, _02309_, _02308_);
  nor (_02310_, _01083_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  nor (_02311_, _01052_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  nand (_02312_, _02311_, _01080_);
  nand (_02313_, _02312_, _23493_);
  nor (_21126_, _02313_, _02310_);
  nor (_02314_, _22479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  nor (_02315_, _22482_, _21586_);
  nor (_21127_, _02315_, _02314_);
  nor (_02316_, _23786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  nor (_02317_, _23789_, _21414_);
  nor (_21129_, _02317_, _02316_);
  nor (_02318_, _23786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  nor (_02319_, _23789_, _21526_);
  nor (_21130_, _02319_, _02318_);
  nor (_02320_, _22490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  nor (_02321_, _22492_, _21451_);
  nor (_21131_, _02321_, _02320_);
  nor (_02322_, _24159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  nor (_02323_, _24161_, _21474_);
  nor (_21134_, _02323_, _02322_);
  nor (_02324_, _24159_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  nor (_02325_, _24161_, _21586_);
  nor (_21135_, _02325_, _02324_);
  nor (_02326_, _23786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7]);
  nor (_02327_, _23789_, _21626_);
  nor (_21136_, _02327_, _02326_);
  nor (_02328_, _01183_, _21530_);
  nor (_02330_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  not (_02331_, _02328_);
  nor (_02332_, _02331_, _21451_);
  nor (_21140_, _02332_, _02330_);
  not (_02333_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_02334_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_02335_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nand (_02337_, _02335_, _02334_);
  nor (_02338_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  not (_02340_, _02338_);
  nor (_02341_, _02340_, _02337_);
  not (_02343_, _02341_);
  not (_02344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_02345_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nand (_02346_, _02345_, _02344_);
  nor (_02347_, _02346_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nand (_02348_, _02347_, _01134_);
  nor (_02349_, _02348_, _02343_);
  nor (_02350_, _02349_, _01142_);
  nor (_02351_, _02350_, _02333_);
  nand (_02352_, _01134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  not (_02353_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_02354_, _01134_, _02353_);
  nand (_02356_, _02354_, _01141_);
  nand (_02357_, _02356_, _02352_);
  nor (_02358_, _02357_, _02351_);
  nor (_02359_, _02358_, _01130_);
  not (_02360_, _01130_);
  nand (_02361_, _01055_, ABINPUT[3]);
  nor (_02362_, _02361_, _02360_);
  nor (_02363_, _02362_, _02359_);
  nor (_21141_, _02363_, rst);
  nor (_25044_[0], _21585_, rst);
  not (_02365_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nand (_02366_, _01137_, _02365_);
  nor (_02367_, _01137_, _02365_);
  nor (_02368_, _02367_, rst);
  nand (_02369_, _02368_, _02366_);
  nor (_21142_, _02369_, _01130_);
  nor (_21143_, _21473_, rst);
  nor (_21144_, _21553_, rst);
  nor (_02370_, _21645_, _21589_);
  nor (_02371_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  not (_02372_, _02370_);
  nor (_02373_, _02372_, _21474_);
  nor (_21145_, _02373_, _02371_);
  nor (_02374_, _23791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  nor (_02375_, _23793_, _21504_);
  nor (_21147_, _02375_, _02374_);
  nor (_02376_, _23791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  nor (_02377_, _23793_, _21451_);
  nor (_21148_, _02377_, _02376_);
  nor (_21149_, _21525_, rst);
  nor (_25044_[4], _21413_, rst);
  nand (_02379_, _02367_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_02380_, _02367_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_02381_, _02380_, rst);
  nand (_02382_, _02381_, _02379_);
  nor (_21150_, _02382_, _01130_);
  nor (_02383_, _01183_, _21821_);
  nor (_02384_, _02383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  not (_02385_, _02383_);
  nor (_02386_, _02385_, _21554_);
  nor (_21151_, _02386_, _02384_);
  not (_02387_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor (_02388_, _21308_, _21268_);
  nor (_02389_, _00917_, _00007_);
  nand (_02390_, _02389_, _02388_);
  nor (_02391_, _02390_, _00909_);
  nor (_02392_, _02391_, _02387_);
  nor (_02393_, _01127_, _00927_);
  not (_02394_, _02393_);
  not (_02395_, _02390_);
  nand (_02397_, _02395_, _00931_);
  nand (_02398_, _02397_, _02394_);
  nor (_02399_, _02398_, _02392_);
  nand (_02400_, _02393_, _24867_);
  nand (_02402_, _02400_, _23493_);
  nor (_21152_, _02402_, _02399_);
  nor (_21153_, _21450_, rst);
  nor (_21154_, _21503_, rst);
  not (_02403_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_02404_, _01075_, _02403_);
  not (_02405_, _02404_);
  nor (_02407_, _01072_, _01052_);
  not (_02408_, _02407_);
  nor (_02410_, _02408_, _02405_);
  nor (_02411_, _02410_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  nand (_02412_, _02404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not (_02413_, _02412_);
  nor (_02414_, _02413_, _01072_);
  nor (_02415_, _01066_, _01058_);
  nor (_02416_, _02415_, _01052_);
  not (_02418_, _02416_);
  nor (_02419_, _02418_, _02414_);
  nor (_02420_, _02419_, rst);
  not (_02421_, _02420_);
  nor (_21155_, _02421_, _02411_);
  nor (_02422_, _21899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  nor (_02423_, _21902_, _21526_);
  nor (_21156_, _02423_, _02422_);
  nor (_02424_, _22292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  nor (_02426_, _22294_, _21474_);
  nor (_21157_, _02426_, _02424_);
  nor (_02427_, _01183_, _21566_);
  nor (_02429_, _02427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7]);
  not (_02430_, _02427_);
  nor (_02431_, _02430_, _21626_);
  nor (_25323_, _02431_, _02429_);
  nor (_02432_, _22272_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  nor (_02433_, _22274_, _21474_);
  nor (_21158_, _02433_, _02432_);
  nor (_21159_, _00634_, rst);
  nor (_02434_, _23786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  nor (_02436_, _23789_, _21474_);
  nor (_21160_, _02436_, _02434_);
  not (_02437_, _00052_);
  nor (_21161_, _02437_, rst);
  nor (_02439_, _21821_, _21645_);
  nor (_02440_, _02439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  not (_02442_, _02439_);
  nor (_02443_, _02442_, _21451_);
  nor (_21162_, _02443_, _02440_);
  nor (_02444_, _23786_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  nor (_02445_, _23789_, _21586_);
  nor (_21163_, _02445_, _02444_);
  nor (_02446_, _23791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7]);
  nor (_02447_, _23793_, _21626_);
  nor (_21164_, _02447_, _02446_);
  not (_02448_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  not (_02449_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nor (_02450_, _01077_, _02449_);
  nand (_02451_, _02450_, _01067_);
  nand (_02453_, _02451_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_02454_, _02453_, _01081_);
  nor (_02455_, _02454_, _02448_);
  nand (_02456_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nor (_02458_, _02456_, _01079_);
  nor (_02459_, _02458_, _02455_);
  nor (_21165_, _02459_, rst);
  nor (_02461_, _01083_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  nor (_02462_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _01052_);
  nand (_02464_, _02462_, _01080_);
  nand (_02465_, _02464_, _23493_);
  nor (_21166_, _02465_, _02461_);
  nor (_02466_, _01233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  nor (_02467_, _01235_, _21586_);
  nor (_21167_, _02467_, _02466_);
  nand (_02468_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nand (_02469_, _01142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nand (_02470_, _02469_, _02468_);
  nor (_02471_, _02470_, _01130_);
  nor (_02472_, _01059_, _00129_);
  nor (_02473_, _01055_, _24900_);
  nor (_02474_, _02473_, _02472_);
  nand (_02475_, _02474_, _01130_);
  nand (_02476_, _02475_, _23493_);
  nor (_21168_, _02476_, _02471_);
  nand (_02478_, _02393_, _00121_);
  nand (_02479_, _02478_, _23493_);
  nor (_02480_, _00915_, _21308_);
  not (_02481_, _02480_);
  nor (_02482_, _01127_, _02481_);
  not (_02484_, _02482_);
  nor (_02485_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  not (_02486_, _02485_);
  nor (_02487_, _02486_, _01055_);
  nand (_02488_, _02487_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not (_02489_, _02487_);
  nand (_02490_, _02489_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nand (_02491_, _02490_, _02488_);
  nand (_02492_, _02491_, _02484_);
  not (_02493_, _01318_);
  nand (_02494_, _01027_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nand (_02495_, _02494_, _02493_);
  nand (_02496_, _02495_, _02482_);
  nand (_02497_, _02496_, _02492_);
  nor (_02498_, _02497_, _02393_);
  nor (_21169_, _02498_, _02479_);
  nor (_02499_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nand (_02500_, _23553_, _23070_);
  nand (_02501_, _02500_, _23493_);
  nor (_21170_, _02501_, _02499_);
  nor (_02502_, _21741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  nor (_02503_, _21744_, _21504_);
  nor (_21171_, _02503_, _02502_);
  nand (_02505_, _01017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_02507_, _01020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nand (_02508_, _02507_, _02505_);
  nor (_02509_, _02508_, _01030_);
  nor (_02510_, _01032_, ABINPUT[10]);
  nor (_02511_, _02510_, _02509_);
  nor (_02512_, _02511_, _01037_);
  not (_02513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nand (_02514_, _01037_, _02513_);
  nand (_02515_, _02514_, _23493_);
  nor (_21174_, _02515_, _02512_);
  nor (_02516_, _23795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7]);
  nor (_02517_, _23797_, _21626_);
  nor (_21175_, _02517_, _02516_);
  nor (_02518_, _23791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  nor (_02519_, _23793_, _21474_);
  nor (_21176_, _02519_, _02518_);
  nor (_02520_, _23791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  nor (_02521_, _23793_, _21586_);
  nor (_21178_, _02521_, _02520_);
  nor (_02522_, _22403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  nor (_02523_, _22406_, _21504_);
  nor (_25114_, _02523_, _02522_);
  nor (_02524_, _22403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  nor (_02525_, _22406_, _21586_);
  nor (_21179_, _02525_, _02524_);
  nor (_02526_, _23791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  nor (_02527_, _23793_, _21526_);
  nor (_21201_, _02527_, _02526_);
  nor (_02529_, _21873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  nor (_02530_, _21875_, _21451_);
  nor (_21204_, _02530_, _02529_);
  nor (_02532_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  nand (_02533_, _23553_, _24830_);
  nand (_02534_, _02533_, _23493_);
  nor (_21211_, _02534_, _02532_);
  nor (_02535_, _23791_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  nor (_02536_, _23793_, _21554_);
  nor (_21225_, _02536_, _02535_);
  nor (_02537_, _22557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  nor (_02538_, _22559_, _21474_);
  nor (_21228_, _02538_, _02537_);
  nor (_02539_, _22557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  nor (_02540_, _22559_, _21526_);
  nor (_21299_, _02540_, _02539_);
  nor (_02541_, _23795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  nor (_02542_, _23797_, _21554_);
  nor (_21326_, _02542_, _02541_);
  nor (_02543_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  nand (_02544_, _23553_, _00506_);
  nand (_02545_, _02544_, _23493_);
  nor (_21387_, _02545_, _02543_);
  nor (_02546_, _21949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  nor (_02547_, _21952_, _21474_);
  nor (_21399_, _02547_, _02546_);
  nor (_02548_, _23795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  nor (_02549_, _23797_, _21474_);
  nor (_21402_, _02549_, _02548_);
  nor (_02550_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7]);
  nor (_02551_, _22473_, _21626_);
  nor (_21405_, _02551_, _02550_);
  nor (_02552_, _21949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  nor (_02553_, _21952_, _21586_);
  nor (_21408_, _02553_, _02552_);
  nor (_02554_, _23795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  nor (_02555_, _23797_, _21586_);
  nor (_25385_, _02555_, _02554_);
  nor (_02556_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7]);
  nor (_02557_, _22537_, _21626_);
  nor (_21447_, _02557_, _02556_);
  nor (_02558_, _21559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7]);
  nor (_02559_, _21626_, _21561_);
  nor (_25254_, _02559_, _02558_);
  nor (_02560_, _21608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  nor (_02561_, _21610_, _21586_);
  nor (_21457_, _02561_, _02560_);
  nor (_02562_, _21608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  nor (_02563_, _21610_, _21526_);
  nor (_21460_, _02563_, _02562_);
  nor (_02564_, _21608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  nor (_02565_, _21610_, _21414_);
  nor (_21463_, _02565_, _02564_);
  nor (_02567_, _21608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  nor (_02568_, _21610_, _21451_);
  nor (_21471_, _02568_, _02567_);
  nor (_02569_, _21608_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  nor (_02570_, _21610_, _21504_);
  nor (_21489_, _02570_, _02569_);
  nor (_02572_, _21600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  nor (_02573_, _21602_, _21554_);
  nor (_21492_, _02573_, _02572_);
  nor (_02574_, _21600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  nor (_02575_, _21602_, _21526_);
  nor (_21509_, _02575_, _02574_);
  nor (_02576_, _21600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  nor (_02577_, _21602_, _21451_);
  nor (_21516_, _02577_, _02576_);
  nor (_02578_, _21600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7]);
  nor (_02579_, _21626_, _21602_);
  nor (_25252_, _02579_, _02578_);
  nor (_02580_, _21590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  nor (_02581_, _21592_, _21474_);
  nor (_21522_, _02581_, _02580_);
  nor (_02582_, _21590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  nor (_02583_, _21592_, _21554_);
  nor (_21527_, _02583_, _02582_);
  nor (_02584_, _21590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  nor (_02585_, _21592_, _21526_);
  nor (_21539_, _02585_, _02584_);
  nor (_02586_, _21590_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  nor (_02587_, _21592_, _21451_);
  nor (_21543_, _02587_, _02586_);
  nor (_02588_, _23795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  nor (_02589_, _23797_, _21451_);
  nor (_21594_, _02589_, _02588_);
  nor (_02590_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  nor (_02591_, _22783_, _21414_);
  nor (_21625_, _02591_, _02590_);
  nor (_02594_, _23795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  nor (_02595_, _23797_, _21414_);
  nor (_21628_, _02595_, _02594_);
  nor (_02596_, _22490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  nor (_02597_, _22492_, _21504_);
  nor (_21630_, _02597_, _02596_);
  nor (_02598_, _23795_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  nor (_02599_, _23797_, _21526_);
  nor (_21633_, _02599_, _02598_);
  nor (_02600_, _22869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7]);
  nor (_02601_, _22872_, _21626_);
  nor (_21650_, _02601_, _02600_);
  nor (_02602_, _22869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  nor (_02603_, _22872_, _21414_);
  nor (_21676_, _02603_, _02602_);
  nor (_02604_, _23799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  nor (_02606_, _23801_, _21414_);
  nor (_25383_, _02606_, _02604_);
  nor (_02607_, _22869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  nor (_02609_, _22872_, _21474_);
  nor (_21705_, _02609_, _02607_);
  nor (_02610_, _23799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  nor (_02611_, _23801_, _21526_);
  nor (_21710_, _02611_, _02610_);
  nor (_02612_, _01003_, _00018_);
  not (_02613_, _02612_);
  not (_02614_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_02615_, _00950_, _02614_);
  nor (_02616_, _02615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  not (_02618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not (_02619_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_02620_, _02619_, _02618_);
  nand (_02621_, _02620_, _23493_);
  nor (_02623_, _02621_, _02616_);
  nand (_02624_, _02623_, _02613_);
  nor (_02625_, _01029_, _00018_);
  not (_02626_, _02625_);
  not (_02627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not (_02628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_02630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not (_02631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_02632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_02633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  not (_02634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_02635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_02636_, _02635_, _02634_);
  not (_02637_, _02636_);
  nor (_02638_, _02637_, _02633_);
  not (_02639_, _02638_);
  nor (_02640_, _02639_, _02632_);
  not (_02641_, _02640_);
  nor (_02642_, _02641_, _02631_);
  not (_02644_, _02642_);
  nor (_02645_, _02644_, _02630_);
  not (_02646_, _02645_);
  nor (_02647_, _02646_, _02628_);
  not (_02648_, _02647_);
  nor (_02649_, _02648_, _02627_);
  not (_02650_, _02649_);
  nand (_02652_, _02650_, _02615_);
  nand (_02653_, _02652_, _02626_);
  nor (_21715_, _02653_, _02624_);
  nor (_02654_, _23799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  nor (_02655_, _23801_, _21554_);
  nor (_21721_, _02655_, _02654_);
  nor (_02656_, _02619_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nor (_02657_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _02618_);
  nor (_02658_, _02657_, _02656_);
  not (_02659_, _02658_);
  not (_02660_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  not (_02662_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not (_02663_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  not (_02664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  not (_02665_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_02666_, _02665_, _02664_);
  nand (_02667_, _02666_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_02669_, _02667_, _02663_);
  nand (_02670_, _02669_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_02671_, _02670_, _02662_);
  nand (_02672_, _02671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_02673_, _02672_, _02660_);
  not (_02674_, t0_i);
  nand (_02675_, _02674_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff );
  nand (_02677_, _02675_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  not (_02678_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nor (_02679_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nor (_02680_, _02679_, _02678_);
  nand (_02681_, _02680_, _02677_);
  nor (_02682_, _02681_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand (_02683_, _02682_, _02673_);
  nor (_02684_, _02683_, _02648_);
  not (_02685_, _02684_);
  nand (_02686_, _02685_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_02687_, _02684_, _02627_);
  nand (_02689_, _02687_, _02686_);
  nand (_02690_, _02689_, _02659_);
  not (_02691_, _02615_);
  nor (_02693_, _02648_, _02691_);
  nor (_02694_, _02693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  not (_02696_, _02693_);
  nor (_02698_, _02696_, _02627_);
  nor (_02699_, _02698_, _02694_);
  nand (_02700_, _02699_, _02620_);
  nand (_02701_, _02700_, _02690_);
  nor (_02702_, _02670_, _02681_);
  nand (_02704_, _02702_, _02649_);
  nor (_02705_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  not (_02707_, _02705_);
  not (_02708_, _02702_);
  nor (_02709_, _02708_, _02648_);
  nor (_02710_, _02709_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_02711_, _02710_, _02707_);
  nand (_02712_, _02711_, _02704_);
  nand (_02714_, _02712_, _02613_);
  nor (_02715_, _02714_, _02701_);
  nor (_02717_, _02613_, ABINPUT[10]);
  nor (_02718_, _02717_, _02715_);
  nor (_02719_, _02718_, _02625_);
  nand (_02720_, _02625_, _02627_);
  nand (_02722_, _02720_, _23493_);
  nor (_21740_, _02722_, _02719_);
  nand (_02723_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5]);
  nand (_02724_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  nand (_02725_, _02724_, _02723_);
  nand (_02726_, _02725_, _00227_);
  nand (_02727_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  nand (_02728_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5]);
  nand (_02729_, _02728_, _02727_);
  nand (_02730_, _02729_, _01417_);
  nand (_02731_, _02730_, _02726_);
  nand (_02732_, _02731_, _00560_);
  nand (_02734_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  nand (_02735_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  nand (_02736_, _02735_, _02734_);
  nand (_02737_, _02736_, _00227_);
  nand (_02738_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  nand (_02739_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5]);
  nand (_02740_, _02739_, _02738_);
  nand (_02741_, _02740_, _01417_);
  nand (_02743_, _02741_, _02737_);
  nand (_02744_, _02743_, _00561_);
  nand (_02745_, _02744_, _02732_);
  nand (_02746_, _02745_, _00466_);
  nand (_02747_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5]);
  nand (_02748_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5]);
  nand (_02749_, _02748_, _02747_);
  nand (_02750_, _02749_, _01417_);
  nor (_02751_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  nor (_02752_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5]);
  nor (_02753_, _02752_, _02751_);
  nand (_02754_, _02753_, _00227_);
  nand (_02756_, _02754_, _02750_);
  nand (_02757_, _02756_, _00560_);
  nand (_02758_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5]);
  nand (_02759_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  nand (_02760_, _02759_, _02758_);
  nand (_02761_, _02760_, _01417_);
  nor (_02762_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  nor (_02763_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5]);
  nor (_02765_, _02763_, _02762_);
  nand (_02766_, _02765_, _00227_);
  nand (_02768_, _02766_, _02761_);
  nand (_02769_, _02768_, _00561_);
  nand (_02771_, _02769_, _02757_);
  nand (_02772_, _02771_, _00465_);
  nand (_02773_, _02772_, _02746_);
  nand (_02774_, _02773_, _00248_);
  nand (_02775_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5]);
  nand (_02777_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  nand (_02778_, _02777_, _02775_);
  nand (_02779_, _02778_, _01417_);
  nand (_02780_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  nand (_02781_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5]);
  nand (_02782_, _02781_, _02780_);
  nand (_02784_, _02782_, _00227_);
  nand (_02785_, _02784_, _02779_);
  nand (_02787_, _02785_, _00560_);
  nand (_02789_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  nand (_02790_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5]);
  nand (_02792_, _02790_, _02789_);
  nand (_02794_, _02792_, _01417_);
  nand (_02795_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5]);
  nand (_02797_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5]);
  nand (_02798_, _02797_, _02795_);
  nand (_02799_, _02798_, _00227_);
  nand (_02800_, _02799_, _02794_);
  nand (_02801_, _02800_, _00561_);
  nand (_02803_, _02801_, _02787_);
  nand (_02804_, _02803_, _00466_);
  nor (_02805_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5]);
  nor (_02806_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5]);
  nor (_02807_, _02806_, _02805_);
  nand (_02808_, _02807_, _01417_);
  nor (_02810_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5]);
  nor (_02811_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5]);
  nor (_02813_, _02811_, _02810_);
  nand (_02814_, _02813_, _00227_);
  nand (_02815_, _02814_, _02808_);
  nand (_02816_, _02815_, _00560_);
  nor (_02818_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5]);
  nor (_02819_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5]);
  nor (_02820_, _02819_, _02818_);
  nor (_02821_, _02820_, _00227_);
  nor (_02822_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5]);
  nor (_02823_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5]);
  nor (_02824_, _02823_, _02822_);
  nor (_02825_, _02824_, _01417_);
  nor (_02826_, _02825_, _02821_);
  nand (_02827_, _02826_, _00561_);
  nand (_02828_, _02827_, _02816_);
  nand (_02830_, _02828_, _00465_);
  nand (_02831_, _02830_, _02804_);
  nand (_02833_, _02831_, _00247_);
  nand (_02835_, _02833_, _02774_);
  nand (_02836_, _02835_, _00320_);
  nand (_02838_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nand (_02839_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nand (_02840_, _02839_, _02838_);
  nand (_02841_, _02840_, _01417_);
  nand (_02843_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nand (_02845_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nand (_02846_, _02845_, _02843_);
  nand (_02848_, _02846_, _00227_);
  nand (_02849_, _02848_, _02841_);
  nand (_02851_, _02849_, _00560_);
  nand (_02852_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nand (_02854_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nand (_02855_, _02854_, _02852_);
  nand (_02856_, _02855_, _01417_);
  nand (_02858_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5]);
  nand (_02860_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nand (_02861_, _02860_, _02858_);
  nand (_02862_, _02861_, _00227_);
  nand (_02864_, _02862_, _02856_);
  nand (_02865_, _02864_, _00561_);
  nand (_02866_, _02865_, _02851_);
  nand (_02868_, _02866_, _00466_);
  nor (_02869_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_02870_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_02871_, _02870_, _02869_);
  nand (_02873_, _02871_, _01417_);
  nor (_02874_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_02875_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5]);
  nor (_02876_, _02875_, _02874_);
  nand (_02877_, _02876_, _00227_);
  nand (_02878_, _02877_, _02873_);
  nand (_02879_, _02878_, _00560_);
  not (_02880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nand (_02881_, _00650_, _02880_);
  nor (_02882_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_02883_, _02882_, _00227_);
  nand (_02884_, _02883_, _02881_);
  nor (_02885_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_02887_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_02889_, _02887_, _02885_);
  nand (_02890_, _02889_, _00227_);
  nand (_02891_, _02890_, _02884_);
  nand (_02892_, _02891_, _00561_);
  nand (_02893_, _02892_, _02879_);
  nand (_02895_, _02893_, _00465_);
  nand (_02896_, _02895_, _02868_);
  nand (_02897_, _02896_, _00248_);
  nand (_02898_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5]);
  nand (_02899_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  nand (_02900_, _02899_, _02898_);
  nand (_02901_, _02900_, _01417_);
  nand (_02902_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  nand (_02903_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  nand (_02904_, _02903_, _02902_);
  nand (_02905_, _02904_, _00227_);
  nand (_02906_, _02905_, _02901_);
  nand (_02907_, _02906_, _00560_);
  nand (_02908_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5]);
  nand (_02909_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5]);
  nand (_02910_, _02909_, _02908_);
  nand (_02912_, _02910_, _01417_);
  nand (_02913_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  nand (_02914_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  nand (_02915_, _02914_, _02913_);
  nand (_02917_, _02915_, _00227_);
  nand (_02918_, _02917_, _02912_);
  nand (_02920_, _02918_, _00561_);
  nand (_02921_, _02920_, _02907_);
  nand (_02922_, _02921_, _00466_);
  not (_02923_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  nand (_02924_, _00650_, _02923_);
  nor (_02925_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5]);
  nor (_02926_, _02925_, _00227_);
  nand (_02927_, _02926_, _02924_);
  nor (_02928_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  nor (_02929_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  nor (_02930_, _02929_, _02928_);
  nand (_02931_, _02930_, _00227_);
  nand (_02932_, _02931_, _02927_);
  nand (_02933_, _02932_, _00560_);
  nor (_02935_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5]);
  nor (_02936_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  nor (_02937_, _02936_, _02935_);
  nand (_02938_, _02937_, _01417_);
  nor (_02939_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  nor (_02940_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  nor (_02941_, _02940_, _02939_);
  nand (_02942_, _02941_, _00227_);
  nand (_02943_, _02942_, _02938_);
  nand (_02944_, _02943_, _00561_);
  nand (_02945_, _02944_, _02933_);
  nand (_02946_, _02945_, _00465_);
  nand (_02947_, _02946_, _02922_);
  nand (_02948_, _02947_, _00247_);
  nand (_02950_, _02948_, _02897_);
  nand (_02951_, _02950_, _00319_);
  nand (_02952_, _02951_, _02836_);
  nor (_02953_, _02952_, _00386_);
  nand (_02954_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5]);
  nand (_02955_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5]);
  nand (_02956_, _02955_, _02954_);
  nand (_02957_, _02956_, _00227_);
  nand (_02958_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5]);
  nand (_02959_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5]);
  nand (_02960_, _02959_, _02958_);
  nand (_02961_, _02960_, _01417_);
  nand (_02962_, _02961_, _02957_);
  nand (_02963_, _02962_, _00560_);
  nand (_02964_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5]);
  nand (_02965_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5]);
  nand (_02966_, _02965_, _02964_);
  nand (_02967_, _02966_, _00227_);
  nand (_02968_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5]);
  nand (_02969_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5]);
  nand (_02972_, _02969_, _02968_);
  nand (_02973_, _02972_, _01417_);
  nand (_02974_, _02973_, _02967_);
  nand (_02975_, _02974_, _00561_);
  nand (_02976_, _02975_, _02963_);
  nand (_02978_, _02976_, _00466_);
  nand (_02979_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5]);
  nand (_02980_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5]);
  nand (_02981_, _02980_, _02979_);
  nand (_02982_, _02981_, _01417_);
  nor (_02983_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5]);
  nor (_02984_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  nor (_02985_, _02984_, _02983_);
  nand (_02986_, _02985_, _00227_);
  nand (_02987_, _02986_, _02982_);
  nand (_02988_, _02987_, _00560_);
  nand (_02989_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5]);
  nand (_02990_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5]);
  nand (_02991_, _02990_, _02989_);
  nand (_02992_, _02991_, _01417_);
  nor (_02993_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  nor (_02994_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5]);
  nor (_02995_, _02994_, _02993_);
  nand (_02996_, _02995_, _00227_);
  nand (_02997_, _02996_, _02992_);
  nand (_02998_, _02997_, _00561_);
  nand (_02999_, _02998_, _02988_);
  nand (_03000_, _02999_, _00465_);
  nand (_03001_, _03000_, _02978_);
  nand (_03002_, _03001_, _00248_);
  nand (_03004_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  nand (_03006_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5]);
  nand (_03007_, _03006_, _03004_);
  nand (_03008_, _03007_, _01417_);
  nand (_03009_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  nand (_03010_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5]);
  nand (_03011_, _03010_, _03009_);
  nand (_03012_, _03011_, _00227_);
  nand (_03013_, _03012_, _03008_);
  nand (_03015_, _03013_, _00560_);
  nand (_03017_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  nand (_03018_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  nand (_03019_, _03018_, _03017_);
  nand (_03020_, _03019_, _01417_);
  nand (_03021_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5]);
  nand (_03022_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5]);
  nand (_03023_, _03022_, _03021_);
  nand (_03024_, _03023_, _00227_);
  nand (_03025_, _03024_, _03020_);
  nand (_03026_, _03025_, _00561_);
  nand (_03027_, _03026_, _03015_);
  nand (_03028_, _03027_, _00466_);
  nor (_03029_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5]);
  nor (_03030_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5]);
  nor (_03031_, _03030_, _03029_);
  nand (_03032_, _03031_, _01417_);
  nor (_03033_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  nor (_03034_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  nor (_03035_, _03034_, _03033_);
  nand (_03036_, _03035_, _00227_);
  nand (_03037_, _03036_, _03032_);
  nand (_03038_, _03037_, _00560_);
  nor (_03039_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  nor (_03040_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5]);
  nor (_03041_, _03040_, _03039_);
  nor (_03042_, _03041_, _00227_);
  nor (_03043_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  nor (_03044_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5]);
  nor (_03046_, _03044_, _03043_);
  nor (_03047_, _03046_, _01417_);
  nor (_03048_, _03047_, _03042_);
  nand (_03050_, _03048_, _00561_);
  nand (_03051_, _03050_, _03038_);
  nand (_03052_, _03051_, _00465_);
  nand (_03053_, _03052_, _03028_);
  nand (_03054_, _03053_, _00247_);
  nand (_03055_, _03054_, _03002_);
  nand (_03056_, _03055_, _00320_);
  nand (_03058_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5]);
  nand (_03059_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5]);
  nand (_03060_, _03059_, _03058_);
  nand (_03061_, _03060_, _01417_);
  nand (_03062_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5]);
  nand (_03063_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5]);
  nand (_03064_, _03063_, _03062_);
  nand (_03065_, _03064_, _00227_);
  nand (_03066_, _03065_, _03061_);
  nand (_03067_, _03066_, _00560_);
  nand (_03068_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5]);
  nand (_03069_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5]);
  nand (_03070_, _03069_, _03068_);
  nand (_03071_, _03070_, _01417_);
  nand (_03073_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5]);
  nand (_03074_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5]);
  nand (_03075_, _03074_, _03073_);
  nand (_03076_, _03075_, _00227_);
  nand (_03077_, _03076_, _03071_);
  nand (_03078_, _03077_, _00561_);
  nand (_03079_, _03078_, _03067_);
  nand (_03080_, _03079_, _00466_);
  nor (_03081_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5]);
  nor (_03082_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5]);
  nor (_03083_, _03082_, _03081_);
  nand (_03084_, _03083_, _01417_);
  nor (_03085_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5]);
  nor (_03086_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5]);
  nor (_03087_, _03086_, _03085_);
  nand (_03088_, _03087_, _00227_);
  nand (_03089_, _03088_, _03084_);
  nand (_03090_, _03089_, _00560_);
  not (_03092_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  nand (_03093_, _00650_, _03092_);
  nor (_03094_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  nor (_03095_, _03094_, _00227_);
  nand (_03096_, _03095_, _03093_);
  nor (_03097_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  nor (_03098_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  nor (_03099_, _03098_, _03097_);
  nand (_03100_, _03099_, _00227_);
  nand (_03101_, _03100_, _03096_);
  nand (_03102_, _03101_, _00561_);
  nand (_03103_, _03102_, _03090_);
  nand (_03104_, _03103_, _00465_);
  nand (_03105_, _03104_, _03080_);
  nand (_03106_, _03105_, _00248_);
  nand (_03107_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5]);
  nand (_03108_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5]);
  nand (_03109_, _03108_, _03107_);
  nand (_03111_, _03109_, _01417_);
  nand (_03112_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5]);
  nand (_03115_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5]);
  nand (_03116_, _03115_, _03112_);
  nand (_03117_, _03116_, _00227_);
  nand (_03118_, _03117_, _03111_);
  nand (_03120_, _03118_, _00560_);
  nand (_03121_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5]);
  nand (_03123_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5]);
  nand (_03124_, _03123_, _03121_);
  nand (_03125_, _03124_, _01417_);
  nand (_03126_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5]);
  nand (_03128_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5]);
  nand (_03129_, _03128_, _03126_);
  nand (_03131_, _03129_, _00227_);
  nand (_03132_, _03131_, _03125_);
  nand (_03133_, _03132_, _00561_);
  nand (_03134_, _03133_, _03120_);
  nand (_03135_, _03134_, _00466_);
  not (_03136_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5]);
  nand (_03138_, _00650_, _03136_);
  nor (_03139_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5]);
  nor (_03141_, _03139_, _00227_);
  nand (_03142_, _03141_, _03138_);
  nor (_03143_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5]);
  nor (_03144_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5]);
  nor (_03145_, _03144_, _03143_);
  nand (_03146_, _03145_, _00227_);
  nand (_03147_, _03146_, _03142_);
  nand (_03149_, _03147_, _00560_);
  nor (_03151_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5]);
  nor (_03152_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5]);
  nor (_03153_, _03152_, _03151_);
  nand (_03154_, _03153_, _01417_);
  nor (_03155_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5]);
  nor (_03156_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5]);
  nor (_03157_, _03156_, _03155_);
  nand (_03158_, _03157_, _00227_);
  nand (_03159_, _03158_, _03154_);
  nand (_03160_, _03159_, _00561_);
  nand (_03161_, _03160_, _03149_);
  nand (_03162_, _03161_, _00465_);
  nand (_03165_, _03162_, _03135_);
  nand (_03166_, _03165_, _00247_);
  nand (_03168_, _03166_, _03106_);
  nand (_03169_, _03168_, _00319_);
  nand (_03170_, _03169_, _03056_);
  nor (_03171_, _03170_, _01629_);
  nor (_03172_, _03171_, _02953_);
  nor (_03173_, _03172_, _00156_);
  nand (_03174_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5]);
  nand (_03175_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5]);
  nand (_03176_, _03175_, _03174_);
  nand (_03177_, _03176_, _01417_);
  nand (_03178_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  nand (_03179_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  nand (_03180_, _03179_, _03178_);
  nand (_03181_, _03180_, _00227_);
  nand (_03182_, _03181_, _03177_);
  nand (_03184_, _03182_, _00560_);
  nand (_03185_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5]);
  nand (_03186_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  nand (_03188_, _03186_, _03185_);
  nand (_03189_, _03188_, _01417_);
  nand (_03190_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5]);
  nand (_03191_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  nand (_03192_, _03191_, _03190_);
  nand (_03193_, _03192_, _00227_);
  nand (_03194_, _03193_, _03189_);
  nand (_03195_, _03194_, _00561_);
  nand (_03196_, _03195_, _03184_);
  nand (_03197_, _03196_, _00466_);
  nor (_03198_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  nor (_03199_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  nor (_03200_, _03199_, _03198_);
  nand (_03202_, _03200_, _01417_);
  nor (_03203_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5]);
  nor (_03204_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5]);
  nor (_03205_, _03204_, _03203_);
  nand (_03206_, _03205_, _00227_);
  nand (_03207_, _03206_, _03202_);
  nand (_03209_, _03207_, _00560_);
  nor (_03211_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5]);
  nor (_03213_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5]);
  nor (_03214_, _03213_, _03211_);
  nand (_03215_, _03214_, _01417_);
  nor (_03216_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  nor (_03217_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  nor (_03218_, _03217_, _03216_);
  nand (_03220_, _03218_, _00227_);
  nand (_03221_, _03220_, _03215_);
  nand (_03222_, _03221_, _00561_);
  nand (_03224_, _03222_, _03209_);
  nand (_03225_, _03224_, _00465_);
  nand (_03226_, _03225_, _03197_);
  nand (_03227_, _03226_, _00247_);
  nand (_03228_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  nand (_03229_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5]);
  nand (_03230_, _03229_, _03228_);
  nand (_03232_, _03230_, _01417_);
  nand (_03233_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5]);
  nand (_03234_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  nand (_03235_, _03234_, _03233_);
  nand (_03236_, _03235_, _00227_);
  nand (_03237_, _03236_, _03232_);
  nand (_03238_, _03237_, _00560_);
  nand (_03239_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5]);
  nand (_03240_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5]);
  nand (_03241_, _03240_, _03239_);
  nand (_03242_, _03241_, _01417_);
  nand (_03243_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  nand (_03244_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5]);
  nand (_03245_, _03244_, _03243_);
  nand (_03246_, _03245_, _00227_);
  nand (_03247_, _03246_, _03242_);
  nand (_03248_, _03247_, _00561_);
  nand (_03249_, _03248_, _03238_);
  nand (_03250_, _03249_, _00466_);
  nor (_03251_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5]);
  nor (_03252_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5]);
  nor (_03253_, _03252_, _03251_);
  nand (_03254_, _03253_, _00227_);
  nand (_03255_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5]);
  nand (_03257_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5]);
  nand (_03258_, _03257_, _03255_);
  nand (_03259_, _03258_, _01417_);
  nand (_03261_, _03259_, _03254_);
  nand (_03262_, _03261_, _00560_);
  nor (_03263_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  nor (_03264_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5]);
  nor (_03265_, _03264_, _03263_);
  nand (_03266_, _03265_, _00227_);
  nand (_03268_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5]);
  nand (_03269_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  nand (_03270_, _03269_, _03268_);
  nand (_03271_, _03270_, _01417_);
  nand (_03272_, _03271_, _03266_);
  nand (_03273_, _03272_, _00561_);
  nand (_03275_, _03273_, _03262_);
  nand (_03276_, _03275_, _00465_);
  nand (_03277_, _03276_, _03250_);
  nand (_03278_, _03277_, _00248_);
  nand (_03279_, _03278_, _03227_);
  nand (_03280_, _03279_, _00320_);
  nand (_03281_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5]);
  nand (_03283_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5]);
  nand (_03284_, _03283_, _03281_);
  nand (_03285_, _03284_, _01417_);
  nand (_03286_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5]);
  nand (_03287_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  nand (_03288_, _03287_, _03286_);
  nand (_03289_, _03288_, _00227_);
  nand (_03290_, _03289_, _03285_);
  nand (_03291_, _03290_, _00560_);
  nand (_03292_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  nand (_03293_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5]);
  nand (_03294_, _03293_, _03292_);
  nand (_03295_, _03294_, _01417_);
  nand (_03296_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  nand (_03297_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  nand (_03298_, _03297_, _03296_);
  nand (_03299_, _03298_, _00227_);
  nand (_03301_, _03299_, _03295_);
  nand (_03302_, _03301_, _00561_);
  nand (_03303_, _03302_, _03291_);
  nand (_03305_, _03303_, _00466_);
  nor (_03306_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  nor (_03307_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5]);
  nor (_03308_, _03307_, _03306_);
  nand (_03309_, _03308_, _00227_);
  nand (_03311_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  nand (_03312_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  nand (_03313_, _03312_, _03311_);
  nand (_03314_, _03313_, _01417_);
  nand (_03315_, _03314_, _03309_);
  nand (_03316_, _03315_, _00560_);
  nor (_03317_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  nor (_03318_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  nor (_03319_, _03318_, _03317_);
  nand (_03321_, _03319_, _00227_);
  nand (_03322_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  nand (_03323_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5]);
  nand (_03324_, _03323_, _03322_);
  nand (_03326_, _03324_, _01417_);
  nand (_03327_, _03326_, _03321_);
  nand (_03328_, _03327_, _00561_);
  nand (_03330_, _03328_, _03316_);
  nand (_03331_, _03330_, _00465_);
  nand (_03332_, _03331_, _03305_);
  nand (_03333_, _03332_, _00248_);
  nand (_03334_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  nand (_03335_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5]);
  nand (_03336_, _03335_, _03334_);
  nand (_03337_, _03336_, _01417_);
  nand (_03338_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  nand (_03339_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5]);
  nand (_03340_, _03339_, _03338_);
  nand (_03341_, _03340_, _00227_);
  nand (_03342_, _03341_, _03337_);
  nand (_03343_, _03342_, _00560_);
  nand (_03344_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5]);
  nand (_03345_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5]);
  nand (_03346_, _03345_, _03344_);
  nand (_03347_, _03346_, _01417_);
  nand (_03348_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5]);
  nand (_03349_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5]);
  nand (_03350_, _03349_, _03348_);
  nand (_03351_, _03350_, _00227_);
  nand (_03352_, _03351_, _03347_);
  nand (_03353_, _03352_, _00561_);
  nand (_03354_, _03353_, _03343_);
  nand (_03355_, _03354_, _00466_);
  nor (_03357_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5]);
  nor (_03358_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5]);
  nor (_03359_, _03358_, _03357_);
  nand (_03361_, _03359_, _01417_);
  nor (_03362_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5]);
  nor (_03363_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5]);
  nor (_03364_, _03363_, _03362_);
  nand (_03365_, _03364_, _00227_);
  nand (_03366_, _03365_, _03361_);
  nand (_03367_, _03366_, _00560_);
  nor (_03368_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5]);
  nor (_03369_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5]);
  nor (_03370_, _03369_, _03368_);
  nand (_03371_, _03370_, _01417_);
  nor (_03372_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5]);
  nor (_03373_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5]);
  nor (_03374_, _03373_, _03372_);
  nand (_03375_, _03374_, _00227_);
  nand (_03376_, _03375_, _03371_);
  nand (_03377_, _03376_, _00561_);
  nand (_03378_, _03377_, _03367_);
  nand (_03379_, _03378_, _00465_);
  nand (_03380_, _03379_, _03355_);
  nand (_03381_, _03380_, _00247_);
  nand (_03382_, _03381_, _03333_);
  nand (_03383_, _03382_, _00319_);
  nand (_03384_, _03383_, _03280_);
  nor (_03385_, _03384_, _00386_);
  nand (_03386_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  nand (_03388_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  nand (_03389_, _03388_, _03386_);
  nand (_03391_, _03389_, _01417_);
  nand (_03392_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  nand (_03393_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  nand (_03394_, _03393_, _03392_);
  nand (_03395_, _03394_, _00227_);
  nand (_03396_, _03395_, _03391_);
  nand (_03398_, _03396_, _00560_);
  nand (_03399_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  nand (_03400_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5]);
  nand (_03401_, _03400_, _03399_);
  nand (_03402_, _03401_, _01417_);
  nand (_03403_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  nand (_03404_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  nand (_03405_, _03404_, _03403_);
  nand (_03406_, _03405_, _00227_);
  nand (_03407_, _03406_, _03402_);
  nand (_03408_, _03407_, _00561_);
  nand (_03409_, _03408_, _03398_);
  nand (_03410_, _03409_, _00466_);
  nor (_03411_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  nor (_03412_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  nor (_03413_, _03412_, _03411_);
  nand (_03414_, _03413_, _00227_);
  nand (_03415_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  nand (_03416_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  nand (_03417_, _03416_, _03415_);
  nand (_03419_, _03417_, _01417_);
  nand (_03420_, _03419_, _03414_);
  nand (_03421_, _03420_, _00560_);
  nor (_03423_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  nor (_03424_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  nor (_03425_, _03424_, _03423_);
  nand (_03427_, _03425_, _00227_);
  nand (_03428_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  nand (_03429_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  nand (_03431_, _03429_, _03428_);
  nand (_03432_, _03431_, _01417_);
  nand (_03433_, _03432_, _03427_);
  nand (_03434_, _03433_, _00561_);
  nand (_03435_, _03434_, _03421_);
  nand (_03436_, _03435_, _00465_);
  nand (_03437_, _03436_, _03410_);
  nand (_03439_, _03437_, _00248_);
  nand (_03440_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  nand (_03442_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  nand (_03443_, _03442_, _03440_);
  nand (_03445_, _03443_, _01417_);
  nand (_03446_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  nand (_03447_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  nand (_03449_, _03447_, _03446_);
  nand (_03450_, _03449_, _00227_);
  nand (_03451_, _03450_, _03445_);
  nand (_03452_, _03451_, _00560_);
  nand (_03454_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  nand (_03455_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  nand (_03456_, _03455_, _03454_);
  nand (_03458_, _03456_, _01417_);
  nand (_03459_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  nand (_03461_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  nand (_03462_, _03461_, _03459_);
  nand (_03463_, _03462_, _00227_);
  nand (_03464_, _03463_, _03458_);
  nand (_03466_, _03464_, _00561_);
  nand (_03468_, _03466_, _03452_);
  nand (_03469_, _03468_, _00466_);
  nor (_03471_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  nor (_03472_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  nor (_03474_, _03472_, _03471_);
  nand (_03475_, _03474_, _01417_);
  nor (_03476_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  nor (_03477_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5]);
  nor (_03479_, _03477_, _03476_);
  nand (_03480_, _03479_, _00227_);
  nand (_03481_, _03480_, _03475_);
  nand (_03482_, _03481_, _00560_);
  nor (_03483_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  nor (_03484_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  nor (_03485_, _03484_, _03483_);
  nand (_03486_, _03485_, _01417_);
  nor (_03488_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  nor (_03489_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  nor (_03490_, _03489_, _03488_);
  nand (_03491_, _03490_, _00227_);
  nand (_03492_, _03491_, _03486_);
  nand (_03493_, _03492_, _00561_);
  nand (_03494_, _03493_, _03482_);
  nand (_03495_, _03494_, _00465_);
  nand (_03496_, _03495_, _03469_);
  nand (_03497_, _03496_, _00247_);
  nand (_03498_, _03497_, _03439_);
  nand (_03499_, _03498_, _00320_);
  nor (_03500_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5]);
  nor (_03502_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  nor (_03503_, _03502_, _03500_);
  nand (_03504_, _03503_, _01417_);
  nor (_03506_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5]);
  nor (_03507_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  nor (_03508_, _03507_, _03506_);
  nand (_03509_, _03508_, _00227_);
  nand (_03510_, _03509_, _03504_);
  nand (_03511_, _03510_, _00561_);
  nor (_03512_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5]);
  nor (_03513_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5]);
  nor (_03514_, _03513_, _03512_);
  nand (_03515_, _03514_, _01417_);
  nor (_03516_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  nor (_03517_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5]);
  nor (_03518_, _03517_, _03516_);
  nand (_03519_, _03518_, _00227_);
  nand (_03521_, _03519_, _03515_);
  nand (_03522_, _03521_, _00560_);
  nand (_03523_, _03522_, _03511_);
  nand (_03524_, _03523_, _00465_);
  nand (_03525_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5]);
  nand (_03526_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5]);
  nand (_03527_, _03526_, _03525_);
  nand (_03528_, _03527_, _01417_);
  nand (_03529_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5]);
  nand (_03530_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5]);
  nand (_03532_, _03530_, _03529_);
  nand (_03534_, _03532_, _00227_);
  nand (_03535_, _03534_, _03528_);
  nand (_03536_, _03535_, _00561_);
  nand (_03537_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  nand (_03538_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5]);
  nand (_03539_, _03538_, _03537_);
  nand (_03540_, _03539_, _01417_);
  nand (_03541_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  nand (_03543_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  nand (_03544_, _03543_, _03541_);
  nand (_03546_, _03544_, _00227_);
  nand (_03548_, _03546_, _03540_);
  nand (_03549_, _03548_, _00560_);
  nand (_03550_, _03549_, _03536_);
  nand (_03551_, _03550_, _00466_);
  nand (_03552_, _03551_, _03524_);
  nand (_03553_, _03552_, _00247_);
  nor (_03554_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  nor (_03555_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  nor (_03556_, _03555_, _03554_);
  nand (_03557_, _03556_, _00227_);
  nand (_03558_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  nand (_03559_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5]);
  nand (_03560_, _03559_, _03558_);
  nand (_03562_, _03560_, _01417_);
  nand (_03563_, _03562_, _03557_);
  nand (_03564_, _03563_, _00561_);
  nor (_03565_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5]);
  nor (_03566_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5]);
  nor (_03567_, _03566_, _03565_);
  nand (_03568_, _03567_, _00227_);
  nand (_03569_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  nand (_03570_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5]);
  nand (_03571_, _03570_, _03569_);
  nand (_03572_, _03571_, _01417_);
  nand (_03573_, _03572_, _03568_);
  nand (_03574_, _03573_, _00560_);
  nand (_03575_, _03574_, _03564_);
  nand (_03576_, _03575_, _00465_);
  nand (_03579_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  nand (_03580_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  nand (_03581_, _03580_, _03579_);
  nand (_03582_, _03581_, _01417_);
  nand (_03583_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5]);
  nand (_03584_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  nand (_03585_, _03584_, _03583_);
  nand (_03586_, _03585_, _00227_);
  nand (_03587_, _03586_, _03582_);
  nand (_03588_, _03587_, _00561_);
  nand (_03589_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  nand (_03590_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  nand (_03591_, _03590_, _03589_);
  nand (_03592_, _03591_, _01417_);
  nand (_03593_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  nand (_03594_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  nand (_03595_, _03594_, _03593_);
  nand (_03596_, _03595_, _00227_);
  nand (_03598_, _03596_, _03592_);
  nand (_03599_, _03598_, _00560_);
  nand (_03600_, _03599_, _03588_);
  nand (_03602_, _03600_, _00466_);
  nand (_03603_, _03602_, _03576_);
  nand (_03604_, _03603_, _00248_);
  nand (_03605_, _03604_, _03553_);
  nand (_03607_, _03605_, _00319_);
  nand (_03608_, _03607_, _03499_);
  nor (_03609_, _03608_, _01629_);
  nor (_03610_, _03609_, _03385_);
  nor (_03611_, _03610_, _00556_);
  nor (_03613_, _03611_, _03173_);
  nor (_03614_, _03613_, _01416_);
  not (_03615_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  nand (_03616_, _01416_, _03615_);
  nand (_03617_, _03616_, _23493_);
  nor (_21743_, _03617_, _03614_);
  not (_03618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  not (_03619_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  not (_03620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  not (_03621_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_03622_, _03621_, _03620_);
  nand (_03623_, _03622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_03624_, _03623_, _03619_);
  nand (_03625_, _03624_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  not (_03626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  not (_03627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_03628_, _03627_, _03626_);
  nand (_03629_, _03628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_03630_, _03629_, _03625_);
  not (_03631_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  not (_03632_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  not (_03633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_03635_, _03633_, _03632_);
  not (_03636_, _03635_);
  nor (_03638_, _03636_, _03631_);
  nand (_03639_, _03638_, _03630_);
  not (_03641_, _03639_);
  not (_03642_, t1_i);
  nand (_03643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _03642_);
  nand (_03644_, _03643_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  nor (_03646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _02614_);
  not (_03648_, _03646_);
  nor (_03649_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  nor (_03650_, _03649_, _03648_);
  nand (_03652_, _03650_, _03644_);
  not (_03653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not (_03654_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  not (_03656_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_03657_, _03656_, _03654_);
  not (_03659_, _03657_);
  nor (_03660_, _03659_, _03653_);
  not (_03661_, _03660_);
  nor (_03662_, _03661_, _03652_);
  nand (_03664_, _03662_, _03641_);
  not (_03665_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  not (_03666_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nor (_03667_, _03666_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_03668_, _03667_);
  nor (_03669_, _03668_, _03665_);
  not (_03670_, _03669_);
  nor (_03672_, _03670_, _03664_);
  nor (_03673_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_03674_, _03661_, _03665_);
  nand (_03675_, _03674_, _03638_);
  nor (_03676_, _03652_, _03625_);
  not (_03677_, _03676_);
  nor (_03678_, _03677_, _03675_);
  nand (_03679_, _03678_, _03673_);
  not (_03680_, _03679_);
  nor (_03681_, _03680_, _03672_);
  nor (_03682_, _03681_, _03618_);
  not (_03683_, _03681_);
  nor (_03685_, _03683_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_03686_, _03685_, _03682_);
  nor (_03687_, _01012_, _00018_);
  not (_03688_, _03687_);
  nand (_03689_, _03688_, _03686_);
  nor (_03691_, _01010_, _21308_);
  nand (_03692_, _03691_, _00009_);
  nor (_03694_, _03692_, _00010_);
  nand (_03695_, _03694_, ABINPUT[10]);
  nand (_03697_, _03695_, _03689_);
  nand (_03698_, _21351_, _24877_);
  nor (_03700_, _00907_, _03698_);
  nand (_03701_, _03700_, _24861_);
  nor (_03702_, _03701_, _00018_);
  nor (_03703_, _03702_, _03697_);
  nand (_03704_, _03702_, _03618_);
  nand (_03705_, _03704_, _23493_);
  nor (_21746_, _03705_, _03703_);
  nor (_03706_, _22512_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7]);
  nor (_03708_, _22514_, _21626_);
  nor (_21755_, _03708_, _03706_);
  nor (_03709_, _23799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7]);
  nor (_03710_, _23801_, _21626_);
  nor (_25384_, _03710_, _03709_);
  nor (_03711_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  nand (_03712_, _23553_, _00444_);
  nand (_03714_, _03712_, _23493_);
  nor (_21765_, _03714_, _03711_);
  nor (_03717_, _23799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  nor (_03718_, _23801_, _21504_);
  nor (_21770_, _03718_, _03717_);
  nor (_03719_, _21850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  nor (_03720_, _21853_, _21474_);
  nor (_21781_, _03720_, _03719_);
  nor (_03721_, _01129_, _00018_);
  nor (_03722_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nand (_03723_, _03721_, _24900_);
  nand (_03724_, _03723_, _23493_);
  nor (_21793_, _03724_, _03722_);
  nor (_03726_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_03727_, _03721_, _00029_);
  nand (_03728_, _03727_, _23493_);
  nor (_21795_, _03728_, _03726_);
  nor (_03729_, _02660_, _02662_);
  nand (_03730_, _03729_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_03731_, _03730_, _02708_);
  nand (_03732_, _03731_, _02619_);
  nor (_03733_, _03732_, _02639_);
  not (_03734_, _03733_);
  nor (_03735_, _03734_, _02632_);
  nand (_03736_, _03735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_03737_, _03736_, _02630_);
  nor (_03738_, _03737_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_03739_, _03738_, _02658_);
  nand (_03740_, _03739_, _02685_);
  nor (_03741_, _02644_, _02691_);
  not (_03742_, _03741_);
  nor (_03743_, _03742_, _02630_);
  nor (_03744_, _03743_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_03745_, _02696_, _02620_);
  nor (_03746_, _03745_, _03744_);
  nand (_03747_, _02702_, _02638_);
  nor (_03748_, _03747_, _02632_);
  nand (_03750_, _03748_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_03751_, _03750_, _02630_);
  nor (_03752_, _03751_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_03753_, _02709_);
  nand (_03754_, _03753_, _02705_);
  nor (_03755_, _03754_, _03752_);
  nor (_03756_, _03755_, _03746_);
  nand (_03758_, _03756_, _03740_);
  nand (_03759_, _03758_, _02613_);
  nor (_03760_, _21351_, _21308_);
  nand (_03761_, _03760_, _24857_);
  nor (_03763_, _03761_, _00018_);
  nand (_03764_, _03763_, _24861_);
  not (_03765_, _03764_);
  nand (_03766_, _03765_, ABINPUT[9]);
  nand (_03767_, _03766_, _03759_);
  nor (_03768_, _03767_, _02625_);
  nand (_03769_, _02625_, _02628_);
  nand (_03770_, _03769_, _23493_);
  nor (_21797_, _03770_, _03768_);
  nand (_03771_, _03734_, _02632_);
  nor (_03772_, _03735_, _02658_);
  nand (_03773_, _03772_, _03771_);
  nand (_03774_, _02636_, _02615_);
  nor (_03775_, _03774_, _02633_);
  not (_03776_, _03775_);
  nor (_03777_, _03776_, _02632_);
  nand (_03779_, _03776_, _02632_);
  nand (_03781_, _03779_, _02620_);
  nor (_03783_, _03781_, _03777_);
  nor (_03784_, _02708_, _02641_);
  nand (_03785_, _03747_, _02632_);
  nand (_03787_, _03785_, _02705_);
  nor (_03788_, _03787_, _03784_);
  nor (_03790_, _03788_, _03783_);
  nand (_03792_, _03790_, _03773_);
  nand (_03793_, _03792_, _03764_);
  nand (_03794_, _03765_, ABINPUT[6]);
  nand (_03795_, _03794_, _03793_);
  nor (_03796_, _03795_, _02625_);
  nand (_03798_, _02625_, _02632_);
  nand (_03799_, _03798_, _23493_);
  nor (_21800_, _03799_, _03796_);
  nor (_03802_, _01025_, _03698_);
  nand (_03803_, _03802_, _00009_);
  nor (_03804_, _03803_, _00010_);
  not (_03805_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand (_03806_, _02612_, _03805_);
  nor (_03807_, _02708_, _02662_);
  not (_03808_, _03807_);
  nand (_03809_, _03808_, _03805_);
  nand (_03810_, _03807_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nand (_03811_, _03810_, _02707_);
  nand (_03812_, _03811_, _02613_);
  nand (_03814_, _03812_, _03809_);
  nor (_03817_, _02707_, _03805_);
  nand (_03819_, _03731_, _02656_);
  nand (_03821_, _02659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_03822_, _03821_, _03819_);
  nor (_03823_, _03822_, _03817_);
  nand (_03824_, _03823_, _03814_);
  nand (_03825_, _03824_, _03806_);
  nor (_03826_, _03825_, _03804_);
  nor (_03827_, _02626_, _00114_);
  nor (_03828_, _03827_, _03826_);
  nor (_21802_, _03828_, rst);
  not (_03829_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_03830_, _02681_, _02665_);
  nand (_03831_, _03830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_03832_, _03831_, _03829_);
  nand (_03833_, _03832_, _02613_);
  nand (_03834_, _03833_, _02663_);
  nand (_03835_, _03832_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_03836_, _03819_, _02632_);
  nor (_03837_, _03836_, _03835_);
  nand (_03838_, _03837_, _02613_);
  nand (_03839_, _03838_, _03834_);
  nor (_03840_, _03839_, _03804_);
  nor (_03841_, _02626_, _24867_);
  nor (_03842_, _03841_, _03840_);
  nor (_21803_, _03842_, rst);
  nor (_03843_, _01036_, _00018_);
  nor (_03844_, _03652_, _03654_);
  not (_03845_, _03844_);
  nor (_03847_, _03845_, _03639_);
  nand (_03849_, _03847_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_03850_, _03849_, _03667_);
  not (_03851_, _03850_);
  nor (_03852_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_03854_, _03852_);
  nor (_03855_, _03854_, _03625_);
  nand (_03856_, _03855_, _03638_);
  nor (_03857_, _03856_, _03659_);
  nor (_03858_, _03857_, _03667_);
  nor (_03860_, _03858_, _03851_);
  nor (_03862_, _03860_, _03687_);
  nor (_03864_, _03862_, _03843_);
  nor (_03866_, _03864_, _03656_);
  not (_03867_, _03847_);
  nor (_03868_, _03850_, _03867_);
  not (_03869_, _03858_);
  not (_03870_, _03856_);
  nand (_03872_, _03870_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_03874_, _03872_, _03869_);
  nor (_03876_, _03874_, _03868_);
  nor (_03879_, _03876_, _03687_);
  nor (_03881_, _03688_, _24900_);
  nor (_03883_, _03881_, _03879_);
  nor (_03885_, _03883_, _03843_);
  nor (_03886_, _03885_, _03866_);
  nor (_21807_, _03886_, rst);
  nor (_03889_, _03677_, _03626_);
  not (_03890_, _03889_);
  nor (_03891_, _03890_, _03627_);
  nand (_03893_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  not (_03894_, _03893_);
  nor (_03896_, _03894_, _03668_);
  nor (_03897_, _03855_, _03667_);
  nor (_03898_, _03897_, _03896_);
  nor (_03900_, _03898_, _03632_);
  not (_03902_, _03898_);
  nor (_03903_, _03902_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_03905_, _03903_, _03900_);
  nor (_03907_, _03905_, _03687_);
  not (_03909_, _03843_);
  nand (_03910_, _03687_, ABINPUT[3]);
  nand (_03912_, _03910_, _03909_);
  nor (_03913_, _03912_, _03907_);
  nand (_03914_, _03702_, _03632_);
  nand (_03915_, _03914_, _23493_);
  nor (_21809_, _03915_, _03913_);
  not (_03916_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  not (_03917_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_03918_, _03666_, _03917_);
  nor (_03919_, _03918_, _03687_);
  nor (_03921_, _03919_, _03916_);
  not (_03922_, _03702_);
  nor (_03923_, _03652_, _03623_);
  not (_03924_, _03923_);
  nor (_03925_, _03924_, _03619_);
  not (_03926_, _03925_);
  nand (_03927_, _03926_, _03916_);
  nor (_03929_, _03918_, _03676_);
  nand (_03931_, _03929_, _03927_);
  not (_03932_, _03629_);
  nor (_03934_, _03926_, _03916_);
  nand (_03935_, _03934_, _03932_);
  nor (_03937_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _03917_);
  not (_03939_, _03937_);
  nor (_03940_, _03939_, _03935_);
  nand (_03942_, _03940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_03944_, _03942_, _03931_);
  nand (_03945_, _03944_, _03688_);
  nand (_03947_, _03945_, _03922_);
  nor (_03948_, _03947_, _03921_);
  nand (_03950_, _03702_, _24900_);
  nand (_03952_, _03950_, _23493_);
  nor (_21813_, _03952_, _03948_);
  nor (_03953_, _03919_, _03621_);
  not (_03954_, _03652_);
  nor (_03956_, _03954_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_03958_, _03652_, _03621_);
  nor (_03959_, _03918_, _03958_);
  nand (_03960_, _03630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_03961_, _03937_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_03963_, _03961_, _03960_);
  nor (_03965_, _03963_, _03959_);
  nor (_03966_, _03965_, _03956_);
  nand (_03968_, _03966_, _03688_);
  nand (_03970_, _03968_, _03922_);
  nor (_03972_, _03970_, _03953_);
  nand (_03974_, _03702_, _00029_);
  nand (_03975_, _03974_, _23493_);
  nor (_21815_, _03975_, _03972_);
  nor (_03976_, _21652_, _21645_);
  nor (_03977_, _03976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  not (_03978_, _03976_);
  nor (_03979_, _03978_, _21586_);
  nor (_21828_, _03979_, _03977_);
  nor (_03980_, _01083_, _02449_);
  nand (_03981_, _03980_, _23493_);
  nand (_03982_, _02451_, _01079_);
  not (_03984_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  nor (_03985_, rst, _01052_);
  not (_03986_, _03985_);
  nor (_03988_, _03986_, _03984_);
  nand (_03989_, _03988_, _03982_);
  nand (_21833_, _03989_, _03981_);
  nand (_03990_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  nand (_03992_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  nand (_03993_, _03992_, _03990_);
  nand (_03994_, _03993_, _01417_);
  nand (_03995_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  nand (_03996_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1]);
  nand (_03997_, _03996_, _03995_);
  nand (_03998_, _03997_, _00227_);
  nand (_03999_, _03998_, _03994_);
  nand (_04000_, _03999_, _00560_);
  nand (_04001_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1]);
  nand (_04002_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1]);
  nand (_04003_, _04002_, _04001_);
  nand (_04004_, _04003_, _01417_);
  nand (_04005_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1]);
  nand (_04006_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1]);
  nand (_04007_, _04006_, _04005_);
  nand (_04009_, _04007_, _00227_);
  nand (_04010_, _04009_, _04004_);
  nand (_04012_, _04010_, _00561_);
  nand (_04014_, _04012_, _04000_);
  nand (_04015_, _04014_, _00466_);
  nor (_04017_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1]);
  nor (_04018_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1]);
  nor (_04020_, _04018_, _04017_);
  nand (_04022_, _04020_, _01417_);
  nor (_04023_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1]);
  nor (_04026_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1]);
  nor (_04027_, _04026_, _04023_);
  nand (_04029_, _04027_, _00227_);
  nand (_04030_, _04029_, _04022_);
  nand (_04032_, _04030_, _00560_);
  nor (_04033_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1]);
  nor (_04034_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1]);
  nor (_04035_, _04034_, _04033_);
  nand (_04037_, _04035_, _01417_);
  nor (_04038_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1]);
  nor (_04040_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1]);
  nor (_04041_, _04040_, _04038_);
  nand (_04043_, _04041_, _00227_);
  nand (_04045_, _04043_, _04037_);
  nand (_04046_, _04045_, _00561_);
  nand (_04048_, _04046_, _04032_);
  nand (_04049_, _04048_, _00465_);
  nand (_04051_, _04049_, _04015_);
  nor (_04052_, _04051_, _00248_);
  nand (_04053_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  nand (_04055_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  nand (_04057_, _04055_, _04053_);
  nand (_04058_, _04057_, _01417_);
  nand (_04060_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  nand (_04061_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  nand (_04062_, _04061_, _04060_);
  nand (_04063_, _04062_, _00227_);
  nand (_04064_, _04063_, _04058_);
  nand (_04065_, _04064_, _00560_);
  nand (_04067_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1]);
  nand (_04069_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1]);
  nand (_04070_, _04069_, _04067_);
  nand (_04072_, _04070_, _01417_);
  nand (_04073_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  nand (_04075_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  nand (_04076_, _04075_, _04073_);
  nand (_04078_, _04076_, _00227_);
  nand (_04079_, _04078_, _04072_);
  nand (_04081_, _04079_, _00561_);
  nand (_04082_, _04081_, _04065_);
  nand (_04084_, _04082_, _00466_);
  nor (_04085_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1]);
  nor (_04086_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  nor (_04087_, _04086_, _04085_);
  nand (_04088_, _04087_, _00227_);
  nand (_04089_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  nand (_04091_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1]);
  nand (_04092_, _04091_, _04089_);
  nand (_04094_, _04092_, _01417_);
  nand (_04095_, _04094_, _04088_);
  nand (_04096_, _04095_, _00560_);
  nor (_04097_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1]);
  nor (_04098_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1]);
  nor (_04099_, _04098_, _04097_);
  nand (_04101_, _04099_, _00227_);
  nand (_04102_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  nand (_04103_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  nand (_04104_, _04103_, _04102_);
  nand (_04105_, _04104_, _01417_);
  nand (_04107_, _04105_, _04101_);
  nand (_04108_, _04107_, _00561_);
  nand (_04109_, _04108_, _04096_);
  nand (_04110_, _04109_, _00465_);
  nand (_04111_, _04110_, _04084_);
  nor (_04112_, _04111_, _00247_);
  nor (_04113_, _04112_, _04052_);
  nand (_04114_, _04113_, _00320_);
  nand (_04115_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1]);
  nand (_04116_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1]);
  nand (_04117_, _04116_, _04115_);
  nand (_04118_, _04117_, _01417_);
  nand (_04119_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nand (_04120_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nand (_04121_, _04120_, _04119_);
  nand (_04122_, _04121_, _00227_);
  nand (_04123_, _04122_, _04118_);
  nand (_04124_, _04123_, _00560_);
  nand (_04126_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1]);
  nand (_04127_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1]);
  nand (_04129_, _04127_, _04126_);
  nand (_04131_, _04129_, _01417_);
  nand (_04132_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1]);
  nand (_04133_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nand (_04134_, _04133_, _04132_);
  nand (_04135_, _04134_, _00227_);
  nand (_04137_, _04135_, _04131_);
  nand (_04138_, _04137_, _00561_);
  nand (_04139_, _04138_, _04124_);
  nand (_04140_, _04139_, _00466_);
  nor (_04142_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_04143_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_04145_, _04143_, _04142_);
  nand (_04146_, _04145_, _00227_);
  nand (_04147_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1]);
  nand (_04148_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nand (_04149_, _04148_, _04147_);
  nand (_04150_, _04149_, _01417_);
  nand (_04151_, _04150_, _04146_);
  nand (_04152_, _04151_, _00560_);
  nor (_04153_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_04154_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1]);
  nor (_04155_, _04154_, _04153_);
  nand (_04156_, _04155_, _00227_);
  nand (_04157_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nand (_04158_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1]);
  nand (_04159_, _04158_, _04157_);
  nand (_04160_, _04159_, _01417_);
  nand (_04161_, _04160_, _04156_);
  nand (_04162_, _04161_, _00561_);
  nand (_04163_, _04162_, _04152_);
  nand (_04165_, _04163_, _00465_);
  nand (_04166_, _04165_, _04140_);
  nand (_04167_, _04166_, _00248_);
  nand (_04168_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1]);
  nand (_04169_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  nand (_04171_, _04169_, _04168_);
  nand (_04172_, _04171_, _01417_);
  nand (_04173_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  nand (_04174_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1]);
  nand (_04175_, _04174_, _04173_);
  nand (_04176_, _04175_, _00227_);
  nand (_04177_, _04176_, _04172_);
  nand (_04178_, _04177_, _00560_);
  nand (_04179_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  nand (_04180_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  nand (_04181_, _04180_, _04179_);
  nand (_04183_, _04181_, _01417_);
  nand (_04184_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1]);
  nand (_04185_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  nand (_04186_, _04185_, _04184_);
  nand (_04188_, _04186_, _00227_);
  nand (_04189_, _04188_, _04183_);
  nand (_04190_, _04189_, _00561_);
  nand (_04191_, _04190_, _04178_);
  nand (_04192_, _04191_, _00466_);
  not (_04194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  nand (_04195_, _00650_, _04194_);
  nor (_04196_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  nor (_04197_, _04196_, _00227_);
  nand (_04199_, _04197_, _04195_);
  nor (_04200_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  nor (_04201_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1]);
  nor (_04202_, _04201_, _04200_);
  nand (_04203_, _04202_, _00227_);
  nand (_04204_, _04203_, _04199_);
  nand (_04205_, _04204_, _00560_);
  nor (_04206_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1]);
  nor (_04207_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1]);
  nor (_04208_, _04207_, _04206_);
  nand (_04209_, _04208_, _01417_);
  nor (_04210_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1]);
  nor (_04211_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  nor (_04212_, _04211_, _04210_);
  nand (_04213_, _04212_, _00227_);
  nand (_04214_, _04213_, _04209_);
  nand (_04215_, _04214_, _00561_);
  nand (_04216_, _04215_, _04205_);
  nand (_04218_, _04216_, _00465_);
  nand (_04219_, _04218_, _04192_);
  nand (_04220_, _04219_, _00247_);
  nand (_04221_, _04220_, _04167_);
  nand (_04222_, _04221_, _00319_);
  nand (_04224_, _04222_, _04114_);
  nor (_04225_, _04224_, _00386_);
  nand (_04226_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1]);
  nand (_04228_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1]);
  nand (_04229_, _04228_, _04226_);
  nand (_04230_, _04229_, _01417_);
  nand (_04231_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1]);
  nand (_04232_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1]);
  nand (_04233_, _04232_, _04231_);
  nand (_04234_, _04233_, _00227_);
  nand (_04235_, _04234_, _04230_);
  nand (_04237_, _04235_, _00560_);
  nand (_04238_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1]);
  nand (_04239_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1]);
  nand (_04240_, _04239_, _04238_);
  nand (_04241_, _04240_, _01417_);
  nand (_04242_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1]);
  nand (_04243_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1]);
  nand (_04245_, _04243_, _04242_);
  nand (_04246_, _04245_, _00227_);
  nand (_04247_, _04246_, _04241_);
  nand (_04248_, _04247_, _00561_);
  nand (_04249_, _04248_, _04237_);
  nand (_04250_, _04249_, _00466_);
  nor (_04251_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1]);
  nor (_04252_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1]);
  nor (_04253_, _04252_, _04251_);
  nand (_04254_, _04253_, _01417_);
  nor (_04255_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  nor (_04256_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1]);
  nor (_04257_, _04256_, _04255_);
  nand (_04258_, _04257_, _00227_);
  nand (_04259_, _04258_, _04254_);
  nand (_04260_, _04259_, _00560_);
  not (_04261_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  nand (_04262_, _00650_, _04261_);
  nor (_04263_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  nor (_04264_, _04263_, _00227_);
  nand (_04265_, _04264_, _04262_);
  nor (_04266_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  nor (_04267_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  nor (_04268_, _04267_, _04266_);
  nand (_04269_, _04268_, _00227_);
  nand (_04270_, _04269_, _04265_);
  nand (_04271_, _04270_, _00561_);
  nand (_04272_, _04271_, _04260_);
  nand (_04273_, _04272_, _00465_);
  nand (_04274_, _04273_, _04250_);
  nand (_04275_, _04274_, _00248_);
  nand (_04277_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  nand (_04278_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1]);
  nand (_04279_, _04278_, _04277_);
  nand (_04281_, _04279_, _01417_);
  nand (_04282_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1]);
  nand (_04283_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1]);
  nand (_04284_, _04283_, _04282_);
  nand (_04285_, _04284_, _00227_);
  nand (_04286_, _04285_, _04281_);
  nand (_04287_, _04286_, _00560_);
  nand (_04288_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1]);
  nand (_04289_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1]);
  nand (_04290_, _04289_, _04288_);
  nand (_04292_, _04290_, _01417_);
  nand (_04293_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1]);
  nand (_04294_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1]);
  nand (_04295_, _04294_, _04293_);
  nand (_04296_, _04295_, _00227_);
  nand (_04297_, _04296_, _04292_);
  nand (_04299_, _04297_, _00561_);
  nand (_04300_, _04299_, _04287_);
  nand (_04301_, _04300_, _00466_);
  not (_04302_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1]);
  nand (_04303_, _00650_, _04302_);
  nor (_04304_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1]);
  nor (_04305_, _04304_, _00227_);
  nand (_04306_, _04305_, _04303_);
  nor (_04307_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1]);
  nor (_04308_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1]);
  nor (_04309_, _04308_, _04307_);
  nand (_04310_, _04309_, _00227_);
  nand (_04311_, _04310_, _04306_);
  nand (_04312_, _04311_, _00560_);
  nor (_04314_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1]);
  nor (_04315_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1]);
  nor (_04316_, _04315_, _04314_);
  nand (_04317_, _04316_, _01417_);
  nor (_04318_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1]);
  nor (_04319_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1]);
  nor (_04320_, _04319_, _04318_);
  nand (_04321_, _04320_, _00227_);
  nand (_04323_, _04321_, _04317_);
  nand (_04324_, _04323_, _00561_);
  nand (_04325_, _04324_, _04312_);
  nand (_04326_, _04325_, _00465_);
  nand (_04327_, _04326_, _04301_);
  nand (_04328_, _04327_, _00247_);
  nand (_04329_, _04328_, _04275_);
  nand (_04330_, _04329_, _00319_);
  nand (_04331_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1]);
  nand (_04332_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1]);
  nand (_04333_, _04332_, _04331_);
  nand (_04334_, _04333_, _00227_);
  nand (_04335_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1]);
  nand (_04336_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1]);
  nand (_04337_, _04336_, _04335_);
  nand (_04338_, _04337_, _01417_);
  nand (_04339_, _04338_, _04334_);
  nand (_04340_, _04339_, _00560_);
  nand (_04343_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1]);
  nand (_04344_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1]);
  nand (_04345_, _04344_, _04343_);
  nand (_04346_, _04345_, _00227_);
  nand (_04347_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1]);
  nand (_04349_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1]);
  nand (_04350_, _04349_, _04347_);
  nand (_04351_, _04350_, _01417_);
  nand (_04352_, _04351_, _04346_);
  nand (_04353_, _04352_, _00561_);
  nand (_04354_, _04353_, _04340_);
  nand (_04355_, _04354_, _00466_);
  nand (_04356_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1]);
  nand (_04358_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1]);
  nand (_04359_, _04358_, _04356_);
  nand (_04360_, _04359_, _01417_);
  nor (_04361_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1]);
  nor (_04362_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  nor (_04363_, _04362_, _04361_);
  nand (_04364_, _04363_, _00227_);
  nand (_04365_, _04364_, _04360_);
  nand (_04366_, _04365_, _00560_);
  nand (_04367_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  nand (_04368_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  nand (_04369_, _04368_, _04367_);
  nand (_04370_, _04369_, _01417_);
  nor (_04372_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1]);
  nor (_04373_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  nor (_04374_, _04373_, _04372_);
  nand (_04375_, _04374_, _00227_);
  nand (_04377_, _04375_, _04370_);
  nand (_04378_, _04377_, _00561_);
  nand (_04379_, _04378_, _04366_);
  nand (_04380_, _04379_, _00465_);
  nand (_04381_, _04380_, _04355_);
  nand (_04382_, _04381_, _00248_);
  nand (_04383_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1]);
  nand (_04384_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1]);
  nand (_04385_, _04384_, _04383_);
  nand (_04386_, _04385_, _01417_);
  nand (_04387_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  nand (_04388_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  nand (_04389_, _04388_, _04387_);
  nand (_04390_, _04389_, _00227_);
  nand (_04391_, _04390_, _04386_);
  nand (_04392_, _04391_, _00560_);
  nand (_04393_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1]);
  nand (_04394_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1]);
  nand (_04395_, _04394_, _04393_);
  nand (_04396_, _04395_, _01417_);
  nand (_04398_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1]);
  nand (_04400_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1]);
  nand (_04401_, _04400_, _04398_);
  nand (_04402_, _04401_, _00227_);
  nand (_04403_, _04402_, _04396_);
  nand (_04404_, _04403_, _00561_);
  nand (_04405_, _04404_, _04392_);
  nand (_04406_, _04405_, _00466_);
  nor (_04408_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1]);
  nor (_04409_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  nor (_04411_, _04409_, _04408_);
  nand (_04412_, _04411_, _01417_);
  nor (_04413_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1]);
  nor (_04414_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  nor (_04415_, _04414_, _04413_);
  nand (_04417_, _04415_, _00227_);
  nand (_04418_, _04417_, _04412_);
  nand (_04419_, _04418_, _00560_);
  nor (_04420_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1]);
  nor (_04421_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  nor (_04423_, _04421_, _04420_);
  nor (_04424_, _04423_, _00227_);
  nor (_04425_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  nor (_04426_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1]);
  nor (_04427_, _04426_, _04425_);
  nor (_04428_, _04427_, _01417_);
  nor (_04429_, _04428_, _04424_);
  nand (_04431_, _04429_, _00561_);
  nand (_04432_, _04431_, _04419_);
  nand (_04433_, _04432_, _00465_);
  nand (_04434_, _04433_, _04406_);
  nand (_04435_, _04434_, _00247_);
  nand (_04436_, _04435_, _04382_);
  nand (_04437_, _04436_, _00320_);
  nand (_04438_, _04437_, _04330_);
  nor (_04439_, _04438_, _01629_);
  nor (_04440_, _04439_, _04225_);
  nor (_04441_, _04440_, _00156_);
  nand (_04442_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  nand (_04444_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  nand (_04445_, _04444_, _04442_);
  nand (_04446_, _04445_, _01417_);
  nand (_04447_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1]);
  nand (_04448_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1]);
  nand (_04450_, _04448_, _04447_);
  nand (_04451_, _04450_, _00227_);
  nand (_04452_, _04451_, _04446_);
  nand (_04453_, _04452_, _00560_);
  nand (_04454_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1]);
  nand (_04455_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  nand (_04456_, _04455_, _04454_);
  nand (_04457_, _04456_, _01417_);
  nand (_04458_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1]);
  nand (_04459_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  nand (_04460_, _04459_, _04458_);
  nand (_04461_, _04460_, _00227_);
  nand (_04463_, _04461_, _04457_);
  nand (_04464_, _04463_, _00561_);
  nand (_04465_, _04464_, _04453_);
  nand (_04466_, _04465_, _00466_);
  nor (_04468_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1]);
  nor (_04469_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  nor (_04470_, _04469_, _04468_);
  nand (_04472_, _04470_, _01417_);
  nor (_04473_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  nor (_04474_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1]);
  nor (_04475_, _04474_, _04473_);
  nand (_04476_, _04475_, _00227_);
  nand (_04477_, _04476_, _04472_);
  nand (_04478_, _04477_, _00560_);
  nor (_04479_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1]);
  nor (_04480_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1]);
  nor (_04481_, _04480_, _04479_);
  nand (_04482_, _04481_, _01417_);
  nor (_04483_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  nor (_04484_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1]);
  nor (_04485_, _04484_, _04483_);
  nand (_04486_, _04485_, _00227_);
  nand (_04487_, _04486_, _04482_);
  nand (_04488_, _04487_, _00561_);
  nand (_04490_, _04488_, _04478_);
  nand (_04491_, _04490_, _00465_);
  nand (_04492_, _04491_, _04466_);
  nand (_04493_, _04492_, _00247_);
  nand (_04494_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1]);
  nand (_04495_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1]);
  nand (_04497_, _04495_, _04494_);
  nand (_04498_, _04497_, _01417_);
  nand (_04500_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1]);
  nand (_04501_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  nand (_04503_, _04501_, _04500_);
  nand (_04504_, _04503_, _00227_);
  nand (_04505_, _04504_, _04498_);
  nand (_04506_, _04505_, _00560_);
  nand (_04507_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1]);
  nand (_04508_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1]);
  nand (_04509_, _04508_, _04507_);
  nand (_04510_, _04509_, _01417_);
  nand (_04511_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  nand (_04513_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1]);
  nand (_04514_, _04513_, _04511_);
  nand (_04515_, _04514_, _00227_);
  nand (_04516_, _04515_, _04510_);
  nand (_04517_, _04516_, _00561_);
  nand (_04518_, _04517_, _04506_);
  nand (_04519_, _04518_, _00466_);
  nor (_04520_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1]);
  nor (_04521_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1]);
  nor (_04522_, _04521_, _04520_);
  nand (_04523_, _04522_, _00227_);
  nand (_04524_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1]);
  nand (_04525_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1]);
  nand (_04526_, _04525_, _04524_);
  nand (_04527_, _04526_, _01417_);
  nand (_04528_, _04527_, _04523_);
  nand (_04529_, _04528_, _00560_);
  nor (_04530_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1]);
  nor (_04531_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1]);
  nor (_04532_, _04531_, _04530_);
  nand (_04533_, _04532_, _00227_);
  nand (_04535_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1]);
  nand (_04536_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1]);
  nand (_04538_, _04536_, _04535_);
  nand (_04539_, _04538_, _01417_);
  nand (_04540_, _04539_, _04533_);
  nand (_04542_, _04540_, _00561_);
  nand (_04543_, _04542_, _04529_);
  nand (_04545_, _04543_, _00465_);
  nand (_04546_, _04545_, _04519_);
  nand (_04547_, _04546_, _00248_);
  nand (_04549_, _04547_, _04493_);
  nand (_04550_, _04549_, _00320_);
  nand (_04551_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1]);
  nand (_04552_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1]);
  nand (_04553_, _04552_, _04551_);
  nand (_04554_, _04553_, _01417_);
  nand (_04555_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  nand (_04556_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  nand (_04557_, _04556_, _04555_);
  nand (_04558_, _04557_, _00227_);
  nand (_04559_, _04558_, _04554_);
  nand (_04560_, _04559_, _00560_);
  nand (_04561_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  nand (_04562_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1]);
  nand (_04563_, _04562_, _04561_);
  nand (_04564_, _04563_, _01417_);
  nand (_04565_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  nand (_04566_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  nand (_04567_, _04566_, _04565_);
  nand (_04568_, _04567_, _00227_);
  nand (_04570_, _04568_, _04564_);
  nand (_04571_, _04570_, _00561_);
  nand (_04572_, _04571_, _04560_);
  nand (_04573_, _04572_, _00466_);
  nor (_04574_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  nor (_04575_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  nor (_04576_, _04575_, _04574_);
  nand (_04577_, _04576_, _00227_);
  nand (_04578_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  nand (_04579_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  nand (_04580_, _04579_, _04578_);
  nand (_04581_, _04580_, _01417_);
  nand (_04582_, _04581_, _04577_);
  nand (_04583_, _04582_, _00560_);
  nor (_04584_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  nor (_04585_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  nor (_04586_, _04585_, _04584_);
  nand (_04587_, _04586_, _00227_);
  nand (_04588_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  nand (_04589_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1]);
  nand (_04590_, _04589_, _04588_);
  nand (_04591_, _04590_, _01417_);
  nand (_04592_, _04591_, _04587_);
  nand (_04594_, _04592_, _00561_);
  nand (_04595_, _04594_, _04583_);
  nand (_04596_, _04595_, _00465_);
  nand (_04597_, _04596_, _04573_);
  nand (_04598_, _04597_, _00248_);
  nand (_04599_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1]);
  nand (_04600_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1]);
  nand (_04601_, _04600_, _04599_);
  nand (_04602_, _04601_, _01417_);
  nand (_04603_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1]);
  nand (_04604_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1]);
  nand (_04605_, _04604_, _04603_);
  nand (_04606_, _04605_, _00227_);
  nand (_04607_, _04606_, _04602_);
  nand (_04608_, _04607_, _00560_);
  nand (_04609_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  nand (_04610_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1]);
  nand (_04611_, _04610_, _04609_);
  nand (_04613_, _04611_, _01417_);
  nand (_04614_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1]);
  nand (_04615_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1]);
  nand (_04617_, _04615_, _04614_);
  nand (_04618_, _04617_, _00227_);
  nand (_04619_, _04618_, _04613_);
  nand (_04620_, _04619_, _00561_);
  nand (_04621_, _04620_, _04608_);
  nand (_04622_, _04621_, _00466_);
  nor (_04623_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1]);
  nor (_04624_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1]);
  nor (_04625_, _04624_, _04623_);
  nand (_04626_, _04625_, _01417_);
  nor (_04627_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1]);
  nor (_04628_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1]);
  nor (_04630_, _04628_, _04627_);
  nand (_04631_, _04630_, _00227_);
  nand (_04632_, _04631_, _04626_);
  nand (_04634_, _04632_, _00560_);
  nor (_04636_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1]);
  nor (_04637_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1]);
  nor (_04638_, _04637_, _04636_);
  nand (_04639_, _04638_, _01417_);
  nor (_04640_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1]);
  nor (_04641_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1]);
  nor (_04642_, _04641_, _04640_);
  nand (_04643_, _04642_, _00227_);
  nand (_04644_, _04643_, _04639_);
  nand (_04645_, _04644_, _00561_);
  nand (_04646_, _04645_, _04634_);
  nand (_04647_, _04646_, _00465_);
  nand (_04649_, _04647_, _04622_);
  nand (_04650_, _04649_, _00247_);
  nand (_04651_, _04650_, _04598_);
  nand (_04652_, _04651_, _00319_);
  nand (_04653_, _04652_, _04550_);
  nor (_04654_, _04653_, _00386_);
  nand (_04655_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  nand (_04656_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  nand (_04657_, _04656_, _04655_);
  nand (_04658_, _04657_, _01417_);
  nand (_04659_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  nand (_04660_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  nand (_04661_, _04660_, _04659_);
  nand (_04662_, _04661_, _00227_);
  nand (_04663_, _04662_, _04658_);
  nand (_04664_, _04663_, _00560_);
  nand (_04665_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  nand (_04666_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  nand (_04667_, _04666_, _04665_);
  nand (_04668_, _04667_, _01417_);
  nand (_04669_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1]);
  nand (_04670_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  nand (_04671_, _04670_, _04669_);
  nand (_04672_, _04671_, _00227_);
  nand (_04673_, _04672_, _04668_);
  nand (_04674_, _04673_, _00561_);
  nand (_04675_, _04674_, _04664_);
  nand (_04676_, _04675_, _00466_);
  nor (_04677_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  nor (_04678_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  nor (_04679_, _04678_, _04677_);
  nand (_04680_, _04679_, _00227_);
  nand (_04682_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  nand (_04683_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  nand (_04684_, _04683_, _04682_);
  nand (_04685_, _04684_, _01417_);
  nand (_04686_, _04685_, _04680_);
  nand (_04688_, _04686_, _00560_);
  nor (_04690_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  nor (_04691_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  nor (_04692_, _04691_, _04690_);
  nand (_04694_, _04692_, _00227_);
  nand (_04695_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  nand (_04696_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  nand (_04698_, _04696_, _04695_);
  nand (_04699_, _04698_, _01417_);
  nand (_04700_, _04699_, _04694_);
  nand (_04702_, _04700_, _00561_);
  nand (_04703_, _04702_, _04688_);
  nand (_04704_, _04703_, _00465_);
  nand (_04705_, _04704_, _04676_);
  nand (_04706_, _04705_, _00248_);
  nand (_04707_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  nand (_04708_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  nand (_04709_, _04708_, _04707_);
  nand (_04710_, _04709_, _01417_);
  nand (_04711_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  nand (_04712_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  nand (_04713_, _04712_, _04711_);
  nand (_04714_, _04713_, _00227_);
  nand (_04715_, _04714_, _04710_);
  nand (_04716_, _04715_, _00560_);
  nand (_04717_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  nand (_04718_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  nand (_04720_, _04718_, _04717_);
  nand (_04722_, _04720_, _01417_);
  nand (_04723_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  nand (_04724_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  nand (_04726_, _04724_, _04723_);
  nand (_04727_, _04726_, _00227_);
  nand (_04728_, _04727_, _04722_);
  nand (_04729_, _04728_, _00561_);
  nand (_04730_, _04729_, _04716_);
  nand (_04732_, _04730_, _00466_);
  nor (_04733_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  nor (_04734_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  nor (_04735_, _04734_, _04733_);
  nand (_04736_, _04735_, _01417_);
  nor (_04737_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  nor (_04738_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  nor (_04739_, _04738_, _04737_);
  nand (_04740_, _04739_, _00227_);
  nand (_04741_, _04740_, _04736_);
  nand (_04742_, _04741_, _00560_);
  nor (_04743_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  nor (_04744_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  nor (_04745_, _04744_, _04743_);
  nand (_04746_, _04745_, _01417_);
  nor (_04748_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  nor (_04749_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  nor (_04750_, _04749_, _04748_);
  nand (_04752_, _04750_, _00227_);
  nand (_04754_, _04752_, _04746_);
  nand (_04755_, _04754_, _00561_);
  nand (_04756_, _04755_, _04742_);
  nand (_04757_, _04756_, _00465_);
  nand (_04759_, _04757_, _04732_);
  nand (_04760_, _04759_, _00247_);
  nand (_04761_, _04760_, _04706_);
  nand (_04762_, _04761_, _00320_);
  nor (_04763_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1]);
  nor (_04764_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  nor (_04765_, _04764_, _04763_);
  nand (_04766_, _04765_, _01417_);
  nor (_04767_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1]);
  nor (_04768_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  nor (_04769_, _04768_, _04767_);
  nand (_04770_, _04769_, _00227_);
  nand (_04772_, _04770_, _04766_);
  nand (_04773_, _04772_, _00561_);
  nor (_04774_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1]);
  nor (_04775_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1]);
  nor (_04776_, _04775_, _04774_);
  nand (_04777_, _04776_, _01417_);
  nor (_04778_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  nor (_04779_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  nor (_04780_, _04779_, _04778_);
  nand (_04781_, _04780_, _00227_);
  nand (_04782_, _04781_, _04777_);
  nand (_04783_, _04782_, _00560_);
  nand (_04784_, _04783_, _04773_);
  nand (_04785_, _04784_, _00465_);
  nand (_04786_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1]);
  nand (_04787_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1]);
  nand (_04788_, _04787_, _04786_);
  nand (_04789_, _04788_, _01417_);
  nand (_04790_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  nand (_04791_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1]);
  nand (_04793_, _04791_, _04790_);
  nand (_04795_, _04793_, _00227_);
  nand (_04796_, _04795_, _04789_);
  nand (_04797_, _04796_, _00561_);
  nand (_04798_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  nand (_04799_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  nand (_04800_, _04799_, _04798_);
  nand (_04801_, _04800_, _01417_);
  nand (_04802_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1]);
  nand (_04803_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  nand (_04804_, _04803_, _04802_);
  nand (_04805_, _04804_, _00227_);
  nand (_04806_, _04805_, _04801_);
  nand (_04807_, _04806_, _00560_);
  nand (_04808_, _04807_, _04797_);
  nand (_04810_, _04808_, _00466_);
  nand (_04811_, _04810_, _04785_);
  nand (_04812_, _04811_, _00247_);
  nor (_04814_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  nor (_04815_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  nor (_04817_, _04815_, _04814_);
  nand (_04818_, _04817_, _00227_);
  nand (_04819_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  nand (_04820_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  nand (_04821_, _04820_, _04819_);
  nand (_04822_, _04821_, _01417_);
  nand (_04823_, _04822_, _04818_);
  nand (_04824_, _04823_, _00561_);
  nor (_04825_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  nor (_04826_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1]);
  nor (_04827_, _04826_, _04825_);
  nand (_04828_, _04827_, _00227_);
  nand (_04829_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1]);
  nand (_04830_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  nand (_04831_, _04830_, _04829_);
  nand (_04832_, _04831_, _01417_);
  nand (_04833_, _04832_, _04828_);
  nand (_04834_, _04833_, _00560_);
  nand (_04835_, _04834_, _04824_);
  nand (_04836_, _04835_, _00465_);
  nand (_04838_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  nand (_04839_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  nand (_04840_, _04839_, _04838_);
  nand (_04841_, _04840_, _01417_);
  nand (_04842_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1]);
  nand (_04843_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  nand (_04844_, _04843_, _04842_);
  nand (_04846_, _04844_, _00227_);
  nand (_04847_, _04846_, _04841_);
  nand (_04848_, _04847_, _00561_);
  nand (_04850_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  nand (_04851_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  nand (_04852_, _04851_, _04850_);
  nand (_04853_, _04852_, _01417_);
  nand (_04854_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  nand (_04855_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  nand (_04856_, _04855_, _04854_);
  nand (_04857_, _04856_, _00227_);
  nand (_04858_, _04857_, _04853_);
  nand (_04859_, _04858_, _00560_);
  nand (_04860_, _04859_, _04848_);
  nand (_04861_, _04860_, _00466_);
  nand (_04862_, _04861_, _04836_);
  nand (_04863_, _04862_, _00248_);
  nand (_04864_, _04863_, _04812_);
  nand (_04866_, _04864_, _00319_);
  nand (_04867_, _04866_, _04762_);
  nor (_04868_, _04867_, _01629_);
  nor (_04869_, _04868_, _04654_);
  nor (_04870_, _04869_, _00556_);
  nor (_04872_, _04870_, _04441_);
  nor (_04873_, _04872_, _01416_);
  not (_04874_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  nand (_04875_, _01416_, _04874_);
  nand (_04876_, _04875_, _23493_);
  nor (_25454_[1], _04876_, _04873_);
  nor (_04877_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand (_04878_, _03721_, _00006_);
  nand (_04879_, _04878_, _23493_);
  nor (_21841_, _04879_, _04877_);
  nand (_04880_, _02683_, _02635_);
  nor (_04881_, _03732_, _02635_);
  nor (_04882_, _04881_, _02658_);
  nand (_04883_, _04882_, _04880_);
  nor (_04884_, _02691_, _02635_);
  nand (_04885_, _02691_, _02635_);
  nand (_04886_, _04885_, _02620_);
  nor (_04887_, _04886_, _04884_);
  nor (_04888_, _02708_, _02635_);
  nand (_04889_, _02708_, _02635_);
  nand (_04891_, _04889_, _02705_);
  nor (_04892_, _04891_, _04888_);
  nor (_04893_, _04892_, _04887_);
  nand (_04894_, _04893_, _04883_);
  nor (_04895_, _04894_, _02612_);
  nand (_04896_, _02612_, _00029_);
  nand (_04897_, _04896_, _02626_);
  nor (_04898_, _04897_, _04895_);
  nor (_04899_, _02626_, _02635_);
  nor (_04900_, _04899_, _04898_);
  nor (_21845_, _04900_, rst);
  nor (_04901_, _02681_, _02612_);
  nor (_04902_, _04901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  not (_04903_, _02670_);
  nand (_04904_, _02656_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_04905_, _04904_, _03730_);
  nand (_04906_, _04905_, _04903_);
  nand (_04907_, _04906_, _03830_);
  nor (_04908_, _04907_, _02612_);
  nor (_04909_, _04908_, _04902_);
  nor (_04910_, _04909_, _02625_);
  nand (_04911_, _02625_, _00029_);
  nand (_04912_, _04911_, _23493_);
  nor (_21848_, _04912_, _04910_);
  nor (_04913_, _03677_, _03632_);
  nand (_04914_, _04913_, _03932_);
  nand (_04915_, _04914_, _03633_);
  nor (_04916_, _04914_, _03633_);
  nor (_04917_, _04916_, _03668_);
  nand (_04918_, _04917_, _04915_);
  not (_04919_, _04913_);
  nand (_04920_, _04919_, _03633_);
  nand (_04921_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_04922_, _03677_, _03636_);
  not (_04923_, _04922_);
  nand (_04924_, _04923_, _03673_);
  nand (_04925_, _04924_, _04921_);
  nand (_04926_, _04925_, _04920_);
  nand (_04927_, _04926_, _04918_);
  nand (_04928_, _04927_, _03688_);
  nand (_04929_, _03694_, ABINPUT[4]);
  nand (_04930_, _04929_, _04928_);
  nor (_04931_, _04930_, _03702_);
  nand (_04933_, _03702_, _03633_);
  nand (_04934_, _04933_, _23493_);
  nor (_21851_, _04934_, _04931_);
  not (_04935_, _03919_);
  nor (_04936_, _03958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nand (_04937_, _03958_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  not (_04938_, _04937_);
  nor (_04939_, _04938_, _04936_);
  nor (_04940_, _04939_, _04935_);
  nor (_04941_, _03919_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_04942_, _04941_, _04940_);
  not (_04943_, _03940_);
  nor (_04944_, _04943_, _03633_);
  nand (_04945_, _04944_, _03688_);
  nand (_04946_, _04945_, _03909_);
  nor (_04947_, _04946_, _04942_);
  nand (_04948_, _03702_, _00006_);
  nand (_04949_, _04948_, _23493_);
  nor (_21854_, _04949_, _04947_);
  nor (_04950_, _21567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1]);
  nor (_04951_, _21569_, _21474_);
  nor (_21886_, _04951_, _04950_);
  nor (_04952_, _22551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1]);
  nor (_04953_, _22555_, _21474_);
  nor (_21888_, _04953_, _04952_);
  nor (_04954_, _22551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  nor (_04955_, _22555_, _21554_);
  nor (_21890_, _04955_, _04954_);
  nor (_04957_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  nand (_04958_, _23553_, _24175_);
  nand (_04959_, _04958_, _23493_);
  nor (_21896_, _04959_, _04957_);
  nor (_04960_, _21567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  nor (_04961_, _21569_, _21526_);
  nor (_21898_, _04961_, _04960_);
  nor (_04962_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  nand (_04963_, _23553_, _00290_);
  nand (_04964_, _04963_, _23493_);
  nor (_21908_, _04964_, _04962_);
  nor (_04965_, _21567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  nor (_04966_, _21569_, _21414_);
  nor (_21909_, _04966_, _04965_);
  nand (_04967_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nand (_04968_, _01142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nand (_04969_, _04968_, _04967_);
  nor (_04970_, _04969_, _01130_);
  nor (_04971_, _01059_, _00114_);
  nor (_04972_, _01055_, _00129_);
  nor (_04973_, _04972_, _04971_);
  nand (_04974_, _04973_, _01130_);
  nand (_04975_, _04974_, _23493_);
  nor (_21912_, _04975_, _04970_);
  nor (_04976_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  nand (_04977_, _23553_, _00370_);
  nand (_04978_, _04977_, _23493_);
  nor (_21916_, _04978_, _04976_);
  nor (_04980_, _24877_, _21268_);
  not (_04981_, _04980_);
  nor (_04982_, _04981_, _21774_);
  not (_04983_, _04982_);
  nor (_04985_, _04983_, _24858_);
  nand (_04986_, _04985_, ABINPUT[3]);
  not (_04987_, _04985_);
  nand (_04988_, _04987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nand (_04989_, _04988_, _04986_);
  nand (_04990_, _04989_, _24861_);
  nor (_04991_, _24858_, _21507_);
  nand (_04992_, _04991_, _04982_);
  nand (_04994_, _04992_, _04988_);
  nand (_04995_, _04994_, _00914_);
  nand (_04996_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nand (_04997_, _04996_, _04995_);
  nor (_04998_, _04997_, rst);
  nand (_21918_, _04998_, _04990_);
  nor (_04999_, _24129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  nor (_05000_, _24131_, _21504_);
  nor (_21921_, _05000_, _04999_);
  nor (_05001_, _01127_, _24903_);
  nand (_05002_, _05001_, ABINPUT[3]);
  not (_05003_, _05001_);
  nand (_05004_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nand (_05005_, _05004_, _05002_);
  nand (_05006_, _05005_, _24861_);
  not (_05007_, _05004_);
  nor (_05008_, _05003_, _21507_);
  nor (_05009_, _05008_, _05007_);
  nor (_05010_, _05009_, _00915_);
  nand (_05011_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nand (_05012_, _05011_, _23493_);
  nor (_05013_, _05012_, _05010_);
  nand (_21925_, _05013_, _05006_);
  nor (_05014_, _00018_, _24877_);
  not (_05015_, _01010_);
  nand (_05016_, _05015_, _05014_);
  nand (_05017_, _05016_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_05018_, _01010_, _21507_);
  nand (_05019_, _05018_, _05014_);
  nand (_05020_, _05019_, _05017_);
  nand (_05021_, _05020_, _00914_);
  not (_05023_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nor (_05024_, _00018_, _24903_);
  nor (_05025_, _05024_, _05023_);
  not (_05026_, _05024_);
  nor (_05027_, _05026_, _00129_);
  nor (_05028_, _05027_, _05025_);
  nor (_05029_, _05028_, _00010_);
  nand (_05030_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nand (_05031_, _05030_, _23493_);
  nor (_05032_, _05031_, _05029_);
  nand (_21927_, _05032_, _05021_);
  nor (_05033_, _21873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  nor (_05034_, _21875_, _21414_);
  nor (_21936_, _05034_, _05033_);
  nor (_05035_, _21567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7]);
  nor (_05037_, _21626_, _21569_);
  nor (_21941_, _05037_, _05035_);
  nand (_05038_, _04985_, ABINPUT[4]);
  nand (_05040_, _04987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nand (_05041_, _05040_, _05038_);
  nand (_05042_, _05041_, _24861_);
  nand (_05043_, _04982_, _00011_);
  nand (_05044_, _05043_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_05045_, _00020_, _21507_);
  nand (_05046_, _05045_, _04982_);
  nand (_05047_, _05046_, _05044_);
  nand (_05048_, _05047_, _00914_);
  nand (_05049_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nand (_05050_, _05049_, _05048_);
  nor (_05051_, _05050_, rst);
  nand (_21950_, _05051_, _05042_);
  nor (_05052_, _01025_, _21351_);
  nand (_05053_, _05052_, _05014_);
  nand (_05054_, _05053_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  not (_05055_, _05052_);
  nor (_05056_, _05055_, _21507_);
  nand (_05057_, _05056_, _05014_);
  nand (_05058_, _05057_, _05054_);
  nand (_05059_, _05058_, _00914_);
  not (_05060_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nor (_05061_, _05024_, _05060_);
  nor (_05062_, _05026_, _00114_);
  nor (_05063_, _05062_, _05061_);
  nor (_05064_, _05063_, _00010_);
  nand (_05065_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nand (_05066_, _05065_, _23493_);
  nor (_05067_, _05066_, _05064_);
  nand (_21953_, _05067_, _05059_);
  nor (_05068_, _24129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5]);
  nor (_05069_, _24131_, _21451_);
  nor (_25382_, _05069_, _05068_);
  nor (_05070_, _23799_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  nor (_05071_, _23801_, _21586_);
  nor (_22089_, _05071_, _05070_);
  nand (_05072_, _05024_, _24900_);
  nor (_05073_, _05024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nor (_05074_, _05073_, _00010_);
  nand (_05075_, _05074_, _05072_);
  not (_05076_, _05014_);
  nor (_05077_, _01001_, _05076_);
  nor (_05078_, _05077_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand (_05079_, _05077_, _21507_);
  nand (_05080_, _05079_, _00914_);
  nor (_05081_, _05080_, _05078_);
  nand (_05082_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand (_05083_, _05082_, _23493_);
  nor (_05084_, _05083_, _05081_);
  nand (_22093_, _05084_, _05075_);
  nand (_05085_, _05026_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nand (_05086_, _05024_, ABINPUT[0]);
  nand (_05087_, _05086_, _05085_);
  nand (_05088_, _05087_, _00914_);
  not (_05090_, _05085_);
  nor (_05091_, _05026_, _00029_);
  nor (_05092_, _05091_, _05090_);
  nor (_05093_, _05092_, _00010_);
  nand (_05094_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nand (_05095_, _05094_, _23493_);
  nor (_05096_, _05095_, _05093_);
  nand (_22097_, _05096_, _05088_);
  nor (_05097_, _01127_, _24877_);
  nand (_05098_, _05097_, _00908_);
  nand (_05099_, _05098_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nand (_05100_, _05097_, _00931_);
  nand (_05101_, _05100_, _05099_);
  nand (_05102_, _05101_, _00914_);
  nor (_05103_, _05003_, _24867_);
  not (_05104_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_05105_, _05001_, _05104_);
  nor (_05107_, _05105_, _05103_);
  nor (_05108_, _05107_, _00010_);
  nand (_05109_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nand (_05110_, _05109_, _23493_);
  nor (_05111_, _05110_, _05108_);
  nand (_22104_, _05111_, _05102_);
  nor (_05112_, _24877_, _24897_);
  not (_05113_, _05112_);
  nor (_05114_, _05113_, _21774_);
  not (_05115_, _05114_);
  nor (_05116_, _05115_, _24858_);
  nand (_05117_, _05116_, ABINPUT[9]);
  not (_05118_, _05116_);
  nand (_05119_, _05118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nand (_05120_, _05119_, _05117_);
  nand (_05121_, _05120_, _24861_);
  not (_05122_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nor (_05123_, _05055_, _05115_);
  nor (_05124_, _05123_, _05122_);
  not (_05125_, _05056_);
  nor (_05126_, _05125_, _05115_);
  nor (_05127_, _05126_, _05124_);
  nor (_05128_, _05127_, _00915_);
  nand (_05129_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nand (_05130_, _05129_, _23493_);
  nor (_05131_, _05130_, _05128_);
  nand (_22107_, _05131_, _05121_);
  nand (_05132_, _05116_, ABINPUT[4]);
  nand (_05133_, _05118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nand (_05134_, _05133_, _05132_);
  nand (_05135_, _05134_, _24861_);
  not (_05136_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_05137_, _05115_, _00020_);
  nor (_05138_, _05137_, _05136_);
  not (_05140_, _05045_);
  nor (_05142_, _05140_, _05115_);
  nor (_05143_, _05142_, _05138_);
  nor (_05144_, _05143_, _00915_);
  nand (_05145_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nand (_05146_, _05145_, _23493_);
  nor (_05147_, _05146_, _05144_);
  nand (_22110_, _05147_, _05135_);
  nor (_05148_, _21850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  nor (_05150_, _21853_, _21554_);
  nor (_22112_, _05150_, _05148_);
  nand (_05151_, _04985_, ABINPUT[8]);
  nand (_05152_, _04987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand (_05153_, _05152_, _05151_);
  nand (_05154_, _05153_, _24861_);
  nand (_05156_, _04982_, _05015_);
  nand (_05158_, _05156_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand (_05159_, _05018_, _04982_);
  nand (_05160_, _05159_, _05158_);
  nand (_05161_, _05160_, _00914_);
  nand (_05162_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand (_05164_, _05162_, _05161_);
  nor (_05166_, _05164_, rst);
  nand (_22120_, _05166_, _05154_);
  nor (_05168_, _21559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  nor (_05169_, _21586_, _21561_);
  nor (_22129_, _05169_, _05168_);
  nor (_05170_, _21559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  nor (_05171_, _21561_, _21554_);
  nor (_22157_, _05171_, _05170_);
  nor (_05173_, _21869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7]);
  nor (_05174_, _21871_, _21626_);
  nor (_22163_, _05174_, _05173_);
  nor (_05175_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  nand (_05176_, _23553_, _00062_);
  nand (_05177_, _05176_, _23493_);
  nor (_22177_, _05177_, _05175_);
  nor (_05178_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  not (_05179_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand (_05180_, _23553_, _05179_);
  nand (_05181_, _05180_, _23493_);
  nor (_25042_[24], _05181_, _05178_);
  nor (_05182_, _21869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  nor (_05183_, _21871_, _21504_);
  nor (_22185_, _05183_, _05182_);
  nor (_05184_, _21873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  nor (_05185_, _21875_, _21526_);
  nor (_22218_, _05185_, _05184_);
  nor (_05186_, _24129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  nor (_05187_, _24131_, _21586_);
  nor (_22237_, _05187_, _05186_);
  nand (_05188_, _24769_, _23044_);
  nand (_05189_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_05190_, _05189_, _05188_);
  nor (_05191_, _05190_, _23518_);
  nor (_25021_[2], _05191_, rst);
  nor (_05192_, _22551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  nor (_05193_, _22555_, _21526_);
  nor (_22244_, _05193_, _05192_);
  nor (_05194_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  not (_05195_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_05197_, _23553_, _05195_);
  nand (_05198_, _05197_, _23493_);
  nor (_22247_, _05198_, _05194_);
  nor (_05199_, _21559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  nor (_05201_, _21561_, _21526_);
  nor (_22254_, _05201_, _05199_);
  nor (_05202_, _21531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1]);
  nor (_05203_, _21533_, _21474_);
  nor (_25255_, _05203_, _05202_);
  nor (_05204_, _24129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  nor (_05205_, _24131_, _21526_);
  nor (_22267_, _05205_, _05204_);
  nor (_05206_, _24129_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  nor (_05208_, _24131_, _21554_);
  nor (_25381_, _05208_, _05206_);
  nand (_05209_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor (_05210_, _05209_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  nand (_05211_, _05210_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor (_22304_, _05211_, rst);
  nor (_05212_, _00531_, _00461_);
  not (_05213_, _05212_);
  nor (_05215_, _00647_, _00052_);
  not (_05216_, _05215_);
  nor (_05217_, _05216_, _05213_);
  nor (_05219_, _00385_, _00556_);
  not (_05220_, _05219_);
  nor (_05221_, _05220_, _00317_);
  not (_05222_, _05221_);
  nor (_05223_, _05222_, _00225_);
  nand (_05224_, _05223_, _05217_);
  not (_05225_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  nor (_05226_, _05225_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_05227_, _05226_);
  nor (_05228_, _05227_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not (_05229_, _05228_);
  nor (_05230_, _05229_, _05224_);
  nor (_05231_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_05232_, _05231_, _00246_);
  nand (_05233_, _05232_, _00317_);
  nor (_05234_, _05233_, _05220_);
  nand (_05235_, _05234_, _05217_);
  nor (_05236_, _00634_, _02437_);
  nor (_05237_, _00384_, _00556_);
  nand (_05238_, _05237_, _00317_);
  not (_05239_, _05238_);
  nand (_05240_, _05239_, _00246_);
  not (_05241_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  nor (_05242_, _05227_, _05241_);
  nand (_05243_, _05242_, _05212_);
  nor (_05244_, _05243_, _05240_);
  nand (_05245_, _05244_, _05236_);
  nand (_05246_, _05245_, _05235_);
  nor (_05247_, _05246_, _05230_);
  nor (_05248_, _05247_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_05250_, _00634_, _24856_);
  nor (_05251_, _00647_, _21320_);
  nor (_05252_, _05251_, _05250_);
  nor (_05253_, _02437_, _24855_);
  nor (_05254_, _00052_, _21285_);
  nor (_05255_, _05254_, _05253_);
  nand (_05256_, _05255_, _05252_);
  nor (_05257_, _00641_, _21308_);
  nor (_05258_, _00461_, _24877_);
  nor (_05259_, _05258_, _05257_);
  nor (_05260_, _00531_, _21351_);
  nor (_05261_, _00671_, _00905_);
  nor (_05262_, _05261_, _05260_);
  not (_05263_, _05262_);
  nor (_05264_, _05263_, _05259_);
  not (_05265_, _05264_);
  nor (_05266_, _05265_, _05256_);
  not (_05267_, _05266_);
  nor (_05269_, _00246_, _21268_);
  nor (_05270_, _00225_, _24897_);
  nor (_05272_, _05270_, _05269_);
  nor (_05273_, _00317_, _21337_);
  nor (_05274_, _00318_, _21336_);
  nor (_05275_, _05274_, _05273_);
  nor (_05276_, _05275_, _05272_);
  nor (_05277_, _00385_, _21365_);
  nor (_05278_, _00384_, _21377_);
  nor (_05279_, _05278_, _05277_);
  nor (_05280_, _05279_, _00657_);
  nand (_05281_, _05280_, _05276_);
  nor (_05282_, _05281_, _05267_);
  nand (_05283_, _05282_, _00912_);
  nor (_05284_, _21227_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  not (_05285_, _05284_);
  nor (_05286_, _05285_, _05283_);
  not (_05287_, _05286_);
  nor (_05288_, _05241_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_05289_, _05288_, _05225_);
  nor (_05290_, _05289_, _05224_);
  nor (_05291_, _05272_, _05259_);
  nor (_05293_, _05279_, _05275_);
  not (_05294_, _05293_);
  nor (_05295_, _05294_, _00657_);
  nand (_05296_, _05295_, _05291_);
  nand (_05297_, _05236_, _00531_);
  nand (_05298_, _05297_, _00916_);
  nor (_05299_, _05298_, _05296_);
  nor (_05300_, _05299_, _05290_);
  nand (_05301_, _05300_, _05287_);
  nor (_05302_, _05301_, _05248_);
  nor (_05303_, _00647_, _02437_);
  nand (_05304_, _05303_, _05244_);
  nand (_05305_, _05304_, _23493_);
  nor (_22309_, _05305_, _05302_);
  nor (_05306_, _24110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  nor (_05307_, _24112_, _21414_);
  nor (_22340_, _05307_, _05306_);
  nor (_05308_, _23545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  nor (_05309_, _23547_, _21526_);
  nor (_22345_, _05309_, _05308_);
  nor (_05310_, _24110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  nor (_05311_, _24112_, _21526_);
  nor (_22350_, _05311_, _05310_);
  nor (_05312_, _21531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  nor (_05313_, _21554_, _21533_);
  nor (_22375_, _05313_, _05312_);
  nor (_05314_, _21782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5]);
  nor (_05315_, _21784_, _21451_);
  nor (_25218_, _05315_, _05314_);
  nor (_05317_, _21782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  nor (_05318_, _21784_, _21504_);
  nor (_22391_, _05318_, _05317_);
  nor (_05320_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand (_05321_, _23553_, _00283_);
  nand (_05322_, _05321_, _23493_);
  nor (_22400_, _05322_, _05320_);
  nor (_05323_, _22454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  nor (_05324_, _22456_, _21526_);
  nor (_22405_, _05324_, _05323_);
  nor (_05326_, _22490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  nor (_05328_, _22492_, _21414_);
  nor (_22419_, _05328_, _05326_);
  nor (_05329_, _24110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  nor (_05330_, _24112_, _21504_);
  nor (_22433_, _05330_, _05329_);
  nor (_05331_, _24110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5]);
  nor (_05332_, _24112_, _21451_);
  nor (_22436_, _05332_, _05331_);
  nor (_05333_, _23833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7]);
  nor (_05334_, _23835_, _21626_);
  nor (_22460_, _05334_, _05333_);
  nor (_05335_, _21531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  nor (_05336_, _21533_, _21414_);
  nor (_25257_, _05336_, _05335_);
  nor (_05337_, _21782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  nor (_05338_, _21784_, _21526_);
  nor (_22469_, _05338_, _05337_);
  nor (_05340_, _21531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  nor (_05341_, _21533_, _21504_);
  nor (_22472_, _05341_, _05340_);
  nor (_05342_, _21782_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  nor (_05343_, _21784_, _21414_);
  nor (_22480_, _05343_, _05342_);
  nor (_05344_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  not (_05345_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_05346_, _23553_, _05345_);
  nand (_05347_, _05346_, _23493_);
  nor (_22518_, _05347_, _05344_);
  nor (_05348_, _21869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5]);
  nor (_05349_, _21871_, _21451_);
  nor (_22522_, _05349_, _05348_);
  nor (_05350_, _22396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  nor (_05351_, _22398_, _21504_);
  nor (_22530_, _05351_, _05350_);
  nor (_05353_, _24110_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1]);
  nor (_05355_, _24112_, _21474_);
  nor (_22552_, _05355_, _05353_);
  nor (_05356_, _21645_, _21374_);
  nor (_05357_, _05356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7]);
  not (_05358_, _05356_);
  nor (_05360_, _05358_, _21626_);
  nor (_22575_, _05360_, _05357_);
  nor (_05361_, _21483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  nor (_05362_, _21586_, _21485_);
  nor (_22580_, _05362_, _05361_);
  nor (_05363_, _23044_, _21279_);
  not (_05364_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  nor (_05365_, _23153_, _05364_);
  nor (_05366_, _23050_, _24830_);
  nor (_05367_, _23076_, _24835_);
  nor (_05368_, _05367_, _05366_);
  not (_05369_, _05368_);
  nor (_05370_, _23073_, _05195_);
  nor (_05371_, _23107_, _23257_);
  nor (_05372_, _05371_, _05370_);
  nor (_05373_, _23067_, _23259_);
  nor (_05374_, _23058_, _23233_);
  nor (_05375_, _05374_, _05373_);
  nand (_05376_, _05375_, _05372_);
  nor (_05377_, _05376_, _05369_);
  nor (_05378_, _05377_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_05379_, _05378_, _05365_);
  nor (_05380_, _05379_, _23490_);
  nor (_05381_, _05380_, _05363_);
  nor (_22589_, _05381_, rst);
  nor (_05382_, _21483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1]);
  nor (_05383_, _21485_, _21474_);
  nor (_22597_, _05383_, _05382_);
  nor (_05384_, _21483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  nor (_05385_, _21526_, _21485_);
  nor (_25259_, _05385_, _05384_);
  nor (_05386_, _22403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  nor (_05387_, _22406_, _21554_);
  nor (_22610_, _05387_, _05386_);
  nor (_05388_, _22500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1]);
  nor (_05389_, _22502_, _21474_);
  nor (_22618_, _05389_, _05388_);
  nor (_05390_, _21483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  nor (_05391_, _21485_, _21414_);
  nor (_22643_, _05391_, _05390_);
  nor (_05393_, _22450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  nor (_05394_, _22452_, _21554_);
  nor (_22687_, _05394_, _05393_);
  nor (_05395_, _23806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  nor (_05397_, _23808_, _21586_);
  nor (_22691_, _05397_, _05395_);
  nor (_05398_, _01083_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  nor (_05400_, _01052_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  nand (_05401_, _05400_, _01080_);
  nand (_05403_, _05401_, _23493_);
  nor (_22694_, _05403_, _05398_);
  nor (_05404_, _21816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  nor (_05405_, _21818_, _21526_);
  nor (_25205_, _05405_, _05404_);
  nor (_05406_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  nor (_05407_, _22563_, _21504_);
  nor (_25077_, _05407_, _05406_);
  nor (_05408_, _23810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7]);
  nor (_05409_, _23812_, _21626_);
  nor (_22711_, _05409_, _05408_);
  nor (_05411_, _22465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  nor (_05412_, _22467_, _21586_);
  nor (_22715_, _05412_, _05411_);
  nor (_05413_, _02439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  nor (_05415_, _02442_, _21586_);
  nor (_22720_, _05415_, _05413_);
  nor (_05418_, _01142_, _02344_);
  not (_05419_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor (_05420_, _01143_, _05419_);
  nor (_05422_, _05420_, _05418_);
  nor (_05424_, _05422_, _01130_);
  nand (_05425_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _02387_);
  nand (_05427_, _05425_, _01059_);
  nor (_05428_, _05427_, _02360_);
  nor (_05430_, _05428_, _05424_);
  nor (_22722_, _05430_, rst);
  nand (_05431_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nand (_05432_, _01142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  nand (_05434_, _05432_, _05431_);
  nor (_05435_, _05434_, _01130_);
  nor (_05436_, _01055_, ABINPUT[10]);
  nand (_05437_, _05436_, _01130_);
  nand (_05438_, _05437_, _23493_);
  nor (_22727_, _05438_, _05435_);
  nor (_05439_, _21816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  nor (_05440_, _21818_, _21554_);
  nor (_22729_, _05440_, _05439_);
  nor (_05441_, _23806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  nor (_05442_, _23808_, _21414_);
  nor (_22737_, _05442_, _05441_);
  nor (_05443_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  nor (_05445_, _22473_, _21586_);
  nor (_22742_, _05445_, _05443_);
  nor (_05446_, _23806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  nor (_05447_, _23808_, _21526_);
  nor (_22748_, _05447_, _05446_);
  nor (_05448_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1]);
  nor (_05449_, _22508_, _21474_);
  nor (_22753_, _05449_, _05448_);
  nor (_05450_, _21816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  nor (_05452_, _21818_, _21586_);
  nor (_22755_, _05452_, _05450_);
  nor (_05453_, _01183_, _21652_);
  nor (_05454_, _05453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  not (_05455_, _05453_);
  nor (_05456_, _05455_, _21504_);
  nor (_22774_, _05456_, _05454_);
  nor (_05457_, _22465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7]);
  nor (_05458_, _22467_, _21626_);
  nor (_22777_, _05458_, _05457_);
  nor (_05459_, _05453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5]);
  nor (_05460_, _05455_, _21451_);
  nor (_25336_, _05460_, _05459_);
  nor (_05461_, _05453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  nor (_05462_, _05455_, _21414_);
  nor (_22788_, _05462_, _05461_);
  nor (_05463_, _23806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  nor (_05464_, _23808_, _21554_);
  nor (_22809_, _05464_, _05463_);
  nor (_05465_, _21850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7]);
  nor (_05467_, _21853_, _21626_);
  nor (_22814_, _05467_, _05465_);
  nor (_05468_, _23810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  nor (_05469_, _23812_, _21526_);
  nor (_22850_, _05469_, _05468_);
  nor (_05470_, _23810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  nor (_05471_, _23812_, _21554_);
  nor (_22859_, _05471_, _05470_);
  nor (_05472_, _23810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  nor (_05473_, _23812_, _21414_);
  nor (_22868_, _05473_, _05472_);
  nor (_05474_, _23810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  nor (_05475_, _23812_, _21504_);
  nor (_22871_, _05475_, _05474_);
  nor (_05476_, _23810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5]);
  nor (_05477_, _23812_, _21451_);
  nor (_22875_, _05477_, _05476_);
  nor (_05478_, _22479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  nor (_05479_, _22482_, _21414_);
  nor (_22880_, _05479_, _05478_);
  nor (_05481_, _21483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5]);
  nor (_05482_, _21485_, _21451_);
  nor (_22888_, _05482_, _05481_);
  nor (_05483_, _21483_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7]);
  nor (_05484_, _21626_, _21485_);
  nor (_22906_, _05484_, _05483_);
  nor (_05485_, _24094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  nor (_05486_, _24096_, _21414_);
  nor (_22916_, _05486_, _05485_);
  nor (_05487_, _24094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  nor (_05488_, _24096_, _21504_);
  nor (_22926_, _05488_, _05487_);
  nor (_05489_, _24094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5]);
  nor (_05490_, _24096_, _21451_);
  nor (_22935_, _05490_, _05489_);
  nor (_05492_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  nor (_05493_, _22280_, _21504_);
  nor (_22944_, _05493_, _05492_);
  nor (_05496_, _24094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7]);
  nor (_05497_, _24096_, _21626_);
  nor (_22959_, _05497_, _05496_);
  nor (_05498_, _23810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  nor (_05499_, _23812_, _21586_);
  nor (_22964_, _05499_, _05498_);
  nand (_05500_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nand (_05501_, _23493_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_22979_, _05501_, _05500_);
  nor (_05502_, _01383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  nor (_05503_, _01385_, _21526_);
  nor (_22985_, _05503_, _05502_);
  nor (_05505_, _23865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7]);
  nor (_05506_, _23868_, _21626_);
  nor (_23019_, _05506_, _05505_);
  nor (_05507_, _24094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  nor (_05508_, _24096_, _21586_);
  nor (_25369_, _05508_, _05507_);
  nor (_05509_, _02439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7]);
  nor (_05511_, _02442_, _21626_);
  nor (_23024_, _05511_, _05509_);
  nor (_05512_, _22021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  nor (_05513_, _22023_, _21586_);
  nor (_23033_, _05513_, _05512_);
  nor (_05516_, _01184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  nor (_05517_, _01186_, _21504_);
  nor (_23053_, _05517_, _05516_);
  nor (_05519_, _21689_, _21645_);
  nor (_05520_, _05519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  not (_05521_, _05519_);
  nor (_05522_, _05521_, _21504_);
  nor (_23071_, _05522_, _05520_);
  nor (_05526_, _01184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5]);
  nor (_05528_, _01186_, _21451_);
  nor (_23089_, _05528_, _05526_);
  nor (_05529_, _24094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  nor (_05530_, _24096_, _21554_);
  nor (_23093_, _05530_, _05529_);
  nor (_05531_, _24094_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1]);
  nor (_05532_, _24096_, _21474_);
  nor (_25370_, _05532_, _05531_);
  nor (_05533_, _22479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  nor (_05534_, _22482_, _21554_);
  nor (_23136_, _05534_, _05533_);
  nor (_05535_, _23865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1]);
  nor (_05536_, _23868_, _21474_);
  nor (_23142_, _05536_, _05535_);
  nor (_05537_, _22838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7]);
  nor (_05539_, _22840_, _21626_);
  nor (_23158_, _05539_, _05537_);
  nor (_05540_, _23865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  nor (_05541_, _23868_, _21586_);
  nor (_23171_, _05541_, _05540_);
  nor (_05543_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1]);
  nor (_05544_, _22783_, _21474_);
  nor (_25127_, _05544_, _05543_);
  nor (_05545_, _23865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  nor (_05546_, _23868_, _21526_);
  nor (_23196_, _05546_, _05545_);
  nor (_05547_, _23865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  nor (_05548_, _23868_, _21414_);
  nor (_23205_, _05548_, _05547_);
  nor (_05549_, _21850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  nor (_05550_, _21853_, _21504_);
  nor (_25197_, _05550_, _05549_);
  nor (_05551_, _05453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1]);
  nor (_05553_, _05455_, _21474_);
  nor (_23252_, _05553_, _05551_);
  nor (_05554_, _22838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  nor (_05555_, _22840_, _21586_);
  nor (_23260_, _05555_, _05554_);
  nor (_05556_, _21822_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  nor (_05557_, _21824_, _21554_);
  nor (_23267_, _05557_, _05556_);
  nor (_05558_, _00907_, _21351_);
  not (_05559_, _05558_);
  nor (_05560_, _05559_, _21308_);
  nor (_05561_, _00915_, _00018_);
  nand (_05562_, _05561_, _05560_);
  nor (_05563_, _05562_, _21507_);
  nor (_05564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_05565_, _05564_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  not (_05566_, _05565_);
  not (_05567_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_05568_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_05569_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_05571_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_05572_, _05571_, _05569_);
  not (_05573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor (_05574_, _05573_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_05575_, _05574_, _05572_);
  nor (_05577_, _05575_, _05568_);
  nor (_05579_, _05577_, _05567_);
  not (_05580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor (_05581_, _05580_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_05582_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_05583_, _05571_, _05582_);
  nor (_05584_, _05583_, _05581_);
  nor (_05585_, _05584_, _05568_);
  not (_05586_, _05585_);
  not (_05587_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nor (_05588_, _05587_, _05571_);
  nand (_05589_, _05571_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  not (_05590_, _05589_);
  nor (_05591_, _05590_, _05588_);
  not (_05592_, _05591_);
  nor (_05593_, _05592_, _05586_);
  nand (_05594_, _05593_, _05579_);
  nand (_05595_, _05594_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nand (_05596_, _05595_, _05566_);
  nand (_05597_, _05596_, _05562_);
  nor (_05598_, _00927_, _00018_);
  not (_05599_, _05598_);
  nand (_05600_, _05599_, _05597_);
  nor (_05601_, _05600_, _05563_);
  nand (_05602_, _05598_, _00106_);
  nand (_05603_, _05602_, _23493_);
  nor (_23270_, _05603_, _05601_);
  nor (_05604_, _23817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  nor (_05605_, _23819_, _21414_);
  nor (_23274_, _05605_, _05604_);
  not (_05606_, _05500_);
  not (_05607_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  not (_05608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  nor (_05609_, _05608_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_05610_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  not (_05611_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  nor (_05612_, _05611_, _05571_);
  nor (_05614_, _05612_, _05610_);
  not (_05615_, _05614_);
  nor (_05616_, _05615_, _05609_);
  nor (_05617_, _05616_, _05568_);
  not (_05619_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nand (_05620_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nor (_05622_, _05620_, _05619_);
  not (_05623_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  not (_05624_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  not (_05625_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  nor (_05626_, _05625_, _05624_);
  not (_05627_, _05626_);
  nor (_05628_, _05627_, _05623_);
  not (_05629_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nand (_05630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nor (_05631_, _05630_, _05629_);
  nor (_05632_, _05631_, _05628_);
  not (_05633_, _05632_);
  nor (_05634_, _05633_, _05622_);
  not (_05635_, _05634_);
  not (_05636_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_05637_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_05638_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_05639_, _05638_, _05637_);
  not (_05641_, _05639_);
  nor (_05642_, _05641_, _05636_);
  not (_05644_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_05645_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_05646_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor (_05647_, _05646_, _05645_);
  not (_05648_, _05647_);
  nor (_05649_, _05648_, _05644_);
  nor (_05650_, _05649_, _05642_);
  not (_05651_, _05650_);
  not (_05652_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nand (_05653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nor (_05654_, _05653_, _05652_);
  nor (_05655_, _05654_, _05651_);
  not (_05656_, _05655_);
  nor (_05657_, _05656_, _05635_);
  nor (_05658_, _05657_, _05617_);
  nor (_05659_, _05610_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  nor (_05660_, _05641_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  nor (_05661_, _05648_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nor (_05663_, _05661_, _05660_);
  nor (_05664_, _05653_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor (_05665_, _05620_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  nor (_05666_, _05627_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_05667_, _05630_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_05668_, _05667_, _05666_);
  not (_05669_, _05668_);
  nor (_05670_, _05669_, _05665_);
  not (_05671_, _05670_);
  nor (_05672_, _05671_, _05664_);
  nand (_05673_, _05672_, _05663_);
  nand (_05674_, _05673_, _05659_);
  not (_05675_, _05674_);
  nor (_05676_, _05675_, _05658_);
  not (_05677_, _05676_);
  nor (_05678_, _05677_, _05607_);
  not (_05679_, _05658_);
  nor (_05680_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _05571_);
  nor (_05681_, _05607_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_05682_, _05681_, _05680_);
  nor (_05684_, _05682_, _05679_);
  nor (_05686_, _05684_, _05678_);
  nor (_05687_, _05686_, _05606_);
  not (_05688_, _05682_);
  nor (_05690_, _05688_, _05500_);
  nor (_05691_, _05690_, _05687_);
  nor (_23281_, _05691_, rst);
  nor (_05693_, _05453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  nor (_05694_, _05455_, _21586_);
  nor (_23291_, _05694_, _05693_);
  nor (_05696_, _01183_, _21631_);
  nor (_05698_, _05696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7]);
  not (_05699_, _05696_);
  nor (_05700_, _05699_, _21626_);
  nor (_23311_, _05700_, _05698_);
  nor (_05701_, _01184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  nor (_05702_, _01186_, _21586_);
  nor (_23314_, _05702_, _05701_);
  nor (_05703_, _22490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  nor (_05704_, _22492_, _21526_);
  nor (_23322_, _05704_, _05703_);
  nor (_05706_, _22869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  nor (_05707_, _22872_, _21504_);
  nor (_23325_, _05707_, _05706_);
  nor (_05708_, _01184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1]);
  nor (_05709_, _01186_, _21474_);
  nor (_23336_, _05709_, _05708_);
  nor (_05710_, _01184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  nor (_05711_, _01186_, _21526_);
  nor (_23340_, _05711_, _05710_);
  nor (_05712_, _01184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  nor (_05713_, _01186_, _21554_);
  nor (_23344_, _05713_, _05712_);
  not (_05714_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor (_05715_, _00742_, _05714_);
  nor (_05716_, _00740_, _00106_);
  nor (_05717_, _05716_, _05715_);
  nor (_23357_, _05717_, rst);
  not (_05718_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_05719_, _00738_, _00013_);
  nand (_05721_, _05719_, _24859_);
  not (_05722_, _05721_);
  nor (_05723_, _05722_, _05718_);
  nor (_05724_, _05721_, _00106_);
  nor (_05725_, _05724_, _05723_);
  nor (_23361_, _05725_, rst);
  nor (_05726_, _24858_, _21308_);
  not (_05727_, _00738_);
  nand (_05728_, _05727_, _05726_);
  nor (_05729_, _05728_, _24860_);
  nor (_05730_, _05729_, _00079_);
  not (_05731_, _05726_);
  nor (_05732_, _05731_, _24860_);
  nand (_05733_, _05727_, _05732_);
  nor (_05734_, _05733_, _00106_);
  nor (_05735_, _05734_, _05730_);
  nor (_23363_, _05735_, rst);
  not (_05736_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_05737_, _00020_, _21308_);
  nand (_05738_, _05737_, _05727_);
  nor (_05740_, _05738_, _24860_);
  nor (_05741_, _05740_, _05736_);
  not (_05742_, _05737_);
  nor (_05743_, _05742_, _24860_);
  nand (_05744_, _05743_, _05727_);
  nor (_05745_, _05744_, _00106_);
  nor (_05746_, _05745_, _05741_);
  nor (_23380_, _05746_, rst);
  not (_05747_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  not (_05748_, _00737_);
  nor (_05749_, _05748_, _24849_);
  nand (_05751_, _24902_, _05749_);
  nor (_05753_, _05751_, _24860_);
  nor (_05754_, _05753_, _05747_);
  not (_05755_, _05753_);
  nor (_05756_, _05755_, _00106_);
  nor (_05758_, _05756_, _05754_);
  nor (_23390_, _05758_, rst);
  not (_05760_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor (_05762_, _00847_, _05760_);
  nor (_05764_, _00848_, _00106_);
  nor (_05765_, _05764_, _05762_);
  nor (_25028_[7], _05765_, rst);
  nor (_05766_, _24661_, _00089_);
  nor (_05767_, _24663_, _00106_);
  nor (_05768_, _05767_, _05766_);
  nor (_23395_, _05768_, rst);
  nor (_05770_, _23817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  nor (_05771_, _23819_, _21504_);
  nor (_23399_, _05771_, _05770_);
  not (_05772_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nand (_05773_, _05737_, _05749_);
  nor (_05774_, _05773_, _24860_);
  nor (_05775_, _05774_, _05772_);
  nand (_05777_, _05743_, _05749_);
  nor (_05779_, _05777_, _00106_);
  nor (_05781_, _05779_, _05775_);
  nor (_23401_, _05781_, rst);
  nor (_05784_, _22403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  nor (_05785_, _22406_, _21526_);
  nor (_23406_, _05785_, _05784_);
  nor (_05786_, _05696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  nor (_05787_, _05699_, _21554_);
  nor (_25334_, _05787_, _05786_);
  nor (_05788_, _23557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  nor (_05789_, _23560_, _21554_);
  nor (_23417_, _05789_, _05788_);
  nor (_05790_, _05696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1]);
  nor (_05791_, _05699_, _21474_);
  nor (_23437_, _05791_, _05790_);
  nor (_05793_, _23825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7]);
  nor (_05794_, _23827_, _21626_);
  nor (_23439_, _05794_, _05793_);
  nor (_05795_, _05696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  nor (_05796_, _05699_, _21586_);
  nor (_23446_, _05796_, _05795_);
  nor (_05797_, _22465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  nor (_05798_, _22467_, _21554_);
  nor (_23453_, _05798_, _05797_);
  nor (_05799_, _22465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  nor (_05800_, _22467_, _21414_);
  nor (_25080_, _05800_, _05799_);
  nor (_05801_, _23817_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1]);
  nor (_05802_, _23819_, _21474_);
  nor (_25368_, _05802_, _05801_);
  nor (_05803_, _01383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7]);
  nor (_05804_, _01385_, _21626_);
  nor (_23483_, _05804_, _05803_);
  nor (_05805_, _21690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1]);
  nor (_05806_, _21692_, _21474_);
  nor (_23494_, _05806_, _05805_);
  nand (_05807_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nand (_05808_, _01142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nand (_05809_, _05808_, _05807_);
  nor (_05810_, _05809_, _01130_);
  nor (_05811_, _01059_, _24867_);
  nor (_05812_, _01055_, _00121_);
  nor (_05813_, _05812_, _05811_);
  nand (_05814_, _05813_, _01130_);
  nand (_05815_, _05814_, _23493_);
  nor (_23503_, _05815_, _05810_);
  nor (_05816_, _23825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  nor (_05817_, _23827_, _21526_);
  nor (_23506_, _05817_, _05816_);
  nor (_05818_, _23825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  nor (_05819_, _23827_, _21414_);
  nor (_23511_, _05819_, _05818_);
  nor (_05820_, _05696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  nor (_05821_, _05699_, _21526_);
  nor (_25335_, _05821_, _05820_);
  nor (_05822_, _05696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5]);
  nor (_05823_, _05699_, _21451_);
  nor (_23526_, _05823_, _05822_);
  nor (_05824_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  nor (_05825_, _22508_, _21554_);
  nor (_23530_, _05825_, _05824_);
  nor (_05826_, _05696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  nor (_05827_, _05699_, _21414_);
  nor (_23533_, _05827_, _05826_);
  nor (_05828_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  nand (_05829_, _03721_, _00106_);
  nand (_05830_, _05829_, _23493_);
  nor (_23538_, _05830_, _05828_);
  nor (_05831_, _01194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  nor (_05832_, _01196_, _21526_);
  nor (_23548_, _05832_, _05831_);
  nor (_05834_, _01194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  nor (_05835_, _01196_, _21554_);
  nor (_23550_, _05835_, _05834_);
  nor (_05836_, _21430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  nor (_05837_, _21586_, _21432_);
  nor (_25260_, _05837_, _05836_);
  nor (_05838_, _03937_, _03667_);
  nor (_05839_, _05838_, _03687_);
  not (_05840_, _05839_);
  nand (_05841_, _05840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_05842_, _03891_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_05843_, _05842_, _03894_);
  nand (_05844_, _05843_, _05839_);
  nand (_05845_, _05844_, _05841_);
  nor (_05846_, _04943_, _03618_);
  nand (_05847_, _05846_, _03688_);
  nand (_05848_, _05847_, _03909_);
  nor (_05849_, _05848_, _05845_);
  nand (_05850_, _03702_, _00106_);
  nand (_05851_, _05850_, _23493_);
  nor (_23566_, _05851_, _05849_);
  nor (_23573_, rst, _03642_);
  nor (_05852_, _22551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7]);
  nor (_05853_, _22555_, _21626_);
  nor (_25084_, _05853_, _05852_);
  nor (_05854_, _23825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5]);
  nor (_05855_, _23827_, _21451_);
  nor (_25367_, _05855_, _05854_);
  nor (_05856_, _22454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  nor (_05857_, _22456_, _21586_);
  nor (_25085_, _05857_, _05856_);
  nor (_05858_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand (_05859_, _23553_, _23183_);
  nand (_05860_, _05859_, _23493_);
  nor (_25042_[11], _05860_, _05858_);
  nor (_05861_, _00880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  nor (_05862_, _00882_, _21504_);
  nor (_23605_, _05862_, _05861_);
  nor (_05863_, _23873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7]);
  nor (_05864_, _23875_, _21626_);
  nor (_23618_, _05864_, _05863_);
  nor (_05865_, _23873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  nor (_05866_, _23875_, _21504_);
  nor (_23621_, _05866_, _05865_);
  nor (_05868_, _23825_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  nor (_05869_, _23827_, _21586_);
  nor (_23635_, _05869_, _05868_);
  nor (_05870_, _23873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  nor (_05871_, _23875_, _21526_);
  nor (_23645_, _05871_, _05870_);
  nor (_05872_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5]);
  nor (_05873_, _22280_, _21451_);
  nor (_23649_, _05873_, _05872_);
  nor (_05874_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  nor (_05876_, _22280_, _21526_);
  nor (_23656_, _05876_, _05874_);
  nor (_05878_, _22278_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1]);
  nor (_05879_, _22280_, _21474_);
  nor (_25154_, _05879_, _05878_);
  nor (_23674_, rst, _02674_);
  nor (_05881_, _24050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7]);
  nor (_05883_, _24052_, _21626_);
  nor (_23688_, _05883_, _05881_);
  nor (_05885_, _24050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  nor (_05886_, _24052_, _21504_);
  nor (_25365_, _05886_, _05885_);
  nor (_05887_, _22838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  nor (_05889_, _22840_, _21414_);
  nor (_23699_, _05889_, _05887_);
  nor (_05891_, _01194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  nor (_05892_, _01196_, _21504_);
  nor (_23703_, _05892_, _05891_);
  nor (_05894_, _22292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7]);
  nor (_05895_, _22294_, _21626_);
  nor (_23706_, _05895_, _05894_);
  nor (_05897_, _21430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  nor (_05898_, _21554_, _21432_);
  nor (_23712_, _05898_, _05897_);
  nor (_05899_, _23873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  nor (_05900_, _23875_, _21586_);
  nor (_23715_, _05900_, _05899_);
  nand (_05901_, _02705_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  nand (_05903_, _02656_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_05904_, _05903_, _03731_);
  not (_05905_, _03731_);
  nand (_05907_, _03810_, _02660_);
  nand (_05908_, _05907_, _02707_);
  nand (_05909_, _05908_, _05905_);
  nand (_05910_, _05909_, _05904_);
  nand (_05911_, _05910_, _05901_);
  nor (_05912_, _05911_, _02612_);
  nand (_05913_, _02612_, _02660_);
  nand (_05914_, _05913_, _02626_);
  nor (_05915_, _05914_, _05912_);
  nor (_05917_, _02626_, _00106_);
  nor (_05918_, _05917_, _05915_);
  nor (_23720_, _05918_, rst);
  nor (_05920_, _01194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5]);
  nor (_05921_, _01196_, _21451_);
  nor (_23724_, _05921_, _05920_);
  nor (_05922_, _02625_, rst);
  not (_05923_, _05922_);
  not (_05924_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not (_05925_, _02681_);
  nor (_05926_, _05925_, _05924_);
  not (_05927_, _05926_);
  nand (_05928_, _05927_, _02704_);
  nand (_05929_, _05928_, _02705_);
  nand (_05930_, _02650_, _02619_);
  nand (_05931_, _05930_, _03731_);
  nand (_05932_, _05931_, _05927_);
  nand (_05933_, _05932_, _02707_);
  nand (_05934_, _05933_, _05929_);
  nand (_05935_, _05934_, _02613_);
  nor (_23731_, _05935_, _05923_);
  nor (_05938_, _03652_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nand (_05940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_05942_, _05940_, _05938_);
  nand (_05944_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _03917_);
  nor (_05945_, _05944_, _03954_);
  nor (_05946_, _05945_, _05942_);
  nand (_05947_, _05946_, _04943_);
  nor (_05949_, _05947_, _03682_);
  nor (_05950_, _03702_, _03687_);
  nand (_05951_, _05950_, _23493_);
  nor (_23734_, _05951_, _05949_);
  nor (_05952_, _01183_, _21482_);
  nor (_05953_, _05952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  not (_05954_, _05952_);
  nor (_05955_, _05954_, _21414_);
  nor (_25333_, _05955_, _05953_);
  nor (_05957_, _05952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  nor (_05958_, _05954_, _21526_);
  nor (_25332_, _05958_, _05957_);
  nor (_05960_, _05952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7]);
  nor (_05961_, _05954_, _21626_);
  nor (_23762_, _05961_, _05960_);
  nor (_05962_, _05952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  nor (_05964_, _05954_, _21504_);
  nor (_23765_, _05964_, _05962_);
  nor (_05966_, _24050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1]);
  nor (_05968_, _24052_, _21474_);
  nor (_23773_, _05968_, _05966_);
  nor (_05970_, _01383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5]);
  nor (_05971_, _01385_, _21451_);
  nor (_23780_, _05971_, _05970_);
  nor (_05974_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7]);
  nor (_05975_, _02331_, _21626_);
  nor (_25331_, _05975_, _05974_);
  nor (_05976_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  nor (_05977_, _02331_, _21504_);
  nor (_23787_, _05977_, _05976_);
  nor (_05978_, _24050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  nor (_05979_, _24052_, _21554_);
  nor (_23804_, _05979_, _05978_);
  nor (_05981_, _05356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  nor (_05982_, _05358_, _21554_);
  nor (_23820_, _05982_, _05981_);
  nor (_05983_, _22465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  nor (_05985_, _22467_, _21504_);
  nor (_25082_, _05985_, _05983_);
  nor (_05987_, _24050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  nor (_05988_, _24052_, _21586_);
  nor (_23823_, _05988_, _05987_);
  nand (_05989_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nand (_05990_, _01142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nand (_05991_, _05990_, _05989_);
  nor (_05992_, _05991_, _01130_);
  nor (_05994_, _01059_, _00121_);
  nor (_05995_, _01055_, _00006_);
  nor (_05996_, _05995_, _05994_);
  nand (_05997_, _05996_, _01130_);
  nand (_05998_, _05997_, _23493_);
  nor (_23866_, _05998_, _05992_);
  nor (_06000_, _24050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  nor (_06001_, _24052_, _21414_);
  nor (_23869_, _06001_, _06000_);
  not (_06002_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  not (_06003_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_06005_, _23553_, _06003_);
  not (_06006_, _06005_);
  nor (_06007_, _06006_, _06002_);
  nor (_06008_, _06005_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_06009_, _06008_, _06007_);
  nor (_06010_, _06009_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_06011_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_06013_, _06011_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor (_06014_, _06013_, _06010_);
  not (_06015_, _23553_);
  nor (_06016_, _06015_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_06017_, _06016_, _06005_);
  nor (_06018_, _06017_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_06019_, _06011_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor (_06020_, _06019_, _06018_);
  not (_06021_, _06020_);
  nor (_06022_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_06024_, _06011_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor (_06026_, _06024_, _06022_);
  not (_06027_, _06026_);
  nor (_06028_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_06029_, _06011_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nor (_06031_, _06029_, _06028_);
  nor (_06033_, _06031_, _06027_);
  nand (_06034_, _06033_, _06021_);
  nor (_06036_, _06034_, _06014_);
  nand (_06037_, _06036_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_06038_, _06014_);
  nor (_06039_, _06038_, \oc8051_symbolic_cxrom1.regvalid [13]);
  not (_06040_, _06039_);
  nor (_06041_, _06014_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_06042_, _06041_, _06021_);
  nand (_06043_, _06042_, _06040_);
  not (_06045_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_06047_, _06020_, _06038_);
  not (_06048_, _06047_);
  nor (_06050_, _06048_, _06045_);
  not (_06051_, _06050_);
  nand (_06052_, _06051_, _06043_);
  nand (_06054_, _06052_, _06033_);
  nand (_06055_, _06054_, _06037_);
  not (_06056_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_06057_, _06020_, _06014_);
  not (_06059_, _06057_);
  nor (_06060_, _06059_, _06056_);
  not (_06061_, _06060_);
  nor (_06062_, _06021_, _06038_);
  nand (_06063_, _06062_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nand (_06064_, _06063_, _06061_);
  not (_06065_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_06066_, _06048_, _06065_);
  not (_06067_, _06066_);
  nor (_06068_, _06021_, _06014_);
  nand (_06069_, _06068_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nand (_06071_, _06069_, _06067_);
  nor (_06072_, _06071_, _06064_);
  nor (_06074_, _06031_, _06026_);
  not (_06075_, _06074_);
  nor (_06076_, _06075_, _06072_);
  nor (_06077_, _06038_, \oc8051_symbolic_cxrom1.regvalid [14]);
  not (_06078_, _06077_);
  nor (_06079_, _06014_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_06080_, _06079_, _06021_);
  nand (_06081_, _06080_, _06078_);
  not (_06082_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_06083_, _06048_, _06082_);
  not (_06084_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_06085_, _06059_, _06084_);
  nor (_06086_, _06085_, _06083_);
  nand (_06087_, _06086_, _06081_);
  not (_06089_, _06031_);
  nor (_06091_, _06089_, _06026_);
  nand (_06092_, _06091_, _06087_);
  not (_06093_, _06092_);
  nor (_06094_, _06093_, _06076_);
  not (_06095_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_06096_, _06059_, _06095_);
  not (_06097_, \oc8051_symbolic_cxrom1.regvalid [15]);
  not (_06098_, _06062_);
  nor (_06099_, _06098_, _06097_);
  nor (_06100_, _06099_, _06096_);
  not (_06101_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_06102_, _06048_, _06101_);
  not (_06103_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_06104_, _06068_);
  nor (_06106_, _06104_, _06103_);
  nor (_06108_, _06106_, _06102_);
  nand (_06109_, _06108_, _06100_);
  nor (_06111_, _06089_, _06027_);
  nand (_06112_, _06111_, _06109_);
  nand (_06114_, _06112_, _06094_);
  nor (_06115_, _06114_, _06055_);
  not (_06116_, _06115_);
  nor (_06117_, _06027_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor (_06118_, _06026_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nor (_06119_, _06118_, _06117_);
  nor (_06120_, _06119_, _06089_);
  nor (_06122_, _06027_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor (_06123_, _06026_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_06124_, _06123_, _06122_);
  nor (_06125_, _06124_, _06031_);
  nor (_06126_, _06125_, _06120_);
  nand (_06128_, _06126_, _06021_);
  nor (_06129_, _06031_, _06021_);
  not (_06130_, _06129_);
  not (_06131_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_06133_, _06026_, _06131_);
  not (_06135_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_06136_, _06027_, _06135_);
  nand (_06137_, _06136_, _06133_);
  nor (_06138_, _06137_, _06130_);
  not (_06139_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_06140_, _06026_, _06139_);
  not (_06141_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_06142_, _06027_, _06141_);
  nand (_06143_, _06142_, _06140_);
  nor (_06144_, _06089_, _06021_);
  not (_06145_, _06144_);
  nor (_06147_, _06145_, _06143_);
  nor (_06148_, _06147_, _06138_);
  nand (_06150_, _06148_, _06128_);
  nand (_06151_, _06150_, _06014_);
  nor (_06153_, _06027_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_06155_, _06026_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_06156_, _06155_, _06153_);
  not (_06159_, _06156_);
  nand (_06160_, _06159_, _06089_);
  nor (_06162_, _06027_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor (_06163_, _06026_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nor (_06164_, _06163_, _06162_);
  not (_06165_, _06164_);
  nand (_06166_, _06165_, _06031_);
  nand (_06167_, _06166_, _06160_);
  nor (_06168_, _06167_, _06020_);
  not (_06169_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_06170_, _06026_, _06169_);
  not (_06171_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_06172_, _06027_, _06171_);
  nand (_06173_, _06172_, _06170_);
  nor (_06175_, _06173_, _06130_);
  nor (_06176_, _06175_, _06168_);
  nor (_06177_, _06027_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nor (_06178_, _06026_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nor (_06180_, _06178_, _06177_);
  nand (_06181_, _06180_, _06144_);
  nand (_06183_, _06181_, _06176_);
  nand (_06184_, _06183_, _06038_);
  nand (_06185_, _06184_, _06151_);
  nand (_06186_, _06185_, _06116_);
  nand (_06187_, _06115_, word_in[7]);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _06187_, _06186_);
  nor (_06188_, _22292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  nor (_06189_, _22294_, _21504_);
  nor (_23886_, _06189_, _06188_);
  not (_06191_, _06091_);
  not (_06192_, _06111_);
  nor (_06193_, _06192_, _06021_);
  nor (_06194_, _06193_, _06038_);
  nor (_06195_, _06192_, _06104_);
  nor (_06196_, _06195_, _06194_);
  not (_06197_, _06196_);
  nor (_06199_, _06111_, _06020_);
  nor (_06200_, _06199_, _06193_);
  nor (_06202_, _06200_, _06197_);
  not (_06203_, _06202_);
  nor (_06206_, _06203_, _06095_);
  nor (_06207_, _06196_, \oc8051_symbolic_cxrom1.regvalid [15]);
  not (_06209_, _06200_);
  nor (_06211_, _06209_, _06038_);
  nor (_06212_, _06209_, _06103_);
  nor (_06214_, _06212_, _06211_);
  nor (_06215_, _06214_, _06207_);
  nor (_06217_, _06200_, _06196_);
  not (_06218_, _06217_);
  nor (_06219_, _06218_, _06101_);
  nor (_06220_, _06219_, _06215_);
  not (_06222_, _06220_);
  nor (_06223_, _06222_, _06206_);
  nor (_06225_, _06223_, _06191_);
  not (_06226_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_06227_, _06203_, _06226_);
  nor (_06228_, _06197_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_06229_, _06209_, _06039_);
  not (_06230_, _06229_);
  nor (_06231_, _06230_, _06228_);
  nor (_06234_, _06218_, _06045_);
  nor (_06235_, _06234_, _06231_);
  not (_06237_, _06235_);
  nor (_06238_, _06237_, _06227_);
  nor (_06240_, _06238_, _06075_);
  not (_06241_, _06033_);
  nor (_06243_, _06203_, _06084_);
  nor (_06244_, _06196_, \oc8051_symbolic_cxrom1.regvalid [14]);
  not (_06245_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_06246_, _06209_, _06245_);
  nor (_06247_, _06246_, _06211_);
  nor (_06249_, _06247_, _06244_);
  nor (_06250_, _06218_, _06082_);
  nor (_06252_, _06250_, _06249_);
  not (_06253_, _06252_);
  nor (_06254_, _06253_, _06243_);
  nor (_06255_, _06254_, _06241_);
  nor (_06256_, _06203_, _06056_);
  nor (_06257_, _06197_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_06258_, _06038_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_06260_, _06209_, _06258_);
  not (_06261_, _06260_);
  nor (_06262_, _06261_, _06257_);
  nor (_06264_, _06218_, _06065_);
  nor (_06265_, _06264_, _06262_);
  not (_06267_, _06265_);
  nor (_06268_, _06267_, _06256_);
  nor (_06270_, _06268_, _06192_);
  nor (_06271_, _06270_, _06255_);
  not (_06272_, _06271_);
  nor (_06274_, _06272_, _06240_);
  not (_06275_, _06274_);
  nor (_06277_, _06275_, _06225_);
  not (_06278_, _06277_);
  nor (_06280_, _06091_, _06033_);
  nor (_06281_, _06027_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_06283_, _06026_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor (_06284_, _06283_, _06281_);
  nand (_06286_, _06284_, _06280_);
  not (_06287_, _06280_);
  nor (_06289_, _06027_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nor (_06290_, _06026_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor (_06291_, _06290_, _06289_);
  nand (_06292_, _06291_, _06287_);
  nand (_06293_, _06292_, _06286_);
  nand (_06294_, _06293_, _06217_);
  nor (_06295_, _06027_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nor (_06297_, _06026_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor (_06298_, _06297_, _06295_);
  not (_06300_, _06298_);
  nor (_06302_, _06300_, _06280_);
  nor (_06303_, _06027_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_06304_, _06026_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_06306_, _06304_, _06303_);
  not (_06307_, _06306_);
  nor (_06308_, _06307_, _06287_);
  nor (_06309_, _06308_, _06302_);
  nor (_06310_, _06309_, _06203_);
  nor (_06311_, _06209_, _06014_);
  nor (_06312_, _06027_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nor (_06313_, _06026_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nor (_06314_, _06313_, _06312_);
  nand (_06315_, _06314_, _06287_);
  nor (_06316_, _06027_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_06317_, _06026_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_06319_, _06317_, _06316_);
  nand (_06320_, _06319_, _06280_);
  nand (_06321_, _06320_, _06315_);
  nand (_06322_, _06321_, _06311_);
  nor (_06323_, _06027_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_06325_, _06026_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_06326_, _06325_, _06323_);
  nand (_06327_, _06326_, _06280_);
  nor (_06328_, _06027_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nor (_06329_, _06026_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nor (_06330_, _06329_, _06328_);
  nand (_06332_, _06330_, _06287_);
  nand (_06333_, _06332_, _06327_);
  nand (_06334_, _06333_, _06211_);
  nand (_06335_, _06334_, _06322_);
  nor (_06336_, _06335_, _06310_);
  nand (_06337_, _06336_, _06294_);
  nand (_06338_, _06337_, _06278_);
  nand (_06339_, _06277_, word_in[15]);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _06339_, _06338_);
  nor (_06341_, _06104_, _06089_);
  nor (_06342_, _06144_, _06038_);
  nor (_06343_, _06342_, _06341_);
  not (_06344_, _06343_);
  nor (_06345_, _06344_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_06346_, _06089_, _06020_);
  nor (_06347_, _06346_, _06129_);
  nor (_06348_, _06347_, _06258_);
  not (_06349_, _06348_);
  nor (_06351_, _06349_, _06345_);
  not (_06352_, _06347_);
  nor (_06353_, _06352_, _06343_);
  not (_06355_, _06353_);
  nor (_06356_, _06355_, _06065_);
  nor (_06358_, _06352_, _06344_);
  not (_06359_, _06358_);
  nor (_06361_, _06359_, _06056_);
  nor (_06362_, _06361_, _06356_);
  not (_06363_, _06362_);
  nor (_06364_, _06363_, _06351_);
  nor (_06365_, _06364_, _06191_);
  nor (_06366_, _06359_, _06084_);
  nor (_06367_, _06344_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_06368_, _06347_, _06077_);
  not (_06370_, _06368_);
  nor (_06371_, _06370_, _06367_);
  nor (_06372_, _06355_, _06082_);
  nor (_06373_, _06372_, _06371_);
  not (_06375_, _06373_);
  nor (_06376_, _06375_, _06366_);
  nor (_06377_, _06376_, _06075_);
  nor (_06378_, _06355_, _06101_);
  nor (_06379_, _06343_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_06381_, _06347_, _06038_);
  nor (_06382_, _06347_, _06103_);
  nor (_06384_, _06382_, _06381_);
  nor (_06385_, _06384_, _06379_);
  nor (_06387_, _06359_, _06095_);
  nor (_06388_, _06387_, _06385_);
  not (_06390_, _06388_);
  nor (_06391_, _06390_, _06378_);
  nor (_06392_, _06391_, _06241_);
  nor (_06393_, _06355_, _06045_);
  nor (_06394_, _06343_, \oc8051_symbolic_cxrom1.regvalid [13]);
  not (_06395_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_06396_, _06347_, _06395_);
  nor (_06397_, _06396_, _06381_);
  nor (_06398_, _06397_, _06394_);
  nor (_06400_, _06359_, _06226_);
  nor (_06401_, _06400_, _06398_);
  not (_06403_, _06401_);
  nor (_06404_, _06403_, _06393_);
  nor (_06405_, _06404_, _06192_);
  nor (_06406_, _06405_, _06392_);
  not (_06407_, _06406_);
  nor (_06409_, _06407_, _06377_);
  not (_06410_, _06409_);
  nor (_06411_, _06410_, _06365_);
  nand (_06412_, _06411_, word_in[23]);
  not (_06413_, _06411_);
  nor (_06414_, _06164_, _06031_);
  nor (_06415_, _06156_, _06089_);
  nor (_06417_, _06415_, _06414_);
  nand (_06418_, _06417_, _06347_);
  not (_06419_, _06346_);
  nor (_06420_, _06173_, _06419_);
  not (_06421_, _06180_);
  nor (_06423_, _06421_, _06130_);
  nor (_06424_, _06423_, _06420_);
  nand (_06425_, _06424_, _06418_);
  nand (_06426_, _06425_, _06343_);
  nand (_06427_, _06124_, _06031_);
  nand (_06428_, _06119_, _06089_);
  nand (_06429_, _06428_, _06427_);
  nand (_06430_, _06429_, _06347_);
  nor (_06431_, _06419_, _06137_);
  nor (_06433_, _06143_, _06130_);
  nor (_06434_, _06433_, _06431_);
  nand (_06436_, _06434_, _06430_);
  nand (_06437_, _06436_, _06344_);
  nand (_06439_, _06437_, _06426_);
  nand (_06440_, _06439_, _06413_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _06440_, _06412_);
  nor (_06442_, _06074_, _06021_);
  nor (_06443_, _06075_, _06020_);
  nor (_06444_, _06443_, _06442_);
  not (_06445_, _06444_);
  not (_06446_, _06442_);
  nor (_06447_, _06446_, _06038_);
  nor (_06448_, _06442_, _06014_);
  nor (_06449_, _06448_, _06447_);
  nor (_06450_, _06449_, _06103_);
  not (_06451_, _06449_);
  nor (_06452_, _06451_, _06097_);
  nor (_06454_, _06452_, _06450_);
  nor (_06455_, _06454_, _06445_);
  nor (_06457_, _06449_, _06095_);
  nor (_06458_, _06451_, _06101_);
  nor (_06460_, _06458_, _06457_);
  nor (_06461_, _06460_, _06444_);
  nor (_06462_, _06461_, _06455_);
  nor (_06464_, _06462_, _06075_);
  nor (_06465_, _06449_, _06226_);
  nor (_06466_, _06451_, _06045_);
  nor (_06468_, _06466_, _06465_);
  nor (_06471_, _06468_, _06444_);
  nor (_06473_, _06451_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_06474_, _06445_, _06041_);
  not (_06476_, _06474_);
  nor (_06477_, _06476_, _06473_);
  nor (_06479_, _06477_, _06471_);
  nor (_06481_, _06479_, _06191_);
  nor (_06482_, _06449_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_06483_, _06445_, _06258_);
  not (_06485_, _06483_);
  nor (_06487_, _06485_, _06482_);
  nor (_06489_, _06449_, _06056_);
  nor (_06490_, _06451_, _06065_);
  nor (_06491_, _06490_, _06489_);
  nor (_06492_, _06491_, _06444_);
  nor (_06493_, _06492_, _06487_);
  nor (_06494_, _06493_, _06241_);
  nor (_06495_, _06449_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_06497_, _06445_, _06077_);
  not (_06498_, _06497_);
  nor (_06499_, _06498_, _06495_);
  nor (_06501_, _06449_, _06084_);
  nor (_06502_, _06451_, _06082_);
  nor (_06504_, _06502_, _06501_);
  nor (_06505_, _06504_, _06444_);
  nor (_06506_, _06505_, _06499_);
  nor (_06507_, _06506_, _06192_);
  nor (_06508_, _06507_, _06494_);
  not (_06509_, _06508_);
  nor (_06510_, _06509_, _06481_);
  not (_06512_, _06510_);
  nor (_06513_, _06512_, _06464_);
  not (_06514_, _06513_);
  nand (_06516_, _06330_, _06280_);
  nand (_06517_, _06326_, _06287_);
  nand (_06519_, _06517_, _06516_);
  nand (_06520_, _06519_, _06444_);
  nand (_06522_, _06284_, _06287_);
  nand (_06524_, _06291_, _06280_);
  nand (_06526_, _06524_, _06522_);
  nand (_06527_, _06526_, _06445_);
  nand (_06529_, _06527_, _06520_);
  nand (_06531_, _06529_, _06449_);
  nand (_06533_, _06314_, _06280_);
  nand (_06534_, _06319_, _06287_);
  nand (_06535_, _06534_, _06533_);
  nand (_06536_, _06535_, _06444_);
  nand (_06538_, _06306_, _06287_);
  nand (_06539_, _06298_, _06280_);
  nand (_06541_, _06539_, _06538_);
  nand (_06543_, _06541_, _06445_);
  nand (_06544_, _06543_, _06536_);
  nand (_06546_, _06544_, _06451_);
  nand (_06547_, _06546_, _06531_);
  nand (_06549_, _06547_, _06514_);
  nand (_06551_, _06513_, word_in[31]);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _06551_, _06549_);
  nor (_06553_, _22454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  nor (_06555_, _22456_, _21554_);
  nor (_25086_, _06555_, _06553_);
  nor (_06556_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand (_06557_, _23553_, _23048_);
  nand (_06558_, _06557_, _23493_);
  nor (_23916_, _06558_, _06556_);
  nor (_06561_, _21777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  nor (_06562_, _21779_, _21414_);
  nor (_25219_, _06562_, _06561_);
  nor (_06563_, _24050_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  nor (_06564_, _24052_, _21526_);
  nor (_25364_, _06564_, _06563_);
  nor (_06566_, _06514_, rst);
  not (_06568_, _06566_);
  nor (_06569_, _06568_, _06451_);
  not (_06570_, _06569_);
  nor (_06571_, _06570_, _06445_);
  not (_06572_, _06571_);
  nor (_06573_, _06572_, _06075_);
  not (_06574_, _06573_);
  nor (_06575_, _06413_, rst);
  nand (_06576_, _06575_, _06381_);
  nor (_06577_, _06576_, _06241_);
  nor (_06578_, _06278_, rst);
  not (_06579_, _06578_);
  nor (_06581_, _06579_, _06209_);
  nand (_06583_, _06581_, _06197_);
  nor (_06585_, _06583_, _06191_);
  nor (_06587_, _06192_, _06098_);
  not (_06589_, _06587_);
  nor (_06590_, _06116_, rst);
  not (_06591_, _06590_);
  nor (_06592_, _06591_, _06589_);
  nor (_06593_, _06592_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  not (_06595_, _06592_);
  nor (_06596_, _06595_, word_in[7]);
  nor (_06597_, _06596_, _06593_);
  nor (_06598_, _06597_, _06585_);
  not (_06599_, _06585_);
  nor (_06600_, _06339_, rst);
  nor (_06601_, _06600_, _06599_);
  nor (_06603_, _06601_, _06598_);
  nor (_06604_, _06603_, _06577_);
  not (_06605_, _06577_);
  nor (_06606_, _06412_, rst);
  nor (_06607_, _06606_, _06605_);
  nor (_06608_, _06607_, _06604_);
  nand (_06609_, _06608_, _06574_);
  nor (_06610_, _06551_, rst);
  nand (_06611_, _06610_, _06573_);
  nand (_25008_[7], _06611_, _06609_);
  not (_06612_, _06443_);
  nor (_06613_, _06612_, _06014_);
  not (_06614_, _06447_);
  nand (_06615_, _06614_, _06056_);
  nor (_06616_, _06615_, _06613_);
  nor (_24964_[0], _06616_, rst);
  nor (_06617_, _06358_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_24964_[1], _06617_, rst);
  not (_06618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  not (_06619_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nand (_06620_, _06619_, _06618_);
  nor (_06621_, _06620_, _00930_);
  nor (_06622_, _02481_, _00008_);
  nand (_06624_, _06622_, _24904_);
  nand (_06625_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nor (_06626_, _05559_, _21507_);
  not (_06627_, _06626_);
  nand (_06628_, _06627_, _06625_);
  nor (_06629_, _06628_, _06624_);
  nor (_06630_, _06629_, _06621_);
  nor (_06631_, _06630_, _00928_);
  nand (_06633_, _00928_, _00106_);
  nand (_06634_, _06633_, _23493_);
  nor (_23986_, _06634_, _06631_);
  nor (_06635_, _05952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1]);
  nor (_06636_, _05954_, _21474_);
  nor (_23988_, _06636_, _06635_);
  nor (_06637_, _00955_, _00943_);
  nand (_06638_, _06637_, _00996_);
  nor (_06639_, _06638_, _00983_);
  nor (_06640_, _06639_, _01240_);
  nand (_06641_, _01240_, _06619_);
  nand (_06642_, _06641_, _23493_);
  nor (_23995_, _06642_, _06640_);
  nor (_06643_, _05952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  nor (_06644_, _05954_, _21586_);
  nor (_24001_, _06644_, _06643_);
  nor (_06645_, _00981_, _00955_);
  nor (_06646_, _06645_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  not (_06647_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor (_06648_, _00944_, _06647_);
  nor (_06650_, _06648_, _00985_);
  nor (_06651_, _06650_, _06646_);
  nor (_06652_, _06651_, _00991_);
  nand (_06653_, _00991_, _06647_);
  nand (_06654_, _06653_, _01006_);
  nor (_06655_, _06654_, _06652_);
  nor (_06657_, _01013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor (_06658_, _06657_, _01239_);
  nor (_06659_, _06658_, _06655_);
  nand (_06660_, _01013_, _00106_);
  nand (_06661_, _06660_, _23493_);
  nor (_24007_, _06661_, _06659_);
  nand (_06663_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor (_06664_, _06663_, _00985_);
  not (_06666_, _00973_);
  nand (_06667_, _06666_, _00954_);
  nand (_06668_, _06667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor (_06669_, _06667_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor (_06670_, _06669_, _00991_);
  nand (_06671_, _06670_, _06668_);
  nor (_06673_, _06671_, _06664_);
  nand (_06674_, _00991_, _02513_);
  nand (_06675_, _06674_, _01006_);
  nor (_06676_, _06675_, _06673_);
  nor (_06678_, _01013_, ABINPUT[10]);
  nor (_06679_, _06678_, _01239_);
  nor (_06680_, _06679_, _06676_);
  nand (_06682_, _01013_, _00959_);
  nand (_06683_, _06682_, _23493_);
  nor (_24009_, _06683_, _06680_);
  nor (_06684_, _06145_, _06038_);
  nor (_06685_, _06059_, _06031_);
  nor (_06686_, _06685_, _06587_);
  not (_06687_, _06686_);
  nor (_06688_, _06191_, _06059_);
  nor (_06689_, _06688_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_06690_, _06689_, _06687_);
  nor (_06691_, _06690_, _06036_);
  nor (_06692_, _06691_, _06684_);
  nor (_06693_, _06613_, _06587_);
  nor (_06694_, _06191_, _06098_);
  not (_06695_, _06690_);
  nand (_06696_, _06027_, _06084_);
  nand (_06698_, _06696_, _06685_);
  nand (_06699_, _06698_, _06695_);
  nand (_06700_, _06699_, _06694_);
  nand (_06701_, _06700_, _06693_);
  nor (_06702_, _06701_, _06692_);
  nor (_24964_[2], _06702_, rst);
  not (_06703_, _00983_);
  nor (_06704_, _00955_, _00942_);
  nand (_06705_, _06704_, _01239_);
  nor (_06706_, _06705_, _06703_);
  not (_06708_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  nand (_06709_, _06705_, _06708_);
  nand (_06710_, _06709_, _23493_);
  nor (_24024_, _06710_, _06706_);
  nor (_06711_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  nor (_06712_, _02331_, _21586_);
  nor (_24037_, _06712_, _06711_);
  nor (_06714_, _01042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor (_06715_, _01044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nor (_06716_, _06715_, _06714_);
  nor (_06718_, _06716_, _01037_);
  nand (_06719_, _01037_, _00106_);
  nand (_06720_, _06719_, _23493_);
  nor (_24040_, _06720_, _06718_);
  not (_06721_, _06036_);
  nor (_06723_, _06192_, _06059_);
  not (_06725_, _06723_);
  nand (_06727_, _06725_, _06095_);
  nand (_06729_, _06727_, _06203_);
  nor (_06731_, _06721_, _06095_);
  nor (_06733_, _06731_, _06688_);
  nand (_06734_, _06733_, _06729_);
  nand (_06735_, _06734_, _06359_);
  nand (_06736_, _06735_, _06721_);
  not (_06738_, _06613_);
  nand (_06739_, _06727_, _06684_);
  nand (_06740_, _06739_, _06738_);
  nor (_06741_, _06740_, _06736_);
  nor (_24964_[3], _06741_, rst);
  nor (_06742_, _21430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  nor (_06743_, _21432_, _21414_);
  nor (_24047_, _06743_, _06742_);
  nor (_06745_, _01233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7]);
  nor (_06746_, _01235_, _21626_);
  nor (_24056_, _06746_, _06745_);
  not (_06747_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not (_06748_, _06448_);
  nor (_06750_, _06748_, _06111_);
  nor (_06751_, _06750_, _06747_);
  nor (_06752_, _06075_, _06104_);
  not (_06753_, _06752_);
  nand (_06754_, _06199_, _06038_);
  not (_06755_, _06754_);
  nand (_06756_, _06755_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nand (_06757_, _06756_, _06753_);
  nor (_06758_, _06757_, _06751_);
  nor (_06759_, _06758_, _06057_);
  nand (_06760_, _06287_, _06057_);
  not (_06761_, _06760_);
  not (_06762_, _06685_);
  nor (_06763_, _06762_, _06747_);
  nor (_06765_, _06763_, _06761_);
  nand (_06766_, _06765_, _06725_);
  nor (_06767_, _06766_, _06759_);
  nor (_24964_[4], _06767_, rst);
  nor (_06768_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  nor (_06769_, _02331_, _21526_);
  nor (_25330_, _06769_, _06768_);
  nor (_06770_, _22450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  nor (_06771_, _22452_, _21526_);
  nor (_25088_, _06771_, _06770_);
  nor (_06772_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  nor (_06773_, _02331_, _21554_);
  nor (_25329_, _06773_, _06772_);
  nor (_06774_, _22450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  nor (_06775_, _22452_, _21586_);
  nor (_24093_, _06775_, _06774_);
  nor (_06777_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7]);
  nor (_06778_, _22569_, _21626_);
  nor (_24099_, _06778_, _06777_);
  nor (_06780_, _06194_, _06068_);
  nor (_06781_, _06104_, _06241_);
  nor (_06782_, _06781_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_06783_, _06074_, _06104_);
  nor (_06784_, _06783_, _06194_);
  nor (_06785_, _06784_, _06782_);
  nor (_06786_, _06721_, _06395_);
  not (_06787_, _06786_);
  nand (_06789_, _06787_, _06753_);
  nor (_06791_, _06789_, _06785_);
  nor (_06792_, _06791_, _06780_);
  not (_06793_, _06782_);
  nand (_06794_, _06793_, _06587_);
  nand (_06796_, _06613_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_06797_, _06786_, _06688_);
  nand (_06798_, _06797_, _06796_);
  nor (_06800_, _06798_, _06723_);
  nand (_06802_, _06800_, _06794_);
  nor (_06803_, _06802_, _06792_);
  nor (_24964_[5], _06803_, rst);
  nor (_06804_, _01233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  nor (_06805_, _01235_, _21526_);
  nor (_24114_, _06805_, _06804_);
  nor (_06806_, _01233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  nor (_06807_, _01235_, _21554_);
  nor (_24116_, _06807_, _06806_);
  nor (_06809_, _01233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1]);
  nor (_06810_, _01235_, _21474_);
  nor (_24124_, _06810_, _06809_);
  nor (_06811_, _01233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  nor (_06812_, _01235_, _21414_);
  nor (_24139_, _06812_, _06811_);
  nor (_06814_, _01233_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5]);
  nor (_06815_, _01235_, _21451_);
  nor (_24141_, _06815_, _06814_);
  nor (_06816_, _06754_, _06245_);
  nor (_06817_, _06816_, _06723_);
  nand (_06818_, _06817_, _06753_);
  not (_06819_, _06781_);
  nand (_06820_, _06145_, _06038_);
  nor (_06821_, _06191_, _06104_);
  not (_06822_, _06821_);
  nand (_06823_, _06027_, _06038_);
  nor (_06824_, _06057_, _06245_);
  nand (_06825_, _06824_, _06823_);
  nand (_06826_, _06825_, _06822_);
  nand (_06827_, _06826_, _06820_);
  nand (_06829_, _06827_, _06819_);
  nor (_06830_, _06829_, _06818_);
  nor (_24964_[6], _06830_, rst);
  nor (_06831_, _01183_, _21558_);
  nor (_06833_, _06831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5]);
  not (_06834_, _06831_);
  nor (_06836_, _06834_, _21451_);
  nor (_24182_, _06836_, _06833_);
  nor (_06838_, _06038_, _06103_);
  nor (_06839_, _06725_, _06103_);
  nor (_06841_, _06839_, _06752_);
  nand (_06842_, _06755_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand (_06844_, _06842_, _06841_);
  nor (_06845_, _06844_, _06341_);
  nand (_06846_, _06845_, _06819_);
  nor (_06847_, _06846_, _06838_);
  nor (_24964_[7], _06847_, rst);
  nor (_06848_, _06831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  nor (_06849_, _06834_, _21414_);
  nor (_25324_, _06849_, _06848_);
  nor (_06850_, _06831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7]);
  nor (_06851_, _06834_, _21626_);
  nor (_25326_, _06851_, _06850_);
  nor (_06853_, _21430_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  nor (_06854_, _21504_, _21432_);
  nor (_24228_, _06854_, _06853_);
  nor (_06856_, _06748_, _06065_);
  not (_06858_, _06783_);
  nor (_06859_, _06612_, _06038_);
  not (_06860_, _06859_);
  nand (_06861_, _06860_, _06065_);
  nand (_06862_, _06861_, _06014_);
  nand (_06864_, _06862_, _06858_);
  nor (_06865_, _06864_, _06856_);
  nor (_24964_[8], _06865_, rst);
  nor (_06868_, _06831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  nor (_06869_, _06834_, _21586_);
  nor (_24237_, _06869_, _06868_);
  nor (_06871_, _22557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5]);
  nor (_06873_, _22559_, _21451_);
  nor (_24259_, _06873_, _06871_);
  nor (_06874_, _06831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  nor (_06875_, _06834_, _21554_);
  nor (_24262_, _06875_, _06874_);
  nor (_06876_, _22403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  nor (_06877_, _22406_, _21414_);
  nor (_24270_, _06877_, _06876_);
  nor (_06878_, _06443_, _06038_);
  nand (_06879_, _06038_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nand (_06880_, _06034_, _06045_);
  nand (_06881_, _06880_, _06014_);
  nand (_06882_, _06881_, _06879_);
  nand (_06883_, _06882_, _06878_);
  nor (_06884_, _06752_, _06723_);
  nand (_06885_, _06760_, _06884_);
  nand (_06886_, _06885_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_06887_, _06738_, _06045_);
  nand (_06888_, _06781_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nand (_06889_, _06888_, _06822_);
  nor (_06890_, _06889_, _06887_);
  nand (_06891_, _06890_, _06886_);
  nor (_06892_, _06891_, _06859_);
  nand (_06893_, _06892_, _06883_);
  nor (_06894_, _06893_, _06195_);
  nor (_24964_[9], _06894_, rst);
  nor (_06895_, _02427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  nor (_06896_, _02430_, _21554_);
  nor (_24281_, _06896_, _06895_);
  nor (_06897_, _02427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1]);
  nor (_06898_, _02430_, _21474_);
  nor (_24285_, _06898_, _06897_);
  nor (_06900_, _02427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  nor (_06901_, _02430_, _21586_);
  nor (_25320_, _06901_, _06900_);
  nor (_06902_, _02427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5]);
  nor (_06903_, _02430_, _21451_);
  nor (_24311_, _06903_, _06902_);
  nor (_06904_, _02427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  nor (_06905_, _02430_, _21414_);
  nor (_25321_, _06905_, _06904_);
  nor (_06906_, _02427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  nor (_06907_, _02430_, _21526_);
  nor (_24321_, _06907_, _06906_);
  not (_06908_, t2_i);
  nor (_24323_, rst, _06908_);
  nor (_06909_, _06034_, _06038_);
  not (_06910_, _06909_);
  nand (_06911_, _06910_, _06860_);
  nor (_06912_, _06347_, _06014_);
  not (_06913_, _06912_);
  nor (_06914_, _06913_, _06082_);
  not (_06915_, _06195_);
  nand (_06916_, _06762_, _06822_);
  nand (_06918_, _06916_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand (_06919_, _06918_, _06915_);
  nor (_06920_, _06919_, _06914_);
  nor (_06922_, _06381_, _06694_);
  nand (_06923_, _06922_, _06589_);
  nor (_06924_, _06760_, _06082_);
  nand (_06925_, _06613_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_06926_, _06191_, _06048_);
  not (_06927_, _06926_);
  nand (_06928_, _06927_, _06925_);
  nor (_06929_, _06928_, _06924_);
  nand (_06931_, _06859_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand (_06932_, _06195_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand (_06933_, _06932_, _06931_);
  nand (_06934_, _06311_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_06935_, _06026_, _06020_);
  nor (_06936_, _06935_, _06082_);
  nand (_06937_, _06936_, _06014_);
  nand (_06938_, _06937_, _06934_);
  nor (_06939_, _06938_, _06933_);
  nand (_06940_, _06939_, _06929_);
  nand (_06941_, _06940_, _06923_);
  nand (_06942_, _06941_, _06920_);
  nor (_06943_, _06942_, _06911_);
  nor (_24964_[10], _06943_, rst);
  nor (_06945_, _01183_, _21864_);
  nor (_06946_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1]);
  not (_06947_, _06945_);
  nor (_06948_, _06947_, _21474_);
  nor (_24334_, _06948_, _06946_);
  nor (_06949_, _21632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1]);
  nor (_06950_, _21635_, _21474_);
  nor (_24339_, _06950_, _06949_);
  nor (_06951_, _01198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  nor (_06952_, _01200_, _21526_);
  nor (_24341_, _06952_, _06951_);
  nor (_06954_, _01198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  nor (_06955_, _01200_, _21554_);
  nor (_25319_, _06955_, _06954_);
  nor (_06956_, _22500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  nor (_06957_, _22502_, _21504_);
  nor (_24347_, _06957_, _06956_);
  nor (_06958_, _01198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1]);
  nor (_06959_, _01200_, _21474_);
  nor (_24354_, _06959_, _06958_);
  not (_06960_, t2ex_i);
  nor (_24356_, rst, _06960_);
  nand (_06961_, _06960_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  nor (_24358_, _06961_, rst);
  nor (_06962_, _02383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1]);
  nor (_06963_, _02385_, _21474_);
  nor (_25310_, _06963_, _06962_);
  nor (_06964_, _01198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  nor (_06966_, _01200_, _21414_);
  nor (_24371_, _06966_, _06964_);
  nor (_06967_, _01198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  nor (_06968_, _01200_, _21504_);
  nor (_24374_, _06968_, _06967_);
  nor (_06969_, _01198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5]);
  nor (_06970_, _01200_, _21451_);
  nor (_24377_, _06970_, _06969_);
  nor (_06971_, _01183_, _21374_);
  nor (_06972_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  not (_06973_, _06971_);
  nor (_06974_, _06973_, _21504_);
  nor (_24388_, _06974_, _06972_);
  nand (_06975_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _06908_);
  nor (_24392_, _06975_, rst);
  nor (_06976_, _06192_, _06048_);
  nor (_06977_, _06976_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_06978_, _06910_, _06101_);
  nor (_06979_, _06978_, _06211_);
  nor (_06980_, _06979_, _06977_);
  not (_06981_, _06311_);
  nor (_06982_, _06981_, _06101_);
  not (_06983_, _06982_);
  nor (_06984_, _06915_, _06101_);
  nor (_06985_, _06984_, _06926_);
  nand (_06986_, _06985_, _06983_);
  nor (_06988_, _06986_, _06980_);
  nor (_06990_, _06988_, _06922_);
  not (_06991_, _06693_);
  nand (_06992_, _06991_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_06993_, _06984_, _06859_);
  nor (_06994_, _06760_, _06101_);
  nor (_06995_, _06994_, _06982_);
  nand (_06996_, _06995_, _06993_);
  nor (_06999_, _06996_, _06909_);
  nand (_07000_, _06999_, _06992_);
  nor (_07001_, _07000_, _06990_);
  nor (_24964_[11], _07001_, rst);
  nor (_07002_, _01183_, _21599_);
  nor (_07003_, _07002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  not (_07004_, _07002_);
  nor (_07005_, _07004_, _21526_);
  nor (_24415_, _07005_, _07003_);
  nor (_07006_, _07002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  nor (_07008_, _07004_, _21554_);
  nor (_24418_, _07008_, _07006_);
  nor (_07009_, _07002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1]);
  nor (_07010_, _07004_, _21474_);
  nor (_25315_, _07010_, _07009_);
  nor (_07011_, _23044_, _21345_);
  not (_07012_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2]);
  nor (_07013_, _23153_, _07012_);
  nor (_07015_, _23050_, _00506_);
  nor (_07016_, _23076_, _23217_);
  nor (_07018_, _07016_, _07015_);
  not (_07019_, _07018_);
  nor (_07020_, _23073_, _05345_);
  nor (_07021_, _23107_, _23215_);
  nor (_07022_, _07021_, _07020_);
  nor (_07023_, _23067_, _23212_);
  nor (_07024_, _23058_, _23210_);
  nor (_07025_, _07024_, _07023_);
  nand (_07026_, _07025_, _07022_);
  nor (_07027_, _07026_, _07019_);
  nor (_07028_, _07027_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_07029_, _07028_, _07013_);
  nor (_07030_, _07029_, _23490_);
  nor (_07031_, _07030_, _07011_);
  nor (_25039_[2], _07031_, rst);
  nor (_07032_, _07002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  nor (_07033_, _07004_, _21504_);
  nor (_25318_, _07033_, _07032_);
  nor (_07034_, _07002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5]);
  nor (_07035_, _07004_, _21451_);
  nor (_25317_, _07035_, _07034_);
  nor (_07037_, _07002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  nor (_07038_, _07004_, _21414_);
  nor (_25316_, _07038_, _07037_);
  nor (_07039_, _06098_, _06241_);
  not (_07040_, _07039_);
  nand (_07041_, _07040_, _06381_);
  nand (_07042_, _07041_, _06910_);
  not (_07043_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_07044_, _06443_, _06036_);
  nor (_07045_, _07044_, _07043_);
  nor (_07046_, _06419_, _06014_);
  nor (_07047_, _07046_, _06068_);
  nand (_07048_, _07047_, _06614_);
  nor (_07049_, _07048_, _07045_);
  nor (_07051_, _07049_, _07043_);
  nor (_07052_, _07051_, _07042_);
  nor (_24964_[12], _07052_, rst);
  nor (_07053_, _02383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  nor (_07054_, _02385_, _21526_);
  nor (_25311_, _07054_, _07053_);
  nor (_07056_, _22500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  nor (_07057_, _22502_, _21554_);
  nor (_25059_, _07057_, _07056_);
  nor (_07058_, _21632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  nor (_07059_, _21635_, _21414_);
  nor (_25261_, _07059_, _07058_);
  nor (_07061_, _21690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5]);
  nor (_07062_, _21692_, _21451_);
  nor (_25266_, _07062_, _07061_);
  nor (_07063_, _21690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7]);
  nor (_07064_, _21692_, _21626_);
  nor (_25268_, _07064_, _07063_);
  nor (_07065_, _02383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7]);
  nor (_07066_, _02385_, _21626_);
  nor (_25314_, _07066_, _07065_);
  nor (_07067_, _02383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  nor (_07068_, _02385_, _21504_);
  nor (_25313_, _07068_, _07067_);
  nor (_07069_, _02383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5]);
  nor (_07071_, _02385_, _21451_);
  nor (_25312_, _07071_, _07069_);
  nor (_07072_, _22227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  nor (_07073_, _22229_, _21504_);
  nor (_25179_, _07073_, _07072_);
  nor (_07074_, _21752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  nor (_07075_, _21754_, _21414_);
  nor (_25236_, _07075_, _07074_);
  nor (_07076_, _06381_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_24964_[13], _07076_, rst);
  nor (_07077_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5]);
  nor (_07079_, _06947_, _21451_);
  nor (_25306_, _07079_, _07077_);
  nor (_07081_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  not (_07082_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand (_07083_, _23553_, _07082_);
  nand (_07085_, _07083_, _23493_);
  nor (_25042_[27], _07085_, _07081_);
  nor (_07086_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  nor (_07087_, _06947_, _21414_);
  nor (_25305_, _07087_, _07086_);
  nor (_07088_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  nor (_07089_, _06947_, _21526_);
  nor (_25304_, _07089_, _07088_);
  nor (_07090_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  nor (_07091_, _06947_, _21554_);
  nor (_25303_, _07091_, _07090_);
  nor (_07093_, _00713_, _00690_);
  nor (_07095_, _23143_, _00704_);
  nor (_07097_, _00698_, _07095_);
  not (_07098_, _07097_);
  nor (_07099_, _07098_, _00702_);
  nand (_07100_, _07099_, _07093_);
  nor (_07101_, _00711_, _23245_);
  nor (_07102_, _00699_, _00687_);
  nand (_07103_, _07102_, _07101_);
  nand (_07104_, _07103_, _07100_);
  nor (_07105_, _23400_, _23320_);
  not (_07106_, _07105_);
  nor (_07107_, _07106_, _00699_);
  nand (_07108_, _07107_, _00693_);
  nor (_07109_, _23302_, _23320_);
  not (_07110_, _07109_);
  nor (_07111_, _07110_, _23143_);
  not (_07112_, _07111_);
  nor (_07113_, _23199_, _23084_);
  not (_07114_, _07113_);
  nor (_07115_, _07114_, _07112_);
  not (_07116_, _07115_);
  nand (_07117_, _07116_, _07108_);
  nor (_07118_, _07117_, _07104_);
  not (_07119_, _07093_);
  nor (_07120_, _07119_, _23084_);
  not (_07121_, _07120_);
  nor (_07122_, _07121_, _07106_);
  nor (_07124_, _23245_, _23170_);
  not (_07125_, _07124_);
  nor (_07126_, _07125_, _00690_);
  not (_07127_, _07126_);
  nand (_07128_, _07127_, _00694_);
  nor (_07129_, _07128_, _07122_);
  nand (_07130_, _07129_, _07118_);
  nor (_07131_, _07106_, _00706_);
  not (_07132_, _07131_);
  nor (_07133_, _07132_, _07119_);
  nor (_07134_, _07125_, _00711_);
  not (_07135_, _07134_);
  nor (_07136_, _23143_, _23084_);
  not (_07138_, _07136_);
  nor (_07139_, _07110_, _07138_);
  not (_07140_, _07139_);
  nor (_07141_, _07140_, _07135_);
  not (_07142_, _07141_);
  nor (_07143_, _07110_, _00697_);
  nand (_07144_, _07143_, _00691_);
  nand (_07145_, _07144_, _07142_);
  nor (_07146_, _07145_, _07133_);
  nand (_07147_, _07146_, _00718_);
  nor (_07148_, _07147_, _07130_);
  not (_07149_, _07095_);
  nor (_07151_, _07149_, _00687_);
  not (_07153_, _07151_);
  nor (_07154_, _07106_, _07149_);
  nor (_07156_, _07154_, _00703_);
  nand (_07157_, _07156_, _07153_);
  nor (_07158_, _07157_, _07143_);
  nor (_07159_, _07158_, _07119_);
  nor (_07160_, _00702_, _23143_);
  nand (_07161_, _07160_, _00695_);
  not (_07162_, _07161_);
  nor (_07163_, _00687_, _00697_);
  not (_07164_, _07163_);
  nor (_07165_, _00711_, _23277_);
  not (_07166_, _07165_);
  nor (_07167_, _07166_, _23084_);
  nor (_07168_, _07167_, _07113_);
  nor (_07169_, _07168_, _07164_);
  nor (_07170_, _07169_, _07162_);
  not (_07171_, _07170_);
  nor (_07172_, _07171_, _07159_);
  nand (_07173_, _07172_, _07148_);
  nand (_07174_, _07173_, _23046_);
  nor (_07175_, _00685_, _23496_);
  nor (_07176_, _07175_, rst);
  nand (_25018_[1], _07176_, _07174_);
  nor (_07177_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  nand (_07178_, _23553_, _24180_);
  nand (_07179_, _07178_, _23493_);
  nor (_25042_[28], _07179_, _07177_);
  nor (_07180_, _21632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5]);
  nor (_07182_, _21635_, _21451_);
  nor (_25262_, _07182_, _07180_);
  nor (_07183_, _02383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  nor (_07184_, _02385_, _21586_);
  nor (_25309_, _07184_, _07183_);
  nor (_07185_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7]);
  nor (_07187_, _06947_, _21626_);
  nor (_25308_, _07187_, _07185_);
  nor (_07188_, _21653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  nor (_07189_, _21655_, _21586_);
  nor (_25269_, _07189_, _07188_);
  nor (_07191_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  nor (_07192_, _06947_, _21504_);
  nor (_25307_, _07192_, _07191_);
  nor (_07193_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  nand (_07194_, _23553_, _01337_);
  nand (_07195_, _07194_, _23493_);
  nor (_25042_[29], _07195_, _07193_);
  nor (_07197_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  nand (_07198_, _23553_, _02288_);
  nand (_07200_, _07198_, _23493_);
  nor (_25042_[30], _07200_, _07197_);
  not (_07201_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nand (_07202_, _06192_, _06062_);
  nand (_07203_, _07202_, _07201_);
  nor (_07204_, _07203_, _06976_);
  nor (_24964_[14], _07204_, rst);
  nor (_07206_, _21632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7]);
  nor (_07207_, _21635_, _21626_);
  nor (_25263_, _07207_, _07206_);
  nor (_07208_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5]);
  nor (_07209_, _06973_, _21451_);
  nor (_25301_, _07209_, _07208_);
  nor (_07210_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  nor (_07211_, _22569_, _21504_);
  nor (_25058_, _07211_, _07210_);
  nor (_07212_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  nor (_07213_, _06973_, _21414_);
  nor (_25300_, _07213_, _07212_);
  nor (_07215_, _22162_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  nor (_07216_, _22165_, _21414_);
  nor (_25071_, _07216_, _07215_);
  nor (_07217_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7]);
  nor (_07218_, _06973_, _21626_);
  nor (_25302_, _07218_, _07217_);
  nor (_07219_, _06945_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  nor (_07220_, _06947_, _21586_);
  nor (_24639_, _07220_, _07219_);
  nor (_07221_, _21690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  nor (_07222_, _21692_, _21586_);
  nor (_25264_, _07222_, _07221_);
  nor (_07224_, _21690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  nor (_07225_, _21692_, _21526_);
  nor (_25265_, _07225_, _07224_);
  nor (_07226_, _01183_, _21658_);
  nor (_07227_, _07226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  not (_07228_, _07226_);
  nor (_07229_, _07228_, _21504_);
  nor (_24656_, _07229_, _07227_);
  nor (_07230_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  nor (_07231_, _06973_, _21586_);
  nor (_24658_, _07231_, _07230_);
  nor (_07232_, _07226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7]);
  nor (_07233_, _07228_, _21626_);
  nor (_24660_, _07233_, _07232_);
  nor (_07234_, _21741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  nor (_07235_, _21744_, _21586_);
  nor (_24664_, _07235_, _07234_);
  nor (_07236_, _06062_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_24964_[15], _07236_, rst);
  nor (_07238_, _22693_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7]);
  nor (_07239_, _22696_, _21626_);
  nor (_24772_, _07239_, _07238_);
  nor (_07240_, _22396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7]);
  nor (_07241_, _22398_, _21626_);
  nor (_24787_, _07241_, _07240_);
  nor (_07243_, _05519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1]);
  nor (_07244_, _05521_, _21474_);
  nor (_24806_, _07244_, _07243_);
  nor (_07246_, _02416_, _02403_);
  nor (_07248_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nand (_07249_, _02407_, _02405_);
  nor (_07251_, _07249_, _07248_);
  nor (_07252_, _07251_, _07246_);
  nor (_24825_, _07252_, rst);
  nor (_07254_, _02407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nand (_07255_, _02416_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nand (_07256_, _07255_, _23493_);
  nor (_24846_, _07256_, _07254_);
  not (_07257_, _06694_);
  not (_07258_, _06575_);
  nor (_07259_, _07258_, _07257_);
  not (_07260_, _07259_);
  nor (_07261_, _06579_, _06589_);
  not (_07262_, _07261_);
  not (_07263_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_07264_, _06591_, _06738_);
  not (_07265_, _07264_);
  nand (_07266_, _07265_, _07263_);
  not (_07267_, word_in[0]);
  nand (_07268_, _07264_, _07267_);
  nand (_07270_, _07268_, _07266_);
  nand (_07271_, _07270_, _07262_);
  not (_07272_, word_in[8]);
  nand (_07273_, _07261_, _07272_);
  nand (_07274_, _07273_, _07271_);
  nand (_07275_, _07274_, _07260_);
  nor (_07276_, _06568_, _06445_);
  nor (_07277_, _07276_, _06569_);
  nor (_07278_, _06568_, _06241_);
  nand (_07280_, _07278_, _07277_);
  not (_07281_, _07280_);
  nor (_07283_, _07260_, word_in[16]);
  nor (_07284_, _07283_, _07281_);
  nand (_07285_, _07284_, _07275_);
  nand (_07286_, _07281_, word_in[24]);
  nand (_25005_[0], _07286_, _07285_);
  nor (_07287_, _07264_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_07288_, _07265_, word_in[1]);
  nor (_07289_, _07288_, _07287_);
  nand (_07290_, _07289_, _07262_);
  nand (_07291_, _06277_, word_in[9]);
  nor (_07292_, _07291_, rst);
  nand (_07293_, _07292_, _06587_);
  nand (_07294_, _07293_, _07290_);
  nor (_07295_, _07294_, _07259_);
  nor (_07296_, _07260_, word_in[17]);
  nor (_07297_, _07296_, _07295_);
  nand (_07298_, _07297_, _07280_);
  nand (_07299_, _07281_, word_in[25]);
  nand (_25005_[1], _07299_, _07298_);
  not (_07300_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand (_07301_, _07265_, _07300_);
  not (_07303_, word_in[2]);
  nand (_07304_, _07264_, _07303_);
  nand (_07305_, _07304_, _07301_);
  nand (_07306_, _07305_, _07262_);
  not (_07307_, word_in[10]);
  nand (_07308_, _07261_, _07307_);
  nand (_07309_, _07308_, _07306_);
  nand (_07310_, _07309_, _07260_);
  nor (_07311_, _07260_, word_in[18]);
  nor (_07312_, _07311_, _07281_);
  nand (_07313_, _07312_, _07310_);
  nand (_07314_, _07281_, word_in[26]);
  nand (_25005_[2], _07314_, _07313_);
  not (_07316_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nand (_07318_, _07265_, _07316_);
  not (_07319_, word_in[3]);
  nand (_07320_, _07264_, _07319_);
  nand (_07322_, _07320_, _07318_);
  nand (_07323_, _07322_, _07262_);
  not (_07324_, word_in[11]);
  nand (_07326_, _07261_, _07324_);
  nand (_07327_, _07326_, _07323_);
  nand (_07328_, _07327_, _07260_);
  nor (_07329_, _07260_, word_in[19]);
  nor (_07330_, _07329_, _07281_);
  nand (_07331_, _07330_, _07328_);
  nand (_07332_, _07281_, word_in[27]);
  nand (_25005_[3], _07332_, _07331_);
  not (_07333_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nand (_07334_, _07265_, _07333_);
  not (_07335_, word_in[4]);
  nand (_07336_, _07264_, _07335_);
  nand (_07337_, _07336_, _07334_);
  nand (_07338_, _07337_, _07262_);
  not (_07339_, word_in[12]);
  nand (_07340_, _07261_, _07339_);
  nand (_07341_, _07340_, _07338_);
  nand (_07342_, _07341_, _07260_);
  nor (_07343_, _07260_, word_in[20]);
  nor (_07344_, _07343_, _07281_);
  nand (_07345_, _07344_, _07342_);
  nand (_07346_, _07281_, word_in[28]);
  nand (_25005_[4], _07346_, _07345_);
  not (_07347_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nand (_07348_, _07265_, _07347_);
  not (_07349_, word_in[5]);
  nand (_07350_, _07264_, _07349_);
  nand (_07351_, _07350_, _07348_);
  nand (_07352_, _07351_, _07262_);
  not (_07353_, word_in[13]);
  nand (_07354_, _07261_, _07353_);
  nand (_07355_, _07354_, _07352_);
  nand (_07356_, _07355_, _07260_);
  nor (_07357_, _07260_, word_in[21]);
  nor (_07358_, _07357_, _07281_);
  nand (_07359_, _07358_, _07356_);
  nand (_07361_, _07281_, word_in[29]);
  nand (_25005_[5], _07361_, _07359_);
  not (_07362_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nand (_07363_, _07265_, _07362_);
  not (_07364_, word_in[6]);
  nand (_07365_, _07264_, _07364_);
  nand (_07366_, _07365_, _07363_);
  nand (_07367_, _07366_, _07262_);
  not (_07368_, word_in[14]);
  nand (_07369_, _07261_, _07368_);
  nand (_07370_, _07369_, _07367_);
  nand (_07372_, _07370_, _07260_);
  nor (_07373_, _07260_, word_in[22]);
  nor (_07374_, _07373_, _07281_);
  nand (_07375_, _07374_, _07372_);
  nand (_07376_, _07281_, word_in[30]);
  nand (_25005_[6], _07376_, _07375_);
  not (_07377_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_07378_, _07265_, _07377_);
  not (_07379_, word_in[7]);
  nand (_07380_, _07264_, _07379_);
  nand (_07381_, _07380_, _07378_);
  nand (_07382_, _07381_, _07262_);
  not (_07383_, word_in[15]);
  nand (_07384_, _07261_, _07383_);
  nand (_07385_, _07384_, _07382_);
  nand (_07386_, _07385_, _07260_);
  nor (_07387_, _07260_, word_in[23]);
  nor (_07388_, _07387_, _07281_);
  nand (_07389_, _07388_, _07386_);
  nand (_07390_, _07281_, word_in[31]);
  nand (_25005_[7], _07390_, _07389_);
  nor (_07392_, _22490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  nor (_07393_, _22492_, _21586_);
  nor (_25065_, _07393_, _07392_);
  nor (_07395_, _06568_, _06191_);
  nand (_07396_, _07395_, _07277_);
  not (_07397_, _07396_);
  nor (_07398_, _07258_, _06192_);
  not (_07399_, _07398_);
  nor (_07400_, _07399_, _06359_);
  nor (_07401_, _06579_, _06075_);
  not (_07402_, _07401_);
  nor (_07403_, _07402_, _06203_);
  nor (_07404_, _06591_, _06721_);
  nor (_07405_, _07404_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  not (_07406_, _07404_);
  nor (_07407_, _07406_, word_in[0]);
  nor (_07408_, _07407_, _07405_);
  nor (_07409_, _07408_, _07403_);
  not (_07410_, _07403_);
  nor (_07411_, _07410_, word_in[8]);
  nor (_07413_, _07411_, _07409_);
  nor (_07414_, _07413_, _07400_);
  not (_07416_, _07400_);
  nor (_07417_, _07416_, word_in[16]);
  nor (_07418_, _07417_, _07414_);
  nor (_07419_, _07418_, _07397_);
  nor (_07421_, _07396_, word_in[24]);
  nor (_24989_, _07421_, _07419_);
  nor (_07422_, _07416_, word_in[17]);
  nor (_07424_, _07404_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_07425_, _07406_, word_in[1]);
  nor (_07426_, _07425_, _07424_);
  nor (_07427_, _07426_, _07403_);
  nor (_07428_, _07410_, word_in[9]);
  nor (_07429_, _07428_, _07427_);
  nor (_07430_, _07429_, _07400_);
  nor (_07431_, _07430_, _07422_);
  nor (_07432_, _07431_, _07397_);
  nor (_07433_, _07396_, word_in[25]);
  nor (_24990_, _07433_, _07432_);
  not (_07435_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand (_07436_, _07406_, _07435_);
  nand (_07437_, _07404_, _07303_);
  nand (_07438_, _07437_, _07436_);
  nand (_07439_, _07438_, _07410_);
  nand (_07440_, _07403_, _07307_);
  nand (_07441_, _07440_, _07439_);
  nand (_07442_, _07441_, _07416_);
  nor (_07443_, _07416_, word_in[18]);
  nor (_07445_, _07443_, _07397_);
  nand (_07446_, _07445_, _07442_);
  nand (_07447_, _07397_, word_in[26]);
  nand (_24991_, _07447_, _07446_);
  not (_07448_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nand (_07449_, _07406_, _07448_);
  nand (_07450_, _07404_, _07319_);
  nand (_07451_, _07450_, _07449_);
  nand (_07452_, _07451_, _07410_);
  nand (_07454_, _07403_, _07324_);
  nand (_07455_, _07454_, _07452_);
  nand (_07457_, _07455_, _07416_);
  nor (_07458_, _07416_, word_in[19]);
  nor (_07459_, _07458_, _07397_);
  nand (_07461_, _07459_, _07457_);
  nand (_07462_, _07397_, word_in[27]);
  nand (_24992_, _07462_, _07461_);
  not (_07463_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nand (_07464_, _07406_, _07463_);
  nand (_07465_, _07404_, _07335_);
  nand (_07467_, _07465_, _07464_);
  nand (_07468_, _07467_, _07410_);
  nand (_07469_, _07403_, _07339_);
  nand (_07470_, _07469_, _07468_);
  nand (_07471_, _07470_, _07416_);
  nor (_07472_, _07416_, word_in[20]);
  nor (_07473_, _07472_, _07397_);
  nand (_07474_, _07473_, _07471_);
  nand (_07475_, _07397_, word_in[28]);
  nand (_24993_, _07475_, _07474_);
  not (_07476_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nand (_07477_, _07406_, _07476_);
  nand (_07478_, _07404_, _07349_);
  nand (_07479_, _07478_, _07477_);
  nand (_07480_, _07479_, _07410_);
  nand (_07481_, _07403_, _07353_);
  nand (_07482_, _07481_, _07480_);
  nand (_07483_, _07482_, _07416_);
  nor (_07484_, _07416_, word_in[21]);
  nor (_07485_, _07484_, _07397_);
  nand (_07488_, _07485_, _07483_);
  nand (_07489_, _07397_, word_in[29]);
  nand (_24994_, _07489_, _07488_);
  nor (_07490_, _21653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  nor (_07491_, _21655_, _21526_);
  nor (_00012_, _07491_, _07490_);
  nor (_07492_, _07416_, word_in[22]);
  nor (_07493_, _07404_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_07494_, _07406_, word_in[6]);
  nor (_07495_, _07494_, _07493_);
  nor (_07496_, _07495_, _07403_);
  nor (_07497_, _07410_, word_in[14]);
  nor (_07498_, _07497_, _07496_);
  nor (_07499_, _07498_, _07400_);
  nor (_07500_, _07499_, _07492_);
  nor (_07501_, _07500_, _07397_);
  nor (_07502_, _07396_, word_in[30]);
  nor (_24995_, _07502_, _07501_);
  not (_07503_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_07505_, _07404_, _07503_);
  nor (_07507_, _06187_, rst);
  not (_07508_, _07507_);
  nor (_07509_, _07508_, _06721_);
  nor (_07510_, _07509_, _07505_);
  nor (_07511_, _07510_, _07403_);
  nor (_07512_, _07410_, _07383_);
  nor (_07513_, _07512_, _07511_);
  nor (_07514_, _07513_, _07400_);
  nand (_07515_, _07400_, _06606_);
  nand (_07516_, _07515_, _07396_);
  nor (_07518_, _07516_, _07514_);
  nor (_07519_, _07396_, word_in[31]);
  nor (_24996_, _07519_, _07518_);
  nor (_07520_, _01083_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  nor (_07522_, _01052_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  nand (_07523_, _07522_, _01080_);
  nand (_07524_, _07523_, _23493_);
  nor (_00044_, _07524_, _07520_);
  nor (_07525_, _21842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  nor (_07526_, _21844_, _21586_);
  nor (_00061_, _07526_, _07525_);
  nor (_07527_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  nor (_07528_, _06973_, _21554_);
  nor (_00065_, _07528_, _07527_);
  nor (_07529_, _21873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  nor (_07530_, _21875_, _21504_);
  nor (_00082_, _07530_, _07529_);
  nor (_07531_, _07258_, _06075_);
  not (_07532_, _07531_);
  nor (_07533_, _07532_, _06359_);
  not (_07535_, _07533_);
  nor (_07536_, _06579_, _06241_);
  not (_07537_, _07536_);
  nor (_07539_, _07537_, _06203_);
  not (_07540_, _07539_);
  not (_07541_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nand (_07542_, _06590_, _06688_);
  nand (_07543_, _07542_, _07541_);
  not (_07544_, _07542_);
  nand (_07545_, _07544_, _07267_);
  nand (_07546_, _07545_, _07543_);
  nand (_07547_, _07546_, _07540_);
  nand (_07548_, _07539_, _07272_);
  nand (_07549_, _07548_, _07547_);
  nand (_07551_, _07549_, _07535_);
  nor (_07552_, _06568_, _06192_);
  nand (_07553_, _07552_, _07277_);
  not (_07554_, _07553_);
  nor (_07555_, _07535_, word_in[16]);
  nor (_07556_, _07555_, _07554_);
  nand (_07558_, _07556_, _07551_);
  nand (_07559_, _07554_, word_in[24]);
  nand (_24997_, _07559_, _07558_);
  nand (_07561_, _07554_, word_in[25]);
  not (_07562_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nand (_07563_, _07542_, _07562_);
  not (_07564_, word_in[1]);
  nand (_07565_, _07544_, _07564_);
  nand (_07566_, _07565_, _07563_);
  nand (_07567_, _07566_, _07540_);
  not (_07568_, word_in[9]);
  nand (_07569_, _07539_, _07568_);
  nand (_07570_, _07569_, _07567_);
  nand (_07571_, _07570_, _07535_);
  nor (_07572_, _07535_, word_in[17]);
  nor (_07573_, _07572_, _07554_);
  nand (_07575_, _07573_, _07571_);
  nand (_24998_, _07575_, _07561_);
  nor (_07576_, _07542_, _07303_);
  not (_07577_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_07578_, _07544_, _07577_);
  nor (_07580_, _07578_, _07576_);
  nor (_07581_, _07580_, _07539_);
  nor (_07582_, _07540_, _07307_);
  nor (_07583_, _07582_, _07581_);
  nor (_07584_, _07583_, _07533_);
  nand (_07585_, _07533_, word_in[18]);
  nand (_07586_, _07585_, _07553_);
  nor (_07587_, _07586_, _07584_);
  nor (_07588_, _07553_, word_in[26]);
  nor (_24999_, _07588_, _07587_);
  nor (_07589_, _21741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  nor (_07590_, _21744_, _21554_);
  nor (_00102_, _07590_, _07589_);
  not (_07591_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nand (_07592_, _07542_, _07591_);
  nand (_07593_, _07544_, _07319_);
  nand (_07594_, _07593_, _07592_);
  nand (_07595_, _07594_, _07540_);
  nand (_07596_, _07539_, _07324_);
  nand (_07597_, _07596_, _07595_);
  nand (_07599_, _07597_, _07535_);
  nor (_07600_, _07535_, word_in[19]);
  nor (_07601_, _07600_, _07554_);
  nand (_07602_, _07601_, _07599_);
  nand (_07603_, _07554_, word_in[27]);
  nand (_25000_, _07603_, _07602_);
  not (_07604_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nand (_07605_, _07542_, _07604_);
  nand (_07606_, _07544_, _07335_);
  nand (_07607_, _07606_, _07605_);
  nand (_07608_, _07607_, _07540_);
  nand (_07609_, _07539_, _07339_);
  nand (_07610_, _07609_, _07608_);
  nand (_07611_, _07610_, _07535_);
  nor (_07612_, _07535_, word_in[20]);
  nor (_07613_, _07612_, _07554_);
  nand (_07614_, _07613_, _07611_);
  nand (_07615_, _07554_, word_in[28]);
  nand (_25001_, _07615_, _07614_);
  nand (_07616_, _07554_, word_in[29]);
  not (_07617_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nand (_07618_, _07542_, _07617_);
  nand (_07619_, _07544_, _07349_);
  nand (_07620_, _07619_, _07618_);
  nand (_07621_, _07620_, _07540_);
  nand (_07622_, _07539_, _07353_);
  nand (_07623_, _07622_, _07621_);
  nand (_07624_, _07623_, _07535_);
  nor (_07626_, _07535_, word_in[21]);
  nor (_07627_, _07626_, _07554_);
  nand (_07628_, _07627_, _07624_);
  nand (_25002_, _07628_, _07616_);
  not (_07629_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nand (_07630_, _07542_, _07629_);
  nand (_07631_, _07544_, _07364_);
  nand (_07632_, _07631_, _07630_);
  nand (_07633_, _07632_, _07540_);
  nand (_07634_, _07539_, _07368_);
  nand (_07635_, _07634_, _07633_);
  nand (_07636_, _07635_, _07535_);
  nor (_07637_, _07535_, word_in[22]);
  nor (_07638_, _07637_, _07554_);
  nand (_07639_, _07638_, _07636_);
  nand (_07640_, _07554_, word_in[30]);
  nand (_25003_, _07640_, _07639_);
  not (_07641_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nor (_07643_, _07544_, _07641_);
  nor (_07644_, _07542_, _07508_);
  nor (_07645_, _07644_, _07643_);
  nor (_07646_, _07645_, _07539_);
  nor (_07647_, _07540_, _07383_);
  nor (_07648_, _07647_, _07646_);
  nor (_07649_, _07648_, _07533_);
  nand (_07650_, _07533_, _06606_);
  nand (_07651_, _07650_, _07553_);
  nor (_07653_, _07651_, _07649_);
  nor (_07654_, _07553_, word_in[31]);
  nor (_25004_, _07654_, _07653_);
  nor (_07655_, _21842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1]);
  nor (_07656_, _21844_, _21474_);
  nor (_00166_, _07656_, _07655_);
  nor (_07657_, _06568_, _06738_);
  not (_07658_, _07657_);
  nor (_07659_, _07258_, _06241_);
  not (_07660_, _07659_);
  nor (_07661_, _07660_, _06359_);
  not (_07662_, _07661_);
  nor (_07663_, _07662_, word_in[16]);
  nor (_07665_, _06579_, _06191_);
  not (_07666_, _07665_);
  nor (_07667_, _07666_, _06203_);
  nand (_07668_, _06115_, word_in[0]);
  nor (_07669_, _07668_, rst);
  nand (_07670_, _07669_, _06723_);
  nor (_07671_, _06591_, _06725_);
  not (_07672_, _07671_);
  nand (_07673_, _07672_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nand (_07674_, _07673_, _07670_);
  nor (_07675_, _07674_, _07667_);
  not (_07676_, _07667_);
  nor (_07677_, _07676_, word_in[8]);
  nor (_07678_, _07677_, _07675_);
  nor (_07679_, _07678_, _07661_);
  nor (_07680_, _07679_, _07663_);
  nand (_07681_, _07680_, _07658_);
  nand (_07682_, _07657_, word_in[24]);
  nand (_25009_[0], _07682_, _07681_);
  nand (_07683_, _07672_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nand (_07684_, _06115_, word_in[1]);
  nor (_07685_, _07684_, rst);
  nand (_07686_, _07685_, _06723_);
  nand (_07687_, _07686_, _07683_);
  nor (_07688_, _07687_, _07667_);
  nor (_07689_, _07676_, word_in[9]);
  nor (_07690_, _07689_, _07688_);
  nor (_07691_, _07690_, _07661_);
  nor (_07692_, _07662_, word_in[17]);
  nor (_07693_, _07692_, _07691_);
  nand (_07694_, _07693_, _07658_);
  nand (_07696_, _07657_, word_in[25]);
  nand (_25009_[1], _07696_, _07694_);
  not (_07697_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_07698_, _07671_, _07697_);
  nand (_07699_, _06590_, word_in[2]);
  nor (_07700_, _07699_, _06725_);
  nor (_07701_, _07700_, _07698_);
  nand (_07703_, _07701_, _07676_);
  nand (_07704_, _07667_, _07307_);
  nand (_07705_, _07704_, _07703_);
  nand (_07706_, _07705_, _07662_);
  nor (_07707_, _07662_, word_in[18]);
  nor (_07708_, _07707_, _07657_);
  nand (_07709_, _07708_, _07706_);
  nand (_07710_, _07657_, word_in[26]);
  nand (_25009_[2], _07710_, _07709_);
  not (_07711_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_07713_, _07671_, _07711_);
  nand (_07715_, _06590_, word_in[3]);
  nor (_07716_, _07715_, _06725_);
  nor (_07718_, _07716_, _07713_);
  nand (_07719_, _07718_, _07676_);
  nand (_07720_, _07667_, _07324_);
  nand (_07721_, _07720_, _07719_);
  nand (_07722_, _07721_, _07662_);
  nor (_07723_, _07662_, word_in[19]);
  nor (_07724_, _07723_, _07657_);
  nand (_07725_, _07724_, _07722_);
  nand (_07726_, _07657_, word_in[27]);
  nand (_25009_[3], _07726_, _07725_);
  not (_07727_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_07728_, _07671_, _07727_);
  nand (_07729_, _06590_, word_in[4]);
  nor (_07731_, _07729_, _06725_);
  nor (_07733_, _07731_, _07728_);
  nand (_07734_, _07733_, _07676_);
  nand (_07735_, _07667_, _07339_);
  nand (_07736_, _07735_, _07734_);
  nand (_07737_, _07736_, _07662_);
  nor (_07738_, _07662_, word_in[20]);
  nor (_07740_, _07738_, _07657_);
  nand (_07741_, _07740_, _07737_);
  nand (_07742_, _07657_, word_in[28]);
  nand (_25009_[4], _07742_, _07741_);
  nand (_07744_, _07672_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nand (_07745_, _06115_, word_in[5]);
  nor (_07746_, _07745_, rst);
  nand (_07747_, _07746_, _06723_);
  nand (_07748_, _07747_, _07744_);
  nand (_07749_, _07748_, _07676_);
  nand (_07750_, _07667_, word_in[13]);
  nand (_07751_, _07750_, _07749_);
  nand (_07752_, _07751_, _07662_);
  nand (_07753_, _07661_, word_in[21]);
  nand (_07754_, _07753_, _07752_);
  nand (_07755_, _07754_, _07658_);
  nand (_07756_, _07657_, word_in[29]);
  nand (_25009_[5], _07756_, _07755_);
  nand (_07758_, _07672_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nand (_07759_, _06115_, word_in[6]);
  nor (_07761_, _07759_, rst);
  nand (_07762_, _07761_, _06723_);
  nand (_07763_, _07762_, _07758_);
  nand (_07764_, _07763_, _07676_);
  nand (_07765_, _07667_, word_in[14]);
  nand (_07766_, _07765_, _07764_);
  nand (_07767_, _07766_, _07662_);
  nand (_07768_, _07661_, word_in[22]);
  nand (_07769_, _07768_, _07767_);
  nand (_07770_, _07769_, _07658_);
  nand (_07771_, _07657_, word_in[30]);
  nand (_25009_[6], _07771_, _07770_);
  nand (_07772_, _06610_, _06613_);
  not (_07773_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nor (_07774_, _07671_, _07773_);
  nor (_07775_, _07508_, _06725_);
  nor (_07776_, _07775_, _07774_);
  nor (_07777_, _07776_, _07667_);
  nor (_07778_, _07676_, _07383_);
  nor (_07779_, _07778_, _07777_);
  nand (_07782_, _07779_, _07662_);
  nor (_07784_, _07662_, _06606_);
  nor (_07785_, _07784_, _07657_);
  nand (_07786_, _07785_, _07782_);
  nand (_25009_[7], _07786_, _07772_);
  nor (_07787_, _21690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  nor (_07788_, _21692_, _21414_);
  nor (_00215_, _07788_, _07787_);
  nand (_07789_, _07276_, _06451_);
  nor (_07791_, _07789_, _06241_);
  not (_07792_, _07791_);
  nand (_07793_, _06411_, word_in[16]);
  nor (_07794_, _07793_, rst);
  nor (_07795_, _06913_, _07258_);
  not (_07796_, _07795_);
  nor (_07797_, _07796_, _06191_);
  nand (_07798_, _07797_, _07794_);
  not (_07799_, _07797_);
  nor (_07800_, _06579_, _06725_);
  not (_07801_, _07800_);
  nor (_07802_, _06591_, _06753_);
  nand (_07803_, _07802_, word_in[0]);
  not (_07804_, _07802_);
  nand (_07805_, _07804_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nand (_07806_, _07805_, _07803_);
  nand (_07807_, _07806_, _07801_);
  nand (_07808_, _07800_, word_in[8]);
  nand (_07809_, _07808_, _07807_);
  nand (_07810_, _07809_, _07799_);
  nand (_07811_, _07810_, _07798_);
  nand (_07812_, _07811_, _07792_);
  nand (_07813_, _06513_, word_in[24]);
  nor (_07814_, _07813_, rst);
  nand (_07815_, _07791_, _07814_);
  nand (_25010_[0], _07815_, _07812_);
  nand (_07816_, _06411_, word_in[17]);
  nor (_07817_, _07816_, rst);
  nand (_07819_, _07797_, _07817_);
  nand (_07820_, _07802_, word_in[1]);
  nand (_07821_, _07804_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nand (_07824_, _07821_, _07820_);
  nand (_07825_, _07824_, _07801_);
  nand (_07826_, _07800_, word_in[9]);
  nand (_07827_, _07826_, _07825_);
  nand (_07829_, _07827_, _07799_);
  nand (_07830_, _07829_, _07819_);
  nand (_07831_, _07830_, _07792_);
  nand (_07832_, _06513_, word_in[25]);
  nor (_07833_, _07832_, rst);
  nand (_07834_, _07791_, _07833_);
  nand (_25010_[1], _07834_, _07831_);
  nand (_07836_, _07802_, word_in[2]);
  nand (_07838_, _07804_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand (_07839_, _07838_, _07836_);
  nand (_07841_, _07839_, _07801_);
  nand (_07842_, _07800_, word_in[10]);
  nand (_07843_, _07842_, _07841_);
  nand (_07845_, _07843_, _07799_);
  nand (_07846_, _06411_, word_in[18]);
  nor (_07847_, _07846_, rst);
  nand (_07850_, _07797_, _07847_);
  nand (_07852_, _07850_, _07845_);
  nand (_07854_, _07852_, _07792_);
  nand (_07855_, _06513_, word_in[26]);
  nor (_07856_, _07855_, rst);
  nand (_07857_, _07791_, _07856_);
  nand (_25010_[2], _07857_, _07854_);
  nor (_07858_, _07804_, _07319_);
  not (_07859_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_07860_, _07802_, _07859_);
  nor (_07861_, _07860_, _07858_);
  nor (_07862_, _07861_, _07800_);
  nor (_07864_, _07801_, _07324_);
  nor (_07866_, _07864_, _07862_);
  nor (_07867_, _07866_, _07797_);
  nand (_07868_, _06411_, word_in[19]);
  nor (_07869_, _07868_, rst);
  nand (_07870_, _07797_, _07869_);
  nand (_07871_, _07870_, _07792_);
  nor (_07872_, _07871_, _07867_);
  nand (_07873_, _06513_, word_in[27]);
  nor (_07874_, _07873_, rst);
  nor (_07875_, _07792_, _07874_);
  nor (_25010_[3], _07875_, _07872_);
  nor (_07877_, _07804_, _07335_);
  not (_07878_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_07879_, _07802_, _07878_);
  nor (_07880_, _07879_, _07877_);
  nor (_07881_, _07880_, _07800_);
  nor (_07882_, _07801_, _07339_);
  nor (_07883_, _07882_, _07881_);
  nor (_07884_, _07883_, _07797_);
  nand (_07885_, _06411_, word_in[20]);
  nor (_07887_, _07885_, rst);
  nand (_07888_, _07797_, _07887_);
  nand (_07889_, _07888_, _07792_);
  nor (_07890_, _07889_, _07884_);
  nand (_07891_, _06513_, word_in[28]);
  nor (_07892_, _07891_, rst);
  nor (_07893_, _07792_, _07892_);
  nor (_25010_[4], _07893_, _07890_);
  nand (_07894_, _06411_, word_in[21]);
  nor (_07896_, _07894_, rst);
  nand (_07897_, _07797_, _07896_);
  nand (_07898_, _07802_, word_in[5]);
  nand (_07899_, _07804_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nand (_07900_, _07899_, _07898_);
  nand (_07901_, _07900_, _07801_);
  nand (_07902_, _07800_, word_in[13]);
  nand (_07903_, _07902_, _07901_);
  nand (_07904_, _07903_, _07799_);
  nand (_07905_, _07904_, _07897_);
  nand (_07906_, _07905_, _07792_);
  nand (_07907_, _06513_, word_in[29]);
  nor (_07908_, _07907_, rst);
  nand (_07909_, _07791_, _07908_);
  nand (_25010_[5], _07909_, _07906_);
  nand (_07910_, _06411_, word_in[22]);
  nor (_07911_, _07910_, rst);
  nand (_07912_, _07797_, _07911_);
  nand (_07914_, _07802_, word_in[6]);
  nand (_07915_, _07804_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nand (_07917_, _07915_, _07914_);
  nand (_07918_, _07917_, _07801_);
  nand (_07919_, _07800_, word_in[14]);
  nand (_07920_, _07919_, _07918_);
  nand (_07921_, _07920_, _07799_);
  nand (_07923_, _07921_, _07912_);
  nand (_07924_, _07923_, _07792_);
  nand (_07925_, _06513_, word_in[30]);
  nor (_07926_, _07925_, rst);
  nand (_07927_, _07791_, _07926_);
  nand (_25010_[6], _07927_, _07924_);
  nor (_07928_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1]);
  nor (_07929_, _06973_, _21474_);
  nor (_00289_, _07929_, _07928_);
  nand (_07931_, _07797_, _06606_);
  nand (_07932_, _07804_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_07934_, _07507_, _06752_);
  nand (_07935_, _07934_, _07932_);
  nand (_07936_, _07935_, _07801_);
  nand (_07937_, _07800_, word_in[15]);
  nand (_07938_, _07937_, _07936_);
  nand (_07939_, _07938_, _07799_);
  nand (_07940_, _07939_, _07931_);
  nand (_07941_, _07940_, _07792_);
  nand (_07942_, _07791_, _06610_);
  nand (_25010_[7], _07942_, _07941_);
  nor (_07943_, _07789_, _06191_);
  not (_07944_, _07943_);
  nor (_07945_, _07796_, _06192_);
  nand (_07946_, _07945_, _07794_);
  nor (_07947_, _07402_, _06981_);
  nand (_07949_, _07947_, _07272_);
  nor (_07950_, _06591_, _06819_);
  nand (_07951_, _07950_, word_in[0]);
  not (_07952_, _07950_);
  nand (_07953_, _07952_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand (_07954_, _07953_, _07951_);
  nor (_07955_, _07954_, _07947_);
  nor (_07957_, _07955_, _07945_);
  nand (_07958_, _07957_, _07949_);
  nand (_07960_, _07958_, _07946_);
  nand (_07962_, _07960_, _07944_);
  nand (_07963_, _07943_, _07814_);
  nand (_25011_[0], _07963_, _07962_);
  nor (_07964_, _07952_, _07564_);
  not (_07965_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_07966_, _07950_, _07965_);
  nor (_07968_, _07966_, _07964_);
  nor (_07969_, _07968_, _07947_);
  not (_07970_, _07947_);
  nor (_07971_, _07970_, _07568_);
  nor (_07972_, _07971_, _07969_);
  nor (_07973_, _07972_, _07945_);
  nand (_07974_, _07945_, _07817_);
  nand (_07975_, _07974_, _07944_);
  nor (_07976_, _07975_, _07973_);
  nor (_07977_, _07944_, _07833_);
  nor (_25011_[1], _07977_, _07976_);
  nand (_07978_, _07947_, _07307_);
  nand (_07979_, _07950_, word_in[2]);
  nand (_07980_, _07952_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand (_07981_, _07980_, _07979_);
  nor (_07982_, _07981_, _07947_);
  nor (_07983_, _07982_, _07945_);
  nand (_07984_, _07983_, _07978_);
  nand (_07985_, _07945_, _07847_);
  nand (_07987_, _07985_, _07984_);
  nand (_07988_, _07987_, _07944_);
  nand (_07990_, _07943_, _07856_);
  nand (_25011_[2], _07990_, _07988_);
  nor (_07991_, _07950_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_07992_, _07952_, word_in[3]);
  nor (_07993_, _07992_, _07991_);
  nor (_07994_, _07993_, _07947_);
  nor (_07995_, _07970_, word_in[11]);
  nor (_07996_, _07995_, _07994_);
  nor (_07997_, _07996_, _07945_);
  not (_07998_, _07945_);
  nor (_08000_, _07998_, _07869_);
  nor (_08001_, _08000_, _07997_);
  nor (_08002_, _08001_, _07943_);
  nor (_08003_, _07944_, _07874_);
  nor (_25011_[3], _08003_, _08002_);
  nor (_08004_, _07952_, _07335_);
  not (_08005_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_08006_, _07950_, _08005_);
  nor (_08008_, _08006_, _08004_);
  nor (_08009_, _08008_, _07947_);
  nor (_08011_, _07970_, _07339_);
  nor (_08012_, _08011_, _08009_);
  nor (_08013_, _08012_, _07945_);
  nand (_08014_, _07945_, _07887_);
  nand (_08016_, _08014_, _07944_);
  nor (_08017_, _08016_, _08013_);
  nor (_08018_, _07944_, _07892_);
  nor (_25011_[4], _08018_, _08017_);
  nor (_08019_, _07952_, _07349_);
  not (_08020_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_08022_, _07950_, _08020_);
  nor (_08023_, _08022_, _08019_);
  nor (_08024_, _08023_, _07947_);
  nor (_08025_, _07970_, _07353_);
  nor (_08026_, _08025_, _08024_);
  nor (_08027_, _08026_, _07945_);
  nand (_08028_, _07945_, _07896_);
  nand (_08029_, _08028_, _07944_);
  nor (_08031_, _08029_, _08027_);
  nor (_08033_, _07944_, _07908_);
  nor (_25011_[5], _08033_, _08031_);
  nand (_08035_, _07945_, _07911_);
  nand (_08037_, _07947_, _07368_);
  nand (_08038_, _07950_, word_in[6]);
  nand (_08039_, _07952_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nand (_08040_, _08039_, _08038_);
  nor (_08041_, _08040_, _07947_);
  nor (_08042_, _08041_, _07945_);
  nand (_08044_, _08042_, _08037_);
  nand (_08045_, _08044_, _08035_);
  nand (_08046_, _08045_, _07944_);
  nand (_08047_, _07943_, _07926_);
  nand (_25011_[6], _08047_, _08046_);
  nand (_08048_, _07945_, _06606_);
  nand (_08049_, _07947_, _07383_);
  nand (_08051_, _07507_, _06781_);
  nand (_08053_, _07952_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_08054_, _08053_, _08051_);
  nor (_08055_, _08054_, _07947_);
  nor (_08056_, _08055_, _07945_);
  nand (_08058_, _08056_, _08049_);
  nand (_08059_, _08058_, _08048_);
  nand (_08060_, _08059_, _07944_);
  nand (_08061_, _07943_, _06610_);
  nand (_25011_[7], _08061_, _08060_);
  nor (_08062_, _21752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5]);
  nor (_08063_, _21754_, _21451_);
  nor (_00396_, _08063_, _08062_);
  nor (_08064_, _07789_, _06192_);
  not (_08065_, _08064_);
  nor (_08066_, _07537_, _06981_);
  nand (_08067_, _08066_, _07272_);
  nor (_08069_, _07796_, _06075_);
  nor (_08070_, _06591_, _06822_);
  nand (_08071_, _08070_, word_in[0]);
  not (_08072_, _08070_);
  nand (_08073_, _08072_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nand (_08074_, _08073_, _08071_);
  nor (_08075_, _08074_, _08066_);
  nor (_08076_, _08075_, _08069_);
  nand (_08077_, _08076_, _08067_);
  nand (_08078_, _08069_, _07794_);
  nand (_08079_, _08078_, _08077_);
  nand (_08080_, _08079_, _08065_);
  nand (_08081_, _08064_, _07814_);
  nand (_25012_[0], _08081_, _08080_);
  nor (_08082_, _22531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  nor (_08083_, _22533_, _21414_);
  nor (_00419_, _08083_, _08082_);
  nor (_08084_, _08070_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_08085_, _08072_, word_in[1]);
  nor (_08087_, _08085_, _08084_);
  nor (_08088_, _08087_, _08066_);
  not (_08090_, _08066_);
  nor (_08091_, _08090_, word_in[9]);
  nor (_08092_, _08091_, _08088_);
  nor (_08093_, _08092_, _08069_);
  not (_08094_, _08069_);
  nor (_08095_, _08094_, _07817_);
  nor (_08096_, _08095_, _08093_);
  nor (_08097_, _08096_, _08064_);
  nor (_08098_, _08065_, _07833_);
  nor (_25012_[1], _08098_, _08097_);
  nor (_08099_, _08072_, _07303_);
  not (_08101_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_08102_, _08070_, _08101_);
  nor (_08103_, _08102_, _08099_);
  nor (_08104_, _08103_, _08066_);
  nor (_08105_, _08090_, _07307_);
  nor (_08106_, _08105_, _08104_);
  nor (_08107_, _08106_, _08069_);
  nand (_08108_, _08069_, _07847_);
  nand (_08109_, _08108_, _08065_);
  nor (_08110_, _08109_, _08107_);
  nor (_08111_, _08065_, _07856_);
  nor (_25012_[2], _08111_, _08110_);
  nor (_08112_, _08070_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_08113_, _08072_, word_in[3]);
  nor (_08114_, _08113_, _08112_);
  nor (_08115_, _08114_, _08066_);
  nor (_08116_, _08090_, word_in[11]);
  nor (_08117_, _08116_, _08115_);
  nor (_08118_, _08117_, _08069_);
  nor (_08119_, _08094_, _07869_);
  nor (_08120_, _08119_, _08118_);
  nor (_08121_, _08120_, _08064_);
  nor (_08122_, _08065_, _07874_);
  nor (_25012_[3], _08122_, _08121_);
  nor (_08123_, _08070_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_08124_, _08072_, word_in[4]);
  nor (_08125_, _08124_, _08123_);
  nor (_08126_, _08125_, _08066_);
  nor (_08127_, _08090_, word_in[12]);
  nor (_08128_, _08127_, _08126_);
  nor (_08129_, _08128_, _08069_);
  nor (_08130_, _08094_, _07887_);
  nor (_08131_, _08130_, _08129_);
  nor (_08132_, _08131_, _08064_);
  nor (_08133_, _08065_, _07892_);
  nor (_25012_[4], _08133_, _08132_);
  nor (_08134_, _08070_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_08135_, _08072_, word_in[5]);
  nor (_08136_, _08135_, _08134_);
  nor (_08137_, _08136_, _08066_);
  nor (_08138_, _08090_, word_in[13]);
  nor (_08139_, _08138_, _08137_);
  nor (_08140_, _08139_, _08069_);
  nor (_08141_, _08094_, _07896_);
  nor (_08142_, _08141_, _08140_);
  nor (_08143_, _08142_, _08064_);
  nor (_08145_, _08065_, _07908_);
  nor (_25012_[5], _08145_, _08143_);
  nor (_08148_, _08072_, _07364_);
  not (_08149_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_08150_, _08070_, _08149_);
  nor (_08152_, _08150_, _08148_);
  nor (_08153_, _08152_, _08066_);
  nor (_08154_, _08090_, _07368_);
  nor (_08156_, _08154_, _08153_);
  nor (_08157_, _08156_, _08069_);
  nand (_08158_, _08069_, _07911_);
  nand (_08159_, _08158_, _08065_);
  nor (_08160_, _08159_, _08157_);
  nor (_08161_, _08065_, _07926_);
  nor (_25012_[6], _08161_, _08160_);
  nand (_08162_, _08066_, _07383_);
  nand (_08164_, _08070_, word_in[7]);
  nand (_08165_, _08072_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_08166_, _08165_, _08164_);
  nor (_08167_, _08166_, _08066_);
  nor (_08169_, _08167_, _08069_);
  nand (_08170_, _08169_, _08162_);
  nand (_08171_, _08069_, _06606_);
  nand (_08172_, _08171_, _08170_);
  nand (_08173_, _08172_, _08065_);
  nand (_08174_, _08064_, _06610_);
  nand (_25012_[7], _08174_, _08173_);
  nor (_08176_, _21690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  nor (_08177_, _21692_, _21504_);
  nor (_25267_, _08177_, _08176_);
  nor (_08178_, _07796_, _06241_);
  not (_08179_, _08178_);
  nor (_08180_, _07666_, _06981_);
  not (_08181_, _08180_);
  not (_08182_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor (_08183_, _06591_, _06915_);
  not (_08184_, _08183_);
  nand (_08185_, _08184_, _08182_);
  nand (_08186_, _08183_, _07267_);
  nand (_08187_, _08186_, _08185_);
  nand (_08189_, _08187_, _08181_);
  nand (_08190_, _08180_, _07272_);
  nand (_08191_, _08190_, _08189_);
  nand (_08192_, _08191_, _08179_);
  nor (_08193_, _06568_, _06753_);
  nor (_08195_, _08179_, _07794_);
  nor (_08196_, _08195_, _08193_);
  nand (_08198_, _08196_, _08192_);
  nand (_08199_, _08193_, _07814_);
  nand (_25013_[0], _08199_, _08198_);
  nand (_08200_, _07833_, _06752_);
  not (_08201_, _08193_);
  nand (_08202_, _08180_, _07568_);
  nand (_08204_, _08183_, word_in[1]);
  nand (_08205_, _08184_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nand (_08207_, _08205_, _08204_);
  nor (_08208_, _08207_, _08180_);
  nor (_08209_, _08208_, _08178_);
  nand (_08210_, _08209_, _08202_);
  nand (_08211_, _08178_, _07817_);
  nand (_08213_, _08211_, _08210_);
  nand (_08214_, _08213_, _08201_);
  nand (_25013_[1], _08214_, _08200_);
  nand (_08216_, _08178_, _07847_);
  nand (_08218_, _08180_, _07307_);
  nand (_08219_, _08183_, word_in[2]);
  nand (_08221_, _08184_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nand (_08222_, _08221_, _08219_);
  nor (_08223_, _08222_, _08180_);
  nor (_08224_, _08223_, _08178_);
  nand (_08225_, _08224_, _08218_);
  nand (_08226_, _08225_, _08216_);
  nand (_08227_, _08226_, _08201_);
  nand (_08228_, _08193_, word_in[26]);
  nand (_25013_[2], _08228_, _08227_);
  nand (_08229_, _08178_, _07869_);
  nand (_08230_, _08180_, _07324_);
  nand (_08231_, _08183_, word_in[3]);
  nand (_08232_, _08184_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nand (_08234_, _08232_, _08231_);
  nor (_08235_, _08234_, _08180_);
  nor (_08237_, _08235_, _08178_);
  nand (_08238_, _08237_, _08230_);
  nand (_08239_, _08238_, _08229_);
  nand (_08240_, _08239_, _08201_);
  nand (_08241_, _08193_, word_in[27]);
  nand (_25013_[3], _08241_, _08240_);
  nand (_08243_, _08180_, _07339_);
  nand (_08245_, _08183_, word_in[4]);
  nand (_08246_, _08184_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nand (_08248_, _08246_, _08245_);
  nor (_08249_, _08248_, _08180_);
  nor (_08250_, _08249_, _08178_);
  nand (_08251_, _08250_, _08243_);
  nand (_08252_, _08178_, _07887_);
  nand (_08253_, _08252_, _08251_);
  nand (_08254_, _08253_, _08201_);
  nand (_08255_, _07892_, _06752_);
  nand (_25013_[4], _08255_, _08254_);
  nand (_08256_, _08178_, _07896_);
  nand (_08257_, _08180_, _07353_);
  nand (_08258_, _08183_, word_in[5]);
  nand (_08259_, _08184_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nand (_08260_, _08259_, _08258_);
  nor (_08261_, _08260_, _08180_);
  nor (_08262_, _08261_, _08178_);
  nand (_08263_, _08262_, _08257_);
  nand (_08264_, _08263_, _08256_);
  nand (_08265_, _08264_, _08201_);
  nand (_08267_, _08193_, word_in[29]);
  nand (_25013_[5], _08267_, _08265_);
  nand (_08269_, _08183_, word_in[6]);
  nand (_08270_, _08184_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nand (_08271_, _08270_, _08269_);
  nand (_08273_, _08271_, _08181_);
  nand (_08275_, _08180_, word_in[14]);
  nand (_08277_, _08275_, _08273_);
  nand (_08278_, _08277_, _08179_);
  nand (_08280_, _08178_, _07911_);
  nand (_08281_, _08280_, _08278_);
  nand (_08282_, _08281_, _08201_);
  nand (_08283_, _08193_, _07926_);
  nand (_25013_[6], _08283_, _08282_);
  nand (_08284_, _08178_, _06606_);
  nand (_08286_, _08180_, _07383_);
  nand (_08287_, _08183_, word_in[7]);
  nand (_08288_, _08184_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_08289_, _08288_, _08287_);
  nor (_08290_, _08289_, _08180_);
  nor (_08291_, _08290_, _08178_);
  nand (_08293_, _08291_, _08286_);
  nand (_08294_, _08293_, _08284_);
  nand (_08295_, _08294_, _08201_);
  nand (_08296_, _08193_, word_in[31]);
  nand (_25013_[7], _08296_, _08295_);
  nor (_08297_, _07258_, _06822_);
  nor (_08298_, _06579_, _06915_);
  nor (_08299_, _06860_, _06591_);
  not (_08300_, _08299_);
  nor (_08302_, _08300_, _07267_);
  not (_08303_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_08304_, _08299_, _08303_);
  nor (_08305_, _08304_, _08302_);
  nor (_08306_, _08305_, _08298_);
  not (_08307_, _08298_);
  nor (_08308_, _08307_, _07272_);
  nor (_08309_, _08308_, _08306_);
  nor (_08310_, _08309_, _08297_);
  nor (_08311_, _06570_, _06444_);
  not (_08312_, _08311_);
  nor (_08313_, _08312_, _06241_);
  not (_08314_, _08313_);
  nand (_08315_, _08297_, word_in[16]);
  nand (_08316_, _08315_, _08314_);
  nor (_08317_, _08316_, _08310_);
  nor (_08318_, _08314_, _07814_);
  nor (_25014_[0], _08318_, _08317_);
  nor (_08319_, _08300_, _07564_);
  not (_08320_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_08321_, _08299_, _08320_);
  nor (_08322_, _08321_, _08319_);
  nor (_08323_, _08322_, _08298_);
  nor (_08325_, _08307_, _07568_);
  nor (_08326_, _08325_, _08323_);
  nor (_08327_, _08326_, _08297_);
  nand (_08328_, _08297_, word_in[17]);
  nand (_08329_, _08328_, _08314_);
  nor (_08330_, _08329_, _08327_);
  nor (_08332_, _08314_, _07833_);
  nor (_25014_[1], _08332_, _08330_);
  nand (_08333_, _08297_, word_in[18]);
  not (_08334_, _08297_);
  nand (_08335_, _08299_, word_in[2]);
  nand (_08336_, _08300_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nand (_08338_, _08336_, _08335_);
  nand (_08339_, _08338_, _08307_);
  nand (_08340_, _08298_, word_in[10]);
  nand (_08341_, _08340_, _08339_);
  nand (_08342_, _08341_, _08334_);
  nand (_08343_, _08342_, _08333_);
  nand (_08346_, _08343_, _08314_);
  nand (_08347_, _08313_, _07856_);
  nand (_25014_[2], _08347_, _08346_);
  nand (_08349_, _08297_, word_in[19]);
  nand (_08350_, _08299_, word_in[3]);
  nand (_08351_, _08300_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nand (_08352_, _08351_, _08350_);
  nand (_08353_, _08352_, _08307_);
  nand (_08354_, _08298_, word_in[11]);
  nand (_08355_, _08354_, _08353_);
  nand (_08357_, _08355_, _08334_);
  nand (_08359_, _08357_, _08349_);
  nand (_08361_, _08359_, _08314_);
  nand (_08362_, _08313_, _07874_);
  nand (_25014_[3], _08362_, _08361_);
  nor (_08364_, _08300_, _07335_);
  not (_08365_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_08366_, _08299_, _08365_);
  nor (_08368_, _08366_, _08364_);
  nor (_08369_, _08368_, _08298_);
  nor (_08370_, _08307_, _07339_);
  nor (_08371_, _08370_, _08369_);
  nor (_08372_, _08371_, _08297_);
  nand (_08374_, _08297_, word_in[20]);
  nand (_08375_, _08374_, _08314_);
  nor (_08376_, _08375_, _08372_);
  nor (_08378_, _08314_, _07892_);
  nor (_25014_[4], _08378_, _08376_);
  nor (_08380_, _08299_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_08382_, _08300_, word_in[5]);
  nor (_08385_, _08382_, _08380_);
  nor (_08387_, _08385_, _08298_);
  nor (_08389_, _08307_, word_in[13]);
  nor (_08390_, _08389_, _08387_);
  nor (_08391_, _08390_, _08297_);
  nor (_08392_, _08334_, word_in[21]);
  nor (_08393_, _08392_, _08391_);
  nor (_08395_, _08393_, _08313_);
  nor (_08396_, _08314_, _07908_);
  nor (_25014_[5], _08396_, _08395_);
  nor (_08397_, _08300_, _07364_);
  not (_08398_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_08399_, _08299_, _08398_);
  nor (_08400_, _08399_, _08397_);
  nor (_08401_, _08400_, _08298_);
  nor (_08402_, _08307_, _07368_);
  nor (_08403_, _08402_, _08401_);
  nor (_08404_, _08403_, _08297_);
  nand (_08405_, _08297_, word_in[22]);
  nand (_08406_, _08405_, _08314_);
  nor (_08408_, _08406_, _08404_);
  nor (_08409_, _08314_, _07926_);
  nor (_25014_[6], _08409_, _08408_);
  nor (_08411_, _08300_, _07379_);
  not (_08412_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_08413_, _08299_, _08412_);
  nor (_08414_, _08413_, _08411_);
  nor (_08415_, _08414_, _08298_);
  nor (_08416_, _08307_, _07383_);
  nor (_08417_, _08416_, _08415_);
  nor (_08418_, _08417_, _08297_);
  nand (_08419_, _06606_, _06821_);
  nand (_08420_, _08419_, _08314_);
  nor (_08421_, _08420_, _08418_);
  nor (_08422_, _08314_, _06610_);
  nor (_25014_[7], _08422_, _08421_);
  nor (_08423_, _07226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1]);
  nor (_08424_, _07228_, _21474_);
  nor (_00614_, _08424_, _08423_);
  nor (_08426_, _22531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5]);
  nor (_08428_, _22533_, _21451_);
  nor (_00630_, _08428_, _08426_);
  nor (_08429_, _07402_, _06218_);
  nor (_08430_, _06910_, _06591_);
  nor (_08431_, _08430_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  not (_08432_, _08430_);
  nor (_08433_, _08432_, word_in[0]);
  nor (_08434_, _08433_, _08431_);
  nor (_08435_, _08434_, _08429_);
  nor (_08436_, _07399_, _06355_);
  not (_08437_, _08436_);
  nand (_08439_, _08429_, _07272_);
  nand (_08441_, _08439_, _08437_);
  nor (_08442_, _08441_, _08435_);
  nor (_08444_, _08312_, _06191_);
  not (_08446_, _08444_);
  nand (_08448_, _08436_, _07794_);
  nand (_08449_, _08448_, _08446_);
  nor (_08451_, _08449_, _08442_);
  nor (_08453_, _08446_, _07814_);
  nor (_25015_[0], _08453_, _08451_);
  nor (_08456_, _08432_, _07564_);
  not (_08457_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_08458_, _08430_, _08457_);
  nor (_08459_, _08458_, _08456_);
  nor (_08460_, _08459_, _08429_);
  not (_08461_, _08429_);
  nor (_08462_, _08461_, _07568_);
  nor (_08463_, _08462_, _08460_);
  nand (_08465_, _08463_, _08437_);
  nor (_08466_, _08437_, _07817_);
  nor (_08467_, _08466_, _08444_);
  nand (_08468_, _08467_, _08465_);
  nand (_08469_, _08444_, _07833_);
  nand (_25015_[1], _08469_, _08468_);
  nor (_08470_, _08432_, _07303_);
  not (_08472_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_08474_, _08430_, _08472_);
  nor (_08475_, _08474_, _08470_);
  nor (_08477_, _08475_, _08429_);
  nor (_08478_, _08461_, _07307_);
  nor (_08479_, _08478_, _08477_);
  nand (_08480_, _08479_, _08437_);
  nor (_08481_, _08437_, _07847_);
  nor (_08483_, _08481_, _08444_);
  nand (_08485_, _08483_, _08480_);
  nand (_08487_, _08444_, _07856_);
  nand (_25015_[2], _08487_, _08485_);
  not (_08488_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nand (_08489_, _08432_, _08488_);
  nand (_08491_, _08430_, _07319_);
  nand (_08492_, _08491_, _08489_);
  nand (_08493_, _08492_, _08461_);
  nand (_08494_, _08429_, _07324_);
  nand (_08495_, _08494_, _08493_);
  nand (_08496_, _08495_, _08437_);
  nor (_08497_, _08437_, _07869_);
  nor (_08499_, _08497_, _08444_);
  nand (_08500_, _08499_, _08496_);
  nand (_08501_, _08444_, _07874_);
  nand (_25015_[3], _08501_, _08500_);
  nor (_08502_, _08430_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_08503_, _08432_, word_in[4]);
  nor (_08504_, _08503_, _08502_);
  nor (_08505_, _08504_, _08429_);
  nand (_08506_, _08429_, _07339_);
  nand (_08508_, _08506_, _08437_);
  nor (_08509_, _08508_, _08505_);
  nand (_08510_, _08436_, _07887_);
  nand (_08511_, _08510_, _08446_);
  nor (_08513_, _08511_, _08509_);
  nor (_08515_, _08446_, _07892_);
  nor (_25015_[4], _08515_, _08513_);
  nor (_08517_, _08432_, _07349_);
  not (_08519_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_08521_, _08430_, _08519_);
  nor (_08523_, _08521_, _08517_);
  nor (_08524_, _08523_, _08429_);
  nor (_08525_, _08461_, _07353_);
  nor (_08526_, _08525_, _08524_);
  nor (_08529_, _08526_, _08436_);
  nand (_08530_, _08436_, _07896_);
  nand (_08531_, _08530_, _08446_);
  nor (_08532_, _08531_, _08529_);
  nor (_08533_, _08446_, _07908_);
  nor (_25015_[5], _08533_, _08532_);
  not (_08535_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nand (_08536_, _08432_, _08535_);
  nand (_08538_, _08430_, _07364_);
  nand (_08539_, _08538_, _08536_);
  nand (_08540_, _08539_, _08461_);
  nand (_08541_, _08429_, _07368_);
  nand (_08542_, _08541_, _08540_);
  nand (_08543_, _08542_, _08437_);
  nor (_08544_, _08437_, _07911_);
  nor (_08545_, _08544_, _08444_);
  nand (_08546_, _08545_, _08543_);
  nand (_08547_, _08444_, _07926_);
  nand (_25015_[6], _08547_, _08546_);
  nor (_08548_, _08432_, _07379_);
  not (_08551_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor (_08552_, _08430_, _08551_);
  nor (_08553_, _08552_, _08548_);
  nor (_08554_, _08553_, _08429_);
  nor (_08555_, _08461_, _07383_);
  nor (_08556_, _08555_, _08554_);
  nor (_08557_, _08556_, _08436_);
  nand (_08558_, _08436_, _06606_);
  nand (_08559_, _08558_, _08446_);
  nor (_08560_, _08559_, _08557_);
  nor (_08561_, _08446_, _06610_);
  nor (_25015_[7], _08561_, _08560_);
  nor (_08562_, _07226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  nor (_08563_, _07228_, _21586_);
  nor (_00679_, _08563_, _08562_);
  nor (_08564_, _07537_, _06218_);
  nor (_08565_, _06927_, _06591_);
  nor (_08567_, _08565_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  not (_08568_, _08565_);
  nor (_08569_, _08568_, word_in[0]);
  nor (_08571_, _08569_, _08567_);
  nor (_08572_, _08571_, _08564_);
  nor (_08573_, _07532_, _06355_);
  not (_08574_, _08573_);
  nand (_08575_, _08564_, _07272_);
  nand (_08576_, _08575_, _08574_);
  nor (_08577_, _08576_, _08572_);
  nor (_08578_, _08312_, _06192_);
  not (_08579_, _08578_);
  nand (_08580_, _08573_, _07794_);
  nand (_08581_, _08580_, _08579_);
  nor (_08582_, _08581_, _08577_);
  nor (_08583_, _08579_, word_in[24]);
  nor (_24965_, _08583_, _08582_);
  not (_08584_, _08564_);
  not (_08586_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nand (_08587_, _08568_, _08586_);
  nand (_08588_, _08565_, _07564_);
  nand (_08590_, _08588_, _08587_);
  nand (_08591_, _08590_, _08584_);
  nand (_08592_, _08564_, _07568_);
  nand (_08593_, _08592_, _08591_);
  nand (_08594_, _08593_, _08574_);
  nor (_08595_, _08574_, _07817_);
  nor (_08596_, _08595_, _08578_);
  nand (_08597_, _08596_, _08594_);
  nand (_08598_, _08578_, _07833_);
  nand (_24966_, _08598_, _08597_);
  nand (_08600_, _08568_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nand (_08602_, _08565_, word_in[2]);
  nand (_08603_, _08602_, _08600_);
  nand (_08604_, _08603_, _08584_);
  nand (_08605_, _08564_, word_in[10]);
  nand (_08606_, _08605_, _08604_);
  nand (_08608_, _08606_, _08574_);
  nand (_08610_, _08573_, _07847_);
  nand (_08611_, _08610_, _08608_);
  nand (_08612_, _08611_, _08579_);
  nand (_08613_, _08578_, word_in[26]);
  nand (_24967_, _08613_, _08612_);
  not (_08615_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nand (_08616_, _08568_, _08615_);
  nand (_08617_, _08565_, _07319_);
  nand (_08618_, _08617_, _08616_);
  nand (_08619_, _08618_, _08584_);
  nand (_08621_, _08564_, _07324_);
  nand (_08622_, _08621_, _08619_);
  nand (_08623_, _08622_, _08574_);
  nor (_08624_, _08574_, _07869_);
  nor (_08625_, _08624_, _08578_);
  nand (_08626_, _08625_, _08623_);
  nand (_08627_, _08578_, _07874_);
  nand (_24968_, _08627_, _08626_);
  nor (_08628_, _08568_, _07335_);
  not (_08629_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_08630_, _08565_, _08629_);
  nor (_08631_, _08630_, _08628_);
  nor (_08632_, _08631_, _08564_);
  nor (_08633_, _08584_, _07339_);
  nor (_08634_, _08633_, _08632_);
  nand (_08636_, _08634_, _08574_);
  nor (_08637_, _08574_, _07887_);
  nor (_08638_, _08637_, _08578_);
  nand (_08639_, _08638_, _08636_);
  nand (_08640_, _08578_, word_in[28]);
  nand (_24969_, _08640_, _08639_);
  nor (_08641_, _08568_, _07349_);
  not (_08642_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_08643_, _08565_, _08642_);
  nor (_08644_, _08643_, _08641_);
  nor (_08645_, _08644_, _08564_);
  nor (_08646_, _08584_, _07353_);
  nor (_08647_, _08646_, _08645_);
  nor (_08648_, _08647_, _08573_);
  nand (_08649_, _08573_, _07896_);
  nand (_08651_, _08649_, _08579_);
  nor (_08653_, _08651_, _08648_);
  nor (_08654_, _08579_, _07908_);
  nor (_24970_, _08654_, _08653_);
  nor (_08655_, _08568_, _07364_);
  not (_08658_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_08659_, _08565_, _08658_);
  nor (_08660_, _08659_, _08655_);
  nor (_08661_, _08660_, _08564_);
  nor (_08663_, _08584_, _07368_);
  nor (_08664_, _08663_, _08661_);
  nor (_08666_, _08664_, _08573_);
  nand (_08667_, _08573_, _07911_);
  nand (_08669_, _08667_, _08579_);
  nor (_08670_, _08669_, _08666_);
  nor (_08671_, _08579_, _07926_);
  nor (_24971_, _08671_, _08670_);
  not (_08672_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nor (_08673_, _08565_, _08672_);
  nor (_08674_, _06927_, _07508_);
  nor (_08675_, _08674_, _08673_);
  nor (_08676_, _08675_, _08564_);
  nor (_08677_, _08584_, _07383_);
  nor (_08679_, _08677_, _08676_);
  nor (_08681_, _08679_, _08573_);
  nand (_08682_, _08573_, _06606_);
  nand (_08683_, _08682_, _08579_);
  nor (_08684_, _08683_, _08681_);
  nor (_08685_, _08579_, _06610_);
  nor (_24972_, _08685_, _08684_);
  not (_08686_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_08687_, _23046_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  nor (_08688_, _08687_, _08686_);
  not (_08690_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_08692_, _08687_);
  nor (_08693_, _08692_, _08690_);
  nor (_08694_, _08693_, _08688_);
  nor (_00735_, _08694_, rst);
  nor (_08695_, _08687_, _08690_);
  not (_08696_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_08697_, _08692_, _08696_);
  nor (_08698_, _08697_, _08695_);
  nor (_00758_, _08698_, rst);
  nor (_08700_, _06860_, _06568_);
  not (_08701_, _08700_);
  nor (_08703_, _07660_, _06355_);
  nor (_08704_, _07666_, _06218_);
  not (_08706_, _06976_);
  nor (_08707_, _08706_, _06591_);
  not (_08708_, _08707_);
  nand (_08709_, _08708_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nand (_08710_, _07669_, _06976_);
  nand (_08711_, _08710_, _08709_);
  nor (_08712_, _08711_, _08704_);
  not (_08713_, _08704_);
  nor (_08714_, _08713_, word_in[8]);
  nor (_08715_, _08714_, _08712_);
  nor (_08716_, _08715_, _08703_);
  not (_08718_, _08703_);
  nor (_08719_, _08718_, _07794_);
  nor (_08720_, _08719_, _08716_);
  nand (_08721_, _08720_, _08701_);
  nand (_08722_, _08700_, word_in[24]);
  nand (_24973_, _08722_, _08721_);
  nand (_08723_, _08703_, _07817_);
  nand (_08724_, _08708_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nand (_08725_, _08707_, _07685_);
  nand (_08726_, _08725_, _08724_);
  nand (_08727_, _08726_, _08713_);
  nand (_08728_, _08704_, word_in[9]);
  nand (_08729_, _08728_, _08727_);
  nand (_08731_, _08729_, _08718_);
  nand (_08732_, _08731_, _08723_);
  nand (_08733_, _08732_, _08701_);
  nand (_08735_, _08700_, word_in[25]);
  nand (_24974_, _08735_, _08733_);
  nand (_08736_, _07856_, _06859_);
  nor (_08737_, _08708_, _07303_);
  not (_08738_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_08739_, _08707_, _08738_);
  nor (_08740_, _08739_, _08737_);
  nor (_08741_, _08740_, _08704_);
  nor (_08742_, _08713_, _07307_);
  nor (_08743_, _08742_, _08741_);
  nand (_08744_, _08743_, _08718_);
  nor (_08745_, _08718_, _07847_);
  nor (_08746_, _08745_, _08700_);
  nand (_08747_, _08746_, _08744_);
  nand (_24975_, _08747_, _08736_);
  not (_08749_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nand (_08750_, _08708_, _08749_);
  nand (_08752_, _08707_, _07319_);
  nand (_08753_, _08752_, _08750_);
  nand (_08755_, _08753_, _08713_);
  nand (_08757_, _08704_, _07324_);
  nand (_08759_, _08757_, _08755_);
  nand (_08760_, _08759_, _08718_);
  nor (_08762_, _08718_, _07869_);
  nor (_08764_, _08762_, _08700_);
  nand (_08766_, _08764_, _08760_);
  nand (_08767_, _08700_, word_in[27]);
  nand (_24976_, _08767_, _08766_);
  not (_08769_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nand (_08770_, _08708_, _08769_);
  nand (_08772_, _08707_, _07335_);
  nand (_08774_, _08772_, _08770_);
  nand (_08776_, _08774_, _08713_);
  nand (_08777_, _08704_, _07339_);
  nand (_08779_, _08777_, _08776_);
  nand (_08781_, _08779_, _08718_);
  nor (_08783_, _08718_, _07887_);
  nor (_08785_, _08783_, _08700_);
  nand (_08787_, _08785_, _08781_);
  nand (_08788_, _08700_, word_in[28]);
  nand (_24977_, _08788_, _08787_);
  nand (_08792_, _07908_, _06859_);
  nor (_08794_, _08708_, _07349_);
  not (_08796_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_08797_, _08707_, _08796_);
  nor (_08798_, _08797_, _08794_);
  nor (_08800_, _08798_, _08704_);
  nor (_08802_, _08713_, _07353_);
  nor (_08803_, _08802_, _08800_);
  nand (_08805_, _08803_, _08718_);
  nor (_08807_, _08718_, _07896_);
  nor (_08809_, _08807_, _08700_);
  nand (_08810_, _08809_, _08805_);
  nand (_24978_, _08810_, _08792_);
  nand (_08811_, _07926_, _06859_);
  not (_08812_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_08813_, _08707_, _08812_);
  nor (_08815_, _08708_, _07364_);
  nor (_08816_, _08815_, _08813_);
  nor (_08818_, _08816_, _08704_);
  nor (_08819_, _08713_, _07368_);
  nor (_08821_, _08819_, _08818_);
  nand (_08823_, _08821_, _08718_);
  nor (_08824_, _08718_, _07911_);
  nor (_08826_, _08824_, _08700_);
  nand (_08828_, _08826_, _08823_);
  nand (_24979_, _08828_, _08811_);
  nor (_08830_, _21741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1]);
  nor (_08832_, _21744_, _21474_);
  nor (_25240_, _08832_, _08830_);
  nand (_08834_, _08703_, _06606_);
  nand (_08835_, _08708_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_08837_, _06976_, _07507_);
  nand (_08838_, _08837_, _08835_);
  nand (_08839_, _08838_, _08713_);
  nand (_08840_, _08704_, word_in[15]);
  nand (_08841_, _08840_, _08839_);
  nand (_08842_, _08841_, _08718_);
  nand (_08844_, _08842_, _08834_);
  nand (_08845_, _08844_, _08701_);
  nand (_08846_, _08700_, word_in[31]);
  nand (_24980_, _08846_, _08845_);
  nor (_08847_, _23557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  nor (_08848_, _23560_, _21504_);
  nor (_00787_, _08848_, _08847_);
  nor (_08849_, _06570_, _06034_);
  not (_08850_, _08849_);
  nor (_08852_, _08706_, _06579_);
  nor (_08854_, _06075_, _06098_);
  nand (_08855_, _08854_, _06590_);
  not (_08857_, _08855_);
  nor (_08858_, _08857_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_08859_, _08855_, word_in[0]);
  nor (_08860_, _08859_, _08858_);
  nor (_08861_, _08860_, _08852_);
  nand (_08863_, _06277_, word_in[8]);
  nor (_08864_, _08863_, rst);
  not (_08865_, _08852_);
  nor (_08867_, _08865_, _08864_);
  nor (_08869_, _08867_, _08861_);
  not (_08870_, _06576_);
  nand (_08871_, _06575_, _06191_);
  nand (_08873_, _08871_, _08870_);
  not (_08874_, _08873_);
  nor (_08876_, _08874_, _08869_);
  nand (_08878_, _08870_, _06091_);
  nor (_08879_, _08878_, _07794_);
  nor (_08880_, _08879_, _08876_);
  nand (_08881_, _08880_, _08850_);
  nand (_08882_, _08849_, _07814_);
  nand (_25006_[0], _08882_, _08881_);
  nor (_08883_, _08857_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_08884_, _08855_, word_in[1]);
  nor (_08885_, _08884_, _08883_);
  nor (_08887_, _08885_, _08852_);
  nor (_08888_, _08865_, _07292_);
  nor (_08890_, _08888_, _08887_);
  nor (_08891_, _08890_, _08874_);
  nor (_08892_, _08873_, _07817_);
  nor (_08893_, _08892_, _08891_);
  nor (_08894_, _08893_, _08849_);
  nor (_08895_, _08850_, word_in[25]);
  nor (_25006_[1], _08895_, _08894_);
  nor (_08896_, _08878_, _07847_);
  nor (_08898_, _08857_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_08899_, _08855_, word_in[2]);
  nor (_08900_, _08899_, _08898_);
  nor (_08901_, _08900_, _08852_);
  nand (_08902_, _06277_, word_in[10]);
  nor (_08903_, _08902_, rst);
  nor (_08904_, _08865_, _08903_);
  nor (_08906_, _08904_, _08901_);
  nor (_08907_, _08906_, _08874_);
  nor (_08908_, _08907_, _08896_);
  nand (_08909_, _08908_, _08850_);
  nand (_08911_, _08849_, _07856_);
  nand (_25006_[2], _08911_, _08909_);
  nor (_08912_, _08857_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_08913_, _08855_, word_in[3]);
  nor (_08915_, _08913_, _08912_);
  nor (_08916_, _08915_, _08852_);
  nand (_08917_, _06277_, word_in[11]);
  nor (_08918_, _08917_, rst);
  nor (_08920_, _08865_, _08918_);
  nor (_08921_, _08920_, _08916_);
  nor (_08923_, _08921_, _08874_);
  nor (_08924_, _08878_, _07869_);
  nor (_08925_, _08924_, _08923_);
  nand (_08926_, _08925_, _08850_);
  nand (_08927_, _08849_, _07874_);
  nand (_25006_[3], _08927_, _08926_);
  nor (_08931_, _08857_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_08932_, _08855_, word_in[4]);
  nor (_08933_, _08932_, _08931_);
  nor (_08934_, _08933_, _08852_);
  nand (_08936_, _06277_, word_in[12]);
  nor (_08937_, _08936_, rst);
  nor (_08939_, _08865_, _08937_);
  nor (_08940_, _08939_, _08934_);
  nor (_08941_, _08940_, _08874_);
  nor (_08942_, _08873_, _07887_);
  nor (_08943_, _08942_, _08941_);
  nor (_08944_, _08943_, _08849_);
  nor (_08945_, _08850_, word_in[28]);
  nor (_25006_[4], _08945_, _08944_);
  nor (_08946_, _08878_, _07896_);
  nor (_08948_, _08857_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_08949_, _08855_, word_in[5]);
  nor (_08951_, _08949_, _08948_);
  nor (_08953_, _08951_, _08852_);
  nand (_08955_, _06277_, word_in[13]);
  nor (_08957_, _08955_, rst);
  nor (_08959_, _08865_, _08957_);
  nor (_08960_, _08959_, _08953_);
  nor (_08961_, _08960_, _08874_);
  nor (_08962_, _08961_, _08946_);
  nand (_08964_, _08962_, _08850_);
  nand (_08966_, _08849_, _07908_);
  nand (_25006_[5], _08966_, _08964_);
  nor (_08968_, _08857_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_08970_, _08855_, word_in[6]);
  nor (_08972_, _08970_, _08968_);
  nor (_08973_, _08972_, _08852_);
  nand (_08974_, _06277_, word_in[14]);
  nor (_08975_, _08974_, rst);
  nor (_08976_, _08865_, _08975_);
  nor (_08978_, _08976_, _08973_);
  nor (_08979_, _08978_, _08874_);
  nor (_08980_, _08873_, _07911_);
  nor (_08982_, _08980_, _08979_);
  nor (_08984_, _08982_, _08849_);
  nor (_08985_, _08850_, word_in[30]);
  nor (_25006_[6], _08985_, _08984_);
  nand (_08987_, _08854_, _07507_);
  nand (_08989_, _08855_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_08991_, _08989_, _08987_);
  nand (_08993_, _08991_, _08865_);
  nand (_08994_, _08852_, _06600_);
  nand (_08996_, _08994_, _08993_);
  nand (_08997_, _08996_, _08873_);
  nand (_08998_, _08874_, _06606_);
  nand (_08999_, _08998_, _08997_);
  nand (_09000_, _08999_, _08850_);
  nand (_09001_, _08849_, word_in[31]);
  nand (_25006_[7], _09001_, _09000_);
  nor (_09002_, _01183_, _21638_);
  nor (_09003_, _09002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7]);
  not (_09004_, _09002_);
  nor (_09006_, _09004_, _21626_);
  nor (_00846_, _09006_, _09003_);
  nor (_09007_, _24380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5]);
  nor (_09009_, _24382_, _21451_);
  nor (_25293_, _09009_, _09007_);
  nor (_09010_, _06572_, _06191_);
  not (_09012_, _09010_);
  nor (_09013_, _06576_, _06192_);
  nor (_09014_, _06583_, _06075_);
  nor (_09015_, _07040_, _06591_);
  nor (_09016_, _09015_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  not (_09017_, _09015_);
  nor (_09018_, _09017_, word_in[0]);
  nor (_09019_, _09018_, _09016_);
  nor (_09020_, _09019_, _09014_);
  not (_09021_, _09014_);
  nor (_09022_, _09021_, _08864_);
  nor (_09023_, _09022_, _09020_);
  nor (_09024_, _09023_, _09013_);
  not (_09025_, _09013_);
  nor (_09026_, _09025_, word_in[16]);
  nor (_09027_, _09026_, _09024_);
  nand (_09028_, _09027_, _09012_);
  nand (_09029_, _09010_, _07814_);
  nand (_24981_, _09029_, _09028_);
  nor (_09030_, _09025_, word_in[17]);
  nor (_09031_, _09015_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_09032_, _09017_, word_in[1]);
  nor (_09033_, _09032_, _09031_);
  nor (_09034_, _09033_, _09014_);
  nor (_09035_, _09021_, _07292_);
  nor (_09036_, _09035_, _09034_);
  nor (_09037_, _09036_, _09013_);
  nor (_09038_, _09037_, _09030_);
  nand (_09039_, _09038_, _09012_);
  nand (_09040_, _09010_, _07833_);
  nand (_24982_, _09040_, _09039_);
  nand (_09041_, _09015_, word_in[2]);
  nand (_09042_, _09017_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand (_09043_, _09042_, _09041_);
  nand (_09044_, _09043_, _09021_);
  nand (_09045_, _09014_, _08903_);
  nand (_09046_, _09045_, _09044_);
  nand (_09047_, _09046_, _09025_);
  nand (_09048_, _09013_, word_in[18]);
  nand (_09049_, _09048_, _09047_);
  nand (_09050_, _09049_, _09012_);
  nand (_09051_, _09010_, _07856_);
  nand (_24983_, _09051_, _09050_);
  nor (_09052_, _09015_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_09053_, _09017_, word_in[3]);
  nor (_09054_, _09053_, _09052_);
  nor (_09055_, _09054_, _09014_);
  nor (_09057_, _09021_, _08918_);
  nor (_09058_, _09057_, _09055_);
  nor (_09060_, _09058_, _09013_);
  nor (_09062_, _09025_, word_in[19]);
  nor (_09063_, _09062_, _09060_);
  nor (_09065_, _09063_, _09010_);
  nor (_09066_, _09012_, _07874_);
  nor (_24984_, _09066_, _09065_);
  nor (_09067_, _09025_, word_in[20]);
  nor (_09068_, _09015_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_09069_, _09017_, word_in[4]);
  nor (_09070_, _09069_, _09068_);
  nor (_09071_, _09070_, _09014_);
  nor (_09072_, _09021_, _08937_);
  nor (_09073_, _09072_, _09071_);
  nor (_09074_, _09073_, _09013_);
  nor (_09075_, _09074_, _09067_);
  nand (_09076_, _09075_, _09012_);
  nand (_09078_, _09010_, _07892_);
  nand (_24985_, _09078_, _09076_);
  nor (_09079_, _09015_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_09080_, _09017_, word_in[5]);
  nor (_09081_, _09080_, _09079_);
  nor (_09082_, _09081_, _09014_);
  nor (_09083_, _09021_, _08957_);
  nor (_09084_, _09083_, _09082_);
  nor (_09085_, _09084_, _09013_);
  nor (_09086_, _09025_, word_in[21]);
  nor (_09087_, _09086_, _09085_);
  nand (_09088_, _09087_, _09012_);
  nand (_09089_, _09010_, _07908_);
  nand (_24986_, _09089_, _09088_);
  nor (_09091_, _09015_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_09092_, _09017_, word_in[6]);
  nor (_09093_, _09092_, _09091_);
  nor (_09094_, _09093_, _09014_);
  nor (_09095_, _09021_, _08975_);
  nor (_09096_, _09095_, _09094_);
  nor (_09097_, _09096_, _09013_);
  nor (_09098_, _09025_, word_in[22]);
  nor (_09099_, _09098_, _09097_);
  nand (_09100_, _09099_, _09012_);
  nand (_09102_, _09010_, _07926_);
  nand (_24987_, _09102_, _09100_);
  nor (_09103_, _09015_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_09104_, _09017_, word_in[7]);
  nor (_09105_, _09104_, _09103_);
  nor (_09106_, _09105_, _09014_);
  nor (_09108_, _09021_, _06600_);
  nor (_09109_, _09108_, _09106_);
  nor (_09110_, _09109_, _09013_);
  nor (_09111_, _09025_, word_in[23]);
  nor (_09112_, _09111_, _09110_);
  nor (_09113_, _09112_, _09010_);
  nor (_09114_, _09012_, _06610_);
  nor (_24988_, _09114_, _09113_);
  nor (_09115_, _06572_, _06192_);
  not (_09116_, _09115_);
  nor (_09117_, _06576_, _06075_);
  nand (_09118_, _09117_, word_in[16]);
  not (_09119_, _09117_);
  nor (_09120_, _06583_, _06241_);
  not (_09121_, _09120_);
  nor (_09122_, _06591_, _07257_);
  nand (_09123_, _09122_, word_in[0]);
  not (_09124_, _09122_);
  nand (_09125_, _09124_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nand (_09127_, _09125_, _09123_);
  nand (_09128_, _09127_, _09121_);
  nand (_09129_, _09120_, _08864_);
  nand (_09130_, _09129_, _09128_);
  nand (_09131_, _09130_, _09119_);
  nand (_09132_, _09131_, _09118_);
  nand (_09133_, _09132_, _09116_);
  nand (_09134_, _09115_, _07814_);
  nand (_25007_[0], _09134_, _09133_);
  nand (_09135_, _09122_, word_in[1]);
  nand (_09136_, _09124_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nand (_09137_, _09136_, _09135_);
  nand (_09138_, _09137_, _09121_);
  nand (_09139_, _09120_, _07292_);
  nand (_09140_, _09139_, _09138_);
  nand (_09141_, _09140_, _09119_);
  nand (_09142_, _09117_, word_in[17]);
  nand (_09143_, _09142_, _09141_);
  nand (_09144_, _09143_, _09116_);
  nand (_09145_, _09115_, _07833_);
  nand (_25007_[1], _09145_, _09144_);
  nand (_09146_, _09122_, word_in[2]);
  nand (_09147_, _09124_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand (_09149_, _09147_, _09146_);
  nand (_09150_, _09149_, _09121_);
  nand (_09151_, _09120_, _08903_);
  nand (_09152_, _09151_, _09150_);
  nand (_09153_, _09152_, _09119_);
  nand (_09154_, _09117_, word_in[18]);
  nand (_09155_, _09154_, _09153_);
  nand (_09156_, _09155_, _09116_);
  nand (_09157_, _09115_, _07856_);
  nand (_25007_[2], _09157_, _09156_);
  nor (_09158_, _09122_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_09159_, _09124_, word_in[3]);
  nor (_09160_, _09159_, _09158_);
  nor (_09161_, _09160_, _09120_);
  nor (_09162_, _09121_, _08918_);
  nor (_09163_, _09162_, _09161_);
  nor (_09164_, _09163_, _09117_);
  nor (_09165_, _09119_, word_in[19]);
  nor (_09166_, _09165_, _09164_);
  nand (_09167_, _09166_, _09116_);
  nand (_09168_, _09115_, _07874_);
  nand (_25007_[3], _09168_, _09167_);
  nor (_09169_, _09119_, word_in[20]);
  nor (_09170_, _09122_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_09171_, _09124_, word_in[4]);
  nor (_09172_, _09171_, _09170_);
  nor (_09173_, _09172_, _09120_);
  nor (_09174_, _09121_, _08937_);
  nor (_09175_, _09174_, _09173_);
  nor (_09176_, _09175_, _09117_);
  nor (_09177_, _09176_, _09169_);
  nor (_09178_, _09177_, _09115_);
  nor (_09179_, _09116_, _07892_);
  nor (_25007_[4], _09179_, _09178_);
  nand (_09180_, _09122_, word_in[5]);
  nand (_09181_, _09124_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nand (_09182_, _09181_, _09180_);
  nand (_09183_, _09182_, _09121_);
  nand (_09184_, _09120_, _08957_);
  nand (_09185_, _09184_, _09183_);
  nand (_09186_, _09185_, _09119_);
  nand (_09187_, _09117_, word_in[21]);
  nand (_09188_, _09187_, _09186_);
  nand (_09189_, _09188_, _09116_);
  nand (_09190_, _09115_, _07908_);
  nand (_25007_[5], _09190_, _09189_);
  nand (_09191_, _09122_, word_in[6]);
  nand (_09192_, _09124_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nand (_09193_, _09192_, _09191_);
  nand (_09194_, _09193_, _09121_);
  nand (_09195_, _09120_, _08975_);
  nand (_09196_, _09195_, _09194_);
  nand (_09197_, _09196_, _09119_);
  nand (_09198_, _09117_, word_in[22]);
  nand (_09199_, _09198_, _09197_);
  nand (_09200_, _09199_, _09116_);
  nand (_09201_, _09115_, _07926_);
  nand (_25007_[6], _09201_, _09200_);
  nor (_09202_, _09122_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nor (_09203_, _09124_, word_in[7]);
  nor (_09204_, _09203_, _09202_);
  nor (_09205_, _09204_, _09120_);
  nor (_09206_, _09121_, _06600_);
  nor (_09207_, _09206_, _09205_);
  nor (_09208_, _09207_, _09117_);
  nor (_09209_, _09119_, word_in[23]);
  nor (_09210_, _09209_, _09208_);
  nor (_09211_, _09210_, _09115_);
  nor (_09212_, _09116_, _06610_);
  nor (_25007_[7], _09212_, _09211_);
  nor (_09213_, _06595_, _07267_);
  not (_09214_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_09215_, _06592_, _09214_);
  nor (_09216_, _09215_, _09213_);
  nor (_09217_, _09216_, _06585_);
  nand (_09218_, _08864_, _06585_);
  nand (_09219_, _09218_, _06605_);
  nor (_09220_, _09219_, _09217_);
  nor (_09221_, _07794_, _06605_);
  nor (_09222_, _09221_, _09220_);
  nand (_09223_, _09222_, _06574_);
  nand (_09224_, _07814_, _06573_);
  nand (_25008_[0], _09224_, _09223_);
  nor (_09225_, _21653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  nor (_09226_, _21655_, _21554_);
  nor (_01008_, _09226_, _09225_);
  nor (_09227_, _06595_, _07564_);
  not (_09228_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_09229_, _06592_, _09228_);
  nor (_09230_, _09229_, _09227_);
  nor (_09231_, _09230_, _06585_);
  nand (_09232_, _07292_, _06585_);
  nand (_09233_, _09232_, _06605_);
  nor (_09234_, _09233_, _09231_);
  nor (_09235_, _07817_, _06605_);
  nor (_09236_, _09235_, _09234_);
  nand (_09237_, _09236_, _06574_);
  nand (_09238_, _07833_, _06573_);
  nand (_25008_[1], _09238_, _09237_);
  nor (_09239_, _06595_, _07303_);
  not (_09240_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_09241_, _06592_, _09240_);
  nor (_09242_, _09241_, _09239_);
  nor (_09243_, _09242_, _06585_);
  nand (_09244_, _08903_, _06585_);
  nand (_09245_, _09244_, _06605_);
  nor (_09246_, _09245_, _09243_);
  nor (_09247_, _07847_, _06605_);
  nor (_09248_, _09247_, _09246_);
  nand (_09249_, _09248_, _06574_);
  nand (_09250_, _07856_, _06573_);
  nand (_25008_[2], _09250_, _09249_);
  nor (_09251_, _06595_, _07319_);
  not (_09252_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_09253_, _06592_, _09252_);
  nor (_09254_, _09253_, _09251_);
  nor (_09255_, _09254_, _06585_);
  nand (_09256_, _08918_, _06585_);
  nand (_09257_, _09256_, _06605_);
  nor (_09258_, _09257_, _09255_);
  nor (_09259_, _07869_, _06605_);
  nor (_09260_, _09259_, _09258_);
  nand (_09261_, _09260_, _06574_);
  nand (_09262_, _07874_, _06573_);
  nand (_25008_[3], _09262_, _09261_);
  nor (_09263_, _06595_, _07335_);
  not (_09264_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_09265_, _06592_, _09264_);
  nor (_09266_, _09265_, _09263_);
  nor (_09267_, _09266_, _06585_);
  nand (_09268_, _08937_, _06585_);
  nand (_09269_, _09268_, _06605_);
  nor (_09270_, _09269_, _09267_);
  nor (_09271_, _07887_, _06605_);
  nor (_09272_, _09271_, _09270_);
  nand (_09273_, _09272_, _06574_);
  nand (_09274_, _07892_, _06573_);
  nand (_25008_[4], _09274_, _09273_);
  nor (_09275_, _06595_, _07349_);
  not (_09276_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_09277_, _06592_, _09276_);
  nor (_09278_, _09277_, _09275_);
  nor (_09279_, _09278_, _06585_);
  nand (_09280_, _08957_, _06585_);
  nand (_09281_, _09280_, _06605_);
  nor (_09282_, _09281_, _09279_);
  nor (_09283_, _07896_, _06605_);
  nor (_09284_, _09283_, _09282_);
  nand (_09285_, _09284_, _06574_);
  nand (_09286_, _07908_, _06573_);
  nand (_25008_[5], _09286_, _09285_);
  nor (_09287_, _06595_, _07364_);
  not (_09288_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_09289_, _06592_, _09288_);
  nor (_09290_, _09289_, _09287_);
  nor (_09291_, _09290_, _06585_);
  nand (_09292_, _08975_, _06585_);
  nand (_09293_, _09292_, _06605_);
  nor (_09294_, _09293_, _09291_);
  nor (_09295_, _07911_, _06605_);
  nor (_09296_, _09295_, _09294_);
  nand (_09297_, _09296_, _06574_);
  nand (_09298_, _07926_, _06573_);
  nand (_25008_[6], _09298_, _09297_);
  nor (_09299_, _21653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  nor (_09300_, _21655_, _21414_);
  nor (_01019_, _09300_, _09299_);
  nor (_09301_, _21777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5]);
  nor (_09302_, _21779_, _21451_);
  nor (_01221_, _09302_, _09301_);
  nor (_09303_, _21777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  nor (_09304_, _21779_, _21526_);
  nor (_01225_, _09304_, _09303_);
  nor (_09305_, _24043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5]);
  nor (_09306_, _24045_, _21451_);
  nor (_25360_, _09306_, _09305_);
  nor (_09307_, _06027_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor (_09308_, _06026_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor (_09309_, _09308_, _09307_);
  nand (_09310_, _09309_, _06031_);
  nor (_09311_, _06027_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_09312_, _06026_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_09313_, _09312_, _09311_);
  nand (_09314_, _09313_, _06089_);
  nand (_09315_, _09314_, _09310_);
  nand (_09316_, _09315_, _06021_);
  nor (_09317_, _06027_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_09318_, _06026_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_09319_, _09318_, _09317_);
  nand (_09320_, _09319_, _06089_);
  nor (_09321_, _06027_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor (_09322_, _06026_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor (_09323_, _09322_, _09321_);
  nand (_09324_, _09323_, _06031_);
  nand (_09325_, _09324_, _09320_);
  nand (_09326_, _09325_, _06020_);
  nand (_09327_, _09326_, _09316_);
  nand (_09328_, _09327_, _06038_);
  nor (_09329_, _06027_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor (_09330_, _06026_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor (_09331_, _09330_, _09329_);
  nand (_09332_, _09331_, _06031_);
  nor (_09333_, _06027_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_09334_, _06026_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_09335_, _09334_, _09333_);
  nand (_09336_, _09335_, _06089_);
  nand (_09337_, _09336_, _09332_);
  nand (_09338_, _09337_, _06021_);
  nor (_09339_, _06027_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_09340_, _06026_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_09341_, _09340_, _09339_);
  nand (_09342_, _09341_, _06089_);
  nor (_09343_, _06027_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_09344_, _06026_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor (_09345_, _09344_, _09343_);
  nand (_09346_, _09345_, _06031_);
  nand (_09347_, _09346_, _09342_);
  nand (_09348_, _09347_, _06020_);
  nand (_09349_, _09348_, _09338_);
  nand (_09350_, _09349_, _06014_);
  nand (_09351_, _09350_, _09328_);
  nand (_09352_, _09351_, _06116_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _09352_, _07668_);
  nor (_09353_, _06027_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_09354_, _06026_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_09355_, _09354_, _09353_);
  nor (_09356_, _09355_, _06089_);
  nor (_09357_, _06027_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_09358_, _06026_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_09359_, _09358_, _09357_);
  nor (_09360_, _09359_, _06031_);
  nor (_09361_, _09360_, _09356_);
  nand (_09362_, _09361_, _06021_);
  nand (_09363_, _06026_, _07965_);
  not (_09364_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nand (_09365_, _06027_, _09364_);
  nand (_09366_, _09365_, _09363_);
  nor (_09367_, _09366_, _06130_);
  not (_09368_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nand (_09369_, _06026_, _09368_);
  not (_09370_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nand (_09371_, _06027_, _09370_);
  nand (_09372_, _09371_, _09369_);
  nor (_09373_, _09372_, _06145_);
  nor (_09374_, _09373_, _09367_);
  nand (_09375_, _09374_, _09362_);
  nand (_09376_, _09375_, _06038_);
  nor (_09377_, _06027_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_09378_, _06026_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_09379_, _09378_, _09377_);
  nand (_09380_, _09379_, _06031_);
  nor (_09381_, _06027_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_09382_, _06026_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_09383_, _09382_, _09381_);
  nand (_09384_, _09383_, _06089_);
  nand (_09385_, _09384_, _09380_);
  nand (_09386_, _09385_, _06021_);
  nor (_09387_, _06027_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_09388_, _06026_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_09389_, _09388_, _09387_);
  nand (_09390_, _09389_, _06089_);
  nor (_09391_, _06027_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_09392_, _06026_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_09393_, _09392_, _09391_);
  nand (_09394_, _09393_, _06031_);
  nand (_09395_, _09394_, _09390_);
  nand (_09396_, _09395_, _06020_);
  nand (_09397_, _09396_, _09386_);
  nand (_09398_, _09397_, _06014_);
  nand (_09399_, _09398_, _09376_);
  nand (_09400_, _09399_, _06116_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _09400_, _07684_);
  nand (_09401_, _06115_, word_in[2]);
  nor (_09402_, _06027_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_09403_, _06026_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_09404_, _09403_, _09402_);
  nor (_09405_, _09404_, _06031_);
  nor (_09406_, _06027_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_09407_, _06026_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_09408_, _09407_, _09406_);
  nor (_09409_, _09408_, _06089_);
  nor (_09410_, _09409_, _09405_);
  nand (_09411_, _09410_, _06021_);
  not (_09413_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand (_09414_, _06026_, _09413_);
  not (_09415_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand (_09416_, _06027_, _09415_);
  nand (_09417_, _09416_, _09414_);
  nor (_09418_, _09417_, _06130_);
  not (_09419_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nand (_09420_, _06026_, _09419_);
  nand (_09421_, _06027_, _08101_);
  nand (_09422_, _09421_, _09420_);
  nor (_09423_, _09422_, _06145_);
  nor (_09424_, _09423_, _09418_);
  nand (_09425_, _09424_, _09411_);
  nand (_09426_, _09425_, _06038_);
  nor (_09427_, _06027_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_09428_, _06026_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_09429_, _09428_, _09427_);
  nor (_09430_, _09429_, _06031_);
  nor (_09431_, _06027_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_09432_, _06026_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_09433_, _09432_, _09431_);
  nor (_09434_, _09433_, _06089_);
  nor (_09435_, _09434_, _09430_);
  nand (_09436_, _09435_, _06021_);
  nor (_09437_, _06027_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_09438_, _06026_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_09439_, _09438_, _09437_);
  nand (_09440_, _09439_, _06089_);
  nor (_09441_, _06027_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_09442_, _06026_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_09443_, _09442_, _09441_);
  nand (_09444_, _09443_, _06031_);
  nand (_09445_, _09444_, _09440_);
  nand (_09446_, _09445_, _06020_);
  nand (_09447_, _09446_, _09436_);
  nand (_09448_, _09447_, _06014_);
  nand (_09449_, _09448_, _09426_);
  nand (_09450_, _09449_, _06116_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _09450_, _09401_);
  nand (_09451_, _06115_, word_in[3]);
  nor (_09452_, _06027_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_09453_, _06026_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_09454_, _09453_, _09452_);
  nor (_09455_, _09454_, _06031_);
  nor (_09456_, _06027_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_09457_, _06026_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_09458_, _09457_, _09456_);
  nor (_09459_, _09458_, _06089_);
  nor (_09460_, _09459_, _09455_);
  nand (_09461_, _09460_, _06021_);
  not (_09462_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nand (_09463_, _06026_, _09462_);
  nand (_09464_, _06027_, _07859_);
  nand (_09465_, _09464_, _09463_);
  nor (_09466_, _09465_, _06130_);
  not (_09467_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nand (_09468_, _06026_, _09467_);
  not (_09469_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nand (_09470_, _06027_, _09469_);
  nand (_09471_, _09470_, _09468_);
  nor (_09472_, _09471_, _06145_);
  nor (_09473_, _09472_, _09466_);
  nand (_09474_, _09473_, _09461_);
  nand (_09475_, _09474_, _06038_);
  nor (_09476_, _06027_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_09477_, _06026_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_09478_, _09477_, _09476_);
  nor (_09479_, _09478_, _06031_);
  nor (_09480_, _06027_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_09481_, _06026_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_09482_, _09481_, _09480_);
  nor (_09483_, _09482_, _06089_);
  nor (_09484_, _09483_, _09479_);
  nand (_09485_, _09484_, _06021_);
  nor (_09486_, _06027_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_09487_, _06026_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_09488_, _09487_, _09486_);
  nand (_09489_, _09488_, _06089_);
  nor (_09490_, _06027_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_09491_, _06026_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_09492_, _09491_, _09490_);
  nand (_09493_, _09492_, _06031_);
  nand (_09494_, _09493_, _09489_);
  nand (_09495_, _09494_, _06020_);
  nand (_09496_, _09495_, _09485_);
  nand (_09497_, _09496_, _06014_);
  nand (_09498_, _09497_, _09475_);
  nand (_09499_, _09498_, _06116_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _09499_, _09451_);
  nand (_09500_, _06115_, word_in[4]);
  nor (_09501_, _06027_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_09502_, _06026_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_09503_, _09502_, _09501_);
  nor (_09504_, _09503_, _06031_);
  nor (_09505_, _06027_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_09506_, _06026_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_09507_, _09506_, _09505_);
  nor (_09508_, _09507_, _06089_);
  nor (_09509_, _09508_, _09504_);
  nand (_09510_, _09509_, _06021_);
  nand (_09511_, _06026_, _08005_);
  nand (_09512_, _06027_, _07878_);
  nand (_09513_, _09512_, _09511_);
  nor (_09514_, _09513_, _06130_);
  not (_09515_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nand (_09516_, _06026_, _09515_);
  not (_09517_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nand (_09518_, _06027_, _09517_);
  nand (_09519_, _09518_, _09516_);
  nor (_09520_, _09519_, _06145_);
  nor (_09521_, _09520_, _09514_);
  nand (_09522_, _09521_, _09510_);
  nand (_09523_, _09522_, _06038_);
  nor (_09524_, _06027_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_09525_, _06026_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_09526_, _09525_, _09524_);
  nor (_09527_, _09526_, _06031_);
  nor (_09529_, _06027_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_09530_, _06026_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_09531_, _09530_, _09529_);
  nor (_09532_, _09531_, _06089_);
  nor (_09533_, _09532_, _09527_);
  nand (_09534_, _09533_, _06021_);
  nor (_09535_, _06027_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_09536_, _06026_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_09537_, _09536_, _09535_);
  nand (_09538_, _09537_, _06089_);
  nor (_09539_, _06027_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_09540_, _06026_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_09541_, _09540_, _09539_);
  nand (_09542_, _09541_, _06031_);
  nand (_09543_, _09542_, _09538_);
  nand (_09544_, _09543_, _06020_);
  nand (_09545_, _09544_, _09534_);
  nand (_09546_, _09545_, _06014_);
  nand (_09547_, _09546_, _09523_);
  nand (_09548_, _09547_, _06116_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _09548_, _09500_);
  nor (_09549_, _06027_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_09550_, _06026_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_09551_, _09550_, _09549_);
  nor (_09552_, _09551_, _06031_);
  nor (_09553_, _06027_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_09554_, _06026_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_09555_, _09554_, _09553_);
  nor (_09556_, _09555_, _06089_);
  nor (_09557_, _09556_, _09552_);
  nand (_09558_, _09557_, _06021_);
  nand (_09559_, _06026_, _08020_);
  not (_09560_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nand (_09561_, _06027_, _09560_);
  nand (_09562_, _09561_, _09559_);
  nor (_09563_, _09562_, _06130_);
  not (_09564_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nand (_09565_, _06026_, _09564_);
  not (_09566_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nand (_09567_, _06027_, _09566_);
  nand (_09568_, _09567_, _09565_);
  nor (_09569_, _09568_, _06145_);
  nor (_09570_, _09569_, _09563_);
  nand (_09571_, _09570_, _09558_);
  nand (_09572_, _09571_, _06038_);
  nor (_09573_, _06027_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_09574_, _06026_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_09575_, _09574_, _09573_);
  nor (_09576_, _09575_, _06031_);
  nor (_09577_, _06027_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_09579_, _06026_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_09580_, _09579_, _09577_);
  nor (_09581_, _09580_, _06089_);
  nor (_09582_, _09581_, _09576_);
  nand (_09583_, _09582_, _06021_);
  nor (_09584_, _06027_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_09585_, _06026_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_09586_, _09585_, _09584_);
  nand (_09587_, _09586_, _06089_);
  nor (_09588_, _06027_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_09589_, _06026_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_09590_, _09589_, _09588_);
  nand (_09591_, _09590_, _06031_);
  nand (_09592_, _09591_, _09587_);
  nand (_09593_, _09592_, _06020_);
  nand (_09594_, _09593_, _09583_);
  nand (_09595_, _09594_, _06014_);
  nand (_09596_, _09595_, _09572_);
  nand (_09597_, _09596_, _06116_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _09597_, _07745_);
  nor (_09598_, _06027_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_09599_, _06026_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_09600_, _09599_, _09598_);
  nor (_09601_, _09600_, _06031_);
  nor (_09602_, _06027_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_09603_, _06026_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_09604_, _09603_, _09602_);
  nor (_09605_, _09604_, _06089_);
  nor (_09606_, _09605_, _09601_);
  nand (_09607_, _09606_, _06021_);
  not (_09608_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nand (_09609_, _06026_, _09608_);
  not (_09610_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nand (_09611_, _06027_, _09610_);
  nand (_09612_, _09611_, _09609_);
  nor (_09613_, _09612_, _06130_);
  not (_09614_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nand (_09615_, _06026_, _09614_);
  nand (_09616_, _06027_, _08149_);
  nand (_09617_, _09616_, _09615_);
  nor (_09618_, _09617_, _06145_);
  nor (_09619_, _09618_, _09613_);
  nand (_09620_, _09619_, _09607_);
  nand (_09621_, _09620_, _06038_);
  nor (_09622_, _06027_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_09623_, _06026_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_09624_, _09623_, _09622_);
  nor (_09625_, _09624_, _06031_);
  nor (_09626_, _06027_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_09627_, _06026_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_09628_, _09627_, _09626_);
  nor (_09629_, _09628_, _06089_);
  nor (_09630_, _09629_, _09625_);
  nand (_09631_, _09630_, _06021_);
  nor (_09632_, _06027_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_09633_, _06026_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_09634_, _09633_, _09632_);
  nand (_09635_, _09634_, _06089_);
  nor (_09636_, _06027_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_09637_, _06026_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_09638_, _09637_, _09636_);
  nand (_09639_, _09638_, _06031_);
  nand (_09640_, _09639_, _09635_);
  nand (_09641_, _09640_, _06020_);
  nand (_09642_, _09641_, _09631_);
  nand (_09643_, _09642_, _06014_);
  nand (_09644_, _09643_, _09621_);
  nand (_09645_, _09644_, _06116_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _09645_, _07759_);
  nor (_09646_, _06027_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nor (_09647_, _06026_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nor (_09648_, _09647_, _09646_);
  nand (_09649_, _09648_, _06287_);
  nor (_09650_, _06027_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_09651_, _06026_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_09652_, _09651_, _09650_);
  nand (_09653_, _09652_, _06280_);
  nand (_09654_, _09653_, _09649_);
  nor (_09655_, _09654_, _06200_);
  nor (_09656_, _06027_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor (_09657_, _06026_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_09658_, _09657_, _09656_);
  nand (_09659_, _09658_, _06287_);
  nor (_09660_, _06027_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_09661_, _06026_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_09662_, _09661_, _09660_);
  nand (_09663_, _09662_, _06280_);
  nand (_09664_, _09663_, _09659_);
  nor (_09665_, _09664_, _06209_);
  nor (_09666_, _09665_, _09655_);
  nand (_09667_, _09666_, _06197_);
  nor (_09668_, _06027_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  nor (_09669_, _06026_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor (_09670_, _09669_, _09668_);
  nand (_09671_, _09670_, _06287_);
  nor (_09672_, _06027_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_09673_, _06026_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_09674_, _09673_, _09672_);
  nand (_09675_, _09674_, _06280_);
  nand (_09676_, _09675_, _09671_);
  nand (_09677_, _09676_, _06209_);
  nor (_09678_, _06027_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor (_09679_, _06026_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor (_09680_, _09679_, _09678_);
  nand (_09681_, _09680_, _06287_);
  nor (_09682_, _06027_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_09683_, _06026_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_09684_, _09683_, _09682_);
  nand (_09685_, _09684_, _06280_);
  nand (_09686_, _09685_, _09681_);
  nand (_09687_, _09686_, _06200_);
  nand (_09688_, _09687_, _09677_);
  nand (_09689_, _09688_, _06196_);
  nand (_09690_, _09689_, _09667_);
  nand (_09691_, _09690_, _06278_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _09691_, _08863_);
  nor (_09692_, _06027_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_09693_, _06026_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_09694_, _09693_, _09692_);
  nand (_09695_, _09694_, _06287_);
  nor (_09696_, _06027_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_09697_, _06026_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_09698_, _09697_, _09696_);
  nand (_09699_, _09698_, _06280_);
  nand (_09700_, _09699_, _09695_);
  nor (_09701_, _09700_, _06209_);
  nor (_09702_, _06027_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_09703_, _06026_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_09704_, _09703_, _09702_);
  nand (_09705_, _09704_, _06287_);
  nor (_09706_, _06027_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_09707_, _06026_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_09708_, _09707_, _09706_);
  nand (_09709_, _09708_, _06280_);
  nand (_09710_, _09709_, _09705_);
  nor (_09711_, _09710_, _06200_);
  nor (_09712_, _09711_, _09701_);
  nand (_09713_, _09712_, _06197_);
  nor (_09714_, _06027_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_09715_, _06026_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_09716_, _09715_, _09714_);
  nand (_09717_, _09716_, _06287_);
  nor (_09718_, _06027_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_09719_, _06026_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_09720_, _09719_, _09718_);
  nand (_09721_, _09720_, _06280_);
  nand (_09722_, _09721_, _09717_);
  nand (_09723_, _09722_, _06209_);
  nor (_09724_, _06027_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_09725_, _06026_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_09727_, _09725_, _09724_);
  nand (_09728_, _09727_, _06287_);
  nor (_09729_, _06027_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_09730_, _06026_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_09731_, _09730_, _09729_);
  nand (_09732_, _09731_, _06280_);
  nand (_09733_, _09732_, _09728_);
  nand (_09734_, _09733_, _06200_);
  nand (_09735_, _09734_, _09723_);
  nand (_09736_, _09735_, _06196_);
  nand (_09737_, _09736_, _09713_);
  nand (_09738_, _09737_, _06278_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _09738_, _07291_);
  nor (_09739_, _06027_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_09740_, _06026_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_09741_, _09740_, _09739_);
  nand (_09742_, _09741_, _06287_);
  nor (_09743_, _06027_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_09744_, _06026_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_09745_, _09744_, _09743_);
  nand (_09746_, _09745_, _06280_);
  nand (_09747_, _09746_, _09742_);
  nor (_09748_, _09747_, _06209_);
  nor (_09749_, _06027_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_09750_, _06026_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_09751_, _09750_, _09749_);
  nand (_09752_, _09751_, _06287_);
  nor (_09753_, _06027_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_09754_, _06026_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_09755_, _09754_, _09753_);
  nand (_09756_, _09755_, _06280_);
  nand (_09757_, _09756_, _09752_);
  nor (_09758_, _09757_, _06200_);
  nor (_09759_, _09758_, _09748_);
  nand (_09760_, _09759_, _06197_);
  nor (_09761_, _06027_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_09762_, _06026_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_09763_, _09762_, _09761_);
  nand (_09764_, _09763_, _06287_);
  nor (_09765_, _06027_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_09766_, _06026_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_09767_, _09766_, _09765_);
  nand (_09768_, _09767_, _06280_);
  nand (_09769_, _09768_, _09764_);
  nand (_09770_, _09769_, _06209_);
  nor (_09771_, _06027_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_09772_, _06026_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_09773_, _09772_, _09771_);
  nand (_09774_, _09773_, _06287_);
  nor (_09775_, _06027_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_09776_, _06026_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_09777_, _09776_, _09775_);
  nand (_09778_, _09777_, _06280_);
  nand (_09779_, _09778_, _09774_);
  nand (_09780_, _09779_, _06200_);
  nand (_09781_, _09780_, _09770_);
  nand (_09782_, _09781_, _06196_);
  nand (_09783_, _09782_, _09760_);
  nand (_09784_, _09783_, _06278_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _09784_, _08902_);
  nor (_09785_, _06027_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_09786_, _06026_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_09787_, _09786_, _09785_);
  nand (_09788_, _09787_, _06287_);
  nor (_09789_, _06027_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_09790_, _06026_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_09791_, _09790_, _09789_);
  nand (_09792_, _09791_, _06280_);
  nand (_09793_, _09792_, _09788_);
  nor (_09794_, _09793_, _06209_);
  nor (_09795_, _06027_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_09796_, _06026_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_09797_, _09796_, _09795_);
  nand (_09798_, _09797_, _06287_);
  nor (_09799_, _06027_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_09800_, _06026_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_09801_, _09800_, _09799_);
  nand (_09802_, _09801_, _06280_);
  nand (_09803_, _09802_, _09798_);
  nor (_09804_, _09803_, _06200_);
  nor (_09805_, _09804_, _09794_);
  nand (_09806_, _09805_, _06197_);
  nor (_09807_, _06027_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_09808_, _06026_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_09809_, _09808_, _09807_);
  nand (_09810_, _09809_, _06287_);
  nor (_09811_, _06027_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_09812_, _06026_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_09813_, _09812_, _09811_);
  nand (_09814_, _09813_, _06280_);
  nand (_09815_, _09814_, _09810_);
  nand (_09816_, _09815_, _06209_);
  nor (_09817_, _06027_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_09818_, _06026_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_09819_, _09818_, _09817_);
  nand (_09820_, _09819_, _06287_);
  nor (_09821_, _06027_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_09822_, _06026_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_09823_, _09822_, _09821_);
  nand (_09824_, _09823_, _06280_);
  nand (_09825_, _09824_, _09820_);
  nand (_09826_, _09825_, _06200_);
  nand (_09827_, _09826_, _09816_);
  nand (_09828_, _09827_, _06196_);
  nand (_09829_, _09828_, _09806_);
  nand (_09830_, _09829_, _06278_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _09830_, _08917_);
  nor (_09831_, _06027_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_09832_, _06026_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_09833_, _09832_, _09831_);
  nand (_09834_, _09833_, _06287_);
  nor (_09835_, _06027_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_09836_, _06026_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_09837_, _09836_, _09835_);
  nand (_09838_, _09837_, _06280_);
  nand (_09839_, _09838_, _09834_);
  nor (_09840_, _09839_, _06200_);
  nor (_09841_, _06027_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_09842_, _06026_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_09843_, _09842_, _09841_);
  nand (_09844_, _09843_, _06287_);
  nor (_09845_, _06027_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_09846_, _06026_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_09847_, _09846_, _09845_);
  nand (_09848_, _09847_, _06280_);
  nand (_09849_, _09848_, _09844_);
  nor (_09850_, _09849_, _06209_);
  nor (_09851_, _09850_, _09840_);
  nand (_09852_, _09851_, _06197_);
  nor (_09853_, _06027_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_09854_, _06026_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_09855_, _09854_, _09853_);
  nand (_09856_, _09855_, _06287_);
  nor (_09857_, _06027_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_09858_, _06026_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_09859_, _09858_, _09857_);
  nand (_09860_, _09859_, _06280_);
  nand (_09861_, _09860_, _09856_);
  nand (_09862_, _09861_, _06209_);
  nor (_09863_, _06027_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_09864_, _06026_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_09865_, _09864_, _09863_);
  nand (_09866_, _09865_, _06287_);
  nor (_09867_, _06027_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_09868_, _06026_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_09869_, _09868_, _09867_);
  nand (_09870_, _09869_, _06280_);
  nand (_09871_, _09870_, _09866_);
  nand (_09872_, _09871_, _06200_);
  nand (_09873_, _09872_, _09862_);
  nand (_09874_, _09873_, _06196_);
  nand (_09875_, _09874_, _09852_);
  nand (_09876_, _09875_, _06278_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _09876_, _08936_);
  nor (_09877_, _06027_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_09878_, _06026_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_09879_, _09878_, _09877_);
  nand (_09880_, _09879_, _06287_);
  nor (_09881_, _06027_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_09882_, _06026_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_09883_, _09882_, _09881_);
  nand (_09884_, _09883_, _06280_);
  nand (_09885_, _09884_, _09880_);
  nor (_09886_, _09885_, _06209_);
  nor (_09887_, _06027_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_09888_, _06026_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_09889_, _09888_, _09887_);
  nand (_09890_, _09889_, _06287_);
  nor (_09891_, _06027_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_09892_, _06026_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_09893_, _09892_, _09891_);
  nand (_09894_, _09893_, _06280_);
  nand (_09895_, _09894_, _09890_);
  nor (_09896_, _09895_, _06200_);
  nor (_09897_, _09896_, _09886_);
  nand (_09898_, _09897_, _06197_);
  nor (_09899_, _06027_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_09900_, _06026_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_09901_, _09900_, _09899_);
  nand (_09902_, _09901_, _06287_);
  nor (_09903_, _06027_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_09904_, _06026_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_09905_, _09904_, _09903_);
  nand (_09906_, _09905_, _06280_);
  nand (_09907_, _09906_, _09902_);
  nand (_09908_, _09907_, _06209_);
  nor (_09909_, _06027_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_09910_, _06026_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_09911_, _09910_, _09909_);
  nand (_09912_, _09911_, _06287_);
  nor (_09913_, _06027_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_09914_, _06026_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_09915_, _09914_, _09913_);
  nand (_09916_, _09915_, _06280_);
  nand (_09917_, _09916_, _09912_);
  nand (_09918_, _09917_, _06200_);
  nand (_09919_, _09918_, _09908_);
  nand (_09920_, _09919_, _06196_);
  nand (_09921_, _09920_, _09898_);
  nand (_09922_, _09921_, _06278_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _09922_, _08955_);
  nor (_09924_, _06027_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_09925_, _06026_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_09926_, _09925_, _09924_);
  nand (_09927_, _09926_, _06287_);
  nor (_09928_, _06027_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_09929_, _06026_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_09930_, _09929_, _09928_);
  nand (_09931_, _09930_, _06280_);
  nand (_09932_, _09931_, _09927_);
  nor (_09933_, _09932_, _06209_);
  nor (_09934_, _06027_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_09935_, _06026_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_09936_, _09935_, _09934_);
  nand (_09937_, _09936_, _06287_);
  nor (_09938_, _06027_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_09939_, _06026_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_09940_, _09939_, _09938_);
  nand (_09941_, _09940_, _06280_);
  nand (_09942_, _09941_, _09937_);
  nor (_09943_, _09942_, _06200_);
  nor (_09944_, _09943_, _09933_);
  nand (_09945_, _09944_, _06197_);
  nor (_09946_, _06027_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_09947_, _06026_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_09948_, _09947_, _09946_);
  nand (_09949_, _09948_, _06287_);
  nor (_09950_, _06027_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_09951_, _06026_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_09952_, _09951_, _09950_);
  nand (_09953_, _09952_, _06280_);
  nand (_09954_, _09953_, _09949_);
  nand (_09955_, _09954_, _06209_);
  nor (_09956_, _06027_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_09957_, _06026_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_09958_, _09957_, _09956_);
  nand (_09959_, _09958_, _06287_);
  nor (_09960_, _06027_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_09961_, _06026_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_09962_, _09961_, _09960_);
  nand (_09963_, _09962_, _06280_);
  nand (_09964_, _09963_, _09959_);
  nand (_09965_, _09964_, _06200_);
  nand (_09966_, _09965_, _09955_);
  nand (_09967_, _09966_, _06196_);
  nand (_09968_, _09967_, _09945_);
  nand (_09969_, _09968_, _06278_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _09969_, _08974_);
  nor (_09970_, _09331_, _06031_);
  nor (_09971_, _09335_, _06089_);
  nor (_09972_, _09971_, _09970_);
  nand (_09973_, _09972_, _06347_);
  nand (_09974_, _09341_, _06031_);
  nand (_09975_, _09345_, _06089_);
  nand (_09976_, _09975_, _09974_);
  nand (_09977_, _09976_, _06352_);
  nand (_09978_, _09977_, _09973_);
  nand (_09979_, _09978_, _06344_);
  nor (_09980_, _09309_, _06031_);
  nor (_09981_, _09313_, _06089_);
  nor (_09982_, _09981_, _09980_);
  nand (_09983_, _09982_, _06347_);
  nand (_09984_, _09319_, _06031_);
  nand (_09985_, _09323_, _06089_);
  nand (_09986_, _09985_, _09984_);
  nand (_09987_, _09986_, _06352_);
  nand (_09988_, _09987_, _09983_);
  nand (_09989_, _09988_, _06343_);
  nand (_09990_, _09989_, _09979_);
  nand (_09991_, _09990_, _06413_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _09991_, _07793_);
  nor (_09992_, _09379_, _06031_);
  nor (_09993_, _09383_, _06089_);
  nor (_09994_, _09993_, _09992_);
  nand (_09995_, _09994_, _06347_);
  nand (_09996_, _09389_, _06031_);
  nand (_09997_, _09393_, _06089_);
  nand (_09998_, _09997_, _09996_);
  nand (_09999_, _09998_, _06352_);
  nand (_10000_, _09999_, _09995_);
  nand (_10001_, _10000_, _06344_);
  nor (_10002_, _09355_, _06031_);
  nor (_10003_, _09359_, _06089_);
  nor (_10004_, _10003_, _10002_);
  nand (_10005_, _10004_, _06347_);
  nor (_10006_, _09366_, _06419_);
  nor (_10007_, _09372_, _06130_);
  nor (_10008_, _10007_, _10006_);
  nand (_10009_, _10008_, _10005_);
  nand (_10010_, _10009_, _06343_);
  nand (_10011_, _10010_, _10001_);
  nand (_10012_, _10011_, _06413_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _10012_, _07816_);
  nor (_10013_, _09433_, _06031_);
  nor (_10014_, _09429_, _06089_);
  nor (_10015_, _10014_, _10013_);
  nand (_10016_, _10015_, _06347_);
  nand (_10017_, _09439_, _06031_);
  nand (_10018_, _09443_, _06089_);
  nand (_10019_, _10018_, _10017_);
  nand (_10020_, _10019_, _06352_);
  nand (_10021_, _10020_, _10016_);
  nand (_10022_, _10021_, _06344_);
  nor (_10023_, _09408_, _06031_);
  nor (_10024_, _09404_, _06089_);
  nor (_10025_, _10024_, _10023_);
  nand (_10026_, _10025_, _06347_);
  nor (_10027_, _09422_, _06130_);
  nor (_10028_, _09417_, _06419_);
  nor (_10029_, _10028_, _10027_);
  nand (_10030_, _10029_, _10026_);
  nand (_10031_, _10030_, _06343_);
  nand (_10032_, _10031_, _10022_);
  nand (_10033_, _10032_, _06413_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _10033_, _07846_);
  nor (_10034_, _09482_, _06031_);
  nor (_10035_, _09478_, _06089_);
  nor (_10036_, _10035_, _10034_);
  nand (_10037_, _10036_, _06347_);
  nand (_10038_, _09488_, _06031_);
  nand (_10039_, _09492_, _06089_);
  nand (_10040_, _10039_, _10038_);
  nand (_10041_, _10040_, _06352_);
  nand (_10042_, _10041_, _10037_);
  nand (_10043_, _10042_, _06344_);
  nor (_10044_, _09458_, _06031_);
  nor (_10045_, _09454_, _06089_);
  nor (_10046_, _10045_, _10044_);
  nand (_10047_, _10046_, _06347_);
  nor (_10048_, _09471_, _06130_);
  nor (_10049_, _09465_, _06419_);
  nor (_10050_, _10049_, _10048_);
  nand (_10051_, _10050_, _10047_);
  nand (_10052_, _10051_, _06343_);
  nand (_10053_, _10052_, _10043_);
  nand (_10054_, _10053_, _06413_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _10054_, _07868_);
  nand (_10055_, _09526_, _06031_);
  nand (_10056_, _09531_, _06089_);
  nand (_10057_, _10056_, _10055_);
  nand (_10058_, _10057_, _06347_);
  nand (_10059_, _09537_, _06031_);
  nand (_10060_, _09541_, _06089_);
  nand (_10061_, _10060_, _10059_);
  nand (_10062_, _10061_, _06352_);
  nand (_10063_, _10062_, _10058_);
  nand (_10064_, _10063_, _06344_);
  nor (_10065_, _09507_, _06031_);
  nor (_10066_, _09503_, _06089_);
  nor (_10067_, _10066_, _10065_);
  nand (_10068_, _10067_, _06347_);
  nor (_10069_, _09519_, _06130_);
  nor (_10070_, _09513_, _06419_);
  nor (_10071_, _10070_, _10069_);
  nand (_10072_, _10071_, _10068_);
  nand (_10073_, _10072_, _06343_);
  nand (_10074_, _10073_, _10064_);
  nand (_10075_, _10074_, _06413_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _10075_, _07885_);
  nand (_10076_, _09575_, _06031_);
  nand (_10077_, _09580_, _06089_);
  nand (_10078_, _10077_, _10076_);
  nand (_10079_, _10078_, _06347_);
  not (_10080_, _09586_);
  nor (_10081_, _10080_, _06419_);
  not (_10082_, _09590_);
  nor (_10083_, _10082_, _06130_);
  nor (_10084_, _10083_, _10081_);
  nand (_10085_, _10084_, _10079_);
  nand (_10086_, _10085_, _06344_);
  nor (_10087_, _09555_, _06031_);
  nor (_10088_, _09551_, _06089_);
  nor (_10089_, _10088_, _10087_);
  nand (_10090_, _10089_, _06347_);
  nor (_10091_, _09568_, _06130_);
  nor (_10092_, _09562_, _06419_);
  nor (_10093_, _10092_, _10091_);
  nand (_10094_, _10093_, _10090_);
  nand (_10095_, _10094_, _06343_);
  nand (_10096_, _10095_, _10086_);
  nand (_10097_, _10096_, _06413_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _10097_, _07894_);
  nor (_10098_, _09628_, _06031_);
  nor (_10099_, _09624_, _06089_);
  nor (_10100_, _10099_, _10098_);
  nand (_10101_, _10100_, _06347_);
  nand (_10102_, _09634_, _06031_);
  nand (_10103_, _09638_, _06089_);
  nand (_10104_, _10103_, _10102_);
  nand (_10105_, _10104_, _06352_);
  nand (_10106_, _10105_, _10101_);
  nand (_10107_, _10106_, _06344_);
  nor (_10108_, _09604_, _06031_);
  nor (_10109_, _09600_, _06089_);
  nor (_10110_, _10109_, _10108_);
  nand (_10111_, _10110_, _06347_);
  nor (_10112_, _09617_, _06130_);
  nor (_10113_, _09612_, _06419_);
  nor (_10114_, _10113_, _10112_);
  nand (_10115_, _10114_, _10111_);
  nand (_10117_, _10115_, _06343_);
  nand (_10118_, _10117_, _10107_);
  nand (_10119_, _10118_, _06413_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _10119_, _07910_);
  nand (_10120_, _09658_, _06280_);
  nand (_10121_, _09662_, _06287_);
  nand (_10122_, _10121_, _10120_);
  nand (_10123_, _10122_, _06444_);
  nand (_10124_, _09652_, _06287_);
  nand (_10125_, _09648_, _06280_);
  nand (_10126_, _10125_, _10124_);
  nand (_10127_, _10126_, _06445_);
  nand (_10128_, _10127_, _10123_);
  nand (_10129_, _10128_, _06449_);
  nand (_10130_, _09680_, _06280_);
  nand (_10131_, _09684_, _06287_);
  nand (_10132_, _10131_, _10130_);
  nand (_10133_, _10132_, _06444_);
  nand (_10134_, _09670_, _06280_);
  nand (_10135_, _09674_, _06287_);
  nand (_10136_, _10135_, _10134_);
  nand (_10137_, _10136_, _06445_);
  nand (_10138_, _10137_, _10133_);
  nand (_10139_, _10138_, _06451_);
  nand (_10140_, _10139_, _10129_);
  nand (_10141_, _10140_, _06514_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _10141_, _07813_);
  nand (_10142_, _09694_, _06280_);
  nand (_10143_, _09698_, _06287_);
  nand (_10144_, _10143_, _10142_);
  nand (_10145_, _10144_, _06444_);
  nand (_10146_, _09704_, _06280_);
  nand (_10147_, _09708_, _06287_);
  nand (_10148_, _10147_, _10146_);
  nand (_10149_, _10148_, _06445_);
  nand (_10150_, _10149_, _10145_);
  nand (_10151_, _10150_, _06449_);
  nand (_10152_, _09727_, _06280_);
  nand (_10153_, _09731_, _06287_);
  nand (_10154_, _10153_, _10152_);
  nand (_10155_, _10154_, _06444_);
  nand (_10156_, _09720_, _06287_);
  nand (_10157_, _09716_, _06280_);
  nand (_10158_, _10157_, _10156_);
  nand (_10159_, _10158_, _06445_);
  nand (_10160_, _10159_, _10155_);
  nand (_10161_, _10160_, _06451_);
  nand (_10162_, _10161_, _10151_);
  nand (_10163_, _10162_, _06514_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _10163_, _07832_);
  nand (_10164_, _09741_, _06280_);
  nand (_10165_, _09745_, _06287_);
  nand (_10166_, _10165_, _10164_);
  nand (_10167_, _10166_, _06444_);
  nand (_10168_, _09755_, _06287_);
  nand (_10169_, _09751_, _06280_);
  nand (_10170_, _10169_, _10168_);
  nand (_10171_, _10170_, _06445_);
  nand (_10172_, _10171_, _10167_);
  nand (_10173_, _10172_, _06449_);
  nand (_10174_, _09773_, _06280_);
  nand (_10175_, _09777_, _06287_);
  nand (_10176_, _10175_, _10174_);
  nand (_10177_, _10176_, _06444_);
  nand (_10178_, _09763_, _06280_);
  nand (_10179_, _09767_, _06287_);
  nand (_10180_, _10179_, _10178_);
  nand (_10181_, _10180_, _06445_);
  nand (_10182_, _10181_, _10177_);
  nand (_10183_, _10182_, _06451_);
  nand (_10184_, _10183_, _10173_);
  nand (_10185_, _10184_, _06514_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _10185_, _07855_);
  nand (_10186_, _09787_, _06280_);
  nand (_10187_, _09791_, _06287_);
  nand (_10188_, _10187_, _10186_);
  nand (_10189_, _10188_, _06444_);
  nand (_10190_, _09801_, _06287_);
  nand (_10191_, _09797_, _06280_);
  nand (_10192_, _10191_, _10190_);
  nand (_10193_, _10192_, _06445_);
  nand (_10194_, _10193_, _10189_);
  nand (_10195_, _10194_, _06449_);
  nand (_10196_, _09819_, _06280_);
  nand (_10197_, _09823_, _06287_);
  nand (_10198_, _10197_, _10196_);
  nand (_10199_, _10198_, _06444_);
  nand (_10200_, _09813_, _06287_);
  nand (_10201_, _09809_, _06280_);
  nand (_10202_, _10201_, _10200_);
  nand (_10203_, _10202_, _06445_);
  nand (_10204_, _10203_, _10199_);
  nand (_10205_, _10204_, _06451_);
  nand (_10206_, _10205_, _10195_);
  nand (_10207_, _10206_, _06514_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _10207_, _07873_);
  nand (_10208_, _09843_, _06280_);
  nand (_10209_, _09847_, _06287_);
  nand (_10210_, _10209_, _10208_);
  nand (_10211_, _10210_, _06444_);
  nand (_10212_, _09837_, _06287_);
  nand (_10213_, _09833_, _06280_);
  nand (_10214_, _10213_, _10212_);
  nand (_10215_, _10214_, _06445_);
  nand (_10216_, _10215_, _10211_);
  nand (_10217_, _10216_, _06449_);
  nand (_10218_, _09865_, _06280_);
  nand (_10219_, _09869_, _06287_);
  nand (_10220_, _10219_, _10218_);
  nand (_10221_, _10220_, _06444_);
  nand (_10222_, _09859_, _06287_);
  nand (_10223_, _09855_, _06280_);
  nand (_10224_, _10223_, _10222_);
  nand (_10225_, _10224_, _06445_);
  nand (_10226_, _10225_, _10221_);
  nand (_10227_, _10226_, _06451_);
  nand (_10228_, _10227_, _10217_);
  nand (_10229_, _10228_, _06514_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _10229_, _07891_);
  nand (_10230_, _09879_, _06280_);
  nand (_10231_, _09883_, _06287_);
  nand (_10232_, _10231_, _10230_);
  nand (_10233_, _10232_, _06444_);
  nand (_10234_, _09893_, _06287_);
  nand (_10235_, _09889_, _06280_);
  nand (_10236_, _10235_, _10234_);
  nand (_10237_, _10236_, _06445_);
  nand (_10238_, _10237_, _10233_);
  nand (_10239_, _10238_, _06449_);
  nand (_10240_, _09911_, _06280_);
  nand (_10242_, _09915_, _06287_);
  nand (_10243_, _10242_, _10240_);
  nand (_10244_, _10243_, _06444_);
  nand (_10245_, _09905_, _06287_);
  nand (_10246_, _09901_, _06280_);
  nand (_10247_, _10246_, _10245_);
  nand (_10248_, _10247_, _06445_);
  nand (_10249_, _10248_, _10244_);
  nand (_10250_, _10249_, _06451_);
  nand (_10251_, _10250_, _10239_);
  nand (_10252_, _10251_, _06514_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _10252_, _07907_);
  nand (_10253_, _09926_, _06280_);
  nand (_10254_, _09930_, _06287_);
  nand (_10255_, _10254_, _10253_);
  nand (_10256_, _10255_, _06444_);
  nand (_10257_, _09940_, _06287_);
  nand (_10258_, _09936_, _06280_);
  nand (_10259_, _10258_, _10257_);
  nand (_10260_, _10259_, _06445_);
  nand (_10261_, _10260_, _10256_);
  nand (_10262_, _10261_, _06449_);
  nand (_10263_, _09958_, _06280_);
  nand (_10264_, _09962_, _06287_);
  nand (_10265_, _10264_, _10263_);
  nand (_10266_, _10265_, _06444_);
  nand (_10267_, _09952_, _06287_);
  nand (_10268_, _09948_, _06280_);
  nand (_10269_, _10268_, _10267_);
  nand (_10270_, _10269_, _06445_);
  nand (_10271_, _10270_, _10266_);
  nand (_10272_, _10271_, _06451_);
  nand (_10273_, _10272_, _10262_);
  nand (_10274_, _10273_, _06514_);
  nand (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _10274_, _07925_);
  nor (_10275_, _23545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  nor (_10276_, _23547_, _21554_);
  nor (_01332_, _10276_, _10275_);
  nor (_10277_, _22454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  nor (_10278_, _22456_, _21414_);
  nor (_01339_, _10278_, _10277_);
  nor (_10279_, _21777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1]);
  nor (_10280_, _21779_, _21474_);
  nor (_01343_, _10280_, _10279_);
  nor (_10281_, _21777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  nor (_10282_, _21779_, _21586_);
  nor (_01349_, _10282_, _10281_);
  nor (_10283_, _24043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7]);
  nor (_10284_, _24045_, _21626_);
  nor (_25362_, _10284_, _10283_);
  nor (_10285_, _24043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  nor (_10286_, _24045_, _21504_);
  nor (_25361_, _10286_, _10285_);
  nor (_10287_, _07226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  nor (_10288_, _07228_, _21414_);
  nor (_01440_, _10288_, _10287_);
  nor (_10289_, _24043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1]);
  nor (_10290_, _24045_, _21474_);
  nor (_25359_, _10290_, _10289_);
  nor (_10291_, _24043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  nor (_10292_, _24045_, _21586_);
  nor (_01454_, _10292_, _10291_);
  not (_10293_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nand (_10294_, _02379_, _10293_);
  nor (_10295_, _02379_, _10293_);
  nor (_10296_, _10295_, rst);
  nand (_10297_, _10296_, _10294_);
  nor (_01458_, _10297_, _01130_);
  nor (_10298_, _22292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  nor (_10299_, _22294_, _21414_);
  nor (_01472_, _10299_, _10298_);
  nor (_10300_, _22292_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  nor (_10301_, _22294_, _21554_);
  nor (_01474_, _10301_, _10300_);
  nor (_10302_, _24043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  nor (_10303_, _24045_, _21526_);
  nor (_01497_, _10303_, _10302_);
  nor (_10304_, _24043_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  nor (_10305_, _24045_, _21554_);
  nor (_01507_, _10305_, _10304_);
  nor (_10306_, _07226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  nor (_10307_, _07228_, _21526_);
  nor (_01512_, _10307_, _10306_);
  nor (_10308_, _07226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  nor (_10309_, _07228_, _21554_);
  nor (_25299_, _10309_, _10308_);
  nor (_10310_, _23829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5]);
  nor (_10311_, _23831_, _21451_);
  nor (_01542_, _10311_, _10310_);
  nor (_10312_, _21653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  nor (_10313_, _21655_, _21504_);
  nor (_01567_, _10313_, _10312_);
  nor (_10314_, _22259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  nor (_10315_, _22261_, _21554_);
  nor (_01569_, _10315_, _10314_);
  nor (_10316_, _23829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  nor (_10317_, _23831_, _21504_);
  nor (_01572_, _10317_, _10316_);
  nor (_10318_, _22259_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  nor (_10319_, _22261_, _21586_);
  nor (_01579_, _10319_, _10318_);
  nor (_10320_, _23829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1]);
  nor (_10321_, _23831_, _21474_);
  nor (_01595_, _10321_, _10320_);
  nor (_10322_, _23829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  nor (_10323_, _23831_, _21526_);
  nor (_01621_, _10323_, _10322_);
  nor (_10324_, _23829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  nor (_10325_, _23831_, _21554_);
  nor (_01648_, _10325_, _10324_);
  nor (_10327_, _23833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  nor (_10328_, _23835_, _21526_);
  nor (_01673_, _10328_, _10327_);
  nor (_10329_, _23833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  nor (_10330_, _23835_, _21554_);
  nor (_25377_, _10330_, _10329_);
  nor (_10331_, _22521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  nor (_10332_, _22524_, _21586_);
  nor (_01695_, _10332_, _10331_);
  nor (_01701_, rst, \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nor (_10333_, _23833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  nor (_10334_, _23835_, _21414_);
  nor (_25378_, _10334_, _10333_);
  nor (_10335_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7]);
  nor (_10336_, _22302_, _21626_);
  nor (_25167_, _10336_, _10335_);
  nor (_10337_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5]);
  nor (_10338_, _22302_, _21451_);
  nor (_01730_, _10338_, _10337_);
  nor (_10339_, _23833_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  nor (_10340_, _23835_, _21586_);
  nor (_01735_, _10340_, _10339_);
  nor (_10341_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5]);
  nor (_10342_, _22473_, _21451_);
  nor (_01744_, _10342_, _10341_);
  nor (_10343_, \oc8051_top_1.oc8051_sfr1.prescaler [1], \oc8051_top_1.oc8051_sfr1.prescaler [0]);
  nand (_10344_, _05209_, _23493_);
  nor (_01761_, _10344_, _10343_);
  nor (_10345_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1]);
  nor (_10346_, _22302_, _21474_);
  nor (_01772_, _10346_, _10345_);
  nor (_10347_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  nor (_10348_, _22302_, _21586_);
  nor (_01785_, _10348_, _10347_);
  nor (_10349_, _21389_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  nor (_10350_, _21586_, _21391_);
  nor (_01788_, _10350_, _10349_);
  nor (_10351_, _22300_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  nor (_10352_, _22302_, _21526_);
  nor (_25165_, _10352_, _10351_);
  nor (_10353_, _23837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  nor (_10354_, _23839_, _21504_);
  nor (_01835_, _10354_, _10353_);
  nor (_10355_, _23837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5]);
  nor (_10356_, _23839_, _21451_);
  nor (_25375_, _10356_, _10355_);
  nor (_10357_, _23837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  nor (_10358_, _23839_, _21586_);
  nor (_01877_, _10358_, _10357_);
  nor (_10359_, _23837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  nor (_10360_, _23839_, _21554_);
  nor (_01886_, _10360_, _10359_);
  nor (_10361_, _09002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1]);
  nor (_10362_, _09004_, _21474_);
  nor (_01903_, _10362_, _10361_);
  nor (_10363_, _23837_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1]);
  nor (_10364_, _23839_, _21474_);
  nor (_01908_, _10364_, _10363_);
  nor (_10365_, _23992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  nor (_10366_, _23994_, _21586_);
  nor (_01938_, _10366_, _10365_);
  nor (_10368_, _23992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1]);
  nor (_10369_, _23994_, _21474_);
  nor (_01955_, _10369_, _10368_);
  nor (_10370_, _23806_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  nor (_10371_, _23808_, _21504_);
  nor (_01977_, _10371_, _10370_);
  nor (_10372_, _09002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  nor (_10373_, _09004_, _21526_);
  nor (_25298_, _10373_, _10372_);
  nor (_10374_, _23992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  nor (_10375_, _23994_, _21414_);
  nor (_25374_, _10375_, _10374_);
  nor (_10376_, _23992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  nor (_10377_, _23994_, _21526_);
  nor (_02012_, _10377_, _10376_);
  nor (_10378_, _22465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5]);
  nor (_10379_, _22467_, _21451_);
  nor (_25081_, _10379_, _10378_);
  nor (_10380_, _23044_, _21302_);
  not (_10381_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  nor (_10382_, _23153_, _10381_);
  nor (_10383_, _23058_, _23183_);
  nor (_10384_, _23067_, _23185_);
  nor (_10385_, _10384_, _10383_);
  nor (_10386_, _23050_, _00444_);
  nor (_10387_, _23107_, _23188_);
  nor (_10388_, _10387_, _10386_);
  nand (_10389_, _10388_, _10385_);
  nor (_10390_, _23073_, _07082_);
  nor (_10391_, _23076_, _23190_);
  nor (_10392_, _10391_, _10390_);
  not (_10393_, _10392_);
  nor (_10394_, _10393_, _10389_);
  nor (_10395_, _10394_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_10396_, _10395_, _10382_);
  nor (_10397_, _10396_, _23490_);
  nor (_10398_, _10397_, _10380_);
  nor (_02018_, _10398_, rst);
  nor (_10399_, _23992_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  nor (_10400_, _23994_, _21504_);
  nor (_02025_, _10400_, _10399_);
  nor (_10401_, _24343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1]);
  nor (_10402_, _24345_, _21474_);
  nor (_02044_, _10402_, _10401_);
  nor (_10403_, _23025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  nor (_10404_, _23027_, _21526_);
  nor (_02050_, _10404_, _10403_);
  nor (_10405_, _24343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  nor (_10406_, _24345_, _21586_);
  nor (_02052_, _10406_, _10405_);
  nor (_10407_, _24343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  nor (_10408_, _24345_, _21504_);
  nor (_02074_, _10408_, _10407_);
  nor (_10409_, _24325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  nor (_10410_, _24327_, _21526_);
  nor (_02077_, _10410_, _10409_);
  not (_10411_, _05210_);
  nand (_10412_, _05209_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  nand (_10413_, _10412_, _10411_);
  nand (_10414_, _10413_, _05211_);
  nor (_25455_[2], _10414_, rst);
  nor (_10415_, _24325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  nor (_10416_, _24327_, _21414_);
  nor (_02083_, _10416_, _10415_);
  nor (_10417_, _24325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  nor (_10418_, _24327_, _21504_);
  nor (_25435_, _10418_, _10417_);
  nor (_10419_, _24343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5]);
  nor (_10420_, _24345_, _21451_);
  nor (_02090_, _10420_, _10419_);
  nor (_10421_, _23025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  nor (_10422_, _23027_, _21554_);
  nor (_25119_, _10422_, _10421_);
  nor (_10423_, _24343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  nor (_10424_, _24345_, _21414_);
  nor (_02103_, _10424_, _10423_);
  nor (_10425_, _24343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  nor (_10426_, _24345_, _21526_);
  nor (_02109_, _10426_, _10425_);
  nor (_10427_, _24331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  nor (_10428_, _24333_, _21526_);
  nor (_02139_, _10428_, _10427_);
  nor (_10429_, _24331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  nor (_10430_, _24333_, _21554_);
  nor (_02145_, _10430_, _10429_);
  nor (_10431_, _24331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1]);
  nor (_10432_, _24333_, _21474_);
  nor (_02147_, _10432_, _10431_);
  nor (_10433_, _24331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  nor (_10434_, _24333_, _21504_);
  nor (_02166_, _10434_, _10433_);
  nor (_10435_, _24331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5]);
  nor (_10436_, _24333_, _21451_);
  nor (_02170_, _10436_, _10435_);
  nor (_10437_, _24331_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  nor (_10438_, _24333_, _21414_);
  nor (_02179_, _10438_, _10437_);
  nor (_10439_, _24027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  nor (_10440_, _24029_, _21504_);
  nor (_25419_, _10440_, _10439_);
  nor (_10442_, _24325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  nor (_10443_, _24327_, _21554_);
  nor (_02220_, _10443_, _10442_);
  nor (_10444_, _22114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  nor (_10445_, _22116_, _21554_);
  nor (_25437_, _10445_, _10444_);
  nor (_10446_, _24325_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7]);
  nor (_10447_, _24327_, _21626_);
  nor (_02227_, _10447_, _10446_);
  nor (_10448_, _22114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  nor (_10449_, _22116_, _21586_);
  nor (_25436_, _10449_, _10448_);
  nor (_10450_, _21816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7]);
  nor (_10451_, _21818_, _21626_);
  nor (_02243_, _10451_, _10450_);
  nor (_10452_, _22114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  nor (_10453_, _22116_, _21504_);
  nor (_02255_, _10453_, _10452_);
  nor (_10454_, _22114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  nor (_10455_, _22116_, _21526_);
  nor (_02260_, _10455_, _10454_);
  nor (_10456_, _22114_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  nor (_10457_, _22116_, _21414_);
  nor (_02267_, _10457_, _10456_);
  nor (_10458_, _21873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7]);
  nor (_10459_, _21875_, _21626_);
  nor (_02270_, _10459_, _10458_);
  nor (_10460_, _05519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  nor (_10461_, _05521_, _21586_);
  nor (_02273_, _10461_, _10460_);
  nor (_10462_, _05453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7]);
  nor (_10463_, _05455_, _21626_);
  nor (_02277_, _10463_, _10462_);
  nor (_10464_, _21899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5]);
  nor (_10465_, _21902_, _21451_);
  nor (_25124_, _10465_, _10464_);
  nor (_10466_, _21810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  nor (_10467_, _21812_, _21586_);
  nor (_02279_, _10467_, _10466_);
  nor (_10468_, _05453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  nor (_10469_, _05455_, _21554_);
  nor (_02282_, _10469_, _10468_);
  nor (_10470_, _01184_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7]);
  nor (_10471_, _01186_, _21626_);
  nor (_02285_, _10471_, _10470_);
  nor (_10472_, _24027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1]);
  nor (_10473_, _24029_, _21474_);
  nor (_02294_, _10473_, _10472_);
  nor (_10474_, _24027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  nor (_10475_, _24029_, _21586_);
  nor (_02297_, _10475_, _10474_);
  nor (_10476_, _24027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  nor (_10477_, _24029_, _21414_);
  nor (_02329_, _10477_, _10476_);
  nor (_10478_, _24027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  nor (_10479_, _24029_, _21526_);
  nor (_02336_, _10479_, _10478_);
  nor (_10480_, _24027_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  nor (_10481_, _24029_, _21554_);
  nor (_02339_, _10481_, _10480_);
  nor (_10482_, _21600_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  nor (_10483_, _21602_, _21586_);
  nor (_02342_, _10483_, _10482_);
  nor (_10484_, _24365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  nor (_10485_, _24367_, _21526_);
  nor (_02364_, _10485_, _10484_);
  nor (_10486_, _24365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  nor (_10487_, _24367_, _21554_);
  nor (_25417_, _10487_, _10486_);
  nor (_10488_, _24365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1]);
  nor (_10489_, _24367_, _21474_);
  nor (_25416_, _10489_, _10488_);
  nor (_10490_, _24365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  nor (_10491_, _24367_, _21586_);
  nor (_25415_, _10491_, _10490_);
  nor (_10492_, _24365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  nor (_10493_, _24367_, _21504_);
  nor (_02401_, _10493_, _10492_);
  nor (_25016_[2], _24799_, rst);
  nor (_10494_, _24365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5]);
  nor (_10495_, _24367_, _21451_);
  nor (_02406_, _10495_, _10494_);
  nor (_10496_, _24365_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  nor (_10497_, _24367_, _21414_);
  nor (_02409_, _10497_, _10496_);
  nor (_10498_, _09002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  nor (_10499_, _09004_, _21554_);
  nor (_02425_, _10499_, _10498_);
  nor (_10500_, _24343_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7]);
  nor (_10501_, _24345_, _21626_);
  nor (_02428_, _10501_, _10500_);
  nor (_10502_, _23829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  nor (_10503_, _23831_, _21586_);
  nor (_02435_, _10503_, _10502_);
  nor (_10504_, _23843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7]);
  nor (_10505_, _23845_, _21626_);
  nor (_02438_, _10505_, _10504_);
  nor (_10506_, _23843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  nor (_10507_, _23845_, _21504_);
  nor (_02441_, _10507_, _10506_);
  nor (_10508_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  nor (_10509_, _22569_, _21526_);
  nor (_02452_, _10509_, _10508_);
  nor (_10510_, _24440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  nor (_10511_, _24442_, _21554_);
  nor (_02457_, _10511_, _10510_);
  nor (_10512_, _21796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5]);
  nor (_10513_, _21799_, _21451_);
  nor (_02460_, _10513_, _10512_);
  nor (_10514_, _24440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1]);
  nor (_10515_, _24442_, _21474_);
  nor (_02463_, _10515_, _10514_);
  nand (_10516_, _23282_, _23283_);
  nor (_10517_, _10516_, _24614_);
  nor (_10518_, _10517_, _24615_);
  nand (_10519_, _10518_, _24613_);
  not (_10520_, _23491_);
  nor (_10521_, _24611_, _10520_);
  nand (_25017_[2], _10521_, _10519_);
  nor (_10522_, _24440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  nor (_10523_, _24442_, _21586_);
  nor (_02477_, _10523_, _10522_);
  nor (_10524_, _21796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  nor (_10525_, _21799_, _21504_);
  nor (_02504_, _10525_, _10524_);
  nor (_10526_, _23843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1]);
  nor (_10527_, _23845_, _21474_);
  nor (_02506_, _10527_, _10526_);
  nor (_10528_, _23843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  nor (_10529_, _23845_, _21414_);
  nor (_02528_, _10529_, _10528_);
  nor (_10530_, _23843_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  nor (_10531_, _23845_, _21526_);
  nor (_02531_, _10531_, _10530_);
  nor (_10532_, _24440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5]);
  nor (_10533_, _24442_, _21451_);
  nor (_02566_, _10533_, _10532_);
  nor (_10534_, _24440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  nor (_10535_, _24442_, _21414_);
  nor (_25413_, _10535_, _10534_);
  nor (_10536_, _24440_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7]);
  nor (_10537_, _24442_, _21626_);
  nor (_02593_, _10537_, _10536_);
  nor (_10538_, _21856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1]);
  nor (_10539_, _21858_, _21474_);
  nor (_25209_, _10539_, _10538_);
  nor (_10540_, _21856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  nor (_10541_, _21858_, _21554_);
  nor (_02605_, _10541_, _10540_);
  nor (_10542_, _00868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  nor (_10543_, _00870_, _21414_);
  nor (_02617_, _10543_, _10542_);
  nor (_10544_, _00868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  nor (_10545_, _00870_, _21526_);
  nor (_02622_, _10545_, _10544_);
  nor (_10546_, _21653_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7]);
  nor (_10547_, _21655_, _21626_);
  nor (_02629_, _10547_, _10546_);
  nor (_10548_, _21796_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7]);
  nor (_10549_, _21799_, _21626_);
  nor (_02643_, _10549_, _10548_);
  nor (_10550_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  nor (_10551_, _24571_, _21586_);
  nor (_02661_, _10551_, _10550_);
  nor (_10552_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1]);
  nor (_10553_, _24609_, _21474_);
  nor (_02668_, _10553_, _10552_);
  nor (_10554_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  nor (_10555_, _24609_, _21526_);
  nor (_25348_, _10555_, _10554_);
  nor (_10556_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5]);
  nor (_10557_, _24609_, _21451_);
  nor (_25349_, _10557_, _10556_);
  nor (_10558_, _24607_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  nor (_10559_, _24609_, _21504_);
  nor (_02676_, _10559_, _10558_);
  nor (_10560_, _24601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5]);
  nor (_10561_, _24603_, _21451_);
  nor (_25342_, _10561_, _10560_);
  nor (_10562_, _24601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  nor (_10563_, _24603_, _21504_);
  nor (_02688_, _10563_, _10562_);
  nor (_10564_, _24593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  nor (_10565_, _24595_, _21586_);
  nor (_02692_, _10565_, _10564_);
  nor (_10566_, _24593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1]);
  nor (_10567_, _24595_, _21474_);
  nor (_02697_, _10567_, _10566_);
  nor (_10568_, _24593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  nor (_10569_, _24595_, _21414_);
  nor (_02703_, _10569_, _10568_);
  nor (_10570_, _24593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5]);
  nor (_10571_, _24595_, _21451_);
  nor (_02706_, _10571_, _10570_);
  nor (_10572_, _24593_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7]);
  nor (_10573_, _24595_, _21626_);
  nor (_02713_, _10573_, _10572_);
  nor (_10574_, _24583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  nor (_10575_, _24585_, _21586_);
  nor (_02716_, _10575_, _10574_);
  nor (_10577_, _24583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  nor (_10578_, _24585_, _21526_);
  nor (_25343_, _10578_, _10577_);
  nor (_10579_, _24583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  nor (_10580_, _24585_, _21414_);
  nor (_02733_, _10580_, _10579_);
  nor (_10581_, _24583_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  nor (_10582_, _24585_, _21504_);
  nor (_25344_, _10582_, _10581_);
  nor (_10583_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  nor (_10584_, _24577_, _21554_);
  nor (_02755_, _10584_, _10583_);
  nor (_10585_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  nor (_10586_, _24577_, _21526_);
  nor (_25346_, _10586_, _10585_);
  nor (_10587_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5]);
  nor (_10588_, _24577_, _21451_);
  nor (_02767_, _10588_, _10587_);
  nor (_10589_, _24575_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7]);
  nor (_10591_, _24577_, _21626_);
  nor (_02770_, _10591_, _10589_);
  nor (_10592_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  nor (_10593_, _24571_, _21554_);
  nor (_02776_, _10593_, _10592_);
  nor (_10594_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  nor (_10595_, _24571_, _21526_);
  nor (_02783_, _10595_, _10594_);
  nor (_10596_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5]);
  nor (_10597_, _24571_, _21451_);
  nor (_02786_, _10597_, _10596_);
  nor (_10598_, _24569_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7]);
  nor (_10599_, _24571_, _21626_);
  nor (_02788_, _10599_, _10598_);
  nor (_10600_, _24559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1]);
  nor (_10601_, _24561_, _21474_);
  nor (_02793_, _10601_, _10600_);
  nor (_10602_, _24559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  nor (_10603_, _24561_, _21526_);
  nor (_02796_, _10603_, _10602_);
  nor (_10604_, _24559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  nor (_10605_, _24561_, _21414_);
  nor (_25351_, _10605_, _10604_);
  nor (_10606_, _24559_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  nor (_10607_, _24561_, _21504_);
  nor (_02802_, _10607_, _10606_);
  nor (_10608_, _24551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1]);
  nor (_10609_, _24553_, _21474_);
  nor (_25352_, _10609_, _10608_);
  nor (_10610_, _24551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  nor (_10611_, _24553_, _21554_);
  nor (_02809_, _10611_, _10610_);
  nor (_10612_, _24551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5]);
  nor (_10613_, _24553_, _21451_);
  nor (_02812_, _10613_, _10612_);
  nor (_10614_, _24551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  nor (_10615_, _24553_, _21504_);
  nor (_02817_, _10615_, _10614_);
  nor (_10616_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  nor (_10617_, _24547_, _21586_);
  nor (_02829_, _10617_, _10616_);
  nor (_10618_, _21856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5]);
  nor (_10619_, _21858_, _21451_);
  nor (_02832_, _10619_, _10618_);
  nor (_10620_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1]);
  nor (_10621_, _24547_, _21474_);
  nor (_02834_, _10621_, _10620_);
  nor (_10622_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  nor (_10623_, _24547_, _21414_);
  nor (_25354_, _10623_, _10622_);
  nor (_10624_, _24545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  nor (_10625_, _24547_, _21504_);
  nor (_02837_, _10625_, _10624_);
  nor (_10626_, _24537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1]);
  nor (_10627_, _24539_, _21474_);
  nor (_25355_, _10627_, _10626_);
  nor (_10628_, _24537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  nor (_10629_, _24539_, _21526_);
  nor (_02844_, _10629_, _10628_);
  nor (_10630_, _24537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5]);
  nor (_10632_, _24539_, _21451_);
  nor (_02847_, _10632_, _10630_);
  nor (_10633_, _24537_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7]);
  nor (_10634_, _24539_, _21626_);
  nor (_02850_, _10634_, _10633_);
  nor (_10635_, _21646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1]);
  nor (_10636_, _21648_, _21474_);
  nor (_02853_, _10636_, _10635_);
  nor (_10637_, _24529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  nor (_10638_, _24531_, _21586_);
  nor (_02857_, _10638_, _10637_);
  nor (_10639_, _24529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  nor (_10640_, _24531_, _21526_);
  nor (_02859_, _10640_, _10639_);
  nor (_10641_, _24529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  nor (_10642_, _24531_, _21414_);
  nor (_02863_, _10642_, _10641_);
  nor (_10643_, _24529_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  nor (_10644_, _24531_, _21504_);
  nor (_02867_, _10644_, _10643_);
  nor (_10645_, _24521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  nor (_10646_, _24523_, _21554_);
  nor (_02872_, _10646_, _10645_);
  nor (_10647_, _24521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  nor (_10648_, _24523_, _21526_);
  nor (_02886_, _10648_, _10647_);
  nor (_10649_, _24521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5]);
  nor (_10650_, _24523_, _21451_);
  nor (_02888_, _10650_, _10649_);
  nor (_10651_, _24521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  nor (_10653_, _24523_, _21504_);
  nor (_02911_, _10653_, _10651_);
  nor (_10654_, _00868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7]);
  nor (_10655_, _00870_, _21626_);
  nor (_02919_, _10655_, _10654_);
  nor (_10656_, _00868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  nor (_10657_, _00870_, _21504_);
  nor (_25337_, _10657_, _10656_);
  nor (_10658_, _00868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5]);
  nor (_10659_, _00870_, _21451_);
  nor (_02934_, _10659_, _10658_);
  nor (_10660_, _24661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7]);
  nor (_10661_, _24663_, _21626_);
  nor (_02971_, _10661_, _10660_);
  nor (_10662_, _24661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  nor (_10663_, _24663_, _21504_);
  nor (_02977_, _10663_, _10662_);
  nor (_10664_, _00868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1]);
  nor (_10665_, _00870_, _21474_);
  nor (_03005_, _10665_, _10664_);
  nor (_10667_, _00868_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  nor (_10668_, _00870_, _21586_);
  nor (_03014_, _10668_, _10667_);
  nor (_10669_, _24661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1]);
  nor (_10670_, _24663_, _21474_);
  nor (_03045_, _10670_, _10669_);
  nor (_10671_, _24661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  nor (_10672_, _24663_, _21586_);
  nor (_03049_, _10672_, _10671_);
  nor (_10673_, _24666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7]);
  nor (_10674_, _24668_, _21626_);
  nor (_03057_, _10674_, _10673_);
  nor (_10675_, _24661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  nor (_10676_, _24663_, _21414_);
  nor (_03072_, _10676_, _10675_);
  nor (_10677_, _24661_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  nor (_10678_, _24663_, _21526_);
  nor (_25328_, _10678_, _10677_);
  nor (_10679_, _21856_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  nor (_10680_, _21858_, _21414_);
  nor (_03110_, _10680_, _10679_);
  nand (_10681_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_10682_, _10681_, _00985_);
  not (_10683_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand (_10684_, _00971_, _00954_);
  nand (_10685_, _10684_, _10683_);
  nand (_10686_, _10685_, _06667_);
  nand (_10687_, _10686_, _00996_);
  nor (_10688_, _10687_, _10682_);
  not (_10689_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nand (_10690_, _00991_, _10689_);
  nand (_10691_, _10690_, _01006_);
  nor (_10692_, _10691_, _10688_);
  nor (_10693_, _01013_, ABINPUT[9]);
  nor (_10694_, _10693_, _01239_);
  nor (_10695_, _10694_, _10692_);
  nand (_10696_, _01013_, _10683_);
  nand (_10697_, _10696_, _23493_);
  nor (_03114_, _10697_, _10695_);
  nor (_10698_, _21646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  nor (_10699_, _21648_, _21554_);
  nor (_03119_, _10699_, _10698_);
  nor (_10700_, _24666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  nor (_10701_, _24668_, _21526_);
  nor (_03122_, _10701_, _10700_);
  nor (_10702_, _24666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  nor (_10703_, _24668_, _21554_);
  nor (_03127_, _10703_, _10702_);
  nor (_10704_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5]);
  nor (_10705_, _22537_, _21451_);
  nor (_03130_, _10705_, _10704_);
  nor (_10706_, _24666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  nor (_10707_, _24668_, _21504_);
  nor (_03137_, _10707_, _10706_);
  nor (_10708_, _24666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5]);
  nor (_10709_, _24668_, _21451_);
  nor (_03148_, _10709_, _10708_);
  nor (_10710_, _24666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  nor (_10711_, _24668_, _21414_);
  nor (_03150_, _10711_, _10710_);
  nor (_10712_, _24670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  nor (_10713_, _24672_, _21414_);
  nor (_25279_, _10713_, _10712_);
  nor (_10714_, _24670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  nor (_10715_, _24672_, _21504_);
  nor (_25280_, _10715_, _10714_);
  nand (_10716_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor (_10717_, _10716_, _00985_);
  nand (_10718_, _00969_, _00954_);
  nand (_10719_, _10718_, _00960_);
  nand (_10720_, _10719_, _10684_);
  nand (_10721_, _10720_, _00996_);
  nor (_10722_, _10721_, _10717_);
  nand (_10723_, _00991_, _01111_);
  nand (_10724_, _10723_, _01006_);
  nor (_10725_, _10724_, _10722_);
  nor (_10726_, _01013_, ABINPUT[8]);
  nor (_10727_, _10726_, _01239_);
  nor (_10728_, _10727_, _10725_);
  nand (_10729_, _01013_, _00960_);
  nand (_10730_, _10729_, _23493_);
  nor (_03164_, _10730_, _10728_);
  nor (_10731_, _24670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5]);
  nor (_10732_, _24672_, _21451_);
  nor (_03167_, _10732_, _10731_);
  nor (_10733_, _21646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  nor (_10734_, _21648_, _21526_);
  nor (_03183_, _10734_, _10733_);
  nor (_10735_, _24666_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  nor (_10736_, _24668_, _21586_);
  nor (_03201_, _10736_, _10735_);
  nor (_10737_, _24670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7]);
  nor (_10738_, _24672_, _21626_);
  nor (_03208_, _10738_, _10737_);
  nor (_10739_, _22521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  nor (_10740_, _22524_, _21414_);
  nor (_03212_, _10740_, _10739_);
  nor (_10741_, _21919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  nor (_10742_, _21922_, _21586_);
  nor (_03219_, _10742_, _10741_);
  nor (_10743_, _00674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  nor (_10744_, _00676_, _21504_);
  nor (_03223_, _10744_, _10743_);
  nor (_10745_, _00674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7]);
  nor (_10746_, _00676_, _21626_);
  nor (_03231_, _10746_, _10745_);
  nor (_10747_, _24670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  nor (_10748_, _24672_, _21554_);
  nor (_03256_, _10748_, _10747_);
  nor (_10749_, _24670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1]);
  nor (_10750_, _24672_, _21474_);
  nor (_03260_, _10750_, _10749_);
  nor (_10751_, _24670_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  nor (_10752_, _24672_, _21586_);
  nor (_03267_, _10752_, _10751_);
  nor (_10753_, _21645_, _21631_);
  nor (_10754_, _10753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  not (_10755_, _10753_);
  nor (_10756_, _10755_, _21586_);
  nor (_03274_, _10756_, _10754_);
  nor (_10758_, _22403_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7]);
  nor (_10759_, _22406_, _21626_);
  nor (_25115_, _10759_, _10758_);
  nor (_10760_, _00674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  nor (_10761_, _00676_, _21586_);
  nor (_03282_, _10761_, _10760_);
  nor (_10762_, _00855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7]);
  nor (_10763_, _00857_, _21626_);
  nor (_03300_, _10763_, _10762_);
  nor (_10764_, _00855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  nor (_10765_, _00857_, _21504_);
  nor (_03304_, _10765_, _10764_);
  nor (_10766_, _22526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  nor (_10767_, _22528_, _21586_);
  nor (_03310_, _10767_, _10766_);
  nor (_10768_, _00674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  nor (_10769_, _00676_, _21526_);
  nor (_03320_, _10769_, _10768_);
  nor (_10770_, _00674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  nor (_10771_, _00676_, _21554_);
  nor (_03325_, _10771_, _10770_);
  nor (_10772_, _00674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1]);
  nor (_10773_, _00676_, _21474_);
  nor (_03329_, _10773_, _10772_);
  nor (_10774_, _00855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1]);
  nor (_10775_, _00857_, _21474_);
  nor (_03356_, _10775_, _10774_);
  nor (_10776_, _21645_, _21607_);
  nor (_10777_, _10776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  not (_10778_, _10776_);
  nor (_10780_, _10778_, _21414_);
  nor (_03360_, _10780_, _10777_);
  nor (_10781_, _00855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  nor (_10782_, _00857_, _21586_);
  nor (_25245_, _10782_, _10781_);
  nor (_10783_, _10776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7]);
  nor (_10784_, _10778_, _21626_);
  nor (_25286_, _10784_, _10783_);
  nor (_10785_, _00855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  nor (_10786_, _00857_, _21414_);
  nor (_03387_, _10786_, _10785_);
  nor (_10787_, _00855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  nor (_10788_, _00857_, _21526_);
  nor (_03390_, _10788_, _10787_);
  nor (_10789_, _00855_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  nor (_10790_, _00857_, _21554_);
  nor (_03397_, _10790_, _10789_);
  nor (_10791_, _24674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  nor (_10792_, _24676_, _21554_);
  nor (_03418_, _10792_, _10791_);
  nor (_10793_, _24674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1]);
  nor (_10794_, _24676_, _21474_);
  nor (_03426_, _10794_, _10793_);
  not (_10795_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor (_10796_, _04981_, _21337_);
  nand (_10797_, _10796_, _21426_);
  nor (_10798_, _10797_, _24858_);
  nor (_10799_, _10798_, _10795_);
  not (_10800_, _04991_);
  nor (_10801_, _10797_, _10800_);
  nor (_10802_, _10801_, _10799_);
  nor (_10803_, _10802_, _00915_);
  nand (_10804_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  not (_10805_, _10799_);
  nand (_10806_, _10798_, ABINPUT[19]);
  nand (_10807_, _10806_, _10805_);
  nand (_10808_, _10807_, _24861_);
  nand (_10809_, _10808_, _10804_);
  nor (_10810_, _10809_, _10803_);
  nor (_03430_, _10810_, rst);
  not (_10811_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_10812_, _10797_, _00020_);
  nor (_10813_, _10812_, _10811_);
  nor (_10814_, _10797_, _05140_);
  nor (_10815_, _10814_, _10813_);
  nor (_10816_, _10815_, _00915_);
  nand (_10817_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  not (_10818_, ABINPUT[20]);
  nand (_10819_, _10798_, _10818_);
  nor (_10820_, _10798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_10821_, _10820_, _00010_);
  nand (_10822_, _10821_, _10819_);
  nand (_10823_, _10822_, _10817_);
  nor (_10824_, _10823_, _10816_);
  nor (_03438_, _10824_, rst);
  not (_10825_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_10826_, _10797_, _00909_);
  nor (_10827_, _10826_, _10825_);
  not (_10828_, _00931_);
  nor (_10829_, _10797_, _10828_);
  nor (_10830_, _10829_, _10827_);
  nor (_10831_, _10830_, _00915_);
  nand (_10832_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not (_10833_, ABINPUT[22]);
  nand (_10834_, _10798_, _10833_);
  nor (_10835_, _10798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_10836_, _10835_, _00010_);
  nand (_10837_, _10836_, _10834_);
  nand (_10838_, _10837_, _10832_);
  nor (_10839_, _10838_, _10831_);
  nor (_03441_, _10839_, rst);
  not (_10840_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nor (_10841_, _10797_, _01027_);
  nor (_10842_, _10841_, _10840_);
  nor (_10843_, _10797_, _02493_);
  nor (_10844_, _10843_, _10842_);
  nor (_10845_, _10844_, _00915_);
  nand (_10846_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  not (_10847_, ABINPUT[21]);
  nand (_10848_, _10798_, _10847_);
  nor (_10850_, _10798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nor (_10851_, _10850_, _00010_);
  nand (_10852_, _10851_, _10848_);
  nand (_10853_, _10852_, _10846_);
  nor (_10854_, _10853_, _10845_);
  nor (_03444_, _10854_, rst);
  not (_10855_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor (_10856_, _10797_, _01010_);
  nor (_10857_, _10856_, _10855_);
  not (_10858_, _05018_);
  nor (_10859_, _10797_, _10858_);
  nor (_10860_, _10859_, _10857_);
  nor (_10861_, _10860_, _00915_);
  nand (_10862_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_10863_, ABINPUT[24]);
  nand (_10864_, _10798_, _10863_);
  nor (_10865_, _10798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nor (_10866_, _10865_, _00010_);
  nand (_10867_, _10866_, _10864_);
  nand (_10868_, _10867_, _10862_);
  nor (_10869_, _10868_, _10861_);
  nor (_03453_, _10869_, rst);
  not (_10870_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor (_10871_, _10797_, _01001_);
  nor (_10872_, _10871_, _10870_);
  not (_10873_, _01093_);
  nor (_10874_, _10797_, _10873_);
  nor (_10875_, _10874_, _10872_);
  nor (_10876_, _10875_, _00915_);
  nand (_10877_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_10878_, ABINPUT[23]);
  nand (_10879_, _10798_, _10878_);
  nor (_10880_, _10798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nor (_10881_, _10880_, _00010_);
  nand (_10882_, _10881_, _10879_);
  nand (_10883_, _10882_, _10877_);
  nor (_10884_, _10883_, _10876_);
  nor (_03457_, _10884_, rst);
  nor (_10885_, _24674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  nor (_10886_, _24676_, _21526_);
  nor (_03460_, _10886_, _10885_);
  nor (_10887_, _21646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  nor (_10888_, _21648_, _21414_);
  nor (_03465_, _10888_, _10887_);
  nor (_10889_, _21816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5]);
  nor (_10890_, _21818_, _21451_);
  nor (_03467_, _10890_, _10889_);
  not (_10891_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor (_10892_, _10797_, _05055_);
  nor (_10893_, _10892_, _10891_);
  nor (_10895_, _10797_, _05125_);
  nor (_10896_, _10895_, _10893_);
  nor (_10897_, _10896_, _00915_);
  nand (_10898_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  not (_10899_, ABINPUT[25]);
  nand (_10900_, _10798_, _10899_);
  nor (_10901_, _10798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nor (_10902_, _10901_, _00010_);
  nand (_10903_, _10902_, _10900_);
  nand (_10904_, _10903_, _10898_);
  nor (_10905_, _10904_, _10897_);
  nor (_03470_, _10905_, rst);
  nor (_10906_, _24674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5]);
  nor (_10907_, _24676_, _21451_);
  nor (_03473_, _10907_, _10906_);
  nor (_10908_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  nor (_10909_, _22221_, _21504_);
  nor (_03478_, _10909_, _10908_);
  nor (_10910_, _24674_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  nor (_10911_, _24676_, _21414_);
  nor (_25228_, _10911_, _10910_);
  nor (_10913_, _03976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  nor (_10914_, _03978_, _21526_);
  nor (_25296_, _10914_, _10913_);
  nor (_10915_, _09002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5]);
  nor (_10916_, _09004_, _21451_);
  nor (_03501_, _10916_, _10915_);
  nor (_10917_, _21919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  nor (_10918_, _21922_, _21526_);
  nor (_03505_, _10918_, _10917_);
  nor (_10919_, _00678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  nor (_10920_, _00681_, _21414_);
  nor (_03531_, _10920_, _10919_);
  nor (_10921_, _21919_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  nor (_10922_, _21922_, _21414_);
  nor (_03533_, _10922_, _10921_);
  nor (_10923_, _00678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  nor (_10924_, _00681_, _21526_);
  nor (_03542_, _10924_, _10923_);
  nor (_10925_, _21646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  nor (_10926_, _21648_, _21504_);
  nor (_03545_, _10926_, _10925_);
  nor (_10927_, _00678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  nor (_10928_, _00681_, _21554_);
  nor (_03547_, _10928_, _10927_);
  nor (_10929_, _00678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5]);
  nor (_10930_, _00681_, _21451_);
  nor (_03561_, _10930_, _10929_);
  nor (_10931_, _00678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7]);
  nor (_10932_, _00681_, _21626_);
  nor (_25216_, _10932_, _10931_);
  nor (_10933_, _00678_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  nor (_10934_, _00681_, _21504_);
  nor (_25215_, _10934_, _10933_);
  nand (_10935_, _00848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  nor (_10936_, _00848_, _24867_);
  not (_10937_, _10936_);
  nand (_03597_, _10937_, _10935_);
  nor (_10938_, _00847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5]);
  nor (_10939_, _00848_, _21451_);
  nor (_03601_, _10939_, _10938_);
  nand (_10940_, _00848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  nor (_10941_, _00848_, _24900_);
  not (_10942_, _10941_);
  nand (_03606_, _10942_, _10940_);
  not (_10943_, _05764_);
  nand (_10944_, _00848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7]);
  nand (_03634_, _10944_, _10943_);
  nor (_10945_, _09002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  nor (_10946_, _09004_, _21414_);
  nor (_03637_, _10946_, _10945_);
  nor (_10947_, _00847_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  nor (_10948_, _00848_, _21504_);
  nor (_03640_, _10948_, _10947_);
  nor (_10949_, _24684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7]);
  nor (_10950_, _24686_, _21626_);
  nor (_03647_, _10950_, _10949_);
  nor (_10951_, _24684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  nor (_10952_, _24686_, _21504_);
  nor (_03651_, _10952_, _10951_);
  nor (_03655_, _00354_, rst);
  nor (_03658_, _00552_, rst);
  nand (_10953_, _00848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1]);
  nor (_10954_, _00848_, _00006_);
  not (_10955_, _10954_);
  nand (_25203_, _10955_, _10953_);
  nand (_10956_, _00848_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  nor (_10957_, _00848_, _00029_);
  not (_10958_, _10957_);
  nand (_03663_, _10958_, _10956_);
  nor (_10959_, _24684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  nor (_10960_, _24686_, _21586_);
  nor (_03684_, _10960_, _10959_);
  nor (_10961_, _21949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  nor (_10962_, _21952_, _21554_);
  nor (_03690_, _10962_, _10961_);
  nor (_10963_, _24684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  nor (_10964_, _24686_, _21526_);
  nor (_03693_, _10964_, _10963_);
  nor (_10965_, _24684_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  nor (_10966_, _24686_, _21554_);
  nor (_03696_, _10966_, _10965_);
  nor (_10967_, _01194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1]);
  nor (_10968_, _01196_, _21474_);
  nor (_03699_, _10968_, _10967_);
  nor (_10969_, rst, _21183_);
  nand (_10970_, _10969_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_10971_, _24410_, _23203_);
  nor (_10972_, _10971_, _24393_);
  not (_10973_, _10972_);
  nor (_10975_, _24410_, _23253_);
  not (_10976_, _10975_);
  nor (_10977_, _23251_, _23359_);
  nor (_10978_, _10977_, _24387_);
  nor (_10979_, _10978_, _24411_);
  nand (_10980_, _10979_, _10976_);
  nor (_10981_, _10980_, _10973_);
  not (_10982_, _00235_);
  nand (_10983_, _23514_, _23410_);
  nand (_10984_, _10983_, _23528_);
  nand (_10985_, _23415_, _23409_);
  nand (_10986_, _10985_, _10984_);
  not (_10987_, _24729_);
  nand (_10988_, _00232_, _23527_);
  nand (_10989_, _10988_, _10987_);
  nor (_10990_, _23415_, _23253_);
  nor (_10991_, _01277_, _23415_);
  nor (_10992_, _10991_, _10990_);
  not (_10993_, _10992_);
  nor (_10994_, _10993_, _10989_);
  nand (_10996_, _10994_, _10986_);
  nor (_10997_, _10996_, _10982_);
  nand (_10998_, _10997_, _10981_);
  nand (_10999_, _10998_, _23491_);
  nand (_25022_[0], _10999_, _10970_);
  nor (_11000_, _01198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  nor (_11001_, _01200_, _21586_);
  nor (_03707_, _11001_, _11000_);
  nor (_11002_, _21913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  nor (_11003_, _21915_, _21554_);
  nor (_25211_, _11003_, _11002_);
  nor (_11004_, _00723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_11005_, _00725_, _21414_);
  nor (_25151_, _11005_, _11004_);
  nor (_11006_, _03976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  nor (_11007_, _03978_, _21414_);
  nor (_03713_, _11007_, _11006_);
  nor (_11008_, _00723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_11009_, _00725_, _21526_);
  nor (_03715_, _11009_, _11008_);
  nor (_11011_, _00723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_11012_, _00725_, _21554_);
  nor (_03716_, _11012_, _11011_);
  nor (_11013_, _00723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7]);
  nor (_11014_, _00725_, _21626_);
  nor (_03749_, _11014_, _11013_);
  nor (_11015_, _00723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_11016_, _00725_, _21504_);
  nor (_03757_, _11016_, _11015_);
  nor (_11017_, _00723_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5]);
  nor (_11018_, _00725_, _21451_);
  nor (_03762_, _11018_, _11017_);
  not (_11019_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_11020_, _00742_, _11019_);
  nor (_11021_, _00740_, _00029_);
  nor (_11022_, _11021_, _11020_);
  nor (_03778_, _11022_, rst);
  nor (_11023_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_11024_, _24692_, _21504_);
  nor (_03780_, _11024_, _11023_);
  nor (_11026_, _00740_, _00006_);
  nor (_11027_, _00742_, _24954_);
  nor (_11028_, _11027_, _11026_);
  nor (_03782_, _11028_, rst);
  nor (_11029_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5]);
  nor (_11030_, _24692_, _21451_);
  nor (_03786_, _11030_, _11029_);
  nor (_11031_, _00740_, _00121_);
  nor (_11032_, _00742_, _00484_);
  nor (_11033_, _11032_, _11031_);
  nor (_03789_, _11033_, rst);
  nor (_11034_, _00742_, _00412_);
  nor (_11035_, _00740_, _24867_);
  nor (_11036_, _11035_, _11034_);
  nor (_03791_, _11036_, rst);
  nor (_11037_, _00740_, _24900_);
  nor (_11038_, _00742_, _00183_);
  nor (_11039_, _11038_, _11037_);
  nor (_03797_, _11039_, rst);
  nor (_11040_, _00742_, _00265_);
  nor (_11042_, _00740_, _00129_);
  nor (_11043_, _11042_, _11040_);
  nor (_03800_, _11043_, rst);
  nor (_11044_, _00740_, _00114_);
  nor (_11045_, _00742_, _00338_);
  nor (_11046_, _11045_, _11044_);
  nor (_03801_, _11046_, rst);
  nor (_11047_, _05722_, _00577_);
  nor (_11048_, _05721_, _00029_);
  nor (_11049_, _11048_, _11047_);
  nor (_03813_, _11049_, rst);
  nor (_11050_, _05722_, _24933_);
  nor (_11051_, _05721_, _00006_);
  nor (_11052_, _11051_, _11050_);
  nor (_03816_, _11052_, rst);
  nor (_11053_, _05722_, _00473_);
  nor (_11054_, _05721_, _00121_);
  nor (_11055_, _11054_, _11053_);
  nor (_03818_, _11055_, rst);
  nor (_11056_, _05722_, _00405_);
  nor (_11058_, _05721_, _24867_);
  nor (_11059_, _11058_, _11056_);
  nor (_03820_, _11059_, rst);
  nor (_11060_, _05722_, _00188_);
  nor (_11061_, _05721_, _24900_);
  nor (_11062_, _11061_, _11060_);
  nor (_25024_[4], _11062_, rst);
  nor (_11063_, _05722_, _00259_);
  nor (_11064_, _05721_, _00129_);
  nor (_11065_, _11064_, _11063_);
  nor (_25024_[5], _11065_, rst);
  nor (_11066_, _05722_, _00326_);
  nor (_11067_, _05721_, _00114_);
  nor (_11068_, _11067_, _11066_);
  nor (_25024_[6], _11068_, rst);
  nor (_11069_, _21949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  nor (_11070_, _21952_, _21414_);
  nor (_03846_, _11070_, _11069_);
  nor (_11071_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1]);
  nor (_11072_, _24692_, _21474_);
  nor (_03848_, _11072_, _11071_);
  nor (_11074_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_11075_, _24692_, _21586_);
  nor (_03853_, _11075_, _11074_);
  nor (_11076_, _05729_, _00572_);
  nor (_11077_, _05733_, _00029_);
  nor (_11078_, _11077_, _11076_);
  nor (_03859_, _11078_, rst);
  nor (_11079_, _05729_, _24923_);
  nor (_11080_, _05733_, _00006_);
  nor (_11081_, _11080_, _11079_);
  nor (_03861_, _11081_, rst);
  nor (_11082_, _05729_, _00490_);
  nor (_11083_, _05733_, _00121_);
  nor (_11084_, _11083_, _11082_);
  nor (_03863_, _11084_, rst);
  nor (_11085_, _05729_, _00400_);
  nor (_11086_, _05733_, _24867_);
  nor (_11087_, _11086_, _11085_);
  nor (_03865_, _11087_, rst);
  nor (_11088_, _05729_, _00196_);
  nor (_11089_, _05733_, _24900_);
  nor (_11090_, _11089_, _11088_);
  nor (_25025_[4], _11090_, rst);
  nor (_11091_, _05729_, _00253_);
  nor (_11092_, _05733_, _00129_);
  nor (_11093_, _11092_, _11091_);
  nor (_25025_[5], _11093_, rst);
  nor (_11094_, _24690_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_11095_, _24692_, _21526_);
  nor (_03871_, _11095_, _11094_);
  nor (_11096_, _05729_, _00343_);
  nor (_11097_, _05733_, _00114_);
  nor (_11098_, _11097_, _11096_);
  nor (_03873_, _11098_, rst);
  nand (_03875_, _00628_, _23493_);
  nand (_03878_, _00047_, _23493_);
  nand (_03880_, _00526_, _23493_);
  nor (_03882_, _00218_, rst);
  nor (_03884_, _00433_, rst);
  nor (_03887_, _00360_, rst);
  nor (_03888_, _00311_, rst);
  nor (_11099_, _05740_, _00569_);
  nor (_11100_, _05744_, _00029_);
  nor (_11101_, _11100_, _11099_);
  nor (_25026_[0], _11101_, rst);
  nor (_11102_, _05740_, _24946_);
  nor (_11103_, _05744_, _00006_);
  nor (_11104_, _11103_, _11102_);
  nor (_03892_, _11104_, rst);
  nor (_11105_, _00727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nor (_11106_, _00730_, _21554_);
  nor (_03895_, _11106_, _11105_);
  nor (_11107_, _00727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nor (_11108_, _00730_, _21526_);
  nor (_03899_, _11108_, _11107_);
  nor (_11109_, _05740_, _00478_);
  nor (_11110_, _05744_, _00121_);
  nor (_11111_, _11110_, _11109_);
  nor (_03901_, _11111_, rst);
  nor (_11112_, _05740_, _00418_);
  nor (_11113_, _05744_, _24867_);
  nor (_11114_, _11113_, _11112_);
  nor (_03904_, _11114_, rst);
  nor (_11115_, _05740_, _00194_);
  nor (_11116_, _05744_, _24900_);
  nor (_11117_, _11116_, _11115_);
  nor (_03906_, _11117_, rst);
  nor (_11118_, _05740_, _00270_);
  nor (_11119_, _05744_, _00129_);
  nor (_11120_, _11119_, _11118_);
  nor (_03908_, _11120_, rst);
  nor (_11121_, _05740_, _00332_);
  nor (_11122_, _05744_, _00114_);
  nor (_11123_, _11122_, _11121_);
  nor (_03911_, _11123_, rst);
  nor (_11124_, _05753_, _00582_);
  nor (_11125_, _05755_, _00029_);
  nor (_11126_, _11125_, _11124_);
  nor (_03928_, _11126_, rst);
  nor (_11127_, _05753_, _24918_);
  nor (_11128_, _05755_, _00006_);
  nor (_11129_, _11128_, _11127_);
  nor (_03930_, _11129_, rst);
  nor (_11130_, _00727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5]);
  nor (_11131_, _00730_, _21451_);
  nor (_03933_, _11131_, _11130_);
  nor (_11132_, _05753_, _00487_);
  nor (_11133_, _05755_, _00121_);
  nor (_11134_, _11133_, _11132_);
  nor (_25027_[2], _11134_, rst);
  nor (_11135_, _05753_, _00398_);
  nor (_11136_, _05755_, _24867_);
  nor (_11137_, _11136_, _11135_);
  nor (_03936_, _11137_, rst);
  nor (_11138_, _05753_, _00201_);
  nor (_11139_, _05755_, _24900_);
  nor (_11140_, _11139_, _11138_);
  nor (_03938_, _11140_, rst);
  nor (_11141_, _05753_, _00263_);
  nor (_11143_, _05755_, _00129_);
  nor (_11144_, _11143_, _11141_);
  nor (_03941_, _11144_, rst);
  nor (_11145_, _05753_, _00341_);
  nor (_11146_, _05755_, _00114_);
  nor (_11147_, _11146_, _11145_);
  nor (_03943_, _11147_, rst);
  nor (_11148_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_11149_, _24698_, _21504_);
  nor (_03946_, _11149_, _11148_);
  nor (_11150_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5]);
  nor (_11151_, _24698_, _21451_);
  nor (_03951_, _11151_, _11150_);
  nor (_11152_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nor (_11153_, _24698_, _21414_);
  nor (_03955_, _11153_, _11152_);
  nor (_11154_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nor (_11155_, _24698_, _21526_);
  nor (_03957_, _11155_, _11154_);
  nor (_11156_, _00847_, _00575_);
  nor (_11158_, _11156_, _10957_);
  nor (_25028_[0], _11158_, rst);
  nor (_11159_, _00847_, _24928_);
  nor (_11160_, _11159_, _10954_);
  nor (_25028_[1], _11160_, rst);
  nor (_11161_, _00847_, _00482_);
  nor (_11162_, _11161_, _00850_);
  nor (_03962_, _11162_, rst);
  nor (_11163_, _00847_, _00410_);
  nor (_11164_, _11163_, _10936_);
  nor (_03964_, _11164_, rst);
  nor (_11165_, _00847_, _00199_);
  nor (_11166_, _11165_, _10941_);
  nor (_03967_, _11166_, rst);
  nor (_11167_, _00847_, _00251_);
  nor (_11168_, _00848_, _00129_);
  nor (_11169_, _11168_, _11167_);
  nor (_03969_, _11169_, rst);
  nor (_11170_, _00847_, _00336_);
  nor (_11171_, _00848_, _00114_);
  nor (_11172_, _11171_, _11170_);
  nor (_03971_, _11172_, rst);
  nor (_11173_, _00727_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nor (_11174_, _00730_, _21586_);
  nor (_03973_, _11174_, _11173_);
  nor (_11175_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7]);
  nor (_11176_, _24698_, _21626_);
  nor (_25093_, _11176_, _11175_);
  nor (_11177_, _00827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5]);
  nor (_11178_, _00829_, _21451_);
  nor (_03983_, _11178_, _11177_);
  nor (_11179_, _00827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7]);
  nor (_11180_, _00829_, _21626_);
  nor (_25073_, _11180_, _11179_);
  nor (_11181_, _00827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_11182_, _00829_, _21504_);
  nor (_03991_, _11182_, _11181_);
  nor (_11183_, _24661_, _00586_);
  nor (_11184_, _24663_, _00029_);
  nor (_11185_, _11184_, _11183_);
  nor (_04008_, _11185_, rst);
  nor (_11186_, _05696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  nor (_11187_, _05699_, _21504_);
  nor (_04011_, _11187_, _11186_);
  nor (_11188_, _24661_, _24951_);
  nor (_11189_, _24663_, _00006_);
  nor (_11190_, _11189_, _11188_);
  nor (_04013_, _11190_, rst);
  nor (_11191_, _24661_, _00476_);
  nor (_11192_, _11191_, _00866_);
  nor (_04016_, _11192_, rst);
  nor (_11193_, _24661_, _00416_);
  nor (_11194_, _24663_, _24867_);
  nor (_11195_, _11194_, _11193_);
  nor (_04019_, _11195_, rst);
  nor (_11196_, _24661_, _00186_);
  nor (_11197_, _24663_, _24900_);
  nor (_11198_, _11197_, _11196_);
  nor (_04021_, _11198_, rst);
  nor (_11199_, _01194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7]);
  nor (_11200_, _01196_, _21626_);
  nor (_04025_, _11200_, _11199_);
  nor (_11201_, _01194_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  nor (_11202_, _01196_, _21414_);
  nor (_04028_, _11202_, _11201_);
  nor (_11203_, _24661_, _00268_);
  nor (_11204_, _24663_, _00129_);
  nor (_11205_, _11204_, _11203_);
  nor (_25029_[5], _11205_, rst);
  nor (_11206_, _24661_, _00329_);
  nor (_11207_, _24663_, _00114_);
  nor (_11208_, _11207_, _11206_);
  nor (_04031_, _11208_, rst);
  nor (_11209_, _05952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5]);
  nor (_11210_, _05954_, _21451_);
  nor (_04036_, _11210_, _11209_);
  nor (_11211_, _05952_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  nor (_11212_, _05954_, _21554_);
  nor (_04039_, _11212_, _11211_);
  nor (_11213_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1]);
  nor (_11214_, _24698_, _21474_);
  nor (_04042_, _11214_, _11213_);
  nor (_11215_, _24696_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nor (_11216_, _24698_, _21586_);
  nor (_04044_, _11216_, _11215_);
  nor (_11217_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1]);
  nor (_11218_, _02331_, _21474_);
  nor (_04047_, _11218_, _11217_);
  nor (_11219_, _02328_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  nor (_11220_, _02331_, _21414_);
  nor (_04050_, _11220_, _11219_);
  not (_11221_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_11222_, _05774_, _11221_);
  nor (_11223_, _05777_, _00029_);
  nor (_11224_, _11223_, _11222_);
  nor (_04054_, _11224_, rst);
  nor (_11225_, _05774_, _24940_);
  nor (_11226_, _05777_, _00006_);
  nor (_11227_, _11226_, _11225_);
  nor (_04056_, _11227_, rst);
  nor (_11229_, _05774_, _00471_);
  nor (_11230_, _05777_, _00121_);
  nor (_11231_, _11230_, _11229_);
  nor (_25030_[2], _11231_, rst);
  nor (_11232_, _05774_, _00403_);
  nor (_11233_, _05777_, _24867_);
  nor (_11234_, _11233_, _11232_);
  nor (_04059_, _11234_, rst);
  nor (_11235_, _05774_, _00181_);
  nor (_11236_, _05777_, _24900_);
  nor (_11237_, _11236_, _11235_);
  nor (_25030_[4], _11237_, rst);
  nor (_11238_, _06831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  nor (_11239_, _06834_, _21504_);
  nor (_25325_, _11239_, _11238_);
  nor (_11240_, _00827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_11241_, _00829_, _21586_);
  nor (_04066_, _11241_, _11240_);
  nor (_11242_, _05774_, _00256_);
  nor (_11243_, _05777_, _00129_);
  nor (_11244_, _11243_, _11242_);
  nor (_04068_, _11244_, rst);
  nor (_11245_, _06831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  nor (_11246_, _06834_, _21526_);
  nor (_04071_, _11246_, _11245_);
  nor (_11247_, _06831_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1]);
  nor (_11248_, _06834_, _21474_);
  nor (_04074_, _11248_, _11247_);
  nor (_11249_, _05774_, _00324_);
  nor (_11250_, _05777_, _00114_);
  nor (_11251_, _11250_, _11249_);
  nor (_04077_, _11251_, rst);
  nor (_11252_, _24702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7]);
  nor (_11253_, _24704_, _21626_);
  nor (_04080_, _11253_, _11252_);
  nor (_11254_, _02427_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  nor (_11255_, _02430_, _21504_);
  nor (_25322_, _11255_, _11254_);
  nor (_11256_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  nor (_11257_, _22783_, _21526_);
  nor (_04090_, _11257_, _11256_);
  nor (_11259_, _07002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7]);
  nor (_11260_, _07004_, _21626_);
  nor (_04093_, _11260_, _11259_);
  nor (_11261_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  nor (_11262_, _22783_, _21554_);
  nor (_25128_, _11262_, _11261_);
  nor (_11263_, _02383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  nor (_11264_, _02385_, _21414_);
  nor (_04100_, _11264_, _11263_);
  nor (_11265_, _00827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_11266_, _00829_, _21526_);
  nor (_04106_, _11266_, _11265_);
  nor (_11267_, _00827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_11268_, _00829_, _21554_);
  nor (_04125_, _11268_, _11267_);
  nor (_11269_, _00827_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1]);
  nor (_11270_, _00829_, _21474_);
  nor (_04128_, _11270_, _11269_);
  nand (_11271_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nor (_11272_, _11271_, _00985_);
  nand (_11273_, _00954_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_11274_, _11273_, _00963_);
  nand (_11275_, _11274_, _01259_);
  nand (_11276_, _11275_, _00996_);
  nor (_11277_, _11276_, _11272_);
  not (_11278_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nand (_11279_, _00991_, _11278_);
  nand (_11280_, _11279_, _01006_);
  nor (_11281_, _11280_, _11277_);
  nor (_11282_, _01013_, ABINPUT[4]);
  nor (_11283_, _11282_, _01239_);
  nor (_11284_, _11283_, _11281_);
  nand (_11285_, _01013_, _00963_);
  nand (_11286_, _11285_, _23493_);
  nor (_04136_, _11286_, _11284_);
  nor (_11287_, _21949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  nor (_11288_, _21952_, _21526_);
  nor (_04141_, _11288_, _11287_);
  nor (_11289_, _03976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  nor (_11291_, _03978_, _21504_);
  nor (_04144_, _11291_, _11289_);
  nor (_11292_, _24702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_11293_, _24704_, _21586_);
  nor (_25061_, _11293_, _11292_);
  nor (_11294_, _24702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1]);
  nor (_11295_, _24704_, _21474_);
  nor (_04170_, _11295_, _11294_);
  nor (_11296_, _24702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_11297_, _24704_, _21414_);
  nor (_25062_, _11297_, _11296_);
  nor (_11298_, _24702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_11299_, _24704_, _21526_);
  nor (_04182_, _11299_, _11298_);
  nor (_11300_, _24702_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_11301_, _24704_, _21554_);
  nor (_04187_, _11301_, _11300_);
  nand (_11302_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nand (_11303_, _01142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nand (_11304_, _11303_, _11302_);
  nor (_11305_, _11304_, _01130_);
  nor (_11306_, _01059_, _00006_);
  nor (_11307_, _01055_, _00029_);
  nor (_11308_, _11307_, _11306_);
  nand (_11309_, _11308_, _01130_);
  nand (_11310_, _11309_, _23493_);
  nor (_04193_, _11310_, _11305_);
  nor (_11311_, _00954_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nand (_11312_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor (_11313_, _11312_, _00983_);
  nor (_11314_, _11313_, _11273_);
  nor (_11315_, _11314_, _11311_);
  nor (_11316_, _11315_, _00991_);
  nand (_11317_, _00991_, _01219_);
  nand (_11318_, _11317_, _01006_);
  nor (_11319_, _11318_, _11316_);
  nor (_11320_, _01013_, ABINPUT[3]);
  nor (_11321_, _11320_, _01239_);
  nor (_11322_, _11321_, _11319_);
  nand (_11323_, _01013_, _00964_);
  nand (_11324_, _11323_, _23493_);
  nor (_04198_, _11324_, _11322_);
  nor (_11325_, _00818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nor (_11326_, _00820_, _21586_);
  nor (_04217_, _11326_, _11325_);
  nor (_11327_, _00818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nor (_11328_, _00820_, _21554_);
  nor (_04223_, _11328_, _11327_);
  nor (_11329_, _03976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5]);
  nor (_11330_, _03978_, _21451_);
  nor (_04227_, _11330_, _11329_);
  nor (_11331_, _00818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1]);
  nor (_11332_, _00820_, _21474_);
  nor (_04236_, _11332_, _11331_);
  nor (_11333_, _00818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nor (_11334_, _00820_, _21414_);
  nor (_25452_, _11334_, _11333_);
  nor (_11335_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand (_11336_, _23553_, _23233_);
  nand (_11337_, _11336_, _23493_);
  nor (_04276_, _11337_, _11335_);
  nor (_11338_, _00818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_11339_, _00820_, _21504_);
  nor (_04280_, _11339_, _11338_);
  nor (_11340_, _00818_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5]);
  nor (_11341_, _00820_, _21451_);
  nor (_25453_, _11341_, _11340_);
  nor (_11342_, _22521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  nor (_11343_, _22524_, _21504_);
  nor (_04291_, _11343_, _11342_);
  nor (_11344_, _00812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nor (_11345_, _00814_, _21526_);
  nor (_04313_, _11345_, _11344_);
  nor (_11346_, _00812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nor (_11347_, _00814_, _21554_);
  nor (_04322_, _11347_, _11346_);
  nor (_11348_, _00812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5]);
  nor (_11349_, _00814_, _21451_);
  nor (_04342_, _11349_, _11348_);
  nor (_11350_, _00812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7]);
  nor (_11351_, _00814_, _21626_);
  nor (_04348_, _11351_, _11350_);
  nor (_11352_, _00812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_11353_, _00814_, _21504_);
  nor (_04357_, _11353_, _11352_);
  nor (_11354_, _22465_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  nor (_11355_, _22467_, _21526_);
  nor (_04371_, _11355_, _11354_);
  nor (_11356_, _24706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nor (_11357_, _24708_, _21504_);
  nor (_04399_, _11357_, _11356_);
  nor (_11358_, _24706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7]);
  nor (_11359_, _24708_, _21626_);
  nor (_04407_, _11359_, _11358_);
  not (_11360_, _05231_);
  nand (_11361_, _11360_, ABINPUT[0]);
  nand (_11362_, _05231_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand (_11363_, _11362_, _11361_);
  nor (_11364_, _04981_, _00911_);
  nand (_11365_, _11364_, _00916_);
  not (_11367_, _11365_);
  nor (_11368_, _11367_, _11363_);
  nand (_11369_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand (_11370_, _11369_, _06627_);
  nor (_11371_, _11370_, _11365_);
  nor (_11372_, _11371_, _11368_);
  nor (_11373_, _11372_, _24865_);
  nand (_11374_, _24865_, _00106_);
  nand (_11375_, _11374_, _23493_);
  nor (_04416_, _11375_, _11373_);
  nor (_11376_, _00812_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nor (_11377_, _00814_, _21586_);
  nor (_04430_, _11377_, _11376_);
  nor (_11378_, _24706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1]);
  nor (_11379_, _24708_, _21474_);
  nor (_04443_, _11379_, _11378_);
  nor (_11380_, _24706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nor (_11381_, _24708_, _21586_);
  nor (_04449_, _11381_, _11380_);
  nor (_11382_, _24706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nor (_11383_, _24708_, _21414_);
  nor (_04462_, _11383_, _11382_);
  nor (_11384_, _21829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5]);
  nor (_11385_, _21831_, _21451_);
  nor (_04467_, _11385_, _11384_);
  nor (_11386_, _24706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nor (_11387_, _24708_, _21526_);
  nor (_04471_, _11387_, _11386_);
  nor (_11388_, _24706_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nor (_11389_, _24708_, _21554_);
  nor (_04489_, _11389_, _11388_);
  nor (_11390_, _00732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nor (_11391_, _00734_, _21554_);
  nor (_04496_, _11391_, _11390_);
  nor (_11392_, _00732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nor (_11393_, _00734_, _21414_);
  nor (_04499_, _11393_, _11392_);
  nor (_11394_, _00732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nor (_11395_, _00734_, _21526_);
  nor (_04502_, _11395_, _11394_);
  nor (_11396_, _00732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nor (_11397_, _00734_, _21504_);
  nor (_04512_, _11397_, _11396_);
  nor (_11398_, _00732_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5]);
  nor (_11399_, _00734_, _21451_);
  nor (_25405_, _11399_, _11398_);
  nor (_11400_, _00797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nor (_11401_, _00799_, _21504_);
  nor (_04534_, _11401_, _11400_);
  nor (_11402_, _22521_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5]);
  nor (_11403_, _22524_, _21451_);
  nor (_04537_, _11403_, _11402_);
  nor (_11404_, _21816_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1]);
  nor (_11405_, _21818_, _21474_);
  nor (_04541_, _11405_, _11404_);
  nor (_11406_, _00797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5]);
  nor (_11407_, _00799_, _21451_);
  nor (_04544_, _11407_, _11406_);
  nor (_11408_, _00797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nor (_11409_, _00799_, _21586_);
  nor (_04593_, _11409_, _11408_);
  nor (_11411_, _00797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nor (_11412_, _00799_, _21526_);
  nor (_04612_, _11412_, _11411_);
  nor (_11413_, _00797_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nor (_11414_, _00799_, _21554_);
  nor (_04616_, _11414_, _11413_);
  nor (_11415_, _24710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nor (_11416_, _24712_, _21526_);
  nor (_04629_, _11416_, _11415_);
  nor (_11418_, _24710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nor (_11419_, _24712_, _21554_);
  nor (_04633_, _11419_, _11418_);
  nor (_11420_, _24710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nor (_11421_, _24712_, _21504_);
  nor (_25376_, _11421_, _11420_);
  nor (_11422_, _24710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5]);
  nor (_11423_, _24712_, _21451_);
  nor (_04648_, _11423_, _11422_);
  nor (_11424_, _03976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7]);
  nor (_11425_, _03978_, _21626_);
  nor (_25297_, _11425_, _11424_);
  nor (_11426_, _22021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  nor (_11427_, _22023_, _21554_);
  nor (_04681_, _11427_, _11426_);
  nor (_11428_, _00788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7]);
  nor (_11429_, _00790_, _21626_);
  nor (_04687_, _11429_, _11428_);
  nor (_11430_, _21842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  nor (_11431_, _21844_, _21526_);
  nor (_04693_, _11431_, _11430_);
  nor (_11433_, _21747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7]);
  nor (_11434_, _21749_, _21626_);
  nor (_04697_, _11434_, _11433_);
  nor (_11435_, _24710_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nor (_11436_, _24712_, _21586_);
  nor (_04701_, _11436_, _11435_);
  nor (_11437_, _00788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nor (_11438_, _00790_, _21554_);
  nor (_04719_, _11438_, _11437_);
  nor (_11439_, _00788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1]);
  nor (_11440_, _00790_, _21474_);
  nor (_04721_, _11440_, _11439_);
  nor (_11441_, _00788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nor (_11442_, _00790_, _21586_);
  nor (_04731_, _11442_, _11441_);
  nor (_11443_, _00788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5]);
  nor (_11444_, _00790_, _21451_);
  nor (_04751_, _11444_, _11443_);
  nor (_11445_, _21747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  nor (_11447_, _21749_, _21504_);
  nor (_04753_, _11447_, _11445_);
  nor (_11448_, _00788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nor (_11449_, _00790_, _21414_);
  nor (_25363_, _11449_, _11448_);
  nor (_11450_, _00788_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nor (_11451_, _00790_, _21526_);
  nor (_04758_, _11451_, _11450_);
  nor (_11452_, _22991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  nor (_11453_, _22993_, _21586_);
  nor (_25111_, _11453_, _11452_);
  nor (_11454_, _00764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5]);
  nor (_11455_, _00766_, _21451_);
  nor (_25347_, _11455_, _11454_);
  nor (_11456_, _00764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nor (_11457_, _00766_, _21414_);
  nor (_04794_, _11457_, _11456_);
  nor (_11458_, _00764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nor (_11459_, _00766_, _21504_);
  nor (_04809_, _11459_, _11458_);
  nor (_11461_, _00764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7]);
  nor (_11462_, _00766_, _21626_);
  nor (_04813_, _11462_, _11461_);
  nor (_11463_, _22991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1]);
  nor (_11464_, _22993_, _21474_);
  nor (_04845_, _11464_, _11463_);
  nor (_11465_, _00740_, ABINPUT[3]);
  nor (_11466_, _00742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nor (_04849_, _11466_, _11465_);
  nor (_11467_, _22500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  nor (_11468_, _22502_, _21414_);
  nor (_04865_, _11468_, _11467_);
  nor (_11469_, _21810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5]);
  nor (_11470_, _21812_, _21451_);
  nor (_04932_, _11470_, _11469_);
  nor (_11471_, _22526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  nor (_11472_, _22528_, _21414_);
  nor (_04979_, _11472_, _11471_);
  nor (_11473_, _05519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7]);
  nor (_11474_, _05521_, _21626_);
  nor (_04984_, _11474_, _11473_);
  nor (_11475_, _22396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5]);
  nor (_11476_, _22398_, _21451_);
  nor (_04993_, _11476_, _11475_);
  not (_11477_, _10981_);
  nand (_11478_, _11477_, _23491_);
  nand (_11479_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_11480_, _23516_, _21183_);
  nand (_11481_, _11480_, _11479_);
  nand (_11482_, _11481_, _23493_);
  nand (_25022_[1], _11482_, _11478_);
  nor (_11483_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nand (_11484_, _23553_, _00611_);
  nand (_11485_, _11484_, _23493_);
  nor (_05022_, _11485_, _11483_);
  nor (_11486_, _22526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  nor (_11487_, _22528_, _21526_);
  nor (_05036_, _11487_, _11486_);
  nor (_11488_, _22531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1]);
  nor (_11489_, _22533_, _21474_);
  nor (_05089_, _11489_, _11488_);
  nor (_11490_, _22991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  nor (_11491_, _22993_, _21526_);
  nor (_05106_, _11491_, _11490_);
  nor (_11492_, _00880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1]);
  nor (_11493_, _00882_, _21474_);
  nor (_05139_, _11493_, _11492_);
  nor (_11494_, _01042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_11495_, _01044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_11496_, _11495_, _11494_);
  nor (_11498_, _11496_, _01037_);
  nand (_11499_, _01037_, _00121_);
  nand (_11500_, _11499_, _23493_);
  nor (_05141_, _11500_, _11498_);
  nor (_11501_, _22531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  nor (_11502_, _22533_, _21554_);
  nor (_05149_, _11502_, _11501_);
  not (_11503_, _24907_);
  not (_11504_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand (_11505_, _04980_, _00918_);
  nor (_11506_, _11505_, _00020_);
  nor (_11507_, _11506_, _11504_);
  nor (_11508_, _11365_, _05140_);
  nor (_11509_, _11508_, _11507_);
  nor (_11510_, _11509_, _11503_);
  nor (_11511_, _24907_, _00006_);
  nor (_11512_, _11511_, _11510_);
  nor (_05155_, _11512_, rst);
  nand (_11513_, ABINPUT[2], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_11514_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_11516_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _11514_);
  nand (_11517_, _11516_, _11513_);
  nor (_11518_, _11517_, _11367_);
  nand (_11519_, _01027_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand (_11520_, _11519_, _02493_);
  nor (_11521_, _11520_, _11365_);
  nor (_11522_, _11521_, _11518_);
  nor (_11523_, _11522_, _24865_);
  nand (_11524_, _24865_, _00121_);
  nand (_11525_, _11524_, _23493_);
  nor (_05157_, _11525_, _11523_);
  nor (_11526_, _11505_, _01001_);
  nor (_11527_, _11526_, _24898_);
  nor (_11528_, _11365_, _10873_);
  nor (_11529_, _11528_, _11527_);
  nor (_11530_, _11529_, _24865_);
  nor (_11531_, _11530_, _24908_);
  nor (_05163_, _11531_, rst);
  not (_11532_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor (_11533_, _11505_, _01010_);
  nor (_11534_, _11533_, _11532_);
  nor (_11535_, _11365_, _10858_);
  nor (_11536_, _11535_, _11534_);
  nor (_11537_, _11536_, _11503_);
  nor (_11538_, _24907_, _00129_);
  nor (_11539_, _11538_, _11537_);
  nor (_05165_, _11539_, rst);
  nor (_11540_, _11505_, _00909_);
  nor (_11541_, _11540_, _24847_);
  nor (_11542_, _11365_, _10828_);
  nor (_11543_, _11542_, _11541_);
  nor (_11544_, _11543_, _24865_);
  nor (_11545_, _11544_, _24869_);
  nor (_05167_, _11545_, rst);
  nand (_11546_, _24865_, _00114_);
  nand (_11547_, _11546_, _23493_);
  nand (_11548_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not (_11549_, _11548_);
  nand (_11550_, _11549_, ABINPUT[1]);
  nand (_11551_, _11548_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_11552_, _11551_, _11550_);
  nand (_11553_, _11552_, _11365_);
  nand (_11554_, _05055_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_11555_, _11554_, _05125_);
  nand (_11556_, _11555_, _11367_);
  nand (_11557_, _11556_, _11553_);
  nor (_11558_, _11557_, _24865_);
  nor (_05172_, _11558_, _11547_);
  nor (_11559_, _03976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  nor (_11560_, _03978_, _21554_);
  nor (_05196_, _11560_, _11559_);
  nor (_11561_, _03976_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1]);
  nor (_11562_, _03978_, _21474_);
  nor (_05207_, _11562_, _11561_);
  nor (_11563_, _21865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  nor (_11564_, _21867_, _21414_);
  nor (_05214_, _11564_, _11563_);
  nor (_11565_, _21864_, _21645_);
  nor (_11566_, _11565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  not (_11567_, _11565_);
  nor (_11568_, _11567_, _21554_);
  nor (_05268_, _11568_, _11566_);
  nor (_11569_, _00667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nor (_11570_, _00669_, _21504_);
  nor (_05316_, _11570_, _11569_);
  nor (_11571_, _00667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5]);
  nor (_11572_, _00669_, _21451_);
  nor (_05319_, _11572_, _11571_);
  nor (_11573_, _01042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_11574_, _01044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_11575_, _11574_, _11573_);
  nor (_11576_, _11575_, _01037_);
  nand (_11577_, _01037_, _00114_);
  nand (_11578_, _11577_, _23493_);
  nor (_05325_, _11578_, _11576_);
  nor (_11579_, _11565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  nor (_11580_, _11567_, _21586_);
  nor (_25276_, _11580_, _11579_);
  nor (_11581_, _00667_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nor (_11582_, _00669_, _21554_);
  nor (_05339_, _11582_, _11581_);
  nor (_11584_, _00740_, ABINPUT[10]);
  nor (_11585_, _00742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7]);
  nor (_05352_, _11585_, _11584_);
  not (_11586_, ABINPUT[18]);
  nor (_11587_, _05229_, _11586_);
  not (_11588_, ABINPUT[26]);
  nor (_11589_, _21337_, _24897_);
  nand (_11590_, _11589_, _21426_);
  nor (_11591_, _11590_, _24903_);
  nand (_11592_, _11591_, _24861_);
  nand (_11593_, _11592_, _05289_);
  not (_11594_, _11593_);
  nor (_11595_, _11594_, _11588_);
  not (_11596_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_11597_, _21365_, _21337_);
  not (_11598_, _11597_);
  nor (_11599_, _11598_, _00917_);
  nand (_11600_, _11599_, _05112_);
  nor (_11601_, _11600_, _05559_);
  nor (_11603_, _11601_, _11596_);
  nor (_11604_, _11600_, _06627_);
  nor (_11605_, _11604_, _11603_);
  nor (_11606_, _11605_, _11593_);
  nor (_11607_, _11606_, _11595_);
  nor (_11608_, _11607_, _05228_);
  nor (_11609_, _11608_, _11587_);
  nor (_05354_, _11609_, rst);
  nor (_11610_, _00740_, ABINPUT[6]);
  nor (_11611_, _00742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nor (_05396_, _11611_, _11610_);
  nor (_11612_, _21913_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1]);
  nor (_11613_, _21915_, _21474_);
  nor (_05399_, _11613_, _11612_);
  nor (_11614_, _00740_, ABINPUT[8]);
  nor (_11615_, _00742_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5]);
  nor (_05402_, _11615_, _11614_);
  nor (_11616_, _22479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1]);
  nor (_11617_, _22482_, _21474_);
  nor (_05414_, _11617_, _11616_);
  nor (_11618_, _01042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor (_11619_, _01044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_11620_, _11619_, _11618_);
  nor (_11621_, _11620_, _01037_);
  nand (_11622_, _01037_, _00129_);
  nand (_11623_, _11622_, _23493_);
  nor (_05416_, _11623_, _11621_);
  nor (_11624_, _00764_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1]);
  nor (_11625_, _00766_, _21474_);
  nor (_05417_, _11625_, _11624_);
  nor (_11626_, _21850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  nor (_11627_, _21853_, _21526_);
  nor (_05421_, _11627_, _11626_);
  nor (_11628_, _21850_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  nor (_11629_, _21853_, _21414_);
  nor (_05423_, _11629_, _11628_);
  nor (_11630_, _24601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  nor (_11631_, _24603_, _21526_);
  nor (_25340_, _11631_, _11630_);
  nor (_11632_, _21810_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1]);
  nor (_11633_, _21812_, _21474_);
  nor (_05426_, _11633_, _11632_);
  nor (_11634_, _24601_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  nor (_11635_, _24603_, _21586_);
  nor (_05429_, _11635_, _11634_);
  nor (_11636_, _01042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_11637_, _01044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_11638_, _11637_, _11636_);
  nor (_11639_, _11638_, _01037_);
  nand (_11640_, _01037_, _24900_);
  nand (_11641_, _11640_, _23493_);
  nor (_05433_, _11641_, _11639_);
  nor (_11642_, _22567_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1]);
  nor (_11643_, _22569_, _21474_);
  nor (_25057_, _11643_, _11642_);
  nor (_11644_, _22484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  nor (_11645_, _22486_, _21504_);
  nor (_05444_, _11645_, _11644_);
  nor (_11646_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  nor (_11647_, _22498_, _21586_);
  nor (_05491_, _11647_, _11646_);
  nor (_11648_, _11593_, _05228_);
  not (_11649_, _11648_);
  not (_11650_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_11651_, _11600_, _24858_);
  nor (_11652_, _11651_, _11650_);
  nor (_11653_, _11600_, _10800_);
  nor (_11654_, _11653_, _11652_);
  nor (_11655_, _11654_, _11649_);
  not (_11656_, ABINPUT[11]);
  nor (_11657_, _05229_, _11656_);
  not (_11658_, ABINPUT[19]);
  nor (_11659_, _05228_, _11658_);
  nand (_11660_, _11659_, _11593_);
  not (_11661_, _11660_);
  nor (_11662_, _11661_, _11657_);
  not (_11663_, _11662_);
  nor (_11664_, _11663_, _11655_);
  nor (_05494_, _11664_, rst);
  nor (_05495_, _00556_, rst);
  nand (_11666_, _05228_, ABINPUT[12]);
  not (_11667_, _11666_);
  nor (_11668_, _11594_, _10818_);
  not (_11669_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_11670_, _11598_, _05113_);
  not (_11671_, _11670_);
  nor (_11672_, _11671_, _00917_);
  not (_11673_, _11672_);
  nor (_11674_, _11649_, _11673_);
  not (_11675_, _11674_);
  nor (_11676_, _11675_, _00011_);
  nor (_11677_, _11676_, _11673_);
  nor (_11678_, _11677_, _11669_);
  nor (_11679_, _11675_, _05140_);
  nor (_11680_, _11679_, _11678_);
  nor (_11681_, _11680_, _11593_);
  nor (_11682_, _11681_, _11668_);
  nor (_11683_, _11682_, _05228_);
  nor (_11684_, _11683_, _11667_);
  nor (_05510_, _11684_, rst);
  not (_11685_, ABINPUT[14]);
  nor (_11686_, _05229_, _11685_);
  not (_11687_, _11600_);
  nand (_11688_, _11687_, _00931_);
  not (_11689_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_11690_, _11600_, _00909_);
  nor (_11691_, _11690_, _11689_);
  nor (_11692_, _11691_, _11593_);
  nand (_11693_, _11692_, _11688_);
  nand (_11694_, _11593_, _10833_);
  nand (_11695_, _11694_, _11693_);
  nor (_11696_, _11695_, _05228_);
  nor (_11697_, _11696_, _11686_);
  nor (_05514_, _11697_, rst);
  nand (_11698_, _05228_, ABINPUT[13]);
  not (_11699_, _11698_);
  nor (_11700_, _11594_, _10847_);
  not (_11701_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_11702_, _11600_, _01027_);
  nor (_11703_, _11702_, _11701_);
  nor (_11704_, _11600_, _02493_);
  nor (_11705_, _11704_, _11703_);
  nor (_11706_, _11705_, _11593_);
  nor (_11707_, _11706_, _11700_);
  nor (_11708_, _11707_, _05228_);
  nor (_11709_, _11708_, _11699_);
  nor (_05515_, _11709_, rst);
  nor (_11710_, _05519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  nor (_11711_, _05521_, _21526_);
  nor (_25295_, _11711_, _11710_);
  not (_11712_, ABINPUT[15]);
  nor (_11713_, _05229_, _11712_);
  nor (_11714_, _11594_, _10878_);
  not (_11715_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_11716_, _11687_, _11715_);
  nor (_11717_, _01000_, _11715_);
  nor (_11718_, _11717_, _01093_);
  nor (_11719_, _11718_, _11675_);
  nor (_11720_, _11719_, _11716_);
  nor (_11721_, _11720_, _11593_);
  nor (_11722_, _11721_, _11714_);
  nor (_11723_, _11722_, _05228_);
  nor (_11724_, _11723_, _11713_);
  nor (_05518_, _11724_, rst);
  not (_11725_, ABINPUT[17]);
  nor (_11726_, _05229_, _11725_);
  nor (_11727_, _05228_, _10899_);
  nand (_11728_, _11727_, _11593_);
  not (_11729_, _11728_);
  nor (_11730_, _11729_, _11726_);
  not (_11731_, _11730_);
  not (_11732_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_11733_, _11600_, _05055_);
  nor (_11734_, _11733_, _11732_);
  nor (_11735_, _11600_, _05125_);
  nor (_11736_, _11735_, _11734_);
  nor (_11737_, _11736_, _11649_);
  nor (_11738_, _11737_, _11731_);
  nor (_05523_, _11738_, rst);
  nor (_11739_, _05229_, ABINPUT[16]);
  nor (_11741_, _11675_, _10858_);
  not (_11742_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_11743_, _11600_, _01010_);
  nor (_11744_, _11743_, _11742_);
  nand (_11745_, _11744_, _11648_);
  nand (_11746_, _05229_, _10863_);
  nand (_11747_, _11746_, _11649_);
  nand (_11748_, _11747_, _11745_);
  nor (_11749_, _11748_, _11741_);
  nor (_11750_, _11749_, _11739_);
  not (_11751_, _11750_);
  nor (_05525_, _11751_, rst);
  nor (_05527_, _24909_, rst);
  nor (_05538_, _00103_, rst);
  nor (_05552_, _00073_, rst);
  nor (_11752_, _23044_, _21210_);
  not (_11753_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  nor (_11754_, _11753_, _23153_);
  nor (_11755_, _23058_, _23385_);
  nor (_11756_, _23067_, _00057_);
  nor (_11758_, _11756_, _11755_);
  nor (_11759_, _23050_, _00062_);
  nor (_11760_, _23107_, _23388_);
  nor (_11761_, _11760_, _11759_);
  nand (_11762_, _11761_, _11758_);
  not (_11763_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nor (_11764_, _23073_, _11763_);
  nor (_11765_, _23076_, _23391_);
  nor (_11766_, _11765_, _11764_);
  not (_11767_, _11766_);
  nor (_11768_, _11767_, _11762_);
  nor (_11769_, _11768_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11770_, _11769_, _11754_);
  nor (_11771_, _11770_, _23490_);
  nor (_11772_, _11771_, _11752_);
  nor (_05570_, _11772_, rst);
  nor (_11773_, _24497_, _23510_);
  not (_11774_, _11773_);
  nor (_11775_, _05558_, _00010_);
  not (_11776_, _11775_);
  nor (_11777_, _11776_, _05296_);
  not (_11778_, _11777_);
  nor (_11779_, _11778_, _11774_);
  not (_11780_, _11779_);
  nor (_11781_, _23407_, _23330_);
  not (_11782_, _11781_);
  nand (_11783_, _11782_, _23472_);
  nand (_11784_, _24386_, _11783_);
  not (_11785_, _11784_);
  nand (_11786_, _24515_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_11787_, _21403_, _21396_);
  nor (_11788_, _21546_, _21544_);
  nor (_11789_, _11788_, _11787_);
  nor (_11790_, _21496_, _21490_);
  nor (_11791_, _21583_, _21578_);
  nor (_11792_, _11791_, _11790_);
  nand (_11793_, _11792_, _11789_);
  nor (_11794_, _21442_, _21437_);
  nor (_11795_, _21461_, _21458_);
  nor (_11796_, _11795_, _11794_);
  not (_11798_, _11796_);
  nor (_11799_, _11798_, _11793_);
  not (_11800_, _11799_);
  not (_11801_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  nor (_11802_, _11801_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  not (_11803_, _11802_);
  nor (_11804_, _21616_, _21614_);
  nand (_11805_, _21519_, _21515_);
  not (_11806_, _11805_);
  nor (_11807_, _11806_, _11804_);
  nand (_11808_, _11807_, _11803_);
  nor (_11809_, _11808_, _11800_);
  nor (_11810_, _11803_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_11811_, _11810_, _11809_);
  nand (_11812_, _11811_, _11773_);
  not (_11813_, _11812_);
  nor (_11814_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_11815_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand (_11816_, _11815_, _11814_);
  nor (_11817_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_11818_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nand (_11819_, _11818_, _11817_);
  nor (_11820_, _11819_, _11816_);
  nand (_11821_, _11820_, _24429_);
  not (_11822_, _24516_);
  nor (_11823_, ABINPUT[32], ABINPUT[31]);
  nor (_11824_, ABINPUT[34], ABINPUT[33]);
  nand (_11825_, _11824_, _11823_);
  nor (_11826_, ABINPUT[28], ABINPUT[27]);
  nor (_11827_, ABINPUT[30], ABINPUT[29]);
  nand (_11829_, _11827_, _11826_);
  nor (_11830_, _11829_, _11825_);
  not (_11831_, _11830_);
  nor (_11832_, _11831_, _11822_);
  nand (_11833_, _11832_, _11774_);
  nand (_11834_, _11833_, _11821_);
  nor (_11835_, _11834_, _11813_);
  nand (_11836_, _11835_, _11786_);
  not (_11837_, _11836_);
  not (_11838_, _24737_);
  nor (_11839_, _11838_, _24495_);
  not (_11840_, _11839_);
  not (_11841_, _24428_);
  nor (_11842_, _24513_, _11841_);
  nor (_11843_, _11842_, _23283_);
  nor (_11844_, _11843_, _11840_);
  nor (_11845_, _11844_, _11837_);
  nor (_11846_, _24468_, _23382_);
  not (_11847_, _11846_);
  nand (_11848_, _10992_, _11847_);
  nor (_11849_, _24468_, _23203_);
  not (_11850_, _11849_);
  not (_11851_, _24463_);
  nor (_11852_, _11851_, _23449_);
  nand (_11853_, _11852_, _24715_);
  nand (_11854_, _11853_, _23431_);
  nand (_11855_, _11854_, _11850_);
  nor (_11856_, _11855_, _11848_);
  nor (_11857_, _11856_, _11836_);
  nor (_11858_, _24397_, _23464_);
  nor (_11859_, _11858_, _24788_);
  nand (_11860_, _11859_, _24510_);
  nor (_11861_, _11860_, _11857_);
  not (_11862_, _11861_);
  nor (_11863_, _11862_, _11845_);
  nor (_11864_, _24511_, _23499_);
  nor (_11865_, _11864_, _11863_);
  nor (_11866_, _11865_, _11785_);
  nor (_11867_, _11649_, _11672_);
  nor (_11868_, _11867_, _24786_);
  nor (_11870_, _11367_, _11360_);
  nand (_11871_, _11870_, _24868_);
  nand (_11872_, _11871_, _24515_);
  not (_11873_, _11872_);
  nor (_11874_, _11873_, _11868_);
  not (_11875_, _11874_);
  nor (_11876_, _11875_, _11866_);
  not (_11877_, _11876_);
  nor (_11878_, _11877_, _05286_);
  nand (_11879_, _11878_, _11780_);
  nand (_11880_, _24512_, _23493_);
  nor (_05576_, _11880_, _11879_);
  nor (_11881_, _22219_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  nor (_11882_, _22221_, _21526_);
  nor (_05613_, _11882_, _11881_);
  nor (_11883_, _05519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  nor (_11884_, _05521_, _21554_);
  nor (_05621_, _11884_, _11883_);
  nor (_11885_, _22531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  nor (_11886_, _22533_, _21526_);
  nor (_25116_, _11886_, _11885_);
  nor (_11887_, _21899_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7]);
  nor (_11888_, _21902_, _21626_);
  nor (_25125_, _11888_, _11887_);
  nor (_11889_, _01083_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  nor (_11890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _01052_);
  nand (_11891_, _11890_, _01080_);
  nand (_11892_, _11891_, _23493_);
  nor (_05643_, _11892_, _11889_);
  nor (_11893_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand (_11894_, _23553_, _23388_);
  nand (_11895_, _11894_, _23493_);
  nor (_05685_, _11895_, _11893_);
  not (_11896_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r );
  nor (_05689_, _11896_, rst);
  nor (_11897_, _05519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5]);
  nor (_11898_, _05521_, _21451_);
  nor (_05692_, _11898_, _11897_);
  nor (_11899_, _06971_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  nor (_11900_, _06973_, _21526_);
  nor (_05695_, _11900_, _11899_);
  nor (_11901_, _07226_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5]);
  nor (_11902_, _07228_, _21451_);
  nor (_05697_, _11902_, _11901_);
  not (_11903_, _11879_);
  nor (_11904_, _24460_, _11782_);
  nand (_11905_, _11904_, _00074_);
  nand (_11906_, _24788_, _23499_);
  nor (_11907_, _11906_, _11586_);
  nor (_11908_, _24512_, _11588_);
  nor (_11910_, _11908_, _11907_);
  nand (_11911_, _11910_, _11905_);
  nor (_11912_, _11848_, _24766_);
  not (_11913_, _11859_);
  nand (_11914_, _11842_, _11850_);
  nor (_11915_, _11914_, _11913_);
  nand (_11916_, _11915_, _11912_);
  nand (_11917_, _11916_, _23499_);
  not (_11918_, _11917_);
  nor (_11919_, _10993_, _11846_);
  nand (_11920_, _11919_, _24497_);
  nand (_11921_, _11920_, _23499_);
  nor (_11922_, _24765_, _24460_);
  nor (_11923_, _11922_, _11904_);
  nand (_11924_, _11923_, _24512_);
  not (_11925_, _11924_);
  nand (_11926_, _11925_, _11921_);
  nor (_11927_, _23528_, _24724_);
  nand (_11928_, _11927_, _23499_);
  not (_11929_, _11928_);
  nor (_11931_, _11929_, _11785_);
  nor (_11932_, _11931_, _11926_);
  not (_11933_, _11932_);
  nor (_11934_, _11933_, _11918_);
  nand (_11935_, _11934_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_11936_, _11931_);
  nor (_11937_, _11912_, _23500_);
  nor (_11938_, _11924_, _11937_);
  nor (_11939_, _24716_, _11838_);
  nor (_11940_, _11939_, _24460_);
  nor (_11941_, _11940_, _11918_);
  nand (_11942_, _11941_, _11938_);
  nor (_11943_, _11942_, _11936_);
  nand (_11944_, _11943_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nand (_11945_, _11944_, _11935_);
  nor (_11946_, _11945_, _11911_);
  nand (_11947_, _11946_, _11903_);
  not (_11948_, _11772_);
  nor (_11949_, _11938_, _11948_);
  nor (_11950_, _11926_, _00074_);
  nor (_11951_, _11950_, _11949_);
  nor (_11952_, _11951_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_11953_, _11952_);
  not (_11954_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_11955_, _02307_);
  nor (_11956_, _11938_, _11955_);
  not (_11957_, _00380_);
  nor (_11958_, _11926_, _11957_);
  nor (_11959_, _11958_, _11956_);
  not (_11960_, _11959_);
  nor (_11961_, _11960_, _11954_);
  nor (_11962_, _11959_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_11963_, _11962_, _11961_);
  not (_11964_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_11965_, _01352_);
  nor (_11966_, _11938_, _11965_);
  not (_11967_, _00301_);
  nor (_11968_, _11926_, _11967_);
  nor (_11969_, _11968_, _11966_);
  not (_11970_, _11969_);
  nor (_11972_, _11970_, _11964_);
  not (_11973_, _11972_);
  nor (_11974_, _11969_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_11975_, _11974_);
  not (_11976_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_11977_, _24191_);
  nor (_11978_, _11938_, _11977_);
  not (_11979_, _00175_);
  nor (_11980_, _11926_, _11979_);
  nor (_11981_, _11980_, _11978_);
  not (_11982_, _11981_);
  nor (_11983_, _11982_, _11976_);
  not (_11984_, _11983_);
  not (_11985_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_11986_, _11926_, _10398_);
  not (_11987_, _11986_);
  nor (_11988_, _11926_, _00456_);
  nor (_11989_, _11988_, _11987_);
  not (_11990_, _11989_);
  nor (_11991_, _11990_, _11985_);
  not (_11992_, _11991_);
  nor (_11993_, _11989_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_11994_, _11993_);
  not (_11995_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_11996_, _07031_);
  nor (_11997_, _11938_, _11996_);
  not (_11998_, _00517_);
  nor (_11999_, _11926_, _11998_);
  nor (_12000_, _11999_, _11997_);
  not (_12001_, _12000_);
  nor (_12002_, _12001_, _11995_);
  not (_12003_, _12002_);
  not (_12004_, _05381_);
  nor (_12005_, _11938_, _12004_);
  not (_12006_, _24841_);
  nor (_12007_, _11926_, _12006_);
  nor (_12008_, _12007_, _12005_);
  nand (_12009_, _12008_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_12010_, _23490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  not (_12011_, _12010_);
  not (_12013_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  nor (_12014_, _23153_, _12013_);
  nor (_12015_, _23058_, _00611_);
  nor (_12016_, _23067_, _00601_);
  nor (_12017_, _12016_, _12015_);
  nor (_12018_, _23050_, _00605_);
  nor (_12019_, _23107_, _00599_);
  nor (_12020_, _12019_, _12018_);
  nand (_12021_, _12020_, _12017_);
  nor (_12022_, _23073_, _05179_);
  nor (_12023_, _23076_, _00607_);
  nor (_12024_, _12023_, _12022_);
  not (_12025_, _12024_);
  nor (_12026_, _12025_, _12021_);
  nor (_12027_, _12026_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12028_, _12027_, _12014_);
  nor (_12029_, _12028_, _23490_);
  nor (_12030_, _12029_, _12011_);
  not (_12031_, _12030_);
  nor (_12032_, _12031_, _11938_);
  nor (_12034_, _11926_, _00620_);
  nor (_12035_, _12034_, _12032_);
  nand (_12036_, _12035_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_12037_, _12036_);
  not (_12038_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_12039_, _11926_, _05381_);
  nand (_12040_, _11938_, _24841_);
  nand (_12041_, _12040_, _12039_);
  nor (_12042_, _12041_, _12038_);
  nor (_12043_, _12008_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_12044_, _12043_, _12042_);
  nand (_12045_, _12044_, _12037_);
  nand (_12046_, _12045_, _12009_);
  nor (_12047_, _12000_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_12048_, _12047_, _12002_);
  nand (_12049_, _12048_, _12046_);
  nand (_12050_, _12049_, _12003_);
  nand (_12051_, _12050_, _11994_);
  nand (_12052_, _12051_, _11992_);
  nor (_12053_, _11981_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_12055_, _12053_, _11983_);
  nand (_12056_, _12055_, _12052_);
  nand (_12057_, _12056_, _11984_);
  nand (_12058_, _12057_, _11975_);
  nand (_12059_, _12058_, _11973_);
  nand (_12060_, _12059_, _11963_);
  not (_12061_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  not (_12062_, _11951_);
  nor (_12063_, _12062_, _12061_);
  nor (_12064_, _12063_, _11961_);
  nand (_12065_, _12064_, _12060_);
  nand (_12066_, _12065_, _11953_);
  nand (_12067_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_12068_, _12067_, _12066_);
  nand (_12069_, _12068_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_12070_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_12071_, _11951_, _12070_);
  not (_12072_, _12071_);
  nor (_12073_, _12072_, _12069_);
  nand (_12074_, _12073_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_12076_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nand (_12077_, _12066_, _12076_);
  not (_12078_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  not (_12079_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand (_12080_, _12079_, _12078_);
  nor (_12081_, _12080_, _12077_);
  nor (_12082_, _12062_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand (_12083_, _12082_, _12081_);
  nor (_12084_, _12083_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  not (_12085_, _12084_);
  nand (_12086_, _12085_, _12074_);
  nor (_12087_, _11951_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_12088_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_12089_, _12062_, _12088_);
  nor (_12090_, _12089_, _12087_);
  nand (_12091_, _12090_, _12086_);
  not (_12092_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_12093_, _12062_, _12092_);
  nand (_12094_, _11951_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_12095_, _12094_, _12093_);
  nor (_12097_, _12095_, _12091_);
  nor (_12098_, _12097_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_12099_, _12097_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_12100_, _11922_, _11918_);
  nor (_12101_, _12100_, _11932_);
  nand (_12102_, _12101_, _12099_);
  nor (_12103_, _12102_, _12098_);
  nor (_12104_, _12103_, _11947_);
  not (_12105_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_12106_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_12107_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_12108_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_12109_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_12110_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_12111_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_12112_, _06002_, _12111_);
  not (_12113_, _12112_);
  nor (_12114_, _12113_, _06003_);
  nand (_12115_, _12114_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_12116_, _12115_, _12110_);
  nand (_12118_, _12116_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_12119_, _12118_, _12109_);
  nand (_12120_, _12119_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_12121_, _12120_, _12108_);
  nand (_12122_, _12121_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_12123_, _12122_, _12107_);
  nand (_12124_, _12123_, _06015_);
  nor (_12125_, _12124_, _12106_);
  not (_12126_, _12125_);
  nor (_12127_, _12126_, _12105_);
  nand (_12128_, _12127_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_12129_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_12130_, _12127_);
  nand (_12131_, _12130_, _12129_);
  nand (_12132_, _12131_, _12128_);
  nand (_12133_, _12132_, _11879_);
  nand (_12134_, _12133_, _23493_);
  nor (_05750_, _12134_, _12104_);
  nor (_12135_, _23038_, rst);
  nand (_12136_, _12135_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_12137_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_12138_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  not (_12139_, _12138_);
  nor (_12140_, _12139_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  not (_12141_, _12140_);
  nor (_12142_, _12141_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_12143_, _12142_);
  nor (_12144_, _12143_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_12145_, _12144_);
  nor (_12146_, _12145_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_12148_, _12146_);
  nor (_12149_, _12148_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_12150_, _12149_);
  nor (_12151_, _12150_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_12152_, _12151_);
  nor (_12153_, _12152_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_12154_, _06003_, _23054_);
  not (_12155_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_12156_, _12155_, _23056_);
  not (_12157_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nor (_12158_, _12157_, _23055_);
  not (_12159_, _12158_);
  nor (_12160_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_12161_, _12160_, _12156_);
  not (_12162_, _12161_);
  nor (_12163_, _12162_, _12159_);
  nor (_12164_, _12163_, _12156_);
  nor (_12165_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_12166_, _12165_, _12154_);
  not (_12167_, _12166_);
  nor (_12169_, _12167_, _12164_);
  nor (_12170_, _12169_, _12154_);
  nand (_12171_, _12170_, _12153_);
  not (_12172_, _12171_);
  nand (_12173_, _12172_, _12137_);
  nor (_12174_, _12173_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_12175_, _12174_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_12176_, _12174_);
  nor (_12177_, _12176_, _12129_);
  nor (_12178_, _12177_, _12175_);
  nand (_12179_, _12173_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_12180_, _12179_, _12176_);
  not (_12181_, _12180_);
  nor (_12182_, _12171_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_12183_, _12182_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_12184_, _12182_);
  nor (_12185_, _12184_, _12106_);
  nor (_12186_, _12185_, _12183_);
  nor (_12187_, _12172_, _12107_);
  nor (_12188_, _12187_, _12182_);
  not (_12189_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_12190_, _12170_);
  nor (_12191_, _12190_, _12152_);
  nor (_12192_, _12191_, _12189_);
  nor (_12193_, _12192_, _12172_);
  not (_12194_, _12193_);
  nor (_12195_, _12190_, _12150_);
  nor (_12196_, _12195_, _12108_);
  nor (_12197_, _12196_, _12191_);
  not (_12198_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_12199_, _12190_, _12148_);
  nor (_12200_, _12199_, _12198_);
  nor (_12201_, _12200_, _12195_);
  not (_12202_, _12201_);
  nor (_12203_, _12190_, _12143_);
  nor (_12204_, _12203_, _12110_);
  nor (_12205_, _12190_, _12145_);
  nor (_12206_, _12205_, _12204_);
  not (_12207_, _12206_);
  not (_12208_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_12209_, _12190_, _12141_);
  nor (_12210_, _12209_, _12208_);
  nor (_12211_, _12210_, _12203_);
  not (_12212_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_12213_, _12190_, _12139_);
  nor (_12214_, _12213_, _12212_);
  nor (_12215_, _12214_, _12209_);
  not (_12216_, _12215_);
  nor (_12217_, _07138_, _00687_);
  nor (_12218_, _07110_, _07149_);
  nor (_12219_, _12218_, _12217_);
  nor (_12220_, _12219_, _07135_);
  nor (_12221_, _12218_, _07102_);
  nor (_12222_, _12221_, _00696_);
  nor (_12223_, _12222_, _12220_);
  nor (_12224_, _00696_, _00687_);
  not (_12225_, _12224_);
  nor (_12226_, _12225_, _07098_);
  nor (_12227_, _00706_, _00687_);
  nor (_12228_, _07111_, _12227_);
  nor (_12229_, _12228_, _07119_);
  nor (_12230_, _12229_, _12226_);
  nand (_12231_, _12230_, _12223_);
  nor (_12232_, _07107_, _00715_);
  nor (_12233_, _12232_, _23199_);
  nor (_12234_, _12233_, _07122_);
  nor (_12235_, _07139_, _07107_);
  nor (_12236_, _12235_, _00696_);
  nor (_12237_, _12225_, _07149_);
  nor (_12238_, _12237_, _12236_);
  nand (_12239_, _12238_, _12234_);
  nor (_12240_, _12239_, _12231_);
  not (_12241_, _00714_);
  not (_12242_, _07102_);
  nor (_12243_, _12242_, _12241_);
  nand (_12244_, _07142_, _07100_);
  nor (_12245_, _12244_, _12243_);
  not (_12246_, _12245_);
  nor (_12247_, _12242_, _07135_);
  not (_12248_, _00693_);
  nor (_12249_, _07106_, _07138_);
  not (_12250_, _12249_);
  nor (_12251_, _12250_, _12248_);
  nor (_12252_, _12251_, _12247_);
  not (_12253_, _12252_);
  nor (_12254_, _12253_, _12246_);
  nor (_12255_, _07101_, _00695_);
  nor (_12256_, _12255_, _12250_);
  nor (_12257_, _07107_, _07151_);
  nor (_12258_, _12257_, _07135_);
  nor (_12259_, _12232_, _07166_);
  nor (_12260_, _12259_, _12258_);
  not (_12261_, _12260_);
  nor (_12262_, _12261_, _12256_);
  nand (_12263_, _12262_, _12254_);
  not (_12264_, _12263_);
  nand (_12265_, _12264_, _12240_);
  nor (_12266_, _07101_, _00691_);
  not (_12267_, _07154_);
  nor (_12268_, _12267_, _23348_);
  nor (_12270_, _12268_, _07131_);
  nor (_12271_, _12270_, _12266_);
  nand (_12272_, _07120_, _00688_);
  not (_12273_, _12272_);
  nor (_12274_, _12273_, _07169_);
  nand (_12275_, _07157_, _07093_);
  nand (_12276_, _12275_, _12274_);
  nor (_12277_, _12276_, _12271_);
  nor (_12278_, _12267_, _12248_);
  not (_12279_, _12278_);
  nor (_12280_, _07110_, _00706_);
  nand (_12281_, _07134_, _12280_);
  nand (_12282_, _12281_, _12279_);
  nor (_12283_, _12242_, _07119_);
  not (_12284_, _00703_);
  nor (_12285_, _12241_, _12284_);
  nor (_12286_, _12285_, _12283_);
  not (_12287_, _12286_);
  nor (_12288_, _12287_, _12282_);
  nor (_12289_, _07115_, _07133_);
  nor (_12290_, _07126_, _07162_);
  nand (_12291_, _12290_, _12289_);
  not (_12292_, _12291_);
  nand (_12293_, _12292_, _12288_);
  not (_12294_, _12217_);
  nor (_12295_, _07107_, _00707_);
  nand (_12296_, _12295_, _12294_);
  nand (_12297_, _12296_, _00714_);
  not (_12298_, _12297_);
  nor (_12299_, _07110_, _00699_);
  nor (_12300_, _07154_, _00701_);
  not (_12301_, _12300_);
  nor (_12302_, _12301_, _12299_);
  nor (_12303_, _12302_, _07135_);
  nor (_12304_, _12303_, _12298_);
  not (_12305_, _12304_);
  nor (_12306_, _12305_, _12293_);
  nand (_12307_, _12306_, _12277_);
  nor (_12308_, _12307_, _12265_);
  nor (_12309_, _12161_, _12158_);
  nor (_12310_, _12309_, _12163_);
  not (_12311_, _12310_);
  nor (_12312_, _12311_, _12308_);
  not (_12313_, _12312_);
  nor (_12314_, _12258_, _07171_);
  nand (_12315_, _12314_, _12252_);
  nor (_12316_, _07119_, _12284_);
  nor (_12317_, _07132_, _12248_);
  nor (_12318_, _12317_, _12316_);
  nor (_12319_, _07119_, _12294_);
  nor (_12320_, _12319_, _12278_);
  nand (_12321_, _12320_, _12318_);
  nor (_12322_, _12321_, _12246_);
  not (_12323_, _12322_);
  nor (_12324_, _12323_, _12315_);
  not (_12325_, _12324_);
  nor (_12326_, _12325_, _12308_);
  nor (_12327_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_12328_, _12327_, _12158_);
  not (_12329_, _12328_);
  nor (_12330_, _12329_, _12326_);
  nand (_12331_, _12311_, _12308_);
  nand (_12332_, _12331_, _12313_);
  not (_12333_, _12332_);
  nand (_12334_, _12333_, _12330_);
  nand (_12335_, _12334_, _12313_);
  nor (_12336_, _12170_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_12337_, _12190_, _06002_);
  nor (_12338_, _12337_, _12336_);
  not (_12339_, _12338_);
  nand (_12341_, _12167_, _12164_);
  not (_12342_, _12341_);
  nor (_12343_, _12342_, _12169_);
  not (_12344_, _12343_);
  nor (_12345_, _12344_, _12339_);
  nand (_12346_, _12345_, _12335_);
  nor (_12347_, _12170_, _12139_);
  nor (_12348_, _12138_, _12112_);
  not (_12349_, _12348_);
  nor (_12350_, _12349_, _12336_);
  nor (_12351_, _12350_, _12347_);
  not (_12352_, _12351_);
  nor (_12353_, _12352_, _12346_);
  nand (_12354_, _12353_, _12216_);
  nor (_12355_, _12354_, _12211_);
  nand (_12356_, _12355_, _12207_);
  nor (_12357_, _12205_, _12109_);
  nor (_12358_, _12357_, _12199_);
  nor (_12359_, _12358_, _12356_);
  nand (_12360_, _12359_, _12202_);
  nor (_12361_, _12360_, _12197_);
  nand (_12362_, _12361_, _12194_);
  nor (_12363_, _12362_, _12188_);
  nand (_12364_, _12363_, _12186_);
  nor (_12365_, _12364_, _12181_);
  not (_12366_, _12365_);
  nand (_12367_, _12366_, _12178_);
  nor (_12368_, _12366_, _12178_);
  nor (_12369_, _12368_, _24824_);
  nand (_12370_, _12369_, _12367_);
  nor (_12371_, _24823_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_12372_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  not (_12373_, _12372_);
  nor (_12374_, _12373_, _12371_);
  nand (_12375_, _12374_, _12370_);
  nand (_05752_, _12375_, _12136_);
  nand (_12376_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _23153_);
  nor (_05757_, _12376_, rst);
  nor (_25035_, _23153_, rst);
  not (_12377_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor (_12379_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nand (_12380_, _12379_, _12377_);
  nor (_12381_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  nor (_12382_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nand (_12383_, _12382_, _12381_);
  nor (_12384_, _12383_, _12380_);
  not (_12385_, _12384_);
  nor (_12386_, _12385_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  not (_12387_, _12386_);
  nor (_12388_, _23490_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_12389_, _12388_, _23153_);
  nor (_12390_, _12389_, _12387_);
  nor (_05759_, _12390_, rst);
  nor (_12391_, _12385_, _11753_);
  nor (_12392_, _12391_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_05761_, _12392_, rst);
  nand (_12393_, _01017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nand (_12394_, _01020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand (_12395_, _12394_, _12393_);
  nor (_12396_, _12395_, _01030_);
  nor (_12397_, _01032_, ABINPUT[5]);
  nor (_12398_, _12397_, _12396_);
  nor (_12399_, _12398_, _01037_);
  nand (_12400_, _01037_, _01264_);
  nand (_12401_, _12400_, _23493_);
  nor (_05763_, _12401_, _12399_);
  nor (_12402_, _23553_, _23490_);
  nor (_12403_, _12308_, _23056_);
  nor (_12404_, _12326_, _23055_);
  not (_12405_, _12403_);
  nand (_12406_, _12308_, _23056_);
  nand (_12407_, _12406_, _12405_);
  not (_12408_, _12407_);
  nand (_12409_, _12408_, _12404_);
  not (_12410_, _12409_);
  nor (_12411_, _12410_, _12403_);
  nor (_12412_, _12411_, _23490_);
  not (_12413_, _12412_);
  nor (_12414_, _12413_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_12415_, _12412_, _23054_);
  nor (_12416_, _12415_, _12414_);
  nor (_12417_, _12416_, _12402_);
  nand (_12418_, _12402_, _23066_);
  nor (_12419_, _12418_, _12324_);
  nand (_12420_, _12419_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_12421_, _12420_, _23038_);
  nor (_12422_, _12421_, _12417_);
  nor (_05769_, _12422_, rst);
  nor (_12423_, _05519_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  nor (_12424_, _05521_, _21414_);
  nor (_05776_, _12424_, _12423_);
  nand (_12425_, _01017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand (_12426_, _01020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nand (_12427_, _12426_, _12425_);
  nor (_12428_, _12427_, _01030_);
  nor (_12429_, _01032_, ABINPUT[4]);
  nor (_12430_, _12429_, _12428_);
  nor (_12431_, _12430_, _01037_);
  nand (_12432_, _01037_, _11278_);
  nand (_12433_, _12432_, _23493_);
  nor (_05778_, _12433_, _12431_);
  nor (_12434_, _23273_, _23167_);
  nand (_12435_, _12434_, _23221_);
  nand (_12436_, _23041_, _23153_);
  nor (_12437_, _12436_, _10520_);
  nand (_12438_, _12437_, _23194_);
  not (_12439_, _23080_);
  nand (_12440_, _23137_, _12439_);
  nor (_12441_, _12440_, _12438_);
  nor (_12442_, _23397_, _23112_);
  nand (_12443_, _12442_, _12441_);
  nor (_05780_, _12443_, _12435_);
  nor (_12444_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_12445_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand (_12446_, _12445_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand (_12447_, _12446_, _23493_);
  nor (_05782_, _12447_, _12444_);
  nor (_05783_, _06011_, rst);
  not (_12448_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  nand (_12449_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  not (_12451_, _12449_);
  nor (_12452_, _12451_, _12448_);
  not (_12453_, _12452_);
  nand (_12454_, _12451_, _12448_);
  nand (_12455_, _12454_, _12453_);
  not (_12456_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  not (_12457_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  nor (_12458_, _12448_, _12457_);
  not (_12459_, _12458_);
  nor (_12460_, _12459_, _12456_);
  nor (_12461_, _12458_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_12462_, _12461_, _12460_);
  nor (_12463_, _12462_, _12451_);
  not (_12464_, _12463_);
  nand (_12465_, _12464_, _12455_);
  nor (_12466_, _12452_, _12457_);
  nor (_12467_, _12453_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  nor (_12468_, _12467_, _12466_);
  nor (_12469_, _12460_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  nor (_05833_, _12469_, rst);
  nand (_12471_, _05833_, _12468_);
  nor (_25041_, _12471_, _12465_);
  nor (_12472_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  nand (_12473_, _23553_, _11763_);
  nand (_12474_, _12473_, _23493_);
  nor (_25042_[31], _12474_, _12472_);
  nor (_12475_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand (_12476_, _23553_, _00057_);
  nand (_12477_, _12476_, _23493_);
  nor (_05867_, _12477_, _12475_);
  nor (_12478_, _10753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  nor (_12479_, _10755_, _21414_);
  nor (_05877_, _12479_, _12478_);
  not (_12480_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nor (_12481_, _12480_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor (_05880_, _12481_, rst);
  nor (_12482_, \oc8051_top_1.oc8051_decoder1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  nand (_12483_, _12482_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  nor (_05884_, _12483_, rst);
  not (_12484_, _05884_);
  nand (_12486_, _05783_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  nand (_05882_, _12486_, _12484_);
  nand (_12487_, _24801_, _23493_);
  nor (_05888_, _12487_, _24805_);
  nor (_12488_, _21865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  nor (_12489_, _21867_, _21526_);
  nor (_05890_, _12489_, _12488_);
  nor (_12490_, _09002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  nor (_12491_, _09004_, _21586_);
  nor (_05893_, _12491_, _12490_);
  nor (_12492_, _21766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  nor (_12493_, _21768_, _21586_);
  nor (_05902_, _12493_, _12492_);
  nor (_12494_, _21766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1]);
  nor (_12495_, _21768_, _21474_);
  nor (_25220_, _12495_, _12494_);
  nor (_12496_, _21766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  nor (_12497_, _21768_, _21554_);
  nor (_05906_, _12497_, _12496_);
  nor (_12498_, _21777_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7]);
  nor (_12500_, _21779_, _21626_);
  nor (_05919_, _12500_, _12498_);
  nor (_12501_, _22140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5]);
  nor (_12502_, _22142_, _21451_);
  nor (_05937_, _12502_, _12501_);
  nor (_12503_, _21766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7]);
  nor (_12504_, _21768_, _21626_);
  nor (_05939_, _12504_, _12503_);
  nor (_12505_, _21893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  nor (_12506_, _21895_, _21586_);
  nor (_05941_, _12506_, _12505_);
  nor (_12507_, _21834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  nor (_12508_, _21836_, _21504_);
  nor (_05943_, _12508_, _12507_);
  nor (_12509_, _21893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1]);
  nor (_12510_, _21895_, _21474_);
  nor (_05948_, _12510_, _12509_);
  nor (_12511_, _22484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  nor (_12512_, _22486_, _21586_);
  nor (_05956_, _12512_, _12511_);
  not (_12514_, _12483_);
  nor (_12515_, _12514_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nand (_12516_, _12514_, _10833_);
  nand (_12517_, _12516_, _23493_);
  nor (_05963_, _12517_, _12515_);
  nor (_12518_, _21766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5]);
  nor (_12519_, _21768_, _21451_);
  nor (_25221_, _12519_, _12518_);
  nor (_12520_, _12514_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nand (_12521_, _12514_, _10847_);
  nand (_12522_, _12521_, _23493_);
  nor (_05965_, _12522_, _12520_);
  nor (_12523_, _21766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  nor (_12524_, _21768_, _21504_);
  nor (_05967_, _12524_, _12523_);
  nor (_12525_, _12514_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nand (_12526_, _12514_, _10818_);
  nand (_12527_, _12526_, _23493_);
  nor (_05969_, _12527_, _12525_);
  nor (_12528_, _21766_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  nor (_12530_, _21768_, _21414_);
  nor (_05972_, _12530_, _12528_);
  nor (_12531_, _12514_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nand (_12532_, _12514_, _11658_);
  nand (_12533_, _12532_, _23493_);
  nor (_05973_, _12533_, _12531_);
  nor (_12534_, _22042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  nor (_12535_, _22044_, _21586_);
  nor (_05984_, _12535_, _12534_);
  nor (_12536_, _22042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1]);
  nor (_12537_, _22044_, _21474_);
  nor (_05986_, _12537_, _12536_);
  nor (_12538_, _21829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  nor (_12539_, _21831_, _21586_);
  nor (_05993_, _12539_, _12538_);
  nor (_12540_, _21893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  nor (_12541_, _21895_, _21504_);
  nor (_25222_, _12541_, _12540_);
  nor (_12542_, _21893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7]);
  nor (_12543_, _21895_, _21626_);
  nor (_06004_, _12543_, _12542_);
  nor (_12544_, _21893_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5]);
  nor (_12545_, _21895_, _21451_);
  nor (_06012_, _12545_, _12544_);
  nor (_12546_, _21834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7]);
  nor (_12547_, _21836_, _21626_);
  nor (_06023_, _12547_, _12546_);
  nor (_12548_, _22042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7]);
  nor (_12549_, _22044_, _21626_);
  nor (_06025_, _12549_, _12548_);
  nor (_12550_, _21887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  nor (_12551_, _21891_, _21586_);
  nor (_06030_, _12551_, _12550_);
  nor (_12552_, _21887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1]);
  nor (_12553_, _21891_, _21474_);
  nor (_06032_, _12553_, _12552_);
  nor (_12554_, _21834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  nor (_12555_, _21836_, _21554_);
  nor (_06044_, _12555_, _12554_);
  nor (_12556_, _22484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1]);
  nor (_12558_, _22486_, _21474_);
  nor (_06046_, _12558_, _12556_);
  nor (_12559_, _22042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  nor (_12560_, _22044_, _21414_);
  nor (_06049_, _12560_, _12559_);
  nor (_12561_, _22042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5]);
  nor (_12562_, _22044_, _21451_);
  nor (_25223_, _12562_, _12561_);
  nor (_12563_, _22551_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  nor (_12564_, _22555_, _21586_);
  nor (_06053_, _12564_, _12563_);
  nor (_12565_, _22042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  nor (_12566_, _22044_, _21504_);
  nor (_25224_, _12566_, _12565_);
  nor (_12567_, _22042_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  nor (_12568_, _22044_, _21526_);
  nor (_06058_, _12568_, _12567_);
  nor (_12569_, _21834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1]);
  nor (_12570_, _21836_, _21474_);
  nor (_06070_, _12570_, _12569_);
  nand (_12571_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6]);
  nand (_12572_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6]);
  nand (_12573_, _12572_, _12571_);
  nand (_12574_, _12573_, _00227_);
  nand (_12575_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6]);
  nand (_12576_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6]);
  nand (_12577_, _12576_, _12575_);
  nand (_12578_, _12577_, _01417_);
  nand (_12579_, _12578_, _12574_);
  nand (_12580_, _12579_, _00560_);
  nand (_12582_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6]);
  nand (_12583_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6]);
  nand (_12584_, _12583_, _12582_);
  nand (_12585_, _12584_, _00227_);
  nand (_12586_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6]);
  nand (_12587_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6]);
  nand (_12588_, _12587_, _12586_);
  nand (_12589_, _12588_, _01417_);
  nand (_12590_, _12589_, _12585_);
  nand (_12591_, _12590_, _00561_);
  nand (_12592_, _12591_, _12580_);
  nand (_12593_, _12592_, _00466_);
  nand (_12594_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6]);
  nand (_12595_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6]);
  nand (_12596_, _12595_, _12594_);
  nand (_12597_, _12596_, _01417_);
  nor (_12598_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6]);
  nor (_12599_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6]);
  nor (_12600_, _12599_, _12598_);
  nand (_12601_, _12600_, _00227_);
  nand (_12603_, _12601_, _12597_);
  nand (_12604_, _12603_, _00560_);
  nand (_12605_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6]);
  nand (_12606_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6]);
  nand (_12607_, _12606_, _12605_);
  nand (_12608_, _12607_, _01417_);
  nor (_12609_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6]);
  nor (_12610_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6]);
  nor (_12611_, _12610_, _12609_);
  nand (_12612_, _12611_, _00227_);
  nand (_12613_, _12612_, _12608_);
  nand (_12614_, _12613_, _00561_);
  nand (_12615_, _12614_, _12604_);
  nand (_12616_, _12615_, _00465_);
  nand (_12617_, _12616_, _12593_);
  nand (_12618_, _12617_, _00248_);
  nand (_12619_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6]);
  nand (_12620_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6]);
  nand (_12621_, _12620_, _12619_);
  nand (_12622_, _12621_, _01417_);
  nand (_12624_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6]);
  nand (_12625_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6]);
  nand (_12626_, _12625_, _12624_);
  nand (_12627_, _12626_, _00227_);
  nand (_12628_, _12627_, _12622_);
  nand (_12629_, _12628_, _00560_);
  nand (_12630_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6]);
  nand (_12631_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6]);
  nand (_12632_, _12631_, _12630_);
  nand (_12633_, _12632_, _01417_);
  nand (_12634_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6]);
  nand (_12635_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6]);
  nand (_12636_, _12635_, _12634_);
  nand (_12637_, _12636_, _00227_);
  nand (_12638_, _12637_, _12633_);
  nand (_12639_, _12638_, _00561_);
  nand (_12640_, _12639_, _12629_);
  nand (_12641_, _12640_, _00466_);
  nor (_12642_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6]);
  nor (_12643_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6]);
  nor (_12645_, _12643_, _12642_);
  nand (_12646_, _12645_, _01417_);
  nor (_12647_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6]);
  nor (_12648_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6]);
  nor (_12649_, _12648_, _12647_);
  nand (_12650_, _12649_, _00227_);
  nand (_12651_, _12650_, _12646_);
  nand (_12652_, _12651_, _00560_);
  nor (_12653_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6]);
  nor (_12654_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6]);
  nor (_12655_, _12654_, _12653_);
  nor (_12656_, _12655_, _00227_);
  nor (_12657_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6]);
  nor (_12658_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6]);
  nor (_12659_, _12658_, _12657_);
  nor (_12660_, _12659_, _01417_);
  nor (_12661_, _12660_, _12656_);
  nand (_12662_, _12661_, _00561_);
  nand (_12663_, _12662_, _12652_);
  nand (_12664_, _12663_, _00465_);
  nand (_12666_, _12664_, _12641_);
  nand (_12667_, _12666_, _00247_);
  nand (_12668_, _12667_, _12618_);
  nand (_12669_, _12668_, _00320_);
  nand (_12670_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6]);
  nand (_12671_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6]);
  nand (_12672_, _12671_, _12670_);
  nand (_12673_, _12672_, _01417_);
  nand (_12674_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6]);
  nand (_12675_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6]);
  nand (_12676_, _12675_, _12674_);
  nand (_12677_, _12676_, _00227_);
  nand (_12678_, _12677_, _12673_);
  nand (_12679_, _12678_, _00560_);
  nand (_12680_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6]);
  nand (_12681_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6]);
  nand (_12682_, _12681_, _12680_);
  nand (_12683_, _12682_, _01417_);
  nand (_12684_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6]);
  nand (_12685_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6]);
  nand (_12686_, _12685_, _12684_);
  nand (_12687_, _12686_, _00227_);
  nand (_12688_, _12687_, _12683_);
  nand (_12689_, _12688_, _00561_);
  nand (_12690_, _12689_, _12679_);
  nand (_12691_, _12690_, _00466_);
  nor (_12692_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6]);
  nor (_12693_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6]);
  nor (_12694_, _12693_, _12692_);
  nand (_12695_, _12694_, _01417_);
  nor (_12697_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6]);
  nor (_12698_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6]);
  nor (_12699_, _12698_, _12697_);
  nand (_12700_, _12699_, _00227_);
  nand (_12701_, _12700_, _12695_);
  nand (_12702_, _12701_, _00560_);
  nor (_12703_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6]);
  nor (_12704_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6]);
  nor (_12705_, _12704_, _12703_);
  nand (_12706_, _12705_, _01417_);
  nor (_12707_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6]);
  nor (_12708_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6]);
  nor (_12709_, _12708_, _12707_);
  nand (_12710_, _12709_, _00227_);
  nand (_12711_, _12710_, _12706_);
  nand (_12712_, _12711_, _00561_);
  nand (_12713_, _12712_, _12702_);
  nand (_12714_, _12713_, _00465_);
  nand (_12715_, _12714_, _12691_);
  nand (_12716_, _12715_, _00248_);
  nand (_12718_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6]);
  nand (_12719_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6]);
  nand (_12720_, _12719_, _12718_);
  nand (_12721_, _12720_, _01417_);
  nand (_12722_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6]);
  nand (_12723_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6]);
  nand (_12724_, _12723_, _12722_);
  nand (_12725_, _12724_, _00227_);
  nand (_12726_, _12725_, _12721_);
  nand (_12727_, _12726_, _00560_);
  nand (_12728_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6]);
  nand (_12729_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6]);
  nand (_12730_, _12729_, _12728_);
  nand (_12731_, _12730_, _01417_);
  nand (_12732_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6]);
  nand (_12733_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6]);
  nand (_12734_, _12733_, _12732_);
  nand (_12735_, _12734_, _00227_);
  nand (_12736_, _12735_, _12731_);
  nand (_12737_, _12736_, _00561_);
  nand (_12738_, _12737_, _12727_);
  nand (_12739_, _12738_, _00466_);
  nor (_12740_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6]);
  nor (_12741_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6]);
  nor (_12742_, _12741_, _12740_);
  nand (_12743_, _12742_, _01417_);
  nor (_12744_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6]);
  nor (_12745_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6]);
  nor (_12746_, _12745_, _12744_);
  nand (_12747_, _12746_, _00227_);
  nand (_12748_, _12747_, _12743_);
  nand (_12749_, _12748_, _00560_);
  nor (_12750_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6]);
  nor (_12751_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6]);
  nor (_12752_, _12751_, _12750_);
  nand (_12753_, _12752_, _01417_);
  nor (_12754_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6]);
  nor (_12755_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6]);
  nor (_12756_, _12755_, _12754_);
  nand (_12757_, _12756_, _00227_);
  nand (_12758_, _12757_, _12753_);
  nand (_12759_, _12758_, _00561_);
  nand (_12760_, _12759_, _12749_);
  nand (_12761_, _12760_, _00465_);
  nand (_12762_, _12761_, _12739_);
  nand (_12763_, _12762_, _00247_);
  nand (_12764_, _12763_, _12716_);
  nand (_12765_, _12764_, _00319_);
  nand (_12766_, _12765_, _12669_);
  nor (_12767_, _12766_, _00386_);
  nand (_12768_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6]);
  nand (_12769_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6]);
  nand (_12770_, _12769_, _12768_);
  nand (_12771_, _12770_, _01417_);
  nand (_12772_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6]);
  nand (_12773_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6]);
  nand (_12774_, _12773_, _12772_);
  nand (_12775_, _12774_, _00227_);
  nand (_12776_, _12775_, _12771_);
  nand (_12777_, _12776_, _00560_);
  nand (_12778_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6]);
  nand (_12779_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6]);
  nand (_12780_, _12779_, _12778_);
  nand (_12781_, _12780_, _01417_);
  nand (_12782_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6]);
  nand (_12783_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6]);
  nand (_12784_, _12783_, _12782_);
  nand (_12785_, _12784_, _00227_);
  nand (_12786_, _12785_, _12781_);
  nand (_12787_, _12786_, _00561_);
  nand (_12788_, _12787_, _12777_);
  nand (_12789_, _12788_, _00466_);
  nor (_12790_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6]);
  nor (_12791_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6]);
  nor (_12792_, _12791_, _12790_);
  nand (_12793_, _12792_, _00227_);
  nand (_12794_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6]);
  nand (_12795_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6]);
  nand (_12796_, _12795_, _12794_);
  nand (_12797_, _12796_, _01417_);
  nand (_12798_, _12797_, _12793_);
  nand (_12799_, _12798_, _00560_);
  nor (_12800_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6]);
  nor (_12801_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6]);
  nor (_12802_, _12801_, _12800_);
  nand (_12803_, _12802_, _00227_);
  nand (_12804_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6]);
  nand (_12805_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6]);
  nand (_12806_, _12805_, _12804_);
  nand (_12807_, _12806_, _01417_);
  nand (_12808_, _12807_, _12803_);
  nand (_12809_, _12808_, _00561_);
  nand (_12810_, _12809_, _12799_);
  nand (_12811_, _12810_, _00465_);
  nand (_12812_, _12811_, _12789_);
  nand (_12813_, _12812_, _00248_);
  nand (_12814_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6]);
  nand (_12815_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6]);
  nand (_12816_, _12815_, _12814_);
  nand (_12817_, _12816_, _01417_);
  nand (_12818_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6]);
  nand (_12819_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6]);
  nand (_12820_, _12819_, _12818_);
  nand (_12821_, _12820_, _00227_);
  nand (_12822_, _12821_, _12817_);
  nand (_12823_, _12822_, _00560_);
  nand (_12824_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6]);
  nand (_12825_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6]);
  nand (_12826_, _12825_, _12824_);
  nand (_12827_, _12826_, _01417_);
  nand (_12829_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6]);
  nand (_12830_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6]);
  nand (_12831_, _12830_, _12829_);
  nand (_12832_, _12831_, _00227_);
  nand (_12833_, _12832_, _12827_);
  nand (_12834_, _12833_, _00561_);
  nand (_12835_, _12834_, _12823_);
  nand (_12836_, _12835_, _00466_);
  nor (_12837_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6]);
  nor (_12838_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6]);
  nor (_12839_, _12838_, _12837_);
  nand (_12840_, _12839_, _01417_);
  nor (_12841_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6]);
  nor (_12842_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  nor (_12843_, _12842_, _12841_);
  nand (_12844_, _12843_, _00227_);
  nand (_12845_, _12844_, _12840_);
  nand (_12846_, _12845_, _00560_);
  nor (_12847_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6]);
  nor (_12848_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6]);
  nor (_12849_, _12848_, _12847_);
  nand (_12850_, _12849_, _01417_);
  nor (_12851_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  nor (_12852_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6]);
  nor (_12853_, _12852_, _12851_);
  nand (_12854_, _12853_, _00227_);
  nand (_12855_, _12854_, _12850_);
  nand (_12856_, _12855_, _00561_);
  nand (_12857_, _12856_, _12846_);
  nand (_12858_, _12857_, _00465_);
  nand (_12859_, _12858_, _12836_);
  nand (_12860_, _12859_, _00247_);
  nand (_12861_, _12860_, _12813_);
  nand (_12862_, _12861_, _00320_);
  nor (_12863_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6]);
  nor (_12864_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6]);
  nor (_12865_, _12864_, _12863_);
  nand (_12866_, _12865_, _01417_);
  nor (_12867_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6]);
  nor (_12868_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6]);
  nor (_12870_, _12868_, _12867_);
  nand (_12871_, _12870_, _00227_);
  nand (_12872_, _12871_, _12866_);
  nand (_12873_, _12872_, _00561_);
  nor (_12874_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6]);
  nor (_12875_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6]);
  nor (_12876_, _12875_, _12874_);
  nand (_12877_, _12876_, _01417_);
  nor (_12878_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6]);
  nor (_12879_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6]);
  nor (_12880_, _12879_, _12878_);
  nand (_12881_, _12880_, _00227_);
  nand (_12882_, _12881_, _12877_);
  nand (_12883_, _12882_, _00560_);
  nand (_12884_, _12883_, _12873_);
  nand (_12885_, _12884_, _00465_);
  nand (_12886_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6]);
  nand (_12887_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6]);
  nand (_12888_, _12887_, _12886_);
  nand (_12889_, _12888_, _01417_);
  nand (_12891_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6]);
  nand (_12892_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6]);
  nand (_12893_, _12892_, _12891_);
  nand (_12894_, _12893_, _00227_);
  nand (_12895_, _12894_, _12889_);
  nand (_12896_, _12895_, _00561_);
  nand (_12897_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6]);
  nand (_12898_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6]);
  nand (_12899_, _12898_, _12897_);
  nand (_12900_, _12899_, _01417_);
  nand (_12901_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6]);
  nand (_12902_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6]);
  nand (_12903_, _12902_, _12901_);
  nand (_12904_, _12903_, _00227_);
  nand (_12905_, _12904_, _12900_);
  nand (_12906_, _12905_, _00560_);
  nand (_12907_, _12906_, _12896_);
  nand (_12908_, _12907_, _00466_);
  nand (_12909_, _12908_, _12885_);
  nand (_12910_, _12909_, _00247_);
  nor (_12912_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6]);
  nor (_12913_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6]);
  nor (_12914_, _12913_, _12912_);
  nand (_12915_, _12914_, _00227_);
  nand (_12916_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6]);
  nand (_12917_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6]);
  nand (_12918_, _12917_, _12916_);
  nand (_12919_, _12918_, _01417_);
  nand (_12920_, _12919_, _12915_);
  nand (_12921_, _12920_, _00561_);
  nor (_12922_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6]);
  nor (_12923_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6]);
  nor (_12924_, _12923_, _12922_);
  nand (_12925_, _12924_, _00227_);
  nand (_12926_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6]);
  nand (_12927_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6]);
  nand (_12928_, _12927_, _12926_);
  nand (_12929_, _12928_, _01417_);
  nand (_12930_, _12929_, _12925_);
  nand (_12931_, _12930_, _00560_);
  nand (_12933_, _12931_, _12921_);
  nand (_12934_, _12933_, _00465_);
  nand (_12935_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6]);
  nand (_12936_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6]);
  nand (_12937_, _12936_, _12935_);
  nand (_12938_, _12937_, _01417_);
  nand (_12939_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6]);
  nand (_12940_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6]);
  nand (_12941_, _12940_, _12939_);
  nand (_12942_, _12941_, _00227_);
  nand (_12943_, _12942_, _12938_);
  nand (_12944_, _12943_, _00561_);
  nand (_12945_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6]);
  nand (_12946_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6]);
  nand (_12947_, _12946_, _12945_);
  nand (_12948_, _12947_, _01417_);
  nand (_12949_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6]);
  nand (_12950_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6]);
  nand (_12951_, _12950_, _12949_);
  nand (_12952_, _12951_, _00227_);
  nand (_12954_, _12952_, _12948_);
  nand (_12955_, _12954_, _00560_);
  nand (_12956_, _12955_, _12944_);
  nand (_12957_, _12956_, _00466_);
  nand (_12958_, _12957_, _12934_);
  nand (_12959_, _12958_, _00248_);
  nand (_12960_, _12959_, _12910_);
  nand (_12961_, _12960_, _00319_);
  nand (_12962_, _12961_, _12862_);
  nor (_12963_, _12962_, _01629_);
  nor (_12964_, _12963_, _12767_);
  nor (_12965_, _12964_, _00156_);
  nand (_12966_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6]);
  nand (_12967_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6]);
  nand (_12968_, _12967_, _12966_);
  nand (_12969_, _12968_, _01417_);
  nand (_12970_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6]);
  nand (_12971_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6]);
  nand (_12972_, _12971_, _12970_);
  nand (_12973_, _12972_, _00227_);
  nand (_12975_, _12973_, _12969_);
  nand (_12976_, _12975_, _00560_);
  nand (_12977_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6]);
  nand (_12978_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6]);
  nand (_12979_, _12978_, _12977_);
  nand (_12980_, _12979_, _01417_);
  nand (_12981_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6]);
  nand (_12982_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6]);
  nand (_12983_, _12982_, _12981_);
  nand (_12984_, _12983_, _00227_);
  nand (_12985_, _12984_, _12980_);
  nand (_12986_, _12985_, _00561_);
  nand (_12987_, _12986_, _12976_);
  nand (_12988_, _12987_, _00466_);
  nor (_12989_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6]);
  nor (_12990_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6]);
  nor (_12991_, _12990_, _12989_);
  nand (_12992_, _12991_, _01417_);
  nor (_12993_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6]);
  nor (_12994_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6]);
  nor (_12995_, _12994_, _12993_);
  nand (_12996_, _12995_, _00227_);
  nand (_12997_, _12996_, _12992_);
  nand (_12998_, _12997_, _00560_);
  nor (_12999_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6]);
  nor (_13000_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6]);
  nor (_13001_, _13000_, _12999_);
  nand (_13002_, _13001_, _01417_);
  nor (_13003_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6]);
  nor (_13004_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6]);
  nor (_13006_, _13004_, _13003_);
  nand (_13007_, _13006_, _00227_);
  nand (_13008_, _13007_, _13002_);
  nand (_13009_, _13008_, _00561_);
  nand (_13010_, _13009_, _12998_);
  nand (_13011_, _13010_, _00465_);
  nand (_13012_, _13011_, _12988_);
  nand (_13013_, _13012_, _00247_);
  nand (_13014_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6]);
  nand (_13015_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6]);
  nand (_13016_, _13015_, _13014_);
  nand (_13017_, _13016_, _01417_);
  nand (_13018_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6]);
  nand (_13019_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6]);
  nand (_13020_, _13019_, _13018_);
  nand (_13021_, _13020_, _00227_);
  nand (_13022_, _13021_, _13017_);
  nand (_13023_, _13022_, _00560_);
  nand (_13024_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6]);
  nand (_13025_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6]);
  nand (_13027_, _13025_, _13024_);
  nand (_13028_, _13027_, _01417_);
  nand (_13029_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6]);
  nand (_13030_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6]);
  nand (_13031_, _13030_, _13029_);
  nand (_13032_, _13031_, _00227_);
  nand (_13033_, _13032_, _13028_);
  nand (_13034_, _13033_, _00561_);
  nand (_13035_, _13034_, _13023_);
  nand (_13036_, _13035_, _00466_);
  nor (_13037_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6]);
  nor (_13038_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6]);
  nor (_13039_, _13038_, _13037_);
  nand (_13040_, _13039_, _00227_);
  nand (_13041_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6]);
  nand (_13042_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6]);
  nand (_13043_, _13042_, _13041_);
  nand (_13044_, _13043_, _01417_);
  nand (_13045_, _13044_, _13040_);
  nand (_13046_, _13045_, _00560_);
  nor (_13047_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6]);
  nor (_13048_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6]);
  nor (_13049_, _13048_, _13047_);
  nand (_13050_, _13049_, _00227_);
  nand (_13051_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6]);
  nand (_13052_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  nand (_13053_, _13052_, _13051_);
  nand (_13054_, _13053_, _01417_);
  nand (_13055_, _13054_, _13050_);
  nand (_13056_, _13055_, _00561_);
  nand (_13058_, _13056_, _13046_);
  nand (_13059_, _13058_, _00465_);
  nand (_13060_, _13059_, _13036_);
  nand (_13061_, _13060_, _00248_);
  nand (_13062_, _13061_, _13013_);
  nand (_13063_, _13062_, _00320_);
  nand (_13064_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  nand (_13065_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  nand (_13066_, _13065_, _13064_);
  nand (_13067_, _13066_, _01417_);
  nand (_13068_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6]);
  nand (_13069_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  nand (_13070_, _13069_, _13068_);
  nand (_13071_, _13070_, _00227_);
  nand (_13072_, _13071_, _13067_);
  nand (_13073_, _13072_, _00560_);
  nand (_13074_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6]);
  nand (_13075_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  nand (_13076_, _13075_, _13074_);
  nand (_13077_, _13076_, _01417_);
  nand (_13078_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  nand (_13079_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  nand (_13080_, _13079_, _13078_);
  nand (_13081_, _13080_, _00227_);
  nand (_13082_, _13081_, _13077_);
  nand (_13083_, _13082_, _00561_);
  nand (_13084_, _13083_, _13073_);
  nand (_13085_, _13084_, _00466_);
  nor (_13086_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6]);
  nor (_13087_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  nor (_13088_, _13087_, _13086_);
  nand (_13089_, _13088_, _00227_);
  nand (_13090_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  nand (_13091_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  nand (_13092_, _13091_, _13090_);
  nand (_13093_, _13092_, _01417_);
  nand (_13094_, _13093_, _13089_);
  nand (_13095_, _13094_, _00560_);
  nor (_13096_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6]);
  nor (_13097_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6]);
  nor (_13098_, _13097_, _13096_);
  nand (_13099_, _13098_, _00227_);
  nand (_13100_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6]);
  nand (_13101_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6]);
  nand (_13102_, _13101_, _13100_);
  nand (_13103_, _13102_, _01417_);
  nand (_13104_, _13103_, _13099_);
  nand (_13105_, _13104_, _00561_);
  nand (_13106_, _13105_, _13095_);
  nand (_13107_, _13106_, _00465_);
  nand (_13109_, _13107_, _13085_);
  nand (_13110_, _13109_, _00248_);
  nand (_13111_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  nand (_13112_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6]);
  nand (_13113_, _13112_, _13111_);
  nand (_13114_, _13113_, _01417_);
  nand (_13115_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6]);
  nand (_13116_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6]);
  nand (_13117_, _13116_, _13115_);
  nand (_13118_, _13117_, _00227_);
  nand (_13119_, _13118_, _13114_);
  nand (_13120_, _13119_, _00560_);
  nand (_13121_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6]);
  nand (_13122_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6]);
  nand (_13123_, _13122_, _13121_);
  nand (_13124_, _13123_, _01417_);
  nand (_13125_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6]);
  nand (_13126_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6]);
  nand (_13127_, _13126_, _13125_);
  nand (_13128_, _13127_, _00227_);
  nand (_13129_, _13128_, _13124_);
  nand (_13130_, _13129_, _00561_);
  nand (_13131_, _13130_, _13120_);
  nand (_13132_, _13131_, _00466_);
  nor (_13133_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6]);
  nor (_13134_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6]);
  nor (_13135_, _13134_, _13133_);
  nand (_13136_, _13135_, _01417_);
  nor (_13137_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6]);
  nor (_13138_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6]);
  nor (_13139_, _13138_, _13137_);
  nand (_13140_, _13139_, _00227_);
  nand (_13141_, _13140_, _13136_);
  nand (_13142_, _13141_, _00560_);
  nor (_13143_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6]);
  nor (_13144_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6]);
  nor (_13145_, _13144_, _13143_);
  nand (_13146_, _13145_, _01417_);
  nor (_13147_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6]);
  nor (_13148_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6]);
  nor (_13149_, _13148_, _13147_);
  nand (_13150_, _13149_, _00227_);
  nand (_13151_, _13150_, _13146_);
  nand (_13152_, _13151_, _00561_);
  nand (_13153_, _13152_, _13142_);
  nand (_13154_, _13153_, _00465_);
  nand (_13155_, _13154_, _13132_);
  nand (_13156_, _13155_, _00247_);
  nand (_13157_, _13156_, _13110_);
  nand (_13158_, _13157_, _00319_);
  nand (_13159_, _13158_, _13063_);
  nor (_13160_, _13159_, _00386_);
  nand (_13161_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  nand (_13162_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6]);
  nand (_13163_, _13162_, _13161_);
  nand (_13164_, _13163_, _01417_);
  nand (_13165_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  nand (_13166_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  nand (_13167_, _13166_, _13165_);
  nand (_13168_, _13167_, _00227_);
  nand (_13169_, _13168_, _13164_);
  nand (_13170_, _13169_, _00560_);
  nand (_13171_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  nand (_13172_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  nand (_13173_, _13172_, _13171_);
  nand (_13174_, _13173_, _01417_);
  nand (_13175_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  nand (_13176_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  nand (_13177_, _13176_, _13175_);
  nand (_13178_, _13177_, _00227_);
  nand (_13179_, _13178_, _13174_);
  nand (_13180_, _13179_, _00561_);
  nand (_13181_, _13180_, _13170_);
  nand (_13182_, _13181_, _00466_);
  nor (_13183_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6]);
  nor (_13184_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6]);
  nor (_13185_, _13184_, _13183_);
  nand (_13186_, _13185_, _00227_);
  nand (_13187_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  nand (_13188_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  nand (_13190_, _13188_, _13187_);
  nand (_13191_, _13190_, _01417_);
  nand (_13192_, _13191_, _13186_);
  nand (_13193_, _13192_, _00560_);
  nor (_13194_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6]);
  nor (_13195_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6]);
  nor (_13196_, _13195_, _13194_);
  nand (_13197_, _13196_, _00227_);
  nand (_13198_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  nand (_13199_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  nand (_13200_, _13199_, _13198_);
  nand (_13201_, _13200_, _01417_);
  nand (_13202_, _13201_, _13197_);
  nand (_13203_, _13202_, _00561_);
  nand (_13204_, _13203_, _13193_);
  nand (_13205_, _13204_, _00465_);
  nand (_13206_, _13205_, _13182_);
  nand (_13207_, _13206_, _00248_);
  nand (_13208_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  nand (_13209_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6]);
  nand (_13210_, _13209_, _13208_);
  nand (_13211_, _13210_, _01417_);
  nand (_13212_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6]);
  nand (_13213_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6]);
  nand (_13214_, _13213_, _13212_);
  nand (_13215_, _13214_, _00227_);
  nand (_13216_, _13215_, _13211_);
  nand (_13217_, _13216_, _00560_);
  nand (_13218_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6]);
  nand (_13219_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6]);
  nand (_13220_, _13219_, _13218_);
  nand (_13221_, _13220_, _01417_);
  nand (_13222_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6]);
  nand (_13223_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6]);
  nand (_13224_, _13223_, _13222_);
  nand (_13225_, _13224_, _00227_);
  nand (_13226_, _13225_, _13221_);
  nand (_13227_, _13226_, _00561_);
  nand (_13228_, _13227_, _13217_);
  nand (_13229_, _13228_, _00466_);
  nor (_13230_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6]);
  nor (_13231_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6]);
  nor (_13232_, _13231_, _13230_);
  nand (_13233_, _13232_, _01417_);
  nor (_13234_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6]);
  nor (_13235_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6]);
  nor (_13236_, _13235_, _13234_);
  nand (_13237_, _13236_, _00227_);
  nand (_13238_, _13237_, _13233_);
  nand (_13239_, _13238_, _00560_);
  nor (_13240_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6]);
  nor (_13241_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6]);
  nor (_13242_, _13241_, _13240_);
  nand (_13243_, _13242_, _01417_);
  nor (_13244_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6]);
  nor (_13245_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6]);
  nor (_13246_, _13245_, _13244_);
  nand (_13247_, _13246_, _00227_);
  nand (_13248_, _13247_, _13243_);
  nand (_13249_, _13248_, _00561_);
  nand (_13251_, _13249_, _13239_);
  nand (_13252_, _13251_, _00465_);
  nand (_13253_, _13252_, _13229_);
  nand (_13254_, _13253_, _00247_);
  nand (_13255_, _13254_, _13207_);
  nand (_13256_, _13255_, _00320_);
  nor (_13257_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6]);
  nor (_13258_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  nor (_13259_, _13258_, _13257_);
  nand (_13260_, _13259_, _01417_);
  nor (_13261_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6]);
  nor (_13262_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6]);
  nor (_13263_, _13262_, _13261_);
  nand (_13264_, _13263_, _00227_);
  nand (_13265_, _13264_, _13260_);
  nand (_13266_, _13265_, _00561_);
  nor (_13267_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6]);
  nor (_13268_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6]);
  nor (_13269_, _13268_, _13267_);
  nand (_13270_, _13269_, _01417_);
  nor (_13271_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6]);
  nor (_13272_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6]);
  nor (_13273_, _13272_, _13271_);
  nand (_13274_, _13273_, _00227_);
  nand (_13275_, _13274_, _13270_);
  nand (_13276_, _13275_, _00560_);
  nand (_13277_, _13276_, _13266_);
  nand (_13278_, _13277_, _00465_);
  nand (_13279_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6]);
  nand (_13280_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6]);
  nand (_13281_, _13280_, _13279_);
  nand (_13282_, _13281_, _01417_);
  nand (_13283_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6]);
  nand (_13284_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6]);
  nand (_13285_, _13284_, _13283_);
  nand (_13286_, _13285_, _00227_);
  nand (_13287_, _13286_, _13282_);
  nand (_13288_, _13287_, _00561_);
  nand (_13289_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  nand (_13290_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  nand (_13291_, _13290_, _13289_);
  nand (_13292_, _13291_, _01417_);
  nand (_13293_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  nand (_13294_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  nand (_13295_, _13294_, _13293_);
  nand (_13296_, _13295_, _00227_);
  nand (_13297_, _13296_, _13292_);
  nand (_13298_, _13297_, _00560_);
  nand (_13299_, _13298_, _13288_);
  nand (_13300_, _13299_, _00466_);
  nand (_13301_, _13300_, _13278_);
  nand (_13302_, _13301_, _00247_);
  nor (_13303_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6]);
  nor (_13304_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6]);
  nor (_13305_, _13304_, _13303_);
  nand (_13306_, _13305_, _00227_);
  nand (_13307_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  nand (_13308_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6]);
  nand (_13309_, _13308_, _13307_);
  nand (_13310_, _13309_, _01417_);
  nand (_13312_, _13310_, _13306_);
  nand (_13313_, _13312_, _00561_);
  nor (_13314_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6]);
  nor (_13315_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6]);
  nor (_13316_, _13315_, _13314_);
  nand (_13317_, _13316_, _00227_);
  nand (_13318_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  nand (_13319_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6]);
  nand (_13320_, _13319_, _13318_);
  nand (_13321_, _13320_, _01417_);
  nand (_13322_, _13321_, _13317_);
  nand (_13323_, _13322_, _00560_);
  nand (_13324_, _13323_, _13313_);
  nand (_13325_, _13324_, _00465_);
  nand (_13326_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  nand (_13327_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  nand (_13328_, _13327_, _13326_);
  nand (_13329_, _13328_, _01417_);
  nand (_13330_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6]);
  nand (_13331_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  nand (_13333_, _13331_, _13330_);
  nand (_13334_, _13333_, _00227_);
  nand (_13335_, _13334_, _13329_);
  nand (_13336_, _13335_, _00561_);
  nand (_13337_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6]);
  nand (_13338_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6]);
  nand (_13339_, _13338_, _13337_);
  nand (_13340_, _13339_, _01417_);
  nand (_13341_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6]);
  nand (_13342_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  nand (_13343_, _13342_, _13341_);
  nand (_13344_, _13343_, _00227_);
  nand (_13345_, _13344_, _13340_);
  nand (_13346_, _13345_, _00560_);
  nand (_13347_, _13346_, _13336_);
  nand (_13348_, _13347_, _00466_);
  nand (_13349_, _13348_, _13325_);
  nand (_13350_, _13349_, _00248_);
  nand (_13351_, _13350_, _13302_);
  nand (_13352_, _13351_, _00319_);
  nand (_13354_, _13352_, _13256_);
  nor (_13355_, _13354_, _01629_);
  nor (_13356_, _13355_, _13160_);
  nor (_13357_, _13356_, _00556_);
  nor (_13358_, _13357_, _12965_);
  nor (_13359_, _13358_, _01416_);
  not (_13360_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  nand (_13361_, _01416_, _13360_);
  nand (_13362_, _13361_, _23493_);
  nor (_06073_, _13362_, _13359_);
  nor (_13363_, _21887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7]);
  nor (_13364_, _21891_, _21626_);
  nor (_06088_, _13364_, _13363_);
  nor (_13365_, _22140_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6]);
  nor (_13366_, _22142_, _21504_);
  nor (_06090_, _13366_, _13365_);
  nor (_13367_, _21887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5]);
  nor (_13368_, _21891_, _21451_);
  nor (_06107_, _13368_, _13367_);
  nor (_13369_, _21887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6]);
  nor (_13370_, _21891_, _21504_);
  nor (_06110_, _13370_, _13369_);
  nor (_13371_, _21887_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  nor (_13372_, _21891_, _21414_);
  nor (_06113_, _13372_, _13371_);
  nor (_13373_, _22484_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7]);
  nor (_13374_, _22486_, _21626_);
  nor (_06121_, _13374_, _13373_);
  nor (_13375_, _24380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  nor (_13376_, _24382_, _21554_);
  nor (_25292_, _13376_, _13375_);
  nor (_13377_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nand (_13378_, _23553_, _00366_);
  nand (_13379_, _13378_, _23493_);
  nor (_25043_[30], _13379_, _13377_);
  nor (_13380_, _22557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7]);
  nor (_13381_, _22559_, _21626_);
  nor (_06127_, _13381_, _13380_);
  nor (_13382_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_13383_, _23553_, _00285_);
  nand (_13384_, _13383_, _23493_);
  nor (_25043_[29], _13384_, _13382_);
  nor (_13385_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand (_13386_, _23553_, _23052_);
  nand (_13387_, _13386_, _23493_);
  nor (_06132_, _13387_, _13385_);
  nor (_13388_, _22054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5]);
  nor (_13389_, _22056_, _21451_);
  nor (_06134_, _13389_, _13388_);
  nor (_13390_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand (_13392_, _23553_, _23185_);
  nand (_13393_, _13392_, _23493_);
  nor (_06146_, _13393_, _13390_);
  nor (_13394_, _22054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6]);
  nor (_13395_, _22056_, _21504_);
  nor (_06149_, _13395_, _13394_);
  nor (_13396_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_13397_, _23553_, _23212_);
  nand (_13398_, _13397_, _23493_);
  nor (_06152_, _13398_, _13396_);
  nor (_13399_, _22054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  nor (_13400_, _22056_, _21414_);
  nor (_06154_, _13400_, _13399_);
  nor (_13401_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_13402_, _23553_, _23259_);
  nand (_13403_, _13402_, _23493_);
  nor (_06158_, _13403_, _13401_);
  nor (_13404_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand (_13405_, _23553_, _00601_);
  nand (_13406_, _13405_, _23493_);
  nor (_06161_, _13406_, _13404_);
  nor (_13407_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand (_13408_, _23553_, _23391_);
  nand (_13409_, _13408_, _23493_);
  nor (_25043_[23], _13409_, _13407_);
  nor (_13410_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand (_13411_, _23553_, _23105_);
  nand (_13412_, _13411_, _23493_);
  nor (_06174_, _13412_, _13410_);
  nor (_13413_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand (_13415_, _23553_, _00292_);
  nand (_13416_, _13415_, _23493_);
  nor (_25043_[21], _13416_, _13413_);
  nor (_13417_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand (_13418_, _23553_, _24183_);
  nand (_13419_, _13418_, _23493_);
  nor (_06179_, _13419_, _13417_);
  nor (_13420_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  nor (_13421_, _22563_, _21414_);
  nor (_25076_, _13421_, _13420_);
  nor (_13422_, _10753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6]);
  nor (_13423_, _10755_, _21504_);
  nor (_06190_, _13423_, _13422_);
  nor (_13424_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand (_13425_, _23553_, _23190_);
  nand (_13426_, _13425_, _23493_);
  nor (_06198_, _13426_, _13424_);
  nor (_13427_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand (_13428_, _23553_, _23217_);
  nand (_13429_, _13428_, _23493_);
  nor (_06201_, _13429_, _13427_);
  nor (_13430_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand (_13431_, _23553_, _24835_);
  nand (_13432_, _13431_, _23493_);
  nor (_06205_, _13432_, _13430_);
  nor (_13433_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand (_13434_, _23553_, _00607_);
  nand (_13435_, _13434_, _23493_);
  nor (_06208_, _13435_, _13433_);
  nor (_13436_, _22054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  nor (_13438_, _22056_, _21554_);
  nor (_06210_, _13438_, _13436_);
  nor (_13439_, _22054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  nor (_13440_, _22056_, _21526_);
  nor (_06213_, _13440_, _13439_);
  nor (_13441_, _22054_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1]);
  nor (_13442_, _22056_, _21474_);
  nor (_06216_, _13442_, _13441_);
  nor (_13443_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_13444_, _23553_, _23286_);
  nand (_13445_, _13444_, _23493_);
  nor (_25043_[15], _13445_, _13443_);
  nor (_13446_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_13447_, _23553_, _23100_);
  nand (_13448_, _13447_, _23493_);
  nor (_06221_, _13448_, _13446_);
  nor (_13449_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_13450_, _23553_, _23124_);
  nand (_13451_, _13450_, _23493_);
  nor (_06224_, _13451_, _13449_);
  nor (_13452_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nand (_13453_, _23553_, _23065_);
  nand (_13454_, _13453_, _23493_);
  nor (_06233_, _13454_, _13452_);
  nor (_13455_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_13456_, _23553_, _00448_);
  nand (_13457_, _13456_, _23493_);
  nor (_06236_, _13457_, _13455_);
  nor (_13458_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand (_13459_, _23553_, _23360_);
  nand (_13460_, _13459_, _23493_);
  nor (_06239_, _13460_, _13458_);
  nor (_13461_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_13462_, _23553_, _23264_);
  nand (_13463_, _13462_, _23493_);
  nor (_06242_, _13463_, _13461_);
  nor (_13464_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_13465_, _23553_, _23156_);
  nand (_13466_, _13465_, _23493_);
  nor (_06248_, _13466_, _13464_);
  nor (_13468_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nand (_13469_, _23553_, _23284_);
  nand (_13470_, _13469_, _23493_);
  nor (_06251_, _13470_, _13468_);
  nor (_13471_, _21938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5]);
  nor (_13472_, _21940_, _21451_);
  nor (_06263_, _13472_, _13471_);
  nor (_13473_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nand (_13474_, _23553_, _23090_);
  nand (_13475_, _13474_, _23493_);
  nor (_06266_, _13475_, _13473_);
  nor (_13476_, _21938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6]);
  nor (_13477_, _21940_, _21504_);
  nor (_06269_, _13477_, _13476_);
  nor (_13478_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nand (_13479_, _23553_, _23122_);
  nand (_13480_, _13479_, _23493_);
  nor (_25043_[5], _13480_, _13478_);
  nor (_13481_, _21938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  nor (_13482_, _21940_, _21414_);
  nor (_06273_, _13482_, _13481_);
  nor (_13483_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand (_13484_, _23553_, _23075_);
  nand (_13485_, _13484_, _23493_);
  nor (_06276_, _13485_, _13483_);
  nor (_13486_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  not (_13487_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_13488_, _23553_, _13487_);
  nand (_13489_, _13488_, _23493_);
  nor (_06279_, _13489_, _13486_);
  nor (_13490_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand (_13491_, _23553_, _23204_);
  nand (_13492_, _13491_, _23493_);
  nor (_06282_, _13492_, _13490_);
  nor (_13493_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand (_13494_, _23553_, _23268_);
  nand (_13495_, _13494_, _23493_);
  nor (_06285_, _13495_, _13493_);
  nor (_13496_, _23553_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nand (_13497_, _23553_, _23154_);
  nand (_13498_, _13497_, _23493_);
  nor (_06288_, _13498_, _13496_);
  nor (_13499_, _21938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  nor (_13500_, _21940_, _21554_);
  nor (_06296_, _13500_, _13499_);
  nor (_13501_, _21938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  nor (_13502_, _21940_, _21526_);
  nor (_06299_, _13502_, _13501_);
  nor (_13503_, _21938_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1]);
  nor (_13504_, _21940_, _21474_);
  nor (_06305_, _13504_, _13503_);
  nor (_13505_, _21882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  nor (_13506_, _21884_, _21526_);
  nor (_25225_, _13506_, _13505_);
  nor (_13507_, _21882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  nor (_13508_, _21884_, _21414_);
  nor (_06318_, _13508_, _13507_);
  nor (_13509_, _21882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  nor (_13510_, _21884_, _21554_);
  nor (_06331_, _13510_, _13509_);
  nor (_13511_, _21882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  nor (_13512_, _21884_, _21586_);
  nor (_06340_, _13512_, _13511_);
  nor (_06350_, _12463_, rst);
  nor (_06354_, _12468_, rst);
  nor (_06357_, _12455_, rst);
  nor (_13513_, _21761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  nor (_13514_, _21763_, _21586_);
  nor (_06360_, _13514_, _13513_);
  nor (_13515_, _21761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1]);
  nor (_13517_, _21763_, _21474_);
  nor (_06369_, _13517_, _13515_);
  nor (_13518_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_13519_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand (_13520_, _13519_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand (_13521_, _13520_, _23493_);
  nor (_06374_, _13521_, _13518_);
  nor (_13522_, _23139_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_13523_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nor (_13524_, _13523_, _06011_);
  nor (_13525_, _13524_, _13522_);
  nor (_25040_[5], _13525_, rst);
  nor (_13526_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_13527_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand (_13528_, _13527_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand (_13529_, _13528_, _23493_);
  nor (_06380_, _13529_, _13526_);
  nor (_13530_, _23197_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_13531_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nor (_13532_, _13531_, _06011_);
  nor (_13533_, _13532_, _13530_);
  nor (_25040_[3], _13533_, rst);
  nor (_13534_, _23223_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_13535_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nor (_13536_, _13535_, _06011_);
  nor (_13537_, _13536_, _13534_);
  nor (_06386_, _13537_, rst);
  nor (_13538_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_13539_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand (_13540_, _13539_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nand (_13541_, _13540_, _23493_);
  nor (_06389_, _13541_, _13538_);
  nor (_13542_, _23557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  nor (_13543_, _23560_, _21414_);
  nor (_06399_, _13543_, _13542_);
  nor (_13544_, _23151_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_13545_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nor (_13546_, _13545_, _06011_);
  nor (_13547_, _13546_, _13544_);
  nor (_06402_, _13547_, rst);
  nor (_13548_, _21882_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7]);
  nor (_13549_, _21884_, _21626_);
  nor (_06408_, _13549_, _13548_);
  nor (_13550_, _22198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  nor (_13551_, _22200_, _21586_);
  nor (_06416_, _13551_, _13550_);
  nor (_13552_, _21761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5]);
  nor (_13553_, _21763_, _21451_);
  nor (_06422_, _13553_, _13552_);
  nor (_13554_, _22198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  nor (_13556_, _22200_, _21554_);
  nor (_25193_, _13556_, _13554_);
  nand (_13557_, _24423_, _23499_);
  not (_13558_, _13557_);
  nor (_13559_, _11943_, _13558_);
  nor (_13560_, _13559_, _11658_);
  nand (_13561_, _12031_, _11904_);
  not (_13562_, _11934_);
  nor (_13563_, _13562_, _00619_);
  nor (_13564_, _24512_, _12157_);
  nor (_13565_, _13564_, _13563_);
  nand (_13566_, _13565_, _13561_);
  nor (_13567_, _13566_, _13560_);
  nor (_13568_, _24460_, _24397_);
  nand (_13569_, _13568_, _24485_);
  nand (_13570_, _13569_, _11917_);
  nand (_13571_, _13570_, _11933_);
  not (_13572_, _13571_);
  nor (_13573_, _12035_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_13574_, _13573_, _12037_);
  nand (_13575_, _13574_, _13572_);
  nand (_13576_, _13575_, _13567_);
  nor (_13577_, _13576_, _11879_);
  nand (_13578_, _11879_, _12157_);
  nand (_13579_, _13578_, _23493_);
  nor (_06432_, _13579_, _13577_);
  nor (_13580_, _13562_, _24841_);
  not (_13581_, _11904_);
  nor (_13582_, _13581_, _05381_);
  nor (_13583_, _13582_, _13580_);
  not (_13584_, _13559_);
  nand (_13585_, _13584_, ABINPUT[20]);
  nand (_13586_, _24432_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nand (_13587_, _13586_, _13585_);
  nor (_13588_, _12044_, _12037_);
  nand (_13589_, _13572_, _12045_);
  nor (_13590_, _13589_, _13588_);
  nor (_13591_, _13590_, _13587_);
  nand (_13592_, _13591_, _13583_);
  nor (_13593_, _13592_, _11879_);
  nand (_13594_, _11879_, _12155_);
  nand (_13595_, _13594_, _23493_);
  nor (_06435_, _13595_, _13593_);
  nor (_13596_, _21873_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  nor (_13597_, _21875_, _21586_);
  nor (_06438_, _13597_, _13596_);
  nor (_13598_, _13562_, _00517_);
  nor (_13599_, _13581_, _07031_);
  nor (_13600_, _13599_, _13598_);
  nand (_13601_, _13584_, ABINPUT[21]);
  nand (_13603_, _24432_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nand (_13604_, _13603_, _13601_);
  nand (_13605_, _12041_, _12038_);
  nand (_13606_, _13605_, _12009_);
  nor (_13607_, _13606_, _12036_);
  nor (_13608_, _13607_, _12042_);
  not (_13609_, _12048_);
  nand (_13610_, _13609_, _13608_);
  nand (_13611_, _13610_, _12049_);
  nor (_13612_, _13611_, _13571_);
  nor (_13613_, _13612_, _13604_);
  nand (_13614_, _13613_, _13600_);
  nor (_13615_, _13614_, _11879_);
  not (_13616_, _06017_);
  nand (_13617_, _11879_, _13616_);
  nand (_13618_, _13617_, _23493_);
  nor (_06441_, _13618_, _13615_);
  nor (_13619_, _13562_, _00455_);
  nor (_13620_, _13609_, _13608_);
  nor (_13621_, _13620_, _12002_);
  nand (_13623_, _11994_, _11992_);
  nand (_13624_, _13623_, _13621_);
  nor (_13625_, _13623_, _13621_);
  nor (_13626_, _13625_, _13571_);
  nand (_13627_, _13626_, _13624_);
  nor (_13628_, _13581_, _10398_);
  nand (_13629_, _13584_, ABINPUT[22]);
  nand (_13630_, _24432_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nand (_13631_, _13630_, _13629_);
  nor (_13632_, _13631_, _13628_);
  nand (_13633_, _13632_, _13627_);
  nor (_13634_, _13633_, _13619_);
  nor (_13635_, _13634_, _11879_);
  not (_13636_, _06009_);
  nor (_13637_, _11903_, _13636_);
  nor (_13638_, _13637_, _13635_);
  nor (_06453_, _13638_, rst);
  nor (_13639_, _12055_, _12052_);
  nand (_13640_, _12101_, _12056_);
  nor (_13641_, _13640_, _13639_);
  nand (_13643_, _13584_, ABINPUT[23]);
  nor (_13644_, _13581_, _24191_);
  nand (_13645_, _11934_, _11979_);
  nand (_13646_, _24811_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nand (_13647_, _13646_, _13645_);
  nor (_13648_, _13647_, _13644_);
  nand (_13649_, _13648_, _13643_);
  nor (_13650_, _13649_, _13641_);
  nor (_13651_, _13650_, _11879_);
  nand (_13652_, _12112_, _06005_);
  not (_13654_, _06007_);
  nand (_13655_, _13654_, _12111_);
  nand (_13656_, _13655_, _13652_);
  nor (_13657_, _13656_, _11903_);
  nor (_13658_, _13657_, _13651_);
  nor (_06456_, _13658_, rst);
  nor (_13659_, _13621_, _11993_);
  nor (_13660_, _13659_, _11991_);
  not (_13661_, _12055_);
  nor (_13662_, _13661_, _13660_);
  nor (_13663_, _13662_, _11983_);
  nand (_13664_, _11975_, _11973_);
  nor (_13665_, _13664_, _13663_);
  nand (_13666_, _13664_, _13663_);
  nand (_13667_, _13666_, _12101_);
  nor (_13668_, _13667_, _13665_);
  nand (_13669_, _13584_, ABINPUT[24]);
  nor (_13670_, _13581_, _01352_);
  nand (_13671_, _11934_, _11967_);
  nand (_13672_, _24811_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nand (_13673_, _13672_, _13671_);
  nor (_13674_, _13673_, _13670_);
  nand (_13675_, _13674_, _13669_);
  nor (_13676_, _13675_, _13668_);
  nor (_13677_, _13676_, _11879_);
  nor (_13678_, _12115_, _23553_);
  not (_13679_, _13678_);
  nand (_13680_, _13652_, _12212_);
  nand (_13681_, _13680_, _13679_);
  nor (_13682_, _13681_, _11903_);
  nor (_13683_, _13682_, _13677_);
  nor (_06459_, _13683_, rst);
  nor (_13684_, _13562_, _00380_);
  nor (_13685_, _13581_, _02307_);
  nor (_13686_, _13685_, _13684_);
  nand (_13687_, _13584_, ABINPUT[25]);
  nand (_13688_, _24432_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nand (_13689_, _13688_, _13687_);
  not (_13690_, _11963_);
  nor (_13691_, _13663_, _11974_);
  nor (_13692_, _13691_, _11972_);
  nand (_13693_, _13692_, _13690_);
  nand (_13694_, _13693_, _12060_);
  nor (_13695_, _13694_, _13571_);
  nor (_13696_, _13695_, _13689_);
  nand (_13697_, _13696_, _13686_);
  nor (_13698_, _13697_, _11879_);
  nor (_13699_, _13679_, _12208_);
  not (_13700_, _13699_);
  nand (_13701_, _13679_, _12208_);
  nand (_13702_, _13701_, _13700_);
  nand (_13703_, _13702_, _11879_);
  nand (_13704_, _13703_, _23493_);
  nor (_06463_, _13704_, _13698_);
  nor (_13705_, _12063_, _11952_);
  nor (_13706_, _13692_, _13690_);
  nor (_13707_, _13706_, _11961_);
  not (_13708_, _13707_);
  nor (_13709_, _13708_, _13705_);
  nand (_13710_, _13708_, _13705_);
  nand (_13711_, _13710_, _12101_);
  nor (_13712_, _13711_, _13709_);
  nor (_13713_, _13559_, _11588_);
  nand (_13714_, _11934_, _00074_);
  nor (_13715_, _13581_, _11772_);
  nor (_13716_, _24512_, _12110_);
  nor (_13717_, _13716_, _13715_);
  nand (_13718_, _13717_, _13714_);
  nor (_13719_, _13718_, _13713_);
  nand (_13720_, _13719_, _11903_);
  nor (_13721_, _13720_, _13712_);
  nor (_13722_, _13700_, _12110_);
  not (_13723_, _13722_);
  nand (_13724_, _13700_, _12110_);
  nand (_13725_, _13724_, _13723_);
  nand (_13726_, _13725_, _11879_);
  nand (_13727_, _13726_, _23493_);
  nor (_25034_[7], _13727_, _13721_);
  nand (_13728_, _11904_, _00620_);
  nor (_13729_, _12066_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not (_13731_, _12064_);
  nor (_13732_, _13731_, _13706_);
  nor (_13733_, _13732_, _11952_);
  nor (_13734_, _13733_, _12076_);
  nor (_13735_, _13734_, _13729_);
  nor (_13736_, _13735_, _12062_);
  nand (_13737_, _13735_, _12062_);
  nand (_13738_, _13737_, _13572_);
  nor (_13739_, _13738_, _13736_);
  not (_13740_, _11943_);
  nor (_13741_, _13740_, _12109_);
  nor (_13742_, _24431_, _11658_);
  nor (_13743_, _13742_, _13741_);
  nor (_13744_, _13562_, _00697_);
  nor (_13745_, _13557_, _11656_);
  nor (_13746_, _13745_, _13744_);
  nand (_13747_, _13746_, _13743_);
  nor (_13748_, _13747_, _13739_);
  nand (_13749_, _13748_, _13728_);
  nor (_13750_, _13749_, _11879_);
  nand (_13751_, _13722_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nand (_13752_, _13723_, _12109_);
  nand (_13753_, _13752_, _13751_);
  nand (_13754_, _13753_, _11879_);
  nand (_13755_, _13754_, _23493_);
  nor (_06467_, _13755_, _13750_);
  nor (_13756_, _12066_, _12076_);
  nand (_13757_, _13756_, _12062_);
  nor (_13758_, _13733_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nand (_13759_, _13758_, _11951_);
  nand (_13761_, _13759_, _13757_);
  nor (_13762_, _13761_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_13763_, _13761_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_13764_, _13763_, _12101_);
  nor (_13765_, _13764_, _13762_);
  nor (_13766_, _13740_, _12198_);
  nor (_13767_, _24431_, _10818_);
  nor (_13768_, _13767_, _13766_);
  nand (_13769_, _11929_, ABINPUT[12]);
  nand (_13770_, _13769_, _13768_);
  nand (_13771_, _11934_, _23115_);
  nand (_13772_, _11904_, _12006_);
  nand (_13773_, _13772_, _13771_);
  nor (_13774_, _13773_, _13770_);
  nand (_13775_, _13774_, _11903_);
  nor (_13776_, _13775_, _13765_);
  nor (_13777_, _12120_, _23553_);
  not (_13778_, _13777_);
  nand (_13779_, _13751_, _12198_);
  nand (_13780_, _13779_, _13778_);
  nand (_13781_, _13780_, _11879_);
  nand (_13782_, _13781_, _23493_);
  nor (_06470_, _13782_, _13776_);
  nor (_13783_, _12077_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_13784_, _13783_, _11951_);
  nand (_13785_, _12068_, _12062_);
  nand (_13786_, _13785_, _13784_);
  nor (_13787_, _13786_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand (_13788_, _13786_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand (_13789_, _13788_, _12101_);
  nor (_13791_, _13789_, _13787_);
  nand (_13792_, _11904_, _11998_);
  nor (_13793_, _24512_, _10847_);
  not (_13794_, ABINPUT[13]);
  nor (_13795_, _11906_, _13794_);
  nor (_13796_, _13795_, _13793_);
  nand (_13797_, _13796_, _13792_);
  nand (_13798_, _11934_, _23400_);
  nand (_13799_, _11943_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nand (_13800_, _13799_, _13798_);
  nor (_13801_, _13800_, _13797_);
  nand (_13802_, _13801_, _11903_);
  nor (_13803_, _13802_, _13791_);
  nor (_13804_, _13778_, _12108_);
  not (_13805_, _13804_);
  nand (_13806_, _13778_, _12108_);
  nand (_13807_, _13806_, _13805_);
  nand (_13808_, _13807_, _11879_);
  nand (_13809_, _13808_, _23493_);
  nor (_06472_, _13809_, _13803_);
  not (_13811_, _12069_);
  nand (_13812_, _13811_, _12062_);
  nand (_13813_, _12081_, _11951_);
  nand (_13814_, _13813_, _13812_);
  nor (_13815_, _13814_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand (_13816_, _13814_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand (_13817_, _13816_, _12101_);
  nor (_13818_, _13817_, _13815_);
  nand (_13819_, _11943_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_13820_, _24512_, _10833_);
  nor (_13821_, _11906_, _11685_);
  nor (_13822_, _13821_, _13820_);
  nand (_13823_, _13822_, _13819_);
  nand (_13824_, _11904_, _00456_);
  nand (_13825_, _11934_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand (_13826_, _13825_, _13824_);
  nor (_13827_, _13826_, _13823_);
  nand (_13828_, _13827_, _11903_);
  nor (_13829_, _13828_, _13818_);
  nand (_13830_, _13804_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand (_13831_, _13805_, _12189_);
  nand (_13832_, _13831_, _13830_);
  nand (_13833_, _13832_, _11879_);
  nand (_13834_, _13833_, _23493_);
  nor (_06475_, _13834_, _13829_);
  not (_13835_, _12073_);
  nand (_13836_, _12083_, _13835_);
  nor (_13837_, _13836_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_13838_, _13836_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_13839_, _13838_, _12101_);
  nor (_13840_, _13839_, _13837_);
  nor (_13841_, _13581_, _00175_);
  nor (_13842_, _11926_, _12107_);
  nand (_13843_, _13842_, _11917_);
  nor (_13844_, _24512_, _10878_);
  nor (_13845_, _11906_, _11712_);
  nor (_13846_, _13845_, _13844_);
  nand (_13847_, _13846_, _13843_);
  nor (_13848_, _13847_, _13841_);
  nand (_13849_, _13848_, _11903_);
  nor (_13850_, _13849_, _13840_);
  nor (_13851_, _12108_, _12189_);
  nand (_13852_, _13851_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_13853_, _13852_, _13778_);
  not (_13854_, _13853_);
  nand (_13855_, _13830_, _12107_);
  nand (_13856_, _13855_, _13854_);
  nand (_13857_, _13856_, _11879_);
  nand (_13858_, _13857_, _23493_);
  nor (_06478_, _13858_, _13850_);
  nor (_13859_, _21757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  nor (_13860_, _21759_, _21586_);
  nor (_06480_, _13860_, _13859_);
  nor (_13861_, _12086_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_13862_, _12086_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_13863_, _13862_, _12101_);
  nor (_13864_, _13863_, _13861_);
  nor (_13865_, _13581_, _00301_);
  nor (_13866_, _11926_, _12106_);
  nand (_13867_, _13866_, _11917_);
  not (_13868_, ABINPUT[16]);
  nor (_13869_, _11906_, _13868_);
  nor (_13870_, _24512_, _10863_);
  nor (_13871_, _13870_, _13869_);
  nand (_13872_, _13871_, _13867_);
  nor (_13873_, _13872_, _13865_);
  nand (_13874_, _13873_, _11903_);
  nor (_13875_, _13874_, _13864_);
  nand (_13876_, _13853_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_13877_, _12124_, _12106_);
  nand (_13879_, _13877_, _13876_);
  nand (_13880_, _13879_, _11879_);
  nand (_13881_, _13880_, _23493_);
  nor (_06484_, _13881_, _13875_);
  nor (_13882_, _21877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7]);
  nor (_13883_, _21880_, _21626_);
  nor (_06486_, _13883_, _13882_);
  nor (_13884_, _13581_, _00380_);
  nand (_13885_, _11943_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_13886_, _24432_, ABINPUT[25]);
  nand (_13887_, _13886_, _13885_);
  nor (_13888_, _13887_, _13884_);
  nand (_13889_, _12091_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_13890_, _12074_);
  nor (_13891_, _12084_, _13890_);
  not (_13892_, _12090_);
  nor (_13893_, _13892_, _13891_);
  nand (_13894_, _13893_, _12092_);
  nand (_13895_, _13894_, _13889_);
  nand (_13896_, _13895_, _13572_);
  nand (_13897_, _13896_, _13888_);
  nor (_13898_, _13562_, _12105_);
  nor (_13899_, _13557_, _11725_);
  nor (_13900_, _13899_, _13898_);
  nand (_13901_, _13900_, _11903_);
  nor (_13902_, _13901_, _13897_);
  nand (_13903_, _13876_, _12105_);
  nand (_13904_, _13903_, _12130_);
  nand (_13905_, _13904_, _11879_);
  nand (_13906_, _13905_, _23493_);
  nor (_06488_, _13906_, _13902_);
  nor (_13907_, _02439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  nor (_13908_, _02442_, _21526_);
  nor (_06496_, _13908_, _13907_);
  nor (_13909_, _21757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  nor (_13910_, _21759_, _21526_);
  nor (_06500_, _13910_, _13909_);
  nor (_13911_, _21757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  nor (_13912_, _21759_, _21554_);
  nor (_06503_, _13912_, _13911_);
  nor (_13913_, _21757_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1]);
  nor (_13914_, _21759_, _21474_);
  nor (_06515_, _13914_, _13913_);
  not (_13915_, _12330_);
  nand (_13916_, _12329_, _12326_);
  nand (_13917_, _13916_, _13915_);
  nand (_13918_, _13917_, _24823_);
  nor (_13919_, _24823_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_13920_, _13919_, _12373_);
  nand (_13921_, _13920_, _13918_);
  nand (_13922_, _12135_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  nand (_06518_, _13922_, _13921_);
  nand (_13923_, _12332_, _13915_);
  nand (_13924_, _13923_, _12334_);
  nand (_13925_, _13924_, _24823_);
  nor (_13926_, _24823_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_13927_, _13926_, _12373_);
  nand (_13928_, _13927_, _13925_);
  nand (_13929_, _12135_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nand (_06521_, _13929_, _13928_);
  nor (_13931_, _12343_, _12335_);
  nand (_13932_, _12343_, _12335_);
  nand (_13933_, _13932_, _24823_);
  nor (_13934_, _13933_, _13931_);
  nand (_13935_, _24824_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_13936_, _13935_, _23038_);
  nor (_13937_, _13936_, _13934_);
  nand (_13938_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _06003_);
  nand (_13939_, _13938_, _23493_);
  nor (_06523_, _13939_, _13937_);
  nand (_13940_, _13932_, _12339_);
  nand (_13941_, _13940_, _12346_);
  nand (_13942_, _13941_, _24823_);
  nor (_13943_, _24823_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_13944_, _13943_, _12373_);
  nand (_13945_, _13944_, _13942_);
  nand (_13946_, _12135_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nand (_06525_, _13946_, _13945_);
  nor (_13947_, _22781_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  nor (_13948_, _22783_, _21586_);
  nor (_25126_, _13948_, _13947_);
  not (_13950_, _12353_);
  nand (_13951_, _12352_, _12346_);
  nand (_13952_, _13951_, _13950_);
  nand (_13953_, _13952_, _24823_);
  nor (_13954_, _24823_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_13955_, _13954_, _12373_);
  nand (_13956_, _13955_, _13953_);
  nand (_13957_, _12135_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nand (_06528_, _13957_, _13956_);
  nor (_13958_, _21877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1]);
  nor (_13959_, _21880_, _21474_);
  nor (_06530_, _13959_, _13958_);
  nand (_13960_, _13950_, _12215_);
  nand (_13961_, _13960_, _12354_);
  nand (_13962_, _13961_, _24823_);
  nor (_13963_, _24823_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_13964_, _13963_, _12373_);
  nand (_13965_, _13964_, _13962_);
  nand (_13966_, _12135_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nand (_06532_, _13966_, _13965_);
  not (_13967_, _12211_);
  not (_13968_, _12354_);
  nor (_13969_, _13968_, _13967_);
  not (_13970_, _12355_);
  nand (_13971_, _13970_, _24823_);
  nor (_13972_, _13971_, _13969_);
  nand (_13973_, _24824_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nand (_13974_, _13973_, _23038_);
  nor (_13975_, _13974_, _13972_);
  nand (_13977_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _12208_);
  nand (_13978_, _13977_, _23493_);
  nor (_06537_, _13978_, _13975_);
  nor (_13979_, _21877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  nor (_13980_, _21880_, _21586_);
  nor (_06540_, _13980_, _13979_);
  nor (_13981_, _12355_, _12207_);
  nand (_13982_, _12356_, _24823_);
  nor (_13983_, _13982_, _13981_);
  nand (_13984_, _24824_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_13985_, _13984_, _23038_);
  nor (_13986_, _13985_, _13983_);
  nand (_13987_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _12110_);
  nand (_13988_, _13987_, _23493_);
  nor (_06542_, _13988_, _13986_);
  nand (_13989_, _12358_, _12356_);
  nand (_13990_, _13989_, _24823_);
  nor (_13991_, _13990_, _12359_);
  nand (_13992_, _24824_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nand (_13993_, _13992_, _23038_);
  nor (_13994_, _13993_, _13991_);
  nand (_13995_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _12109_);
  nand (_13996_, _13995_, _23493_);
  nor (_06545_, _13996_, _13994_);
  nand (_13997_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _12198_);
  nand (_13998_, _13997_, _23493_);
  nor (_13999_, _12359_, _12202_);
  nand (_14000_, _12360_, _24823_);
  nor (_14001_, _14000_, _13999_);
  nand (_14002_, _24824_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_14003_, _14002_, _23038_);
  nor (_14004_, _14003_, _14001_);
  nor (_06548_, _14004_, _13998_);
  nand (_14005_, _12135_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  not (_14006_, _12361_);
  nand (_14007_, _12360_, _12197_);
  nand (_14008_, _14007_, _14006_);
  nand (_14009_, _14008_, _24823_);
  nor (_14010_, _24823_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_14011_, _14010_, _12373_);
  nand (_14012_, _14011_, _14009_);
  nand (_06550_, _14012_, _14005_);
  nand (_14013_, _12135_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand (_14014_, _14006_, _12193_);
  nand (_14015_, _14014_, _12362_);
  nand (_14016_, _14015_, _24823_);
  nor (_14017_, _24823_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_14018_, _14017_, _12373_);
  nand (_14019_, _14018_, _14016_);
  nand (_06552_, _14019_, _14013_);
  nand (_14020_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _12107_);
  nand (_14021_, _14020_, _23493_);
  nand (_14022_, _12362_, _12188_);
  nand (_14023_, _14022_, _24823_);
  nor (_14024_, _14023_, _12363_);
  nand (_14025_, _24824_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_14026_, _14025_, _23038_);
  nor (_14027_, _14026_, _14024_);
  nor (_06554_, _14027_, _14021_);
  not (_14028_, _12186_);
  not (_14029_, _12363_);
  nand (_14030_, _14029_, _14028_);
  nand (_14031_, _14030_, _12364_);
  nand (_14032_, _14031_, _24823_);
  nor (_14033_, _24823_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_14034_, _14033_, _12373_);
  nand (_14035_, _14034_, _14032_);
  nand (_14036_, _12135_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nand (_06559_, _14036_, _14035_);
  not (_14037_, _12364_);
  nor (_14038_, _14037_, _12180_);
  nand (_14039_, _12366_, _24823_);
  nor (_14040_, _14039_, _14038_);
  nand (_14041_, _24824_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_14042_, _14041_, _23038_);
  nor (_14043_, _14042_, _14040_);
  nand (_14044_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _12105_);
  nand (_14045_, _14044_, _23493_);
  nor (_06560_, _14045_, _14043_);
  nor (_14046_, _21877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  nor (_14047_, _21880_, _21414_);
  nor (_25233_, _14047_, _14046_);
  nor (_14048_, _21877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  nor (_14049_, _21880_, _21526_);
  nor (_06567_, _14049_, _14048_);
  nor (_14050_, _21877_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  nor (_14051_, _21880_, _21554_);
  nor (_25232_, _14051_, _14050_);
  nor (_14052_, _12387_, _12013_);
  nor (_14053_, _14052_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  nor (_06580_, _14053_, rst);
  nor (_14054_, _21933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  nor (_14055_, _21935_, _21526_);
  nor (_06582_, _14055_, _14054_);
  nor (_14056_, _12387_, _05364_);
  nor (_14057_, _14056_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  nor (_06584_, _14057_, rst);
  nand (_14058_, _23493_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  nor (_14059_, rst, _07012_);
  nand (_14060_, _14059_, _12386_);
  nand (_06586_, _14060_, _14058_);
  nor (_14061_, _21933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  nor (_14062_, _21935_, _21554_);
  nor (_06588_, _14062_, _14061_);
  nor (_14063_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  nor (_14064_, _22563_, _21526_);
  nor (_06594_, _14064_, _14063_);
  nor (_14065_, _10753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5]);
  nor (_14066_, _10755_, _21451_);
  nor (_06602_, _14066_, _14065_);
  nor (_14067_, _21865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6]);
  nor (_14068_, _21867_, _21504_);
  nor (_06623_, _14068_, _14067_);
  nor (_14069_, _21865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5]);
  nor (_14070_, _21867_, _21451_);
  nor (_25247_, _14070_, _14069_);
  nor (_14071_, _21869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  nor (_14072_, _21871_, _21554_);
  nor (_06656_, _14072_, _14071_);
  nand (_14073_, _01143_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nand (_14075_, _01142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nand (_14076_, _14075_, _14073_);
  nor (_14077_, _14076_, _01130_);
  nor (_14078_, _01059_, _24900_);
  nor (_14079_, _01055_, _24867_);
  nor (_14080_, _14079_, _14078_);
  nand (_14081_, _14080_, _01130_);
  nand (_14082_, _14081_, _23493_);
  nor (_06662_, _14082_, _14077_);
  nor (_14083_, _10753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7]);
  nor (_14084_, _10755_, _21626_);
  nor (_06665_, _14084_, _14083_);
  nor (_14085_, _21632_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6]);
  nor (_14086_, _21635_, _21504_);
  nor (_06677_, _14086_, _14085_);
  nand (_14087_, _01017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand (_14088_, _01020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nand (_14089_, _14088_, _14087_);
  nor (_14090_, _14089_, _01030_);
  nor (_14091_, _01032_, ABINPUT[9]);
  nor (_14092_, _14091_, _14090_);
  nor (_14093_, _14092_, _01037_);
  nand (_14094_, _01037_, _10689_);
  nand (_14095_, _14094_, _23493_);
  nor (_06681_, _14095_, _14093_);
  nor (_14096_, _21761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  nor (_14097_, _21763_, _21526_);
  nor (_06697_, _14097_, _14096_);
  nor (_14098_, _22198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  nor (_14099_, _22200_, _21414_);
  nor (_06707_, _14099_, _14098_);
  nor (_14100_, _21761_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6]);
  nor (_14101_, _21763_, _21504_);
  nor (_06713_, _14101_, _14100_);
  nor (_14102_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6]);
  nor (_14103_, _22130_, _21504_);
  nor (_06717_, _14103_, _14102_);
  nor (_14104_, _24380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  nor (_14105_, _24382_, _21414_);
  nor (_06722_, _14105_, _14104_);
  nand (_14106_, _05674_, _05568_);
  nor (_14107_, _14106_, _05658_);
  nand (_14108_, _05680_, _05606_);
  nand (_14109_, _14108_, _23493_);
  nor (_06724_, _14109_, _14107_);
  nor (_14110_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5]);
  nor (_14111_, _22130_, _21451_);
  nor (_06728_, _14111_, _14110_);
  nor (_14112_, _05634_, _05617_);
  nor (_14113_, _05674_, _05658_);
  not (_14114_, _14113_);
  nor (_14115_, _14114_, _05670_);
  nor (_14116_, _14115_, _14112_);
  nor (_14117_, _05606_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_14118_, _14117_);
  nor (_14119_, _14118_, _14116_);
  not (_14120_, _05659_);
  nor (_14121_, _05663_, _14120_);
  not (_14122_, _05664_);
  nor (_14123_, _14122_, _14120_);
  nor (_14125_, _14123_, _14121_);
  nand (_14126_, _14125_, _05679_);
  not (_14127_, _14112_);
  nor (_14128_, _14127_, _05656_);
  nor (_14129_, _14128_, _14118_);
  nand (_14130_, _14129_, _14126_);
  nand (_14131_, _14130_, _05582_);
  nand (_14132_, _14131_, _23493_);
  nor (_06730_, _14132_, _14119_);
  nor (_14133_, _05606_, _05571_);
  not (_14134_, _14133_);
  nor (_14135_, _14134_, _14116_);
  nor (_14136_, _14134_, _14128_);
  nand (_14137_, _14136_, _14126_);
  nand (_14138_, _14137_, _05580_);
  nand (_14139_, _14138_, _23493_);
  nor (_06732_, _14139_, _14135_);
  nor (_14140_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  nor (_14141_, _22130_, _21414_);
  nor (_06737_, _14141_, _14140_);
  nor (_14142_, _23545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7]);
  nor (_14143_, _23547_, _21626_);
  nor (_06744_, _14143_, _14142_);
  nor (_14144_, _23545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6]);
  nor (_14145_, _23547_, _21504_);
  nor (_06749_, _14145_, _14144_);
  nor (_14146_, _22396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1]);
  nor (_14147_, _22398_, _21474_);
  nor (_06764_, _14147_, _14146_);
  nor (_14148_, _21865_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  nor (_14149_, _21867_, _21586_);
  nor (_06779_, _14149_, _14148_);
  nor (_14150_, _21869_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1]);
  nor (_14151_, _21871_, _21474_);
  nor (_25239_, _14151_, _14150_);
  nor (_14152_, _10753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  nor (_14153_, _10755_, _21526_);
  nor (_06788_, _14153_, _14152_);
  nor (_14154_, _22396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  nor (_14155_, _22398_, _21554_);
  nor (_06790_, _14155_, _14154_);
  nor (_14156_, _10753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  nor (_14157_, _10755_, _21554_);
  nor (_06795_, _14157_, _14156_);
  nor (_14158_, _10753_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1]);
  nor (_14159_, _10755_, _21474_);
  nor (_06799_, _14159_, _14158_);
  not (_14160_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_14161_, _05559_, _02484_);
  nor (_14162_, _14161_, _14160_);
  nand (_14163_, _14161_, ABINPUT[0]);
  nand (_14164_, _14163_, _02394_);
  nor (_14165_, _14164_, _14162_);
  nand (_14166_, _02393_, _00106_);
  nand (_14167_, _14166_, _23493_);
  nor (_06808_, _14167_, _14165_);
  nor (_14168_, _22454_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7]);
  nor (_14169_, _22456_, _21626_);
  nor (_06813_, _14169_, _14168_);
  nor (_14170_, _10776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  nor (_14172_, _10778_, _21554_);
  nor (_06828_, _14172_, _14170_);
  nor (_14173_, _05742_, _01127_);
  nand (_14174_, _14173_, _00912_);
  nor (_14175_, _14174_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  not (_14176_, _01135_);
  nand (_14177_, _14176_, _02333_);
  not (_14178_, _01140_);
  nand (_14179_, _02347_, _14178_);
  nor (_14180_, _14179_, _14177_);
  nand (_14181_, _14180_, _02341_);
  nor (_14182_, _02349_, _01131_);
  nand (_14183_, _14182_, _14181_);
  nor (_14184_, _14183_, _14175_);
  nor (_14185_, _14184_, _14175_);
  nor (_06832_, _14185_, rst);
  nor (_14186_, _05559_, _05076_);
  nand (_14187_, _14186_, _24861_);
  nor (_14188_, _14187_, ABINPUT[10]);
  not (_14189_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_14191_, _14187_, _14189_);
  nand (_14192_, _14191_, _23493_);
  nor (_06835_, _14192_, _14188_);
  nand (_14193_, _01142_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_14194_, _14193_, _01130_);
  nor (_14195_, _02360_, _14160_);
  nor (_14196_, _14195_, _14194_);
  nor (_06837_, _14196_, rst);
  nand (_14197_, _10295_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nor (_14198_, _10295_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nor (_14199_, _14198_, rst);
  nand (_14200_, _14199_, _14197_);
  nor (_06840_, _14200_, _01130_);
  not (_14201_, _02349_);
  nand (_14202_, _14178_, _14176_);
  nand (_14203_, _14202_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nand (_14204_, _14203_, _14181_);
  nor (_14205_, _01134_, _01131_);
  nand (_14206_, _14205_, _14204_);
  nand (_14207_, _14206_, _14201_);
  nand (_14208_, _14207_, _23493_);
  nor (_06843_, _14208_, _01130_);
  nor (_14209_, _05566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  nor (_14210_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _14160_);
  nor (_14211_, _06708_, _01090_);
  nor (_14212_, _14211_, _14210_);
  not (_14213_, _14212_);
  nor (_14214_, _14213_, _14209_);
  nor (_14215_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor (_14216_, _14215_, _14214_);
  nor (_14217_, _14216_, _14214_);
  nor (_14218_, _14217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_14219_, _14216_, _14189_);
  nand (_14220_, _14219_, _23493_);
  nor (_06852_, _14220_, _14218_);
  not (_14221_, _14216_);
  nor (_06855_, _14221_, rst);
  nand (_14222_, _01052_, _03984_);
  nand (_14223_, _14222_, _23493_);
  not (_14224_, _01078_);
  nor (_14226_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nor (_14227_, _14226_, _14224_);
  nor (_14228_, _14227_, _01071_);
  nand (_14229_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  nor (_14230_, _14229_, _01071_);
  nor (_14231_, _14230_, rxd_i);
  nor (_14232_, _14231_, _14228_);
  nor (_14233_, _01083_, _03984_);
  nor (_14234_, _14233_, _14232_);
  nor (_06857_, _14234_, _14223_);
  not (_14235_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_14236_, _01080_, _14235_);
  nand (_14237_, _01052_, _01060_);
  nor (_14238_, _14237_, _01055_);
  nand (_14239_, _14238_, _01072_);
  nand (_14240_, _14239_, _14236_);
  nand (_06863_, _14240_, _03985_);
  nand (_14241_, _02413_, _01073_);
  nor (_14242_, _02408_, _14241_);
  nand (_14243_, _14242_, _23493_);
  nand (_14244_, _02420_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nand (_06866_, _14244_, _14243_);
  nor (_14245_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7]);
  nor (_14246_, _22130_, _21626_);
  nor (_06867_, _14246_, _14245_);
  nand (_14247_, _07248_, _01074_);
  nor (_14248_, _02408_, _14247_);
  nor (_14249_, _14248_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  not (_14250_, rxd_i);
  nand (_14251_, _14248_, _14250_);
  nand (_14253_, _14251_, _23493_);
  nor (_06870_, _14253_, _14249_);
  nor (_14254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _01060_);
  nand (_14255_, _01059_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_14256_, _14255_, _14254_);
  nand (_14257_, _14256_, _01072_);
  nand (_14258_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor (_14259_, _14257_, _14250_);
  nor (_14260_, _14259_, rst);
  nand (_06872_, _14260_, _14258_);
  nor (_14261_, _10776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  nor (_14262_, _10778_, _21526_);
  nor (_25285_, _14262_, _14261_);
  nor (_14263_, _22396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  nor (_14264_, _22398_, _21526_);
  nor (_06917_, _14264_, _14263_);
  nor (_14265_, _02481_, _00018_);
  not (_14266_, _14265_);
  nor (_14267_, _14266_, _05055_);
  nor (_14268_, _14267_, _02614_);
  nand (_14269_, _14265_, _05056_);
  nand (_14270_, _14269_, _05599_);
  nor (_14271_, _14270_, _14268_);
  nand (_14272_, _05598_, _00114_);
  nand (_14273_, _14272_, _23493_);
  nor (_06921_, _14273_, _14271_);
  nor (_14274_, _00008_, _21772_);
  not (_14275_, _14274_);
  nor (_14276_, _14275_, _02481_);
  not (_14277_, _14276_);
  nor (_14278_, _14277_, _05559_);
  nor (_14279_, _14278_, _05610_);
  nor (_14280_, _14275_, _00927_);
  not (_14281_, _14280_);
  nand (_14282_, _14276_, _06626_);
  nand (_14283_, _14282_, _14281_);
  nor (_14284_, _14283_, _14279_);
  nand (_14285_, _14280_, _00106_);
  nand (_14286_, _14285_, _23493_);
  nor (_06930_, _14286_, _14284_);
  nor (_14287_, _10776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6]);
  nor (_14288_, _10778_, _21504_);
  nor (_06944_, _14288_, _14287_);
  nor (_14289_, _10776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5]);
  nor (_14290_, _10778_, _21451_);
  nor (_06953_, _14290_, _14289_);
  not (_14291_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nor (_14292_, _01124_, _21772_);
  nand (_14293_, _14292_, _02480_);
  nor (_14294_, _14293_, _05559_);
  nor (_14295_, _14294_, _14291_);
  nor (_14296_, _14293_, _06627_);
  nor (_14297_, _14296_, _14295_);
  nor (_14298_, _05559_, _04983_);
  nand (_14299_, _14298_, _24861_);
  not (_14300_, _14299_);
  nor (_14301_, _14300_, _14297_);
  nor (_14302_, _14299_, _00106_);
  nor (_14303_, _14302_, _14301_);
  nor (_06965_, _14303_, rst);
  nor (_14304_, _21645_, _21558_);
  nor (_14305_, _14304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5]);
  not (_14306_, _14304_);
  nor (_14307_, _14306_, _21451_);
  nor (_06987_, _14307_, _14305_);
  nor (_14308_, _14304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7]);
  nor (_14309_, _14306_, _21626_);
  nor (_06989_, _14309_, _14308_);
  nor (_14310_, _14304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6]);
  nor (_14311_, _14306_, _21504_);
  nor (_07007_, _14311_, _14310_);
  nor (_14312_, _22021_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  nor (_14313_, _22023_, _21414_);
  nor (_07014_, _14313_, _14312_);
  nand (_14314_, _24617_, _23513_);
  nand (_14315_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nand (_14316_, _14315_, _14314_);
  nand (_14317_, _14316_, _23493_);
  not (_14318_, _23150_);
  nand (_14319_, _23424_, _14318_);
  nand (_14321_, _24490_, _23435_);
  nor (_14322_, _14321_, _14319_);
  nand (_14323_, _14322_, _23411_);
  nand (_14324_, _14323_, _23514_);
  not (_14325_, _24414_);
  nor (_14326_, _14325_, _24406_);
  nor (_14327_, _24489_, _23253_);
  nor (_14328_, _14327_, _24408_);
  not (_14329_, _14328_);
  nor (_14330_, _14329_, _10973_);
  nand (_14331_, _14330_, _14326_);
  not (_14332_, _10988_);
  nor (_14333_, _14332_, _10978_);
  nand (_14334_, _14333_, _10976_);
  nor (_14335_, _23457_, _24483_);
  not (_14336_, _14335_);
  nand (_14337_, _23327_, _23381_);
  nand (_14338_, _14337_, _14336_);
  nor (_14339_, _14338_, _14334_);
  nor (_14340_, _23326_, _23203_);
  nand (_14342_, _24482_, _23088_);
  nor (_14343_, _14342_, _23382_);
  nor (_14344_, _14343_, _14340_);
  nor (_14345_, _24614_, _23457_);
  nand (_14346_, _23405_, _23088_);
  nor (_14347_, _14346_, _23528_);
  nor (_14348_, _14347_, _14345_);
  nand (_14349_, _14348_, _14344_);
  nor (_14350_, _14349_, _23534_);
  nand (_14351_, _14350_, _14339_);
  nor (_14352_, _14351_, _14331_);
  nand (_14353_, _14352_, _14324_);
  nand (_14354_, _14353_, _23491_);
  nand (_25020_[0], _14354_, _14317_);
  nor (_14355_, _10776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1]);
  nor (_14356_, _10778_, _21474_);
  nor (_07050_, _14356_, _14355_);
  nor (_14357_, _10776_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  nor (_14358_, _10778_, _21586_);
  nor (_07060_, _14358_, _14357_);
  nor (_14359_, _14304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  nor (_14360_, _14306_, _21586_);
  nor (_07078_, _14360_, _14359_);
  nor (_14361_, _14304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1]);
  nor (_14362_, _14306_, _21474_);
  nor (_07080_, _14362_, _14361_);
  nand (_14363_, _04985_, ABINPUT[7]);
  nand (_14364_, _04987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand (_14365_, _14364_, _14363_);
  nand (_14366_, _14365_, _24861_);
  nand (_14367_, _04982_, _01000_);
  nand (_14368_, _14367_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand (_14369_, _04982_, _01093_);
  nand (_14370_, _14369_, _14368_);
  nand (_14371_, _14370_, _00914_);
  nand (_14372_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nand (_14373_, _14372_, _14371_);
  nor (_14374_, _14373_, rst);
  nand (_07084_, _14374_, _14366_);
  nand (_14375_, _04985_, ABINPUT[6]);
  nand (_14376_, _04987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nand (_14377_, _14376_, _14375_);
  nand (_14378_, _14377_, _24861_);
  nand (_14379_, _04982_, _00908_);
  nand (_14380_, _14379_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nand (_14381_, _04982_, _00931_);
  nand (_14382_, _14381_, _14380_);
  nand (_14383_, _14382_, _00914_);
  nand (_14384_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nand (_14385_, _14384_, _14383_);
  nor (_14387_, _14385_, rst);
  nand (_07092_, _14387_, _14378_);
  nand (_14388_, _04985_, ABINPUT[5]);
  nand (_14389_, _04987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nand (_14390_, _14389_, _14388_);
  nand (_14391_, _14390_, _24861_);
  nand (_14392_, _04982_, _01026_);
  nand (_14393_, _14392_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nand (_14394_, _04982_, _01318_);
  nand (_14395_, _14394_, _14393_);
  nand (_14396_, _14395_, _00914_);
  nand (_14397_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nand (_14398_, _14397_, _14396_);
  nor (_14399_, _14398_, rst);
  nand (_07094_, _14399_, _14391_);
  nor (_14400_, _22991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6]);
  nor (_14401_, _22993_, _21504_);
  nor (_07096_, _14401_, _14400_);
  nand (_14402_, _04985_, ABINPUT[9]);
  nand (_14403_, _04987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nand (_14404_, _14403_, _14402_);
  nand (_14405_, _14404_, _24861_);
  nand (_14406_, _05052_, _04982_);
  nand (_14407_, _14406_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nand (_14408_, _05056_, _04982_);
  nand (_14409_, _14408_, _14407_);
  nand (_14410_, _14409_, _00914_);
  nand (_14411_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nand (_14412_, _14411_, _14410_);
  nor (_14413_, _14412_, rst);
  nand (_07123_, _14413_, _14405_);
  nor (_14414_, _14304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  nor (_14415_, _14306_, _21526_);
  nor (_07137_, _14415_, _14414_);
  nor (_14416_, _14304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  nor (_14417_, _14306_, _21414_);
  nor (_07152_, _14417_, _14416_);
  nor (_14418_, _22531_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7]);
  nor (_14419_, _22533_, _21626_);
  nor (_07155_, _14419_, _14418_);
  nor (_14420_, _21645_, _21566_);
  nor (_14421_, _14420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  not (_14422_, _14420_);
  nor (_14423_, _14422_, _21554_);
  nor (_07186_, _14423_, _14421_);
  nor (_14424_, _14420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  nor (_14425_, _14422_, _21414_);
  nor (_07196_, _14425_, _14424_);
  nor (_14426_, _14420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  nor (_14427_, _14422_, _21526_);
  nor (_25282_, _14427_, _14426_);
  nor (_14429_, _21728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7]);
  nor (_14430_, _21731_, _21626_);
  nor (_07205_, _14430_, _14429_);
  nand (_14431_, _05116_, ABINPUT[3]);
  nand (_14432_, _05118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nand (_14433_, _14432_, _14431_);
  nand (_14434_, _14433_, _24861_);
  not (_14435_, _14432_);
  nor (_14436_, _05115_, _10800_);
  nor (_14437_, _14436_, _14435_);
  nor (_14438_, _14437_, _00915_);
  nand (_14439_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nand (_14440_, _14439_, _23493_);
  nor (_14441_, _14440_, _14438_);
  nand (_07214_, _14441_, _14434_);
  nor (_14442_, _14420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7]);
  nor (_14443_, _14422_, _21626_);
  nor (_07242_, _14443_, _14442_);
  nand (_14444_, _05116_, ABINPUT[8]);
  nand (_14446_, _05118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nand (_14447_, _14446_, _14444_);
  nand (_14448_, _14447_, _24861_);
  not (_14449_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nor (_14450_, _05115_, _01010_);
  nor (_14451_, _14450_, _14449_);
  nor (_14452_, _10858_, _05115_);
  nor (_14453_, _14452_, _14451_);
  nor (_14454_, _14453_, _00915_);
  nand (_14455_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nand (_14456_, _14455_, _23493_);
  nor (_14457_, _14456_, _14454_);
  nand (_07245_, _14457_, _14448_);
  nand (_14458_, _05116_, ABINPUT[7]);
  nand (_14459_, _05118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nand (_14460_, _14459_, _14458_);
  nand (_14461_, _14460_, _24861_);
  not (_14462_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nor (_14463_, _05115_, _01001_);
  nor (_14464_, _14463_, _14462_);
  nor (_14466_, _05115_, _10873_);
  nor (_14467_, _14466_, _14464_);
  nor (_14468_, _14467_, _00915_);
  nand (_14469_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nand (_14470_, _14469_, _23493_);
  nor (_14471_, _14470_, _14468_);
  nand (_07247_, _14471_, _14461_);
  nand (_14472_, _05116_, ABINPUT[6]);
  nand (_14473_, _05118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nand (_14474_, _14473_, _14472_);
  nand (_14475_, _14474_, _24861_);
  not (_14476_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor (_14477_, _05115_, _00909_);
  nor (_14478_, _14477_, _14476_);
  nor (_14479_, _05115_, _10828_);
  nor (_14480_, _14479_, _14478_);
  nor (_14481_, _14480_, _00915_);
  nand (_14482_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nand (_14483_, _14482_, _23493_);
  nor (_14484_, _14483_, _14481_);
  nand (_07250_, _14484_, _14475_);
  nand (_14485_, _05116_, ABINPUT[5]);
  nand (_14486_, _05118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nand (_14487_, _14486_, _14485_);
  nand (_14488_, _14487_, _24861_);
  not (_14489_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nor (_14490_, _05115_, _01027_);
  nor (_14491_, _14490_, _14489_);
  nor (_14492_, _05115_, _02493_);
  nor (_14493_, _14492_, _14491_);
  nor (_14494_, _14493_, _00915_);
  nand (_14495_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nand (_14496_, _14495_, _23493_);
  nor (_14497_, _14496_, _14494_);
  nand (_07253_, _14497_, _14488_);
  nor (_14498_, _23400_, _23043_);
  not (_14499_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nand (_14500_, _23043_, _14499_);
  nand (_14501_, _14500_, _23493_);
  nor (_25019_[7], _14501_, _14498_);
  nor (_14502_, _14420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6]);
  nor (_14503_, _14422_, _21504_);
  nor (_07269_, _14503_, _14502_);
  nor (_14504_, _14420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5]);
  nor (_14505_, _14422_, _21451_);
  nor (_25283_, _14505_, _14504_);
  nand (_14506_, _05001_, ABINPUT[5]);
  nand (_14507_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nand (_14508_, _14507_, _14506_);
  nand (_14509_, _14508_, _24861_);
  not (_14510_, _05097_);
  nor (_14511_, _14510_, _01027_);
  nand (_14512_, _14511_, _21507_);
  not (_14513_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  not (_14514_, _14511_);
  nand (_14515_, _14514_, _14513_);
  nand (_14516_, _14515_, _14512_);
  nor (_14517_, _14516_, _00915_);
  nand (_14518_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nand (_14519_, _14518_, _23493_);
  nor (_14520_, _14519_, _14517_);
  nand (_07279_, _14520_, _14509_);
  nand (_14521_, _05001_, ABINPUT[4]);
  nand (_14522_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nand (_14523_, _14522_, _14521_);
  nand (_14524_, _14523_, _24861_);
  not (_14525_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_14526_, _14510_, _00020_);
  not (_14527_, _14526_);
  nand (_14528_, _14527_, _14525_);
  nand (_14529_, _14526_, _21507_);
  nand (_14530_, _14529_, _14528_);
  nor (_14531_, _14530_, _00915_);
  nand (_14532_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nand (_14533_, _14532_, _23493_);
  nor (_14534_, _14533_, _14531_);
  nand (_07282_, _14534_, _14524_);
  nor (_14535_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6]);
  nor (_14536_, _02372_, _21504_);
  nor (_25281_, _14536_, _14535_);
  nor (_14537_, _23025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5]);
  nor (_14538_, _23027_, _21451_);
  nor (_07302_, _14538_, _14537_);
  nand (_14539_, _05052_, _05097_);
  nand (_14540_, _14539_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nand (_14541_, _05056_, _05097_);
  nand (_14542_, _14541_, _14540_);
  nand (_14543_, _14542_, _00914_);
  nor (_14544_, _05003_, _00114_);
  not (_14545_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_14547_, _05001_, _14545_);
  nor (_14548_, _14547_, _14544_);
  nor (_14549_, _14548_, _00010_);
  nand (_14550_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nand (_14551_, _14550_, _23493_);
  nor (_14552_, _14551_, _14549_);
  nand (_07315_, _14552_, _14543_);
  nor (_14553_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7]);
  nor (_14554_, _02372_, _21626_);
  nor (_07317_, _14554_, _14553_);
  nand (_14555_, _05097_, _05015_);
  nand (_14556_, _14555_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nand (_14557_, _05018_, _05097_);
  nand (_14558_, _14557_, _14556_);
  nand (_14559_, _14558_, _00914_);
  nor (_14560_, _05003_, _00129_);
  not (_14561_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nor (_14562_, _05001_, _14561_);
  nor (_14563_, _14562_, _14560_);
  nor (_14564_, _14563_, _00010_);
  nand (_14565_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nand (_14566_, _14565_, _23493_);
  nor (_14567_, _14566_, _14564_);
  nand (_07321_, _14567_, _14559_);
  nand (_14568_, _05001_, ABINPUT[7]);
  nand (_14569_, _05003_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nand (_14570_, _14569_, _14568_);
  nand (_14571_, _14570_, _24861_);
  nor (_14572_, _14510_, _01001_);
  nand (_14573_, _14572_, _21507_);
  not (_14574_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  not (_14575_, _14572_);
  nand (_14576_, _14575_, _14574_);
  nand (_14577_, _14576_, _14573_);
  nor (_14578_, _14577_, _00915_);
  nand (_14579_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nand (_14580_, _14579_, _23493_);
  nor (_14581_, _14580_, _14578_);
  nand (_07325_, _14581_, _14571_);
  nor (_14582_, _14420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  nor (_14583_, _14422_, _21586_);
  nor (_07360_, _14583_, _14582_);
  nor (_14584_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  nor (_14585_, _02372_, _21554_);
  nor (_07394_, _14585_, _14584_);
  nand (_14586_, _01026_, _05014_);
  nand (_14587_, _14586_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nand (_14588_, _01318_, _05014_);
  nand (_14589_, _14588_, _14587_);
  nand (_14590_, _14589_, _00914_);
  not (_14591_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nor (_14592_, _05024_, _14591_);
  nor (_14593_, _05026_, _00121_);
  nor (_14594_, _14593_, _14592_);
  nor (_14595_, _14594_, _00010_);
  nand (_14596_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nand (_14597_, _14596_, _23493_);
  nor (_14598_, _14597_, _14595_);
  nand (_07412_, _14598_, _14590_);
  nand (_14599_, _00908_, _05014_);
  nand (_14600_, _14599_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nand (_14601_, _00931_, _05014_);
  nand (_14602_, _14601_, _14600_);
  nand (_14603_, _14602_, _00914_);
  not (_14604_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_14605_, _05024_, _14604_);
  nor (_14606_, _05026_, _24867_);
  nor (_14607_, _14606_, _14605_);
  nor (_14608_, _14607_, _00010_);
  nand (_14609_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nand (_14610_, _14609_, _23493_);
  nor (_14611_, _14610_, _14608_);
  nand (_07415_, _14611_, _14603_);
  not (_14612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_14613_, _00013_, _00018_);
  nor (_14614_, _14613_, _14612_);
  nor (_14615_, _05140_, _05076_);
  nor (_14616_, _14615_, _14614_);
  nor (_14617_, _14616_, _00915_);
  nand (_14618_, _05024_, _00006_);
  nor (_14619_, _05024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_14620_, _14619_, _00010_);
  nand (_14621_, _14620_, _14618_);
  nand (_14622_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nand (_14623_, _14622_, _14621_);
  nor (_14624_, _14623_, _14617_);
  nand (_07420_, _14624_, _23493_);
  nor (_14625_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  nor (_14626_, _02372_, _21414_);
  nor (_07434_, _14626_, _14625_);
  nor (_14628_, _01375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6]);
  nor (_14629_, _01377_, _21504_);
  nor (_07453_, _14629_, _14628_);
  nor (_14630_, _01375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5]);
  nor (_14631_, _01377_, _21451_);
  nor (_07456_, _14631_, _14630_);
  nor (_14632_, _22396_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  nor (_14633_, _22398_, _21586_);
  nor (_07460_, _14633_, _14632_);
  nor (_14634_, _21842_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7]);
  nor (_14635_, _21844_, _21626_);
  nor (_25199_, _14635_, _14634_);
  nor (_14636_, _21728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6]);
  nor (_14637_, _21731_, _21504_);
  nor (_07504_, _14637_, _14636_);
  nand (_14638_, _05577_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_14639_, _14638_);
  nor (_14640_, _05591_, _05568_);
  nor (_14641_, _14640_, _05585_);
  nand (_14642_, _14641_, _14639_);
  nand (_14643_, _14642_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand (_14644_, _14643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nor (_14645_, _05742_, _00018_);
  nand (_14646_, _14645_, _00914_);
  nand (_14647_, _14646_, _14644_);
  not (_14648_, _14646_);
  nand (_14649_, _14648_, ABINPUT[0]);
  nand (_14650_, _14649_, _14647_);
  nor (_14651_, _14650_, _05598_);
  nand (_14652_, _05598_, _00006_);
  nand (_14653_, _14652_, _23493_);
  nor (_07517_, _14653_, _14651_);
  nor (_07521_, _05564_, rst);
  not (_14654_, _01063_);
  nand (_14655_, _01072_, _14654_);
  nand (_14656_, _14250_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nand (_14657_, _14656_, _01064_);
  nand (_14658_, _01065_, _01057_);
  nand (_14659_, _14658_, _14657_);
  nand (_14660_, _14659_, _01070_);
  nor (_14661_, _14660_, _14655_);
  nor (_07534_, _14661_, _03986_);
  nor (_14662_, _01375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  nor (_14663_, _01377_, _21554_);
  nor (_07538_, _14663_, _14662_);
  nor (_14664_, _14266_, _00909_);
  not (_14665_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand (_14666_, _14640_, _05586_);
  nor (_14667_, _14666_, _14638_);
  nor (_14668_, _14667_, _14665_);
  nand (_14669_, _14668_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nor (_14670_, _14669_, _14664_);
  nand (_14671_, _14664_, ABINPUT[0]);
  nand (_14672_, _14671_, _05599_);
  nor (_14673_, _14672_, _14670_);
  nand (_14674_, _05598_, _24867_);
  nand (_14675_, _14674_, _23493_);
  nor (_07550_, _14675_, _14673_);
  nand (_14676_, _14265_, _05015_);
  nor (_14677_, _14676_, _21507_);
  not (_14678_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  nand (_14679_, _14678_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  not (_14680_, _14666_);
  nand (_14681_, _14680_, _05579_);
  nand (_14682_, _14681_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  nand (_14683_, _14682_, _14679_);
  nand (_14684_, _14683_, _14676_);
  nand (_14685_, _14684_, _05599_);
  nor (_14686_, _14685_, _14677_);
  nand (_14687_, _05598_, _00129_);
  nand (_14688_, _14687_, _23493_);
  nor (_07560_, _14688_, _14686_);
  nor (_14689_, _01375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1]);
  nor (_14690_, _01377_, _21474_);
  nor (_25278_, _14690_, _14689_);
  nor (_14691_, _05566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  not (_14692_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_14693_, _06708_, _14692_);
  nor (_14694_, _14693_, _14210_);
  not (_14695_, _14694_);
  nor (_14696_, _14695_, _14691_);
  nor (_14697_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nor (_14698_, _14697_, _14696_);
  nor (_14699_, _14698_, _14696_);
  nor (_14700_, _14699_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_14701_, _14698_, _14189_);
  nand (_14702_, _14701_, _23493_);
  nor (_07574_, _14702_, _14700_);
  not (_14703_, _14698_);
  nor (_07579_, _14703_, rst);
  nor (_14705_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  nor (_14706_, _22130_, _21554_);
  nor (_07598_, _14706_, _14705_);
  nor (_14707_, _01375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  nor (_14708_, _01377_, _21526_);
  nor (_07625_, _14708_, _14707_);
  nor (_14709_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1]);
  nor (_14710_, _22130_, _21474_);
  nor (_25246_, _14710_, _14709_);
  nor (_14711_, _22506_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5]);
  nor (_14713_, _22508_, _21451_);
  nor (_07642_, _14713_, _14711_);
  nor (_14714_, _22127_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  nor (_14715_, _22130_, _21586_);
  nor (_07652_, _14715_, _14714_);
  nor (_14716_, _23557_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5]);
  nor (_14717_, _23560_, _21451_);
  nor (_07664_, _14717_, _14716_);
  nor (_14718_, _02439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6]);
  nor (_14719_, _02442_, _21504_);
  nor (_07702_, _14719_, _14718_);
  nor (_14721_, _21728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1]);
  nor (_14722_, _21731_, _21474_);
  nor (_07712_, _14722_, _14721_);
  nor (_14723_, _21728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  nor (_14724_, _21731_, _21586_);
  nor (_07714_, _14724_, _14723_);
  nor (_14725_, _21834_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  nor (_14726_, _21836_, _21414_);
  nor (_25200_, _14726_, _14725_);
  nor (_07730_, _23175_, rst);
  nor (_14727_, _21659_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7]);
  nor (_14728_, _21661_, _21626_);
  nor (_07732_, _14728_, _14727_);
  nor (_14729_, _22408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5]);
  nor (_14730_, _22410_, _21451_);
  nor (_07743_, _14730_, _14729_);
  nor (_07757_, _23279_, rst);
  nor (_07781_, _23229_, rst);
  nor (_07783_, _24870_, rst);
  nor (_14731_, _21747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1]);
  nor (_14732_, _21749_, _21474_);
  nor (_07790_, _14732_, _14731_);
  nor (_14733_, _01383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  nor (_14734_, _01385_, _21554_);
  nor (_07818_, _14734_, _14733_);
  not (_14735_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nor (_14736_, _14293_, _05055_);
  nor (_14737_, _14736_, _14735_);
  nor (_14738_, _14293_, _05125_);
  nor (_14740_, _14738_, _14737_);
  nor (_14741_, _14740_, _14300_);
  nor (_14742_, _14299_, _00114_);
  nor (_14743_, _14742_, _14741_);
  nor (_07823_, _14743_, rst);
  nor (_14744_, _02439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  nor (_14745_, _02442_, _21554_);
  nor (_07828_, _14745_, _14744_);
  nand (_14746_, _04985_, ABINPUT[10]);
  nand (_14747_, _04987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nand (_14748_, _14747_, _14746_);
  nand (_14749_, _14748_, _24861_);
  not (_14750_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_14751_, _14298_, _14750_);
  nor (_14752_, _06627_, _04983_);
  nor (_14753_, _14752_, _14751_);
  nor (_14754_, _14753_, _00915_);
  nand (_14755_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nand (_14756_, _14755_, _23493_);
  nor (_14757_, _14756_, _14754_);
  nand (_07835_, _14757_, _14749_);
  nor (_14758_, _02439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1]);
  nor (_14759_, _02442_, _21474_);
  nor (_07837_, _14759_, _14758_);
  nor (_14760_, _14293_, _10828_);
  nor (_14761_, _14293_, _00909_);
  nor (_14762_, _14761_, _05652_);
  nor (_14763_, _14762_, _14760_);
  nor (_14764_, _14763_, _14300_);
  nor (_14765_, _14299_, _24867_);
  nor (_14766_, _14765_, _14764_);
  nor (_07840_, _14766_, rst);
  nor (_14767_, _22408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  nor (_14768_, _22410_, _21526_);
  nor (_25110_, _14768_, _14767_);
  nor (_14769_, _14293_, _24858_);
  nor (_14770_, _14769_, _05619_);
  nor (_14771_, _14293_, _10800_);
  nor (_14772_, _14771_, _14770_);
  nor (_14773_, _14772_, _14300_);
  nor (_14774_, _14299_, _00029_);
  nor (_14775_, _14774_, _14773_);
  nor (_07844_, _14775_, rst);
  nor (_14776_, _14293_, _01001_);
  nor (_14777_, _14776_, _05644_);
  nor (_14778_, _14293_, _10873_);
  nor (_14779_, _14778_, _14777_);
  nor (_14780_, _14779_, _14300_);
  nor (_14781_, _14299_, _24900_);
  nor (_14782_, _14781_, _14780_);
  nor (_07849_, _14782_, rst);
  nand (_14783_, _05116_, ABINPUT[10]);
  nand (_14784_, _05118_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nand (_14785_, _14784_, _14783_);
  nand (_14786_, _14785_, _24861_);
  not (_14787_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_14788_, _05559_, _05115_);
  nor (_14789_, _14788_, _14787_);
  nor (_14790_, _06627_, _05115_);
  nor (_14791_, _14790_, _14789_);
  nor (_14792_, _14791_, _00915_);
  nand (_14793_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nand (_14794_, _14793_, _23493_);
  nor (_14795_, _14794_, _14792_);
  nand (_07851_, _14795_, _14786_);
  nor (_14796_, _22408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  nor (_14797_, _22410_, _21414_);
  nor (_07853_, _14797_, _14796_);
  nor (_14798_, _21747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  nor (_14799_, _21749_, _21586_);
  nor (_07863_, _14799_, _14798_);
  nand (_14801_, _05558_, _05097_);
  nand (_14802_, _14801_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nand (_14803_, _06626_, _05097_);
  nand (_14804_, _14803_, _14802_);
  nand (_14805_, _14804_, _00914_);
  nor (_14806_, _05003_, _00106_);
  not (_14807_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_14808_, _05001_, _14807_);
  nor (_14809_, _14808_, _14806_);
  nor (_14810_, _14809_, _00010_);
  nand (_14811_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nand (_14812_, _14811_, _23493_);
  nor (_14813_, _14812_, _14810_);
  nand (_07865_, _14813_, _14805_);
  nor (_14814_, _14293_, _01010_);
  nor (_14815_, _14814_, _05636_);
  nor (_14816_, _14293_, _10858_);
  nor (_14817_, _14816_, _14815_);
  nor (_14818_, _14817_, _14300_);
  nor (_14820_, _14299_, _00129_);
  nor (_14821_, _14820_, _14818_);
  nor (_07876_, _14821_, rst);
  nand (_14822_, _05024_, _00106_);
  nor (_14823_, _05024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_14824_, _14823_, _00010_);
  nand (_14825_, _14824_, _14822_);
  not (_14826_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_14827_, _14186_, _14826_);
  nor (_14828_, _06627_, _05076_);
  nor (_14829_, _14828_, _14827_);
  nor (_14830_, _14829_, _00915_);
  nand (_14831_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nand (_14832_, _14831_, _23493_);
  nor (_14833_, _14832_, _14830_);
  nand (_07886_, _14833_, _14825_);
  nor (_14834_, _02439_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  nor (_14835_, _02442_, _21414_);
  nor (_07895_, _14835_, _14834_);
  nor (_14836_, _21728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  nor (_14837_, _21731_, _21526_);
  nor (_07916_, _14837_, _14836_);
  nor (_14838_, _21728_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  nor (_14839_, _21731_, _21554_);
  nor (_07922_, _14839_, _14838_);
  nor (_14840_, _11565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  nor (_14841_, _11567_, _21414_);
  nor (_07930_, _14841_, _14840_);
  nor (_14842_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  nor (_14843_, _02372_, _21526_);
  nor (_07933_, _14843_, _14842_);
  not (_14845_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  nor (_14846_, _14277_, _05055_);
  nor (_14847_, _14846_, _14845_);
  nand (_14848_, _14276_, _05056_);
  nand (_14849_, _14848_, _14281_);
  nor (_14850_, _14849_, _14847_);
  nand (_14851_, _14280_, _00114_);
  nand (_14852_, _14851_, _23493_);
  nor (_07948_, _14852_, _14850_);
  nor (_14853_, _22434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5]);
  nor (_14854_, _22437_, _21451_);
  nor (_07959_, _14854_, _14853_);
  nor (_14855_, _14293_, _05140_);
  nor (_14856_, _14293_, _00020_);
  nor (_14857_, _14856_, _05623_);
  nor (_14858_, _14857_, _14855_);
  nor (_14859_, _14858_, _14300_);
  nor (_14860_, _14299_, _00006_);
  nor (_14861_, _14860_, _14859_);
  nor (_07961_, _14861_, rst);
  nor (_14862_, _11565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5]);
  nor (_14863_, _11567_, _21451_);
  nor (_07967_, _14863_, _14862_);
  nor (_14864_, _11565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  nor (_14865_, _11567_, _21526_);
  nor (_07986_, _14865_, _14864_);
  nor (_14866_, _01375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7]);
  nor (_14867_, _01377_, _21626_);
  nor (_07989_, _14867_, _14866_);
  nor (_14869_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  nor (_14870_, _22537_, _21554_);
  nor (_25113_, _14870_, _14869_);
  nor (_14871_, _22434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  nor (_14872_, _22437_, _21414_);
  nor (_25102_, _14872_, _14871_);
  nor (_14873_, _22434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  nor (_14874_, _22437_, _21554_);
  nor (_08007_, _14874_, _14873_);
  nor (_14875_, _21829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  nor (_14876_, _21831_, _21414_);
  nor (_08010_, _14876_, _14875_);
  nor (_14877_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1]);
  nor (_14878_, _22537_, _21474_);
  nor (_08015_, _14878_, _14877_);
  nor (_14879_, _21904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  nor (_14880_, _21906_, _21586_);
  nor (_08021_, _14880_, _14879_);
  nor (_14881_, _11565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7]);
  nor (_14882_, _11567_, _21626_);
  nor (_08030_, _14882_, _14881_);
  not (_14884_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  nor (_14885_, _02390_, _01010_);
  nor (_14886_, _14885_, _14884_);
  nand (_14887_, _05018_, _02395_);
  nand (_14888_, _14887_, _02394_);
  nor (_14889_, _14888_, _14886_);
  nand (_14890_, _02393_, _00129_);
  nand (_14891_, _14890_, _23493_);
  nor (_08032_, _14891_, _14889_);
  nor (_14892_, _22434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1]);
  nor (_14893_, _22437_, _21474_);
  nor (_08034_, _14893_, _14892_);
  not (_14894_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nor (_14895_, _05055_, _02390_);
  nor (_14896_, _14895_, _14894_);
  nand (_14897_, _05056_, _02395_);
  nand (_14898_, _14897_, _02394_);
  nor (_14899_, _14898_, _14896_);
  nand (_14900_, _02393_, _00114_);
  nand (_14901_, _14900_, _23493_);
  nor (_08036_, _14901_, _14899_);
  nor (_14902_, _02390_, _01001_);
  nor (_14903_, _14902_, _01060_);
  nand (_14904_, _02395_, _01093_);
  nand (_14905_, _14904_, _02394_);
  nor (_14906_, _14905_, _14903_);
  nand (_14907_, _02393_, _24900_);
  nand (_14908_, _14907_, _23493_);
  nor (_08043_, _14908_, _14906_);
  nor (_14910_, _14277_, _01010_);
  nor (_14911_, _14910_, _05637_);
  nand (_14912_, _14276_, _05018_);
  nand (_14913_, _14912_, _14281_);
  nor (_14914_, _14913_, _14911_);
  nand (_14915_, _14280_, _00129_);
  nand (_14916_, _14915_, _23493_);
  nor (_08050_, _14916_, _14914_);
  nor (_14917_, _22412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1]);
  nor (_14918_, _22414_, _21474_);
  nor (_08052_, _14918_, _14917_);
  nor (_14919_, _22412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  nor (_14920_, _22414_, _21554_);
  nor (_08068_, _14920_, _14919_);
  nor (_14921_, _11565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6]);
  nor (_14922_, _11567_, _21504_);
  nor (_25277_, _14922_, _14921_);
  nor (_14923_, _22412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6]);
  nor (_14924_, _22414_, _21504_);
  nor (_08086_, _14924_, _14923_);
  nor (_14925_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5]);
  nor (_14926_, _02372_, _21451_);
  nor (_08089_, _14926_, _14925_);
  nor (_14927_, _14293_, _01027_);
  nor (_14928_, _14927_, _05629_);
  nor (_14929_, _14293_, _02493_);
  nor (_14930_, _14929_, _14928_);
  nor (_14931_, _14930_, _14300_);
  nor (_14932_, _14299_, _00121_);
  nor (_14933_, _14932_, _14931_);
  nor (_08100_, _14933_, rst);
  not (_14934_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nor (_14935_, _14277_, _00909_);
  nor (_14936_, _14935_, _14934_);
  nand (_14937_, _14276_, _00931_);
  nand (_14938_, _14937_, _14281_);
  nor (_14939_, _14938_, _14936_);
  nand (_14940_, _14280_, _24867_);
  nand (_14941_, _14940_, _23493_);
  nor (_08146_, _14941_, _14939_);
  nor (_14942_, _22412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  nor (_14943_, _22414_, _21414_);
  nor (_08147_, _14943_, _14942_);
  not (_14944_, _00595_);
  nor (_08151_, _14944_, rst);
  nor (_14945_, _14266_, _01027_);
  nor (_14946_, _14945_, _14665_);
  nand (_14947_, _14265_, _01318_);
  nand (_14948_, _14947_, _05599_);
  nor (_14949_, _14948_, _14946_);
  nand (_14950_, _05598_, _00121_);
  nand (_14951_, _14950_, _23493_);
  nor (_08155_, _14951_, _14949_);
  not (_14952_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nor (_14953_, _14277_, _01027_);
  nor (_14954_, _14953_, _14952_);
  nand (_14955_, _14276_, _01318_);
  nand (_14956_, _14955_, _14281_);
  nor (_14957_, _14956_, _14954_);
  nand (_14958_, _14280_, _00121_);
  nand (_14959_, _14958_, _23493_);
  nor (_08163_, _14959_, _14957_);
  nor (_14960_, _22421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  nor (_14961_, _22423_, _21526_);
  nor (_08175_, _14961_, _14960_);
  nor (_14962_, _21829_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7]);
  nor (_14963_, _21831_, _21626_);
  nor (_08194_, _14963_, _14962_);
  nor (_14964_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  nor (_14965_, _22545_, _21414_);
  nor (_08197_, _14965_, _14964_);
  not (_14966_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nor (_14967_, _14266_, _24858_);
  nor (_14968_, _14967_, _14966_);
  nand (_14969_, _14967_, ABINPUT[0]);
  nand (_14970_, _14969_, _05599_);
  nor (_14971_, _14970_, _14968_);
  nand (_14972_, _05598_, _00029_);
  nand (_14973_, _14972_, _23493_);
  nor (_08203_, _14973_, _14971_);
  nor (_08206_, _24962_, rst);
  nor (_14974_, _22421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5]);
  nor (_14975_, _22423_, _21451_);
  nor (_08215_, _14975_, _14974_);
  nor (_14976_, _14420_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1]);
  nor (_14977_, _14422_, _21474_);
  nor (_08217_, _14977_, _14976_);
  nor (_14978_, _11565_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1]);
  nor (_14979_, _11567_, _21474_);
  nor (_08220_, _14979_, _14978_);
  nor (_14980_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  nor (_14981_, _22545_, _21526_);
  nor (_25100_, _14981_, _14980_);
  nor (_14982_, _22421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  nor (_14983_, _22423_, _21414_);
  nor (_08233_, _14983_, _14982_);
  nor (_14984_, _21733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  nor (_14985_, _21735_, _21526_);
  nor (_08236_, _14985_, _14984_);
  nor (_14986_, _21646_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5]);
  nor (_14987_, _21648_, _21451_);
  nor (_08242_, _14987_, _14986_);
  not (_14988_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nor (_14989_, _14277_, _24858_);
  nor (_14990_, _14989_, _14988_);
  nand (_14991_, _14989_, ABINPUT[0]);
  nand (_14992_, _14991_, _14281_);
  nor (_14993_, _14992_, _14990_);
  nand (_14994_, _14280_, _00029_);
  nand (_14995_, _14994_, _23493_);
  nor (_08244_, _14995_, _14993_);
  nor (_14996_, _14277_, _01001_);
  nor (_14997_, _14996_, _05645_);
  nand (_14998_, _14276_, _01093_);
  nand (_14999_, _14998_, _14281_);
  nor (_15000_, _14999_, _14997_);
  nand (_15001_, _14280_, _24900_);
  nand (_15002_, _15001_, _23493_);
  nor (_08266_, _15002_, _15000_);
  nor (_08268_, _00498_, rst);
  nor (_15004_, _22412_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5]);
  nor (_15005_, _22414_, _21451_);
  nor (_08272_, _15005_, _15004_);
  nor (_08274_, _00425_, rst);
  nor (_15006_, _22991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  nor (_15007_, _22993_, _21414_);
  nor (_08276_, _15007_, _15006_);
  nor (_15008_, _14277_, _00020_);
  nor (_15009_, _15008_, _05625_);
  nand (_15010_, _14276_, _05045_);
  nand (_15011_, _15010_, _14281_);
  nor (_15012_, _15011_, _15009_);
  nand (_15013_, _14280_, _00006_);
  nand (_15014_, _15013_, _23493_);
  nor (_08279_, _15014_, _15012_);
  nor (_15015_, _14266_, _01001_);
  nor (_15016_, _15015_, _02678_);
  nand (_15017_, _14265_, _01093_);
  nand (_15018_, _15017_, _05599_);
  nor (_15019_, _15018_, _15016_);
  nand (_15021_, _05598_, _24900_);
  nand (_15022_, _15021_, _23493_);
  nor (_08285_, _15022_, _15019_);
  nor (_15023_, _22421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7]);
  nor (_15024_, _22423_, _21626_);
  nor (_25109_, _15024_, _15023_);
  nor (_15025_, _21733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  nor (_15026_, _21735_, _21554_);
  nor (_08301_, _15026_, _15025_);
  nor (_15027_, _21733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1]);
  nor (_15028_, _21735_, _21474_);
  nor (_25243_, _15028_, _15027_);
  nor (_15029_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7]);
  nor (_15030_, _22545_, _21626_);
  nor (_08324_, _15030_, _15029_);
  nor (_15031_, _22500_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  nor (_15032_, _22502_, _21526_);
  nor (_08331_, _15032_, _15031_);
  nor (_15033_, _22425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6]);
  nor (_15034_, _22427_, _21504_);
  nor (_08337_, _15034_, _15033_);
  not (_15035_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_15036_, _08687_, _15035_);
  not (_15037_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_15038_, _08692_, _15037_);
  nor (_15039_, _15038_, _15036_);
  nor (_08345_, _15039_, rst);
  nor (_08348_, _00207_, rst);
  nor (_15040_, _08687_, _12038_);
  not (_15041_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_15043_, _08692_, _15041_);
  nor (_15044_, _15043_, _15040_);
  nor (_25031_[1], _15044_, rst);
  nor (_15045_, _21747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  nor (_15046_, _21749_, _21414_);
  nor (_25238_, _15046_, _15045_);
  nor (_15047_, _08687_, _11995_);
  not (_15048_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_15049_, _08692_, _15048_);
  nor (_15050_, _15049_, _15047_);
  nor (_08356_, _15050_, rst);
  nor (_15051_, _08687_, _11985_);
  not (_15052_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_15053_, _08692_, _15052_);
  nor (_15054_, _15053_, _15051_);
  nor (_08358_, _15054_, rst);
  nor (_15055_, _08687_, _11976_);
  not (_15056_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_15057_, _08692_, _15056_);
  nor (_15058_, _15057_, _15055_);
  nor (_08360_, _15058_, rst);
  nor (_15059_, _14118_, _14114_);
  nand (_15060_, _14117_, _05658_);
  nand (_15061_, _15060_, _05611_);
  nand (_15062_, _15061_, _23493_);
  nor (_08363_, _15062_, _15059_);
  nor (_15063_, _02370_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  nor (_15064_, _02372_, _21586_);
  nor (_08367_, _15064_, _15063_);
  nor (_15065_, _08687_, _11964_);
  not (_15066_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_15067_, _08692_, _15066_);
  nor (_15068_, _15067_, _15065_);
  nor (_25031_[5], _15068_, rst);
  nor (_15069_, _22949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5]);
  nor (_15070_, _22951_, _21451_);
  nor (_08373_, _15070_, _15069_);
  nor (_15071_, _08687_, _11954_);
  not (_15072_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_15073_, _08692_, _15072_);
  nor (_15075_, _15073_, _15071_);
  nor (_25031_[6], _15075_, rst);
  nor (_15076_, _08687_, _12061_);
  not (_15077_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_15078_, _08692_, _15077_);
  nor (_15079_, _15078_, _15076_);
  nor (_08377_, _15079_, rst);
  nor (_15080_, _08687_, _12076_);
  not (_15081_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_15082_, _08692_, _15081_);
  nor (_15083_, _15082_, _15080_);
  nor (_08379_, _15083_, rst);
  nor (_15084_, _08687_, _12078_);
  not (_15085_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_15086_, _08692_, _15085_);
  nor (_15087_, _15086_, _15084_);
  nor (_08381_, _15087_, rst);
  nor (_15088_, _08687_, _12079_);
  not (_15089_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_15090_, _08692_, _15089_);
  nor (_15091_, _15090_, _15088_);
  nor (_08384_, _15091_, rst);
  nor (_15092_, _08687_, _12070_);
  not (_15093_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_15094_, _08692_, _15093_);
  nor (_15095_, _15094_, _15092_);
  nor (_08386_, _15095_, rst);
  not (_15096_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_15097_, _08687_, _15096_);
  not (_15098_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_15099_, _08692_, _15098_);
  nor (_15100_, _15099_, _15097_);
  nor (_08388_, _15100_, rst);
  nor (_15101_, _08687_, _12088_);
  not (_15102_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_15103_, _08692_, _15102_);
  nor (_15104_, _15103_, _15101_);
  nor (_25031_[13], _15104_, rst);
  nor (_15105_, _08687_, _12092_);
  not (_15106_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_15107_, _08692_, _15106_);
  nor (_15108_, _15107_, _15105_);
  nor (_25031_[14], _15108_, rst);
  nor (_15109_, _22425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5]);
  nor (_15110_, _22427_, _21451_);
  nor (_08394_, _15110_, _15109_);
  nor (_15111_, _21904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5]);
  nor (_15112_, _21906_, _21451_);
  nor (_25202_, _15112_, _15111_);
  nor (_15113_, _22425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  nor (_15114_, _22427_, _21414_);
  nor (_08410_, _15114_, _15113_);
  nor (_25033_[5], _00279_, rst);
  nor (_15115_, _22421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6]);
  nor (_15116_, _22423_, _21504_);
  nor (_25108_, _15116_, _15115_);
  nor (_15117_, _14134_, _14114_);
  nand (_15118_, _14133_, _05658_);
  nand (_15119_, _15118_, _05608_);
  nand (_15120_, _15119_, _23493_);
  nor (_08425_, _15120_, _15117_);
  nor (_15121_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  nor (_15122_, _22545_, _21554_);
  nor (_08438_, _15122_, _15121_);
  nor (_15123_, _08687_, _15037_);
  not (_15124_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_15125_, _08692_, _15124_);
  nor (_15126_, _15125_, _15123_);
  nor (_08440_, _15126_, rst);
  nor (_15127_, _08687_, _15041_);
  not (_15128_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_15129_, _08692_, _15128_);
  nor (_15130_, _15129_, _15127_);
  nor (_08443_, _15130_, rst);
  nor (_15131_, _08687_, _15048_);
  not (_15132_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_15133_, _08692_, _15132_);
  nor (_15134_, _15133_, _15131_);
  nor (_08445_, _15134_, rst);
  nor (_15135_, _08687_, _15052_);
  not (_15136_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_15137_, _08692_, _15136_);
  nor (_15138_, _15137_, _15135_);
  nor (_08447_, _15138_, rst);
  nor (_15139_, _22543_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6]);
  nor (_15140_, _22545_, _21504_);
  nor (_08450_, _15140_, _15139_);
  nor (_15141_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor (_15142_, _15141_, _05665_);
  nor (_15143_, _15142_, _05670_);
  nand (_15145_, _05660_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_15146_, _15145_);
  nor (_15147_, _15146_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  not (_15148_, _05661_);
  nor (_15149_, _15148_, _05571_);
  nor (_15150_, _15149_, _05664_);
  not (_15151_, _15150_);
  nor (_15152_, _15151_, _15147_);
  nand (_15153_, _05664_, _05590_);
  nand (_15154_, _15153_, _05668_);
  nor (_15155_, _15154_, _15152_);
  nor (_15156_, _15155_, _15143_);
  not (_15157_, _05665_);
  nor (_15158_, _15157_, _05589_);
  nor (_15159_, _15158_, _05658_);
  nand (_15160_, _15159_, _05675_);
  nor (_15161_, _15160_, _15156_);
  nor (_15162_, _15141_, _05622_);
  nor (_15163_, _15162_, _05634_);
  not (_15164_, _05642_);
  nor (_15166_, _15164_, _05571_);
  nor (_15167_, _15166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  not (_15168_, _05654_);
  nand (_15169_, _05649_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_15170_, _15169_, _15168_);
  nor (_15171_, _15170_, _15167_);
  nand (_15172_, _05654_, _05590_);
  nand (_15173_, _15172_, _05632_);
  nor (_15174_, _15173_, _15171_);
  nor (_15175_, _15174_, _15163_);
  nand (_15176_, _05622_, _05590_);
  nand (_15177_, _15176_, _05658_);
  nor (_15178_, _15177_, _15175_);
  nor (_15179_, _15178_, _15161_);
  nor (_15180_, _15179_, _05606_);
  not (_15181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor (_15182_, _05676_, _05606_);
  not (_15183_, _15182_);
  nand (_15184_, _15183_, _15181_);
  nand (_15185_, _15184_, _23493_);
  nor (_08452_, _15185_, _15180_);
  nor (_08464_, _00352_, rst);
  nor (_15186_, _22425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7]);
  nor (_15187_, _22427_, _21626_);
  nor (_08471_, _15187_, _15186_);
  nor (_15188_, _21747_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  nor (_15189_, _21749_, _21526_);
  nor (_08473_, _15189_, _15188_);
  nor (_15190_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _05571_);
  nor (_15191_, _15190_, _05622_);
  nor (_15192_, _15191_, _05634_);
  not (_15193_, _05588_);
  nor (_15194_, _15168_, _15193_);
  nand (_15195_, _05642_, _05571_);
  nand (_15196_, _15195_, _05587_);
  not (_15197_, _05649_);
  nor (_15198_, _15197_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_15199_, _15198_, _05654_);
  nand (_15200_, _15199_, _15196_);
  nand (_15201_, _15200_, _05632_);
  nor (_15203_, _15201_, _15194_);
  nor (_15204_, _15203_, _15192_);
  nand (_15205_, _05622_, _05588_);
  nand (_15206_, _15205_, _05658_);
  nor (_15207_, _15206_, _15204_);
  nor (_15208_, _15190_, _05665_);
  nor (_15209_, _15208_, _05670_);
  nor (_15210_, _14122_, _15193_);
  nand (_15211_, _05660_, _05571_);
  nand (_15212_, _15211_, _05587_);
  nor (_15213_, _15148_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_15214_, _15213_, _05664_);
  nand (_15215_, _15214_, _15212_);
  nand (_15216_, _15215_, _05668_);
  nor (_15217_, _15216_, _15210_);
  nor (_15218_, _15217_, _15209_);
  nor (_15219_, _15157_, _15193_);
  nor (_15220_, _15219_, _05658_);
  nand (_15221_, _15220_, _05675_);
  nor (_15222_, _15221_, _15218_);
  nor (_15223_, _15222_, _15207_);
  nor (_15224_, _15223_, _05606_);
  nand (_15225_, _15183_, _05587_);
  nand (_15226_, _15225_, _23493_);
  nor (_08476_, _15226_, _15224_);
  nor (_15227_, _05356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  nor (_15228_, _05358_, _21414_);
  nor (_08482_, _15228_, _15227_);
  nor (_15229_, _22949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  nor (_15230_, _22951_, _21526_);
  nor (_08484_, _15230_, _15229_);
  nor (_15231_, _23025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6]);
  nor (_15232_, _23027_, _21504_);
  nor (_08486_, _15232_, _15231_);
  nor (_15233_, _22421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1]);
  nor (_15234_, _22423_, _21474_);
  nor (_08498_, _15234_, _15233_);
  nor (_15235_, _22949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  nor (_15236_, _22951_, _21414_);
  nor (_25097_, _15236_, _15235_);
  nor (_15237_, _08687_, _15056_);
  not (_15238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_15239_, _08692_, _15238_);
  nor (_15240_, _15239_, _15237_);
  nor (_25032_[4], _15240_, rst);
  nor (_15241_, _22408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1]);
  nor (_15242_, _22410_, _21474_);
  nor (_08507_, _15242_, _15241_);
  nor (_15243_, _22949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6]);
  nor (_15244_, _22951_, _21504_);
  nor (_25098_, _15244_, _15243_);
  nor (_15245_, _05356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  nor (_15246_, _05358_, _21526_);
  nor (_08512_, _15246_, _15245_);
  nor (_15247_, _08687_, _15066_);
  not (_15248_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_15249_, _08692_, _15248_);
  nor (_15250_, _15249_, _15247_);
  nor (_08514_, _15250_, rst);
  nor (_15251_, _08687_, _15072_);
  not (_15252_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_15253_, _08692_, _15252_);
  nor (_15254_, _15253_, _15251_);
  nor (_08516_, _15254_, rst);
  nor (_15255_, _08687_, _15077_);
  not (_15256_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_15257_, _08692_, _15256_);
  nor (_15258_, _15257_, _15255_);
  nor (_08518_, _15258_, rst);
  nor (_15259_, _08687_, _15081_);
  not (_15260_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_15261_, _08692_, _15260_);
  nor (_15262_, _15261_, _15259_);
  nor (_08520_, _15262_, rst);
  nor (_15263_, _08687_, _15085_);
  not (_15264_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_15265_, _08692_, _15264_);
  nor (_15266_, _15265_, _15263_);
  nor (_08522_, _15266_, rst);
  nor (_15267_, _22421_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  nor (_15268_, _22423_, _21586_);
  nor (_08528_, _15268_, _15267_);
  nor (_15269_, _05658_, _05606_);
  nor (_15270_, _15269_, _05571_);
  nand (_15271_, _14117_, _05676_);
  nand (_15272_, _15271_, _23493_);
  nor (_08534_, _15272_, _15270_);
  nor (_15273_, _08687_, _15089_);
  not (_15274_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_15275_, _08692_, _15274_);
  nor (_15276_, _15275_, _15273_);
  nor (_08537_, _15276_, rst);
  nor (_15277_, _08687_, _15093_);
  not (_15278_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_15279_, _08692_, _15278_);
  nor (_15280_, _15279_, _15277_);
  nor (_08550_, _15280_, rst);
  nor (_15281_, _08687_, _15098_);
  not (_15282_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_15283_, _08692_, _15282_);
  nor (_15284_, _15283_, _15281_);
  nor (_25032_[12], _15284_, rst);
  nor (_15285_, _08687_, _15102_);
  not (_15286_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_15287_, _08692_, _15286_);
  nor (_15288_, _15287_, _15285_);
  nor (_25032_[13], _15288_, rst);
  nor (_15289_, _08687_, _15106_);
  not (_15290_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_15291_, _08692_, _15290_);
  nor (_15293_, _15291_, _15289_);
  nor (_25032_[14], _15293_, rst);
  nor (_15294_, _22429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5]);
  nor (_15295_, _22431_, _21451_);
  nor (_25105_, _15295_, _15294_);
  nor (_15296_, _22949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  nor (_15297_, _22951_, _21586_);
  nor (_08566_, _15297_, _15296_);
  nor (_15298_, _05356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6]);
  nor (_15299_, _05358_, _21504_);
  nor (_08570_, _15299_, _15298_);
  nor (_15300_, _05356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5]);
  nor (_15301_, _05358_, _21451_);
  nor (_25275_, _15301_, _15300_);
  nor (_15302_, _01375_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  nor (_15303_, _01377_, _21414_);
  nor (_08585_, _15303_, _15302_);
  nor (_15304_, _15182_, _05569_);
  not (_15305_, _05572_);
  not (_15306_, _05628_);
  nor (_15307_, _15306_, _15305_);
  not (_15308_, _05631_);
  nand (_15309_, _15195_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  nand (_15310_, _15309_, _15199_);
  nand (_15311_, _05654_, _15305_);
  nand (_15312_, _15311_, _15310_);
  nand (_15313_, _15312_, _15308_);
  nor (_15314_, _05571_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  nand (_15315_, _15314_, _05631_);
  nand (_15316_, _15315_, _15313_);
  nor (_15317_, _15316_, _05628_);
  nor (_15318_, _15317_, _15307_);
  nor (_15319_, _15318_, _05622_);
  not (_15320_, _05622_);
  nor (_15321_, _15314_, _15320_);
  nor (_15322_, _15321_, _15319_);
  nor (_15323_, _15322_, _05679_);
  nand (_15324_, _15211_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  nand (_15325_, _15324_, _15214_);
  nand (_15326_, _05664_, _15305_);
  nand (_15327_, _15326_, _15325_);
  nor (_15328_, _15327_, _05667_);
  not (_15329_, _05667_);
  nor (_15330_, _15314_, _15329_);
  nor (_15331_, _15330_, _15328_);
  nor (_15332_, _15331_, _05666_);
  nand (_15333_, _05666_, _05572_);
  nand (_15334_, _15333_, _15157_);
  nor (_15335_, _15334_, _15332_);
  nor (_15336_, _14114_, _05665_);
  nor (_15338_, _15314_, _14114_);
  nor (_15339_, _15338_, _15336_);
  nor (_15340_, _15339_, _15335_);
  nor (_15341_, _15340_, _15323_);
  nor (_15342_, _15341_, _05606_);
  nor (_15343_, _15342_, _15304_);
  nor (_08589_, _15343_, rst);
  nor (_15344_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7]);
  nor (_15345_, _22498_, _21626_);
  nor (_08599_, _15345_, _15344_);
  nor (_15346_, _01083_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  nor (_15347_, _01052_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  nand (_15348_, _15347_, _01080_);
  nand (_15349_, _15348_, _23493_);
  nor (_08601_, _15349_, _15346_);
  nor (_15350_, _22949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7]);
  nor (_15351_, _22951_, _21626_);
  nor (_08607_, _15351_, _15350_);
  nor (_15352_, _22429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6]);
  nor (_15353_, _22431_, _21504_);
  nor (_08609_, _15353_, _15352_);
  nand (_15354_, _05672_, _14121_);
  nor (_15355_, _15354_, _05658_);
  nand (_15356_, _05606_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nand (_15357_, _15168_, _05500_);
  nor (_15358_, _15357_, _05617_);
  nor (_15359_, _05650_, _05635_);
  nand (_15360_, _15359_, _15358_);
  nand (_15361_, _15360_, _15356_);
  nor (_15362_, _15361_, _15355_);
  nor (_08614_, _15362_, rst);
  nor (_15363_, _22547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  nor (_15364_, _22549_, _21554_);
  nor (_08620_, _15364_, _15363_);
  nor (_15365_, _05356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  nor (_15366_, _05358_, _21586_);
  nor (_25273_, _15366_, _15365_);
  nand (_15367_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3]);
  nand (_15368_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3]);
  nand (_15369_, _15368_, _15367_);
  nand (_15370_, _15369_, _01417_);
  nand (_15371_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3]);
  nand (_15372_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3]);
  nand (_15373_, _15372_, _15371_);
  nand (_15374_, _15373_, _00227_);
  nand (_15375_, _15374_, _15370_);
  nand (_15376_, _15375_, _00560_);
  nand (_15377_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3]);
  nand (_15378_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3]);
  nand (_15379_, _15378_, _15377_);
  nand (_15380_, _15379_, _01417_);
  nand (_15381_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3]);
  nand (_15382_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3]);
  nand (_15383_, _15382_, _15381_);
  nand (_15384_, _15383_, _00227_);
  nand (_15385_, _15384_, _15380_);
  nand (_15386_, _15385_, _00561_);
  nand (_15387_, _15386_, _15376_);
  nand (_15388_, _15387_, _00466_);
  nor (_15389_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3]);
  nor (_15390_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3]);
  nor (_15391_, _15390_, _15389_);
  nand (_15392_, _15391_, _01417_);
  nor (_15393_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3]);
  nor (_15394_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3]);
  nor (_15395_, _15394_, _15393_);
  nand (_15396_, _15395_, _00227_);
  nand (_15397_, _15396_, _15392_);
  nand (_15398_, _15397_, _00560_);
  nor (_15399_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3]);
  nor (_15401_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3]);
  nor (_15402_, _15401_, _15399_);
  nand (_15403_, _15402_, _01417_);
  nor (_15404_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3]);
  nor (_15405_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3]);
  nor (_15406_, _15405_, _15404_);
  nand (_15407_, _15406_, _00227_);
  nand (_15408_, _15407_, _15403_);
  nand (_15409_, _15408_, _00561_);
  nand (_15410_, _15409_, _15398_);
  nand (_15411_, _15410_, _00465_);
  nand (_15412_, _15411_, _15388_);
  nand (_15413_, _15412_, _00247_);
  nand (_15414_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3]);
  nand (_15415_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3]);
  nand (_15416_, _15415_, _15414_);
  nand (_15417_, _15416_, _01417_);
  nand (_15418_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3]);
  nand (_15419_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3]);
  nand (_15420_, _15419_, _15418_);
  nand (_15421_, _15420_, _00227_);
  nand (_15422_, _15421_, _15417_);
  nand (_15423_, _15422_, _00560_);
  nand (_15424_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3]);
  nand (_15425_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3]);
  nand (_15426_, _15425_, _15424_);
  nand (_15427_, _15426_, _01417_);
  nand (_15428_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3]);
  nand (_15429_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3]);
  nand (_15430_, _15429_, _15428_);
  nand (_15431_, _15430_, _00227_);
  nand (_15432_, _15431_, _15427_);
  nand (_15433_, _15432_, _00561_);
  nand (_15434_, _15433_, _15423_);
  nand (_15435_, _15434_, _00466_);
  nor (_15436_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3]);
  nor (_15437_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3]);
  nor (_15438_, _15437_, _15436_);
  nand (_15439_, _15438_, _00227_);
  nand (_15440_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3]);
  nand (_15441_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3]);
  nand (_15442_, _15441_, _15440_);
  nand (_15443_, _15442_, _01417_);
  nand (_15444_, _15443_, _15439_);
  nand (_15445_, _15444_, _00560_);
  nor (_15446_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3]);
  nor (_15447_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3]);
  nor (_15448_, _15447_, _15446_);
  nand (_15449_, _15448_, _00227_);
  nand (_15450_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3]);
  nand (_15451_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3]);
  nand (_15452_, _15451_, _15450_);
  nand (_15453_, _15452_, _01417_);
  nand (_15454_, _15453_, _15449_);
  nand (_15455_, _15454_, _00561_);
  nand (_15456_, _15455_, _15445_);
  nand (_15457_, _15456_, _00465_);
  nand (_15458_, _15457_, _15435_);
  nand (_15459_, _15458_, _00248_);
  nand (_15460_, _15459_, _15413_);
  nand (_15461_, _15460_, _00320_);
  nand (_15462_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3]);
  nand (_15463_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3]);
  nand (_15464_, _15463_, _15462_);
  nand (_15465_, _15464_, _01417_);
  nand (_15466_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3]);
  nand (_15467_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3]);
  nand (_15468_, _15467_, _15466_);
  nand (_15469_, _15468_, _00227_);
  nand (_15470_, _15469_, _15465_);
  nand (_15471_, _15470_, _00560_);
  nand (_15472_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3]);
  nand (_15473_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3]);
  nand (_15474_, _15473_, _15472_);
  nand (_15475_, _15474_, _01417_);
  nand (_15476_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3]);
  nand (_15477_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3]);
  nand (_15478_, _15477_, _15476_);
  nand (_15479_, _15478_, _00227_);
  nand (_15480_, _15479_, _15475_);
  nand (_15482_, _15480_, _00561_);
  nand (_15483_, _15482_, _15471_);
  nand (_15484_, _15483_, _00466_);
  nor (_15485_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3]);
  nor (_15486_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3]);
  nor (_15487_, _15486_, _15485_);
  nand (_15488_, _15487_, _00227_);
  nand (_15489_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3]);
  nand (_15490_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3]);
  nand (_15491_, _15490_, _15489_);
  nand (_15492_, _15491_, _01417_);
  nand (_15493_, _15492_, _15488_);
  nand (_15494_, _15493_, _00560_);
  nor (_15495_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3]);
  nor (_15496_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3]);
  nor (_15497_, _15496_, _15495_);
  nand (_15498_, _15497_, _00227_);
  nand (_15499_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3]);
  nand (_15500_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3]);
  nand (_15501_, _15500_, _15499_);
  nand (_15503_, _15501_, _01417_);
  nand (_15504_, _15503_, _15498_);
  nand (_15505_, _15504_, _00561_);
  nand (_15506_, _15505_, _15494_);
  nand (_15507_, _15506_, _00465_);
  nand (_15508_, _15507_, _15484_);
  nand (_15509_, _15508_, _00248_);
  nand (_15510_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3]);
  nand (_15511_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3]);
  nand (_15512_, _15511_, _15510_);
  nand (_15513_, _15512_, _01417_);
  nand (_15514_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3]);
  nand (_15515_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3]);
  nand (_15516_, _15515_, _15514_);
  nand (_15517_, _15516_, _00227_);
  nand (_15518_, _15517_, _15513_);
  nand (_15519_, _15518_, _00560_);
  nand (_15520_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3]);
  nand (_15521_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3]);
  nand (_15522_, _15521_, _15520_);
  nand (_15523_, _15522_, _01417_);
  nand (_15524_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3]);
  nand (_15525_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3]);
  nand (_15526_, _15525_, _15524_);
  nand (_15527_, _15526_, _00227_);
  nand (_15528_, _15527_, _15523_);
  nand (_15529_, _15528_, _00561_);
  nand (_15530_, _15529_, _15519_);
  nand (_15531_, _15530_, _00466_);
  nor (_15532_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3]);
  nor (_15533_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3]);
  nor (_15534_, _15533_, _15532_);
  nand (_15535_, _15534_, _01417_);
  nor (_15536_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3]);
  nor (_15537_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3]);
  nor (_15538_, _15537_, _15536_);
  nand (_15539_, _15538_, _00227_);
  nand (_15540_, _15539_, _15535_);
  nand (_15541_, _15540_, _00560_);
  nor (_15542_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3]);
  nor (_15543_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3]);
  nor (_15544_, _15543_, _15542_);
  nand (_15545_, _15544_, _01417_);
  nor (_15546_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3]);
  nor (_15547_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3]);
  nor (_15548_, _15547_, _15546_);
  nand (_15549_, _15548_, _00227_);
  nand (_15550_, _15549_, _15545_);
  nand (_15551_, _15550_, _00561_);
  nand (_15552_, _15551_, _15541_);
  nand (_15553_, _15552_, _00465_);
  nand (_15554_, _15553_, _15531_);
  nand (_15555_, _15554_, _00247_);
  nand (_15556_, _15555_, _15509_);
  nand (_15557_, _15556_, _00319_);
  nand (_15558_, _15557_, _15461_);
  nor (_15559_, _15558_, _00386_);
  nand (_15560_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3]);
  nand (_15561_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3]);
  nand (_15562_, _15561_, _15560_);
  nand (_15563_, _15562_, _01417_);
  nand (_15564_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3]);
  nand (_15565_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3]);
  nand (_15566_, _15565_, _15564_);
  nand (_15567_, _15566_, _00227_);
  nand (_15568_, _15567_, _15563_);
  nand (_15569_, _15568_, _00560_);
  nand (_15570_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3]);
  nand (_15571_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3]);
  nand (_15572_, _15571_, _15570_);
  nand (_15574_, _15572_, _01417_);
  nand (_15575_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3]);
  nand (_15576_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3]);
  nand (_15577_, _15576_, _15575_);
  nand (_15578_, _15577_, _00227_);
  nand (_15579_, _15578_, _15574_);
  nand (_15580_, _15579_, _00561_);
  nand (_15581_, _15580_, _15569_);
  nand (_15582_, _15581_, _00466_);
  nor (_15583_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3]);
  nor (_15584_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3]);
  nor (_15585_, _15584_, _15583_);
  nand (_15586_, _15585_, _00227_);
  nand (_15587_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3]);
  nand (_15588_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3]);
  nand (_15589_, _15588_, _15587_);
  nand (_15590_, _15589_, _01417_);
  nand (_15591_, _15590_, _15586_);
  nand (_15592_, _15591_, _00560_);
  nor (_15593_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  nor (_15594_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3]);
  nor (_15595_, _15594_, _15593_);
  nand (_15596_, _15595_, _00227_);
  nand (_15597_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3]);
  nand (_15598_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3]);
  nand (_15599_, _15598_, _15597_);
  nand (_15600_, _15599_, _01417_);
  nand (_15601_, _15600_, _15596_);
  nand (_15602_, _15601_, _00561_);
  nand (_15603_, _15602_, _15592_);
  nand (_15604_, _15603_, _00465_);
  nand (_15605_, _15604_, _15582_);
  nand (_15606_, _15605_, _00248_);
  nand (_15607_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3]);
  nand (_15608_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3]);
  nand (_15609_, _15608_, _15607_);
  nand (_15610_, _15609_, _01417_);
  nand (_15611_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3]);
  nand (_15612_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3]);
  nand (_15613_, _15612_, _15611_);
  nand (_15615_, _15613_, _00227_);
  nand (_15616_, _15615_, _15610_);
  nand (_15617_, _15616_, _00560_);
  nand (_15618_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3]);
  nand (_15619_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3]);
  nand (_15620_, _15619_, _15618_);
  nand (_15621_, _15620_, _01417_);
  nand (_15622_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3]);
  nand (_15623_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3]);
  nand (_15624_, _15623_, _15622_);
  nand (_15625_, _15624_, _00227_);
  nand (_15626_, _15625_, _15621_);
  nand (_15627_, _15626_, _00561_);
  nand (_15628_, _15627_, _15617_);
  nand (_15629_, _15628_, _00466_);
  nor (_15630_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3]);
  nor (_15631_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3]);
  nor (_15632_, _15631_, _15630_);
  nand (_15633_, _15632_, _01417_);
  nor (_15634_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3]);
  nor (_15636_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3]);
  nor (_15637_, _15636_, _15634_);
  nand (_15638_, _15637_, _00227_);
  nand (_15639_, _15638_, _15633_);
  nand (_15640_, _15639_, _00560_);
  nor (_15641_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3]);
  nor (_15642_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3]);
  nor (_15643_, _15642_, _15641_);
  nand (_15644_, _15643_, _01417_);
  nor (_15645_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3]);
  nor (_15646_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3]);
  nor (_15647_, _15646_, _15645_);
  nand (_15648_, _15647_, _00227_);
  nand (_15649_, _15648_, _15644_);
  nand (_15650_, _15649_, _00561_);
  nand (_15651_, _15650_, _15640_);
  nand (_15652_, _15651_, _00465_);
  nand (_15653_, _15652_, _15629_);
  nand (_15654_, _15653_, _00247_);
  nand (_15655_, _15654_, _15606_);
  nand (_15656_, _15655_, _00320_);
  nor (_15657_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3]);
  nor (_15658_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3]);
  nor (_15659_, _15658_, _15657_);
  nand (_15660_, _15659_, _01417_);
  nor (_15661_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3]);
  nor (_15662_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3]);
  nor (_15663_, _15662_, _15661_);
  nand (_15664_, _15663_, _00227_);
  nand (_15665_, _15664_, _15660_);
  nand (_15666_, _15665_, _00561_);
  nor (_15667_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3]);
  nor (_15668_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3]);
  nor (_15669_, _15668_, _15667_);
  nand (_15670_, _15669_, _01417_);
  nor (_15671_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3]);
  nor (_15672_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3]);
  nor (_15673_, _15672_, _15671_);
  nand (_15674_, _15673_, _00227_);
  nand (_15675_, _15674_, _15670_);
  nand (_15676_, _15675_, _00560_);
  nand (_15677_, _15676_, _15666_);
  nand (_15678_, _15677_, _00465_);
  nand (_15679_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3]);
  nand (_15680_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3]);
  nand (_15681_, _15680_, _15679_);
  nand (_15682_, _15681_, _01417_);
  nand (_15683_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3]);
  nand (_15684_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3]);
  nand (_15685_, _15684_, _15683_);
  nand (_15686_, _15685_, _00227_);
  nand (_15687_, _15686_, _15682_);
  nand (_15688_, _15687_, _00561_);
  nand (_15689_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3]);
  nand (_15690_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3]);
  nand (_15691_, _15690_, _15689_);
  nand (_15692_, _15691_, _01417_);
  nand (_15693_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3]);
  nand (_15694_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3]);
  nand (_15695_, _15694_, _15693_);
  nand (_15696_, _15695_, _00227_);
  nand (_15697_, _15696_, _15692_);
  nand (_15698_, _15697_, _00560_);
  nand (_15699_, _15698_, _15688_);
  nand (_15700_, _15699_, _00466_);
  nand (_15701_, _15700_, _15678_);
  nand (_15702_, _15701_, _00247_);
  nor (_15703_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3]);
  nor (_15704_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3]);
  nor (_15705_, _15704_, _15703_);
  nand (_15706_, _15705_, _00227_);
  nand (_15707_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3]);
  nand (_15708_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3]);
  nand (_15709_, _15708_, _15707_);
  nand (_15710_, _15709_, _01417_);
  nand (_15711_, _15710_, _15706_);
  nand (_15712_, _15711_, _00561_);
  nor (_15713_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3]);
  nor (_15714_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3]);
  nor (_15715_, _15714_, _15713_);
  nand (_15716_, _15715_, _00227_);
  nand (_15717_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3]);
  nand (_15718_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3]);
  nand (_15719_, _15718_, _15717_);
  nand (_15720_, _15719_, _01417_);
  nand (_15721_, _15720_, _15716_);
  nand (_15722_, _15721_, _00560_);
  nand (_15723_, _15722_, _15712_);
  nand (_15724_, _15723_, _00465_);
  nand (_15725_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3]);
  nand (_15726_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3]);
  nand (_15727_, _15726_, _15725_);
  nand (_15728_, _15727_, _01417_);
  nand (_15729_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3]);
  nand (_15730_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3]);
  nand (_15731_, _15730_, _15729_);
  nand (_15732_, _15731_, _00227_);
  nand (_15733_, _15732_, _15728_);
  nand (_15734_, _15733_, _00561_);
  nand (_15735_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3]);
  nand (_15737_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3]);
  nand (_15738_, _15737_, _15735_);
  nand (_15739_, _15738_, _01417_);
  nand (_15740_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3]);
  nand (_15741_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3]);
  nand (_15742_, _15741_, _15740_);
  nand (_15743_, _15742_, _00227_);
  nand (_15744_, _15743_, _15739_);
  nand (_15745_, _15744_, _00560_);
  nand (_15746_, _15745_, _15734_);
  nand (_15747_, _15746_, _00466_);
  nand (_15748_, _15747_, _15724_);
  nand (_15749_, _15748_, _00248_);
  nand (_15750_, _15749_, _15702_);
  nand (_15751_, _15750_, _00319_);
  nand (_15752_, _15751_, _15656_);
  nor (_15753_, _15752_, _01629_);
  nor (_15754_, _15753_, _15559_);
  nor (_15755_, _15754_, _00156_);
  nand (_15756_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3]);
  nand (_15757_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3]);
  nand (_15758_, _15757_, _15756_);
  nand (_15759_, _15758_, _01417_);
  nand (_15760_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  nand (_15761_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3]);
  nand (_15762_, _15761_, _15760_);
  nand (_15763_, _15762_, _00227_);
  nand (_15764_, _15763_, _15759_);
  nand (_15765_, _15764_, _00560_);
  nand (_15766_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3]);
  nand (_15767_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3]);
  nand (_15768_, _15767_, _15766_);
  nand (_15769_, _15768_, _01417_);
  nand (_15770_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3]);
  nand (_15771_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3]);
  nand (_15772_, _15771_, _15770_);
  nand (_15773_, _15772_, _00227_);
  nand (_15774_, _15773_, _15769_);
  nand (_15775_, _15774_, _00561_);
  nand (_15776_, _15775_, _15765_);
  nand (_15778_, _15776_, _00466_);
  nor (_15779_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3]);
  nor (_15780_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3]);
  nor (_15781_, _15780_, _15779_);
  nand (_15782_, _15781_, _01417_);
  nor (_15783_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3]);
  nor (_15784_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3]);
  nor (_15785_, _15784_, _15783_);
  nand (_15786_, _15785_, _00227_);
  nand (_15787_, _15786_, _15782_);
  nand (_15789_, _15787_, _00560_);
  nor (_15790_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3]);
  nor (_15791_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3]);
  nor (_15792_, _15791_, _15790_);
  nand (_15793_, _15792_, _01417_);
  nor (_15794_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3]);
  nor (_15795_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3]);
  nor (_15796_, _15795_, _15794_);
  nand (_15797_, _15796_, _00227_);
  nand (_15798_, _15797_, _15793_);
  nand (_15799_, _15798_, _00561_);
  nand (_15800_, _15799_, _15789_);
  nand (_15801_, _15800_, _00465_);
  nand (_15802_, _15801_, _15778_);
  nand (_15803_, _15802_, _00247_);
  nand (_15804_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3]);
  nand (_15805_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3]);
  nand (_15806_, _15805_, _15804_);
  nand (_15807_, _15806_, _01417_);
  nand (_15808_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3]);
  nand (_15809_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3]);
  nand (_15810_, _15809_, _15808_);
  nand (_15811_, _15810_, _00227_);
  nand (_15812_, _15811_, _15807_);
  nand (_15813_, _15812_, _00560_);
  nand (_15814_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3]);
  nand (_15815_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3]);
  nand (_15816_, _15815_, _15814_);
  nand (_15817_, _15816_, _01417_);
  nand (_15818_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3]);
  nand (_15819_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3]);
  nand (_15820_, _15819_, _15818_);
  nand (_15821_, _15820_, _00227_);
  nand (_15822_, _15821_, _15817_);
  nand (_15823_, _15822_, _00561_);
  nand (_15824_, _15823_, _15813_);
  nand (_15825_, _15824_, _00466_);
  nor (_15826_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3]);
  nor (_15827_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3]);
  nor (_15828_, _15827_, _15826_);
  nand (_15829_, _15828_, _00227_);
  nand (_15830_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3]);
  nand (_15831_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3]);
  nand (_15832_, _15831_, _15830_);
  nand (_15833_, _15832_, _01417_);
  nand (_15834_, _15833_, _15829_);
  nand (_15835_, _15834_, _00560_);
  nor (_15836_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3]);
  nor (_15837_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3]);
  nor (_15838_, _15837_, _15836_);
  nand (_15839_, _15838_, _00227_);
  nand (_15840_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3]);
  nand (_15841_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3]);
  nand (_15842_, _15841_, _15840_);
  nand (_15843_, _15842_, _01417_);
  nand (_15844_, _15843_, _15839_);
  nand (_15845_, _15844_, _00561_);
  nand (_15846_, _15845_, _15835_);
  nand (_15847_, _15846_, _00465_);
  nand (_15848_, _15847_, _15825_);
  nand (_15849_, _15848_, _00248_);
  nand (_15850_, _15849_, _15803_);
  nand (_15851_, _15850_, _00320_);
  nand (_15852_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  nand (_15853_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  nand (_15854_, _15853_, _15852_);
  nand (_15855_, _15854_, _01417_);
  nand (_15856_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3]);
  nand (_15857_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3]);
  nand (_15858_, _15857_, _15856_);
  nand (_15859_, _15858_, _00227_);
  nand (_15860_, _15859_, _15855_);
  nand (_15861_, _15860_, _00560_);
  nand (_15862_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3]);
  nand (_15863_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3]);
  nand (_15864_, _15863_, _15862_);
  nand (_15865_, _15864_, _01417_);
  nand (_15866_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  nand (_15867_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3]);
  nand (_15868_, _15867_, _15866_);
  nand (_15869_, _15868_, _00227_);
  nand (_15870_, _15869_, _15865_);
  nand (_15871_, _15870_, _00561_);
  nand (_15872_, _15871_, _15861_);
  nand (_15873_, _15872_, _00466_);
  nor (_15874_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3]);
  nor (_15875_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3]);
  nor (_15876_, _15875_, _15874_);
  nand (_15877_, _15876_, _00227_);
  nand (_15878_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3]);
  nand (_15879_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3]);
  nand (_15880_, _15879_, _15878_);
  nand (_15881_, _15880_, _01417_);
  nand (_15882_, _15881_, _15877_);
  nand (_15883_, _15882_, _00560_);
  nor (_15884_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3]);
  nor (_15885_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3]);
  nor (_15886_, _15885_, _15884_);
  nand (_15887_, _15886_, _00227_);
  nand (_15888_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3]);
  nand (_15889_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3]);
  nand (_15890_, _15889_, _15888_);
  nand (_15891_, _15890_, _01417_);
  nand (_15892_, _15891_, _15887_);
  nand (_15893_, _15892_, _00561_);
  nand (_15894_, _15893_, _15883_);
  nand (_15895_, _15894_, _00465_);
  nand (_15896_, _15895_, _15873_);
  nand (_15897_, _15896_, _00248_);
  nand (_15898_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3]);
  nand (_15899_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3]);
  nand (_15900_, _15899_, _15898_);
  nand (_15901_, _15900_, _01417_);
  nand (_15902_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3]);
  nand (_15903_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3]);
  nand (_15904_, _15903_, _15902_);
  nand (_15905_, _15904_, _00227_);
  nand (_15906_, _15905_, _15901_);
  nand (_15907_, _15906_, _00560_);
  nand (_15908_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3]);
  nand (_15909_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3]);
  nand (_15910_, _15909_, _15908_);
  nand (_15911_, _15910_, _01417_);
  nand (_15912_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3]);
  nand (_15913_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3]);
  nand (_15914_, _15913_, _15912_);
  nand (_15915_, _15914_, _00227_);
  nand (_15916_, _15915_, _15911_);
  nand (_15917_, _15916_, _00561_);
  nand (_15918_, _15917_, _15907_);
  nand (_15919_, _15918_, _00466_);
  nor (_15920_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3]);
  nor (_15921_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3]);
  nor (_15922_, _15921_, _15920_);
  nand (_15923_, _15922_, _01417_);
  nor (_15924_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3]);
  nor (_15925_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3]);
  nor (_15926_, _15925_, _15924_);
  nand (_15927_, _15926_, _00227_);
  nand (_15928_, _15927_, _15923_);
  nand (_15929_, _15928_, _00560_);
  nor (_15930_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3]);
  nor (_15931_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3]);
  nor (_15932_, _15931_, _15930_);
  nand (_15933_, _15932_, _01417_);
  nor (_15934_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3]);
  nor (_15935_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3]);
  nor (_15936_, _15935_, _15934_);
  nand (_15937_, _15936_, _00227_);
  nand (_15938_, _15937_, _15933_);
  nand (_15939_, _15938_, _00561_);
  nand (_15940_, _15939_, _15929_);
  nand (_15941_, _15940_, _00465_);
  nand (_15942_, _15941_, _15919_);
  nand (_15943_, _15942_, _00247_);
  nand (_15944_, _15943_, _15897_);
  nand (_15945_, _15944_, _00319_);
  nand (_15946_, _15945_, _15851_);
  nor (_15947_, _15946_, _00386_);
  nand (_15948_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3]);
  nand (_15949_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3]);
  nand (_15950_, _15949_, _15948_);
  nand (_15951_, _15950_, _01417_);
  nand (_15952_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3]);
  nand (_15953_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3]);
  nand (_15954_, _15953_, _15952_);
  nand (_15955_, _15954_, _00227_);
  nand (_15956_, _15955_, _15951_);
  nand (_15957_, _15956_, _00560_);
  nand (_15958_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3]);
  nand (_15960_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3]);
  nand (_15961_, _15960_, _15958_);
  nand (_15962_, _15961_, _01417_);
  nand (_15963_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3]);
  nand (_15964_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3]);
  nand (_15965_, _15964_, _15963_);
  nand (_15966_, _15965_, _00227_);
  nand (_15967_, _15966_, _15962_);
  nand (_15968_, _15967_, _00561_);
  nand (_15969_, _15968_, _15957_);
  nand (_15970_, _15969_, _00466_);
  nor (_15971_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  nor (_15972_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  nor (_15973_, _15972_, _15971_);
  nand (_15974_, _15973_, _00227_);
  nand (_15975_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3]);
  nand (_15976_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3]);
  nand (_15977_, _15976_, _15975_);
  nand (_15978_, _15977_, _01417_);
  nand (_15979_, _15978_, _15974_);
  nand (_15980_, _15979_, _00560_);
  nor (_15981_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3]);
  nor (_15982_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3]);
  nor (_15983_, _15982_, _15981_);
  nand (_15984_, _15983_, _00227_);
  nand (_15985_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3]);
  nand (_15986_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3]);
  nand (_15987_, _15986_, _15985_);
  nand (_15988_, _15987_, _01417_);
  nand (_15989_, _15988_, _15984_);
  nand (_15991_, _15989_, _00561_);
  nand (_15992_, _15991_, _15980_);
  nand (_15993_, _15992_, _00465_);
  nand (_15994_, _15993_, _15970_);
  nand (_15995_, _15994_, _00248_);
  nand (_15996_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3]);
  nand (_15997_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3]);
  nand (_15998_, _15997_, _15996_);
  nand (_15999_, _15998_, _01417_);
  nand (_16000_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3]);
  nand (_16001_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3]);
  nand (_16002_, _16001_, _16000_);
  nand (_16003_, _16002_, _00227_);
  nand (_16004_, _16003_, _15999_);
  nand (_16005_, _16004_, _00560_);
  nand (_16006_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3]);
  nand (_16007_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3]);
  nand (_16008_, _16007_, _16006_);
  nand (_16009_, _16008_, _01417_);
  nand (_16010_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3]);
  nand (_16012_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3]);
  nand (_16013_, _16012_, _16010_);
  nand (_16014_, _16013_, _00227_);
  nand (_16015_, _16014_, _16009_);
  nand (_16016_, _16015_, _00561_);
  nand (_16017_, _16016_, _16005_);
  nand (_16018_, _16017_, _00466_);
  nor (_16019_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3]);
  nor (_16020_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3]);
  nor (_16021_, _16020_, _16019_);
  nand (_16022_, _16021_, _01417_);
  nor (_16023_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3]);
  nor (_16024_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3]);
  nor (_16025_, _16024_, _16023_);
  nand (_16026_, _16025_, _00227_);
  nand (_16027_, _16026_, _16022_);
  nand (_16028_, _16027_, _00560_);
  nor (_16029_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3]);
  nor (_16030_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3]);
  nor (_16031_, _16030_, _16029_);
  nand (_16033_, _16031_, _01417_);
  nor (_16034_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  nor (_16035_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3]);
  nor (_16036_, _16035_, _16034_);
  nand (_16037_, _16036_, _00227_);
  nand (_16038_, _16037_, _16033_);
  nand (_16039_, _16038_, _00561_);
  nand (_16040_, _16039_, _16028_);
  nand (_16041_, _16040_, _00465_);
  nand (_16042_, _16041_, _16018_);
  nand (_16043_, _16042_, _00247_);
  nand (_16044_, _16043_, _15995_);
  nand (_16045_, _16044_, _00320_);
  nor (_16046_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3]);
  nor (_16047_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3]);
  nor (_16048_, _16047_, _16046_);
  nand (_16049_, _16048_, _01417_);
  nor (_16050_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3]);
  nor (_16051_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3]);
  nor (_16052_, _16051_, _16050_);
  nand (_16054_, _16052_, _00227_);
  nand (_16055_, _16054_, _16049_);
  nand (_16056_, _16055_, _00561_);
  nor (_16057_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3]);
  nor (_16058_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3]);
  nor (_16059_, _16058_, _16057_);
  nand (_16060_, _16059_, _01417_);
  nor (_16061_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3]);
  nor (_16062_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3]);
  nor (_16063_, _16062_, _16061_);
  nand (_16064_, _16063_, _00227_);
  nand (_16065_, _16064_, _16060_);
  nand (_16066_, _16065_, _00560_);
  nand (_16067_, _16066_, _16056_);
  nand (_16068_, _16067_, _00465_);
  nand (_16069_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3]);
  nand (_16070_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3]);
  nand (_16071_, _16070_, _16069_);
  nand (_16072_, _16071_, _01417_);
  nand (_16073_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3]);
  nand (_16075_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3]);
  nand (_16076_, _16075_, _16073_);
  nand (_16077_, _16076_, _00227_);
  nand (_16078_, _16077_, _16072_);
  nand (_16079_, _16078_, _00561_);
  nand (_16080_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3]);
  nand (_16081_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3]);
  nand (_16082_, _16081_, _16080_);
  nand (_16083_, _16082_, _01417_);
  nand (_16084_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3]);
  nand (_16085_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3]);
  nand (_16086_, _16085_, _16084_);
  nand (_16087_, _16086_, _00227_);
  nand (_16088_, _16087_, _16083_);
  nand (_16089_, _16088_, _00560_);
  nand (_16090_, _16089_, _16079_);
  nand (_16091_, _16090_, _00466_);
  nand (_16092_, _16091_, _16068_);
  nand (_16093_, _16092_, _00247_);
  nor (_16094_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3]);
  nor (_16095_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3]);
  nor (_16096_, _16095_, _16094_);
  nand (_16097_, _16096_, _00227_);
  nand (_16098_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3]);
  nand (_16099_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3]);
  nand (_16100_, _16099_, _16098_);
  nand (_16101_, _16100_, _01417_);
  nand (_16102_, _16101_, _16097_);
  nand (_16103_, _16102_, _00561_);
  nor (_16104_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3]);
  nor (_16105_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3]);
  nor (_16106_, _16105_, _16104_);
  nand (_16107_, _16106_, _00227_);
  nand (_16108_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3]);
  nand (_16109_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3]);
  nand (_16110_, _16109_, _16108_);
  nand (_16111_, _16110_, _01417_);
  nand (_16112_, _16111_, _16107_);
  nand (_16113_, _16112_, _00560_);
  nand (_16114_, _16113_, _16103_);
  nand (_16115_, _16114_, _00465_);
  nand (_16116_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3]);
  nand (_16117_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3]);
  nand (_16118_, _16117_, _16116_);
  nand (_16119_, _16118_, _01417_);
  nand (_16120_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3]);
  nand (_16121_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3]);
  nand (_16122_, _16121_, _16120_);
  nand (_16123_, _16122_, _00227_);
  nand (_16124_, _16123_, _16119_);
  nand (_16125_, _16124_, _00561_);
  nand (_16126_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3]);
  nand (_16127_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3]);
  nand (_16128_, _16127_, _16126_);
  nand (_16129_, _16128_, _01417_);
  nand (_16130_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3]);
  nand (_16131_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3]);
  nand (_16132_, _16131_, _16130_);
  nand (_16133_, _16132_, _00227_);
  nand (_16134_, _16133_, _16129_);
  nand (_16136_, _16134_, _00560_);
  nand (_16137_, _16136_, _16125_);
  nand (_16138_, _16137_, _00466_);
  nand (_16139_, _16138_, _16115_);
  nand (_16140_, _16139_, _00248_);
  nand (_16141_, _16140_, _16093_);
  nand (_16142_, _16141_, _00319_);
  nand (_16143_, _16142_, _16045_);
  nor (_16144_, _16143_, _01629_);
  nor (_16145_, _16144_, _15947_);
  nor (_16146_, _16145_, _00556_);
  nor (_16147_, _16146_, _15755_);
  nor (_16148_, _16147_, _01416_);
  not (_16149_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  nand (_16150_, _01416_, _16149_);
  nand (_16151_, _16150_, _23493_);
  nor (_08635_, _16151_, _16148_);
  nor (_16152_, _22425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1]);
  nor (_16153_, _22427_, _21474_);
  nor (_25106_, _16153_, _16152_);
  nor (_16155_, _22547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  nor (_16156_, _22549_, _21414_);
  nor (_25094_, _16156_, _16155_);
  nor (_16157_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6]);
  nor (_16158_, _22473_, _21504_);
  nor (_08650_, _16158_, _16157_);
  nor (_16159_, _22425_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  nor (_16160_, _22427_, _21586_);
  nor (_08652_, _16160_, _16159_);
  nor (_16161_, _22490_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1]);
  nor (_16162_, _22492_, _21474_);
  nor (_08657_, _16162_, _16161_);
  nor (_08662_, _14058_, _05500_);
  nor (_16163_, _22547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1]);
  nor (_16164_, _22549_, _21474_);
  nor (_08665_, _16164_, _16163_);
  nor (_16165_, _22949_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1]);
  nor (_16166_, _22951_, _21474_);
  nor (_08668_, _16166_, _16165_);
  nor (_16167_, _05356_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1]);
  nor (_16168_, _05358_, _21474_);
  nor (_25274_, _16168_, _16167_);
  nand (_16169_, _23493_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  nor (_08678_, _16169_, _05500_);
  nor (_16170_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3]);
  nor (_16171_, _22498_, _21526_);
  nor (_08680_, _16171_, _16170_);
  nor (_16172_, _12387_, _10381_);
  nor (_16173_, _16172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_08689_, _16173_, rst);
  nor (_16174_, _05500_, _12377_);
  nor (_16175_, _16174_, _15182_);
  nor (_08691_, _16175_, rst);
  nand (_16176_, _05663_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nand (_16177_, _16176_, _14122_);
  nor (_16178_, _16177_, _05667_);
  nor (_16179_, _16178_, _05666_);
  nand (_16180_, _16179_, _15336_);
  nand (_16181_, _15168_, _15308_);
  not (_16182_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_16183_, _05651_, _16182_);
  nor (_16184_, _16183_, _16181_);
  nor (_16185_, _16184_, _05628_);
  nor (_16186_, _05679_, _05622_);
  nand (_16187_, _16186_, _16185_);
  nand (_16188_, _16187_, _16180_);
  nor (_16189_, _16188_, _05606_);
  nand (_16190_, _05606_, _16182_);
  nand (_16191_, _16190_, _23493_);
  nor (_08699_, _16191_, _16189_);
  nor (_16192_, _22535_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  nor (_16193_, _22537_, _21586_);
  nor (_08702_, _16193_, _16192_);
  nor (_16194_, _22547_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7]);
  nor (_16195_, _22549_, _21626_);
  nor (_08705_, _16195_, _16194_);
  nor (_08717_, _00619_, rst);
  not (_16196_, _15336_);
  nor (_16197_, _05660_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_16198_, _16197_, _05661_);
  nor (_16199_, _16198_, _05664_);
  nor (_16200_, _16199_, _05667_);
  nor (_16201_, _16200_, _05666_);
  nor (_16202_, _16201_, _16196_);
  not (_16203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nand (_16204_, _15164_, _16203_);
  nand (_16205_, _16204_, _15197_);
  nand (_16206_, _16205_, _15168_);
  nand (_16207_, _16206_, _15308_);
  nand (_16208_, _16207_, _15306_);
  nand (_16209_, _16208_, _16186_);
  nand (_16210_, _16209_, _05500_);
  nor (_16211_, _16210_, _16202_);
  nand (_16212_, _05606_, _16203_);
  nand (_16213_, _16212_, _23493_);
  nor (_08730_, _16213_, _16211_);
  nor (_16214_, _22991_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7]);
  nor (_16215_, _22993_, _21626_);
  nor (_25112_, _16215_, _16214_);
  not (_16216_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  nor (_16217_, _05500_, _16216_);
  nor (_16218_, _16217_, _15182_);
  nor (_08734_, _16218_, rst);
  nor (_16219_, _01383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  nor (_16220_, _01385_, _21414_);
  nor (_25272_, _16220_, _16219_);
  nor (_16221_, _22922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3]);
  nor (_16222_, _22924_, _21526_);
  nor (_08748_, _16222_, _16221_);
  nand (_16223_, _04935_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_16225_, _16223_, _03702_);
  nand (_16226_, _03924_, _03619_);
  nor (_16227_, _03918_, _03925_);
  nand (_16228_, _16227_, _16226_);
  nor (_16229_, _03939_, _03845_);
  nand (_16230_, _16229_, _03630_);
  nand (_16231_, _16230_, _16228_);
  nand (_16232_, _16231_, _05950_);
  nand (_16233_, _03843_, ABINPUT[6]);
  nand (_16234_, _16233_, _16232_);
  nor (_16235_, _16234_, _16225_);
  nor (_08751_, _16235_, rst);
  not (_16236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand (_16237_, _04938_, _03919_);
  nand (_16238_, _16237_, _16236_);
  nand (_16239_, _03919_, _03923_);
  nand (_16240_, _16239_, _16238_);
  nor (_16241_, _16240_, _03702_);
  nand (_16242_, _03702_, ABINPUT[5]);
  nand (_16243_, _03937_, _03894_);
  nor (_16245_, _16243_, _03631_);
  nand (_16246_, _16245_, _05950_);
  nand (_16247_, _16246_, _16242_);
  nor (_16248_, _16247_, _16241_);
  nor (_08754_, _16248_, rst);
  nor (_16249_, _22434_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7]);
  nor (_16250_, _22437_, _21626_);
  nor (_08756_, _16250_, _16249_);
  nor (_16251_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6]);
  nor (_16252_, _22448_, _21504_);
  nor (_08761_, _16252_, _16251_);
  nand (_16253_, _05840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_16254_, _16253_, _03702_);
  not (_16255_, _05838_);
  nor (_16256_, _03889_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_16257_, _16256_, _03891_);
  nand (_16258_, _16257_, _16255_);
  nand (_16259_, _03940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_16260_, _16259_, _16258_);
  nand (_16261_, _16260_, _05950_);
  nand (_16262_, _03702_, ABINPUT[9]);
  nand (_16263_, _16262_, _16261_);
  nor (_16264_, _16263_, _16254_);
  nor (_08763_, _16264_, rst);
  nand (_16265_, _05840_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_16266_, _16265_, _03702_);
  nor (_16267_, _03676_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_16268_, _16267_, _05838_);
  nand (_16269_, _16268_, _03890_);
  nand (_16270_, _03940_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand (_16272_, _16270_, _16269_);
  nand (_16273_, _16272_, _05950_);
  nand (_16274_, _03702_, ABINPUT[8]);
  nand (_16275_, _16274_, _16273_);
  nor (_16276_, _16275_, _16266_);
  nor (_08765_, _16276_, rst);
  nor (_16277_, _04923_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_16278_, _16277_, _03667_);
  nor (_16279_, _16278_, _04917_);
  nand (_16280_, _16279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand (_16281_, _16280_, _03654_);
  not (_16282_, _16280_);
  nand (_16283_, _16282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_16284_, _16283_, _16281_);
  nor (_16285_, _16284_, _03687_);
  nand (_16286_, _03687_, ABINPUT[6]);
  nand (_16287_, _16286_, _03909_);
  nor (_16288_, _16287_, _16285_);
  nand (_16289_, _03702_, _03654_);
  nand (_16290_, _16289_, _23493_);
  nor (_08768_, _16290_, _16288_);
  nor (_16292_, _03688_, ABINPUT[5]);
  nor (_16293_, _16279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_16294_, _16293_, _16282_);
  nor (_16295_, _16294_, _03687_);
  nor (_16296_, _16295_, _16292_);
  nor (_16297_, _16296_, _03702_);
  nand (_16298_, _03702_, _03631_);
  nand (_16299_, _16298_, _23493_);
  nor (_08771_, _16299_, _16297_);
  nand (_16300_, _03860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand (_16301_, _16300_, _03665_);
  not (_16302_, _16300_);
  nand (_16303_, _16302_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_16304_, _16303_, _16301_);
  nor (_16305_, _16304_, _03687_);
  nand (_16306_, _03687_, ABINPUT[9]);
  nand (_16307_, _16306_, _03909_);
  nor (_16308_, _16307_, _16305_);
  nand (_16309_, _03702_, _03665_);
  nand (_16310_, _16309_, _23493_);
  nor (_08773_, _16310_, _16308_);
  nor (_16311_, _03864_, _03653_);
  nor (_16312_, _03688_, _00129_);
  nand (_16313_, _03860_, _03653_);
  nor (_16314_, _16313_, _03687_);
  nor (_16315_, _16314_, _16312_);
  nor (_16316_, _16315_, _03843_);
  nor (_16317_, _16316_, _16311_);
  nor (_08775_, _16317_, rst);
  not (_16319_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  not (_16320_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nand (_16321_, _16320_, _16319_);
  nor (_16322_, _16321_, _02482_);
  nand (_16323_, _00020_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_16324_, _16323_, _05140_);
  nor (_16325_, _16324_, _02390_);
  nor (_16326_, _16325_, _16322_);
  nor (_16327_, _16326_, _02393_);
  nand (_16328_, _02393_, _00006_);
  nand (_16329_, _16328_, _23493_);
  nor (_08778_, _16329_, _16327_);
  nor (_16330_, _02613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_16331_, _03819_, _02633_);
  not (_16332_, _03832_);
  nor (_16333_, _16332_, _02612_);
  not (_16334_, _03831_);
  nor (_16335_, _16334_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_16336_, _16335_, _16333_);
  nor (_16337_, _16336_, _16331_);
  nor (_16338_, _16337_, _16330_);
  nor (_16339_, _16338_, _02625_);
  nand (_16340_, _02625_, _00121_);
  nand (_16341_, _16340_, _23493_);
  nor (_08780_, _16341_, _16339_);
  nor (_16342_, _03830_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_16343_, _16342_, _16334_);
  nor (_16344_, _03819_, _02634_);
  nor (_16345_, _16344_, _16343_);
  nor (_16346_, _16345_, _03765_);
  nor (_16347_, _03764_, _02664_);
  nor (_16348_, _16347_, _16346_);
  nor (_16349_, _16348_, _03804_);
  nor (_16350_, _02626_, _00006_);
  nor (_16351_, _16350_, _16349_);
  nor (_08782_, _16351_, rst);
  nor (_16352_, _03819_, _02630_);
  nor (_16353_, _02708_, _02705_);
  not (_16354_, _16353_);
  nor (_16355_, _16354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor (_16356_, _16355_, _16352_);
  nor (_16357_, _16356_, _02612_);
  nor (_16358_, _16354_, _02612_);
  nor (_16359_, _16358_, _02662_);
  nor (_16360_, _16359_, _16357_);
  nor (_16361_, _16360_, _02625_);
  nor (_16362_, _02626_, _00129_);
  nor (_16363_, _16362_, _16361_);
  nor (_08784_, _16363_, rst);
  not (_16364_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_16365_, _02708_, _02612_);
  nor (_16366_, _16365_, _16364_);
  nor (_16367_, _03819_, _02631_);
  nor (_16368_, _03835_, _02702_);
  nor (_16369_, _16368_, _16367_);
  nor (_16370_, _16369_, _02612_);
  nor (_16371_, _16370_, _16366_);
  nor (_16372_, _16371_, _02625_);
  nor (_16373_, _02626_, _24900_);
  nor (_16374_, _16373_, _16372_);
  nor (_08786_, _16374_, rst);
  not (_16375_, _02683_);
  nand (_16376_, _16375_, _02636_);
  nand (_16377_, _16376_, _02633_);
  nor (_16378_, _03733_, _02658_);
  nand (_16379_, _16378_, _16377_);
  not (_16380_, _02620_);
  nand (_16381_, _03774_, _02633_);
  nand (_16382_, _16381_, _03776_);
  nor (_16383_, _16382_, _16380_);
  nor (_16385_, _02708_, _02637_);
  nor (_16386_, _16385_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_16387_, _03747_, _02705_);
  nor (_16388_, _16387_, _16386_);
  nor (_16389_, _16388_, _16383_);
  nand (_16390_, _16389_, _16379_);
  nand (_16391_, _16390_, _03764_);
  nand (_16392_, _03765_, ABINPUT[5]);
  nand (_16393_, _16392_, _16391_);
  nand (_16394_, _16393_, _05922_);
  nor (_16395_, _02626_, rst);
  nand (_16396_, _16395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_08789_, _16396_, _16394_);
  nor (_16397_, _04881_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_16398_, _16397_, _02658_);
  nand (_16399_, _16398_, _16376_);
  nor (_16400_, _04884_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_16401_, _03774_, _02620_);
  nor (_16402_, _16401_, _16400_);
  nor (_16403_, _04888_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_16405_, _16385_);
  nand (_16406_, _16405_, _02705_);
  nor (_16407_, _16406_, _16403_);
  nor (_16408_, _16407_, _16402_);
  nand (_16409_, _16408_, _16399_);
  nand (_16410_, _16409_, _03764_);
  nand (_16411_, _03765_, ABINPUT[4]);
  nand (_16412_, _16411_, _16410_);
  nand (_16413_, _16412_, _05922_);
  nand (_16414_, _16395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_08791_, _16414_, _16413_);
  nand (_16415_, _03736_, _02630_);
  nor (_16416_, _03737_, _02658_);
  nand (_16417_, _16416_, _16415_);
  nand (_16418_, _03742_, _02630_);
  nor (_16419_, _03743_, _16380_);
  nand (_16420_, _16419_, _16418_);
  nand (_16421_, _03750_, _02630_);
  nor (_16422_, _03751_, _02707_);
  nand (_16423_, _16422_, _16421_);
  nand (_16424_, _16423_, _16420_);
  nor (_16425_, _16424_, _02612_);
  nand (_16426_, _16425_, _16417_);
  nor (_16427_, _02613_, ABINPUT[8]);
  nor (_16428_, _16427_, _05923_);
  nand (_16429_, _16428_, _16426_);
  nand (_16430_, _16395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_08793_, _16430_, _16429_);
  nand (_16431_, _02612_, _24900_);
  nor (_16432_, _03777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_16433_, _16432_, _03741_);
  nand (_16434_, _16433_, _02620_);
  nor (_16435_, _03735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_16436_, _03736_, _02659_);
  nor (_16437_, _16436_, _16435_);
  nor (_16438_, _03784_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_16439_, _03750_, _02705_);
  nor (_16440_, _16439_, _16438_);
  nor (_16441_, _16440_, _16437_);
  nand (_16442_, _16441_, _16434_);
  nor (_16444_, _16442_, _02612_);
  nor (_16445_, _16444_, _05923_);
  nand (_16446_, _16445_, _16431_);
  nand (_16447_, _16395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_08795_, _16447_, _16446_);
  nor (_16448_, _01383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6]);
  nor (_16449_, _01385_, _21504_);
  nor (_08799_, _16449_, _16448_);
  nor (_16450_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  nand (_16451_, _03721_, _00121_);
  nand (_16452_, _16451_, _23493_);
  nor (_08801_, _16452_, _16450_);
  nor (_16453_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  nand (_16454_, _03721_, _00114_);
  nand (_16455_, _16454_, _23493_);
  nor (_08804_, _16455_, _16453_);
  nor (_16456_, _03721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nand (_16457_, _03721_, _00129_);
  nand (_16458_, _16457_, _23493_);
  nor (_08806_, _16458_, _16456_);
  nor (_08808_, _24841_, rst);
  nand (_16459_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2]);
  nand (_16460_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2]);
  nand (_16461_, _16460_, _16459_);
  nand (_16462_, _16461_, _01417_);
  nand (_16463_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2]);
  nand (_16464_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2]);
  nand (_16465_, _16464_, _16463_);
  nand (_16466_, _16465_, _00227_);
  nand (_16467_, _16466_, _16462_);
  nand (_16468_, _16467_, _00560_);
  nand (_16469_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2]);
  nand (_16470_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2]);
  nand (_16471_, _16470_, _16469_);
  nand (_16472_, _16471_, _01417_);
  nand (_16473_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2]);
  nand (_16474_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2]);
  nand (_16475_, _16474_, _16473_);
  nand (_16476_, _16475_, _00227_);
  nand (_16477_, _16476_, _16472_);
  nand (_16479_, _16477_, _00561_);
  nand (_16480_, _16479_, _16468_);
  nand (_16481_, _16480_, _00466_);
  nor (_16482_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2]);
  nor (_16483_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2]);
  nor (_16484_, _16483_, _16482_);
  nand (_16485_, _16484_, _01417_);
  nor (_16486_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2]);
  nor (_16487_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2]);
  nor (_16488_, _16487_, _16486_);
  nand (_16489_, _16488_, _00227_);
  nand (_16490_, _16489_, _16485_);
  nand (_16491_, _16490_, _00560_);
  nor (_16492_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2]);
  nor (_16493_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2]);
  nor (_16494_, _16493_, _16492_);
  nand (_16495_, _16494_, _01417_);
  nor (_16496_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2]);
  nor (_16497_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2]);
  nor (_16498_, _16497_, _16496_);
  nand (_16499_, _16498_, _00227_);
  nand (_16500_, _16499_, _16495_);
  nand (_16501_, _16500_, _00561_);
  nand (_16502_, _16501_, _16491_);
  nand (_16503_, _16502_, _00465_);
  nand (_16504_, _16503_, _16481_);
  nand (_16505_, _16504_, _00247_);
  nand (_16506_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2]);
  nand (_16507_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2]);
  nand (_16508_, _16507_, _16506_);
  nand (_16509_, _16508_, _01417_);
  nand (_16510_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2]);
  nand (_16511_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2]);
  nand (_16512_, _16511_, _16510_);
  nand (_16513_, _16512_, _00227_);
  nand (_16514_, _16513_, _16509_);
  nand (_16515_, _16514_, _00560_);
  nand (_16516_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2]);
  nand (_16517_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2]);
  nand (_16518_, _16517_, _16516_);
  nand (_16520_, _16518_, _01417_);
  nand (_16521_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2]);
  nand (_16522_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2]);
  nand (_16523_, _16522_, _16521_);
  nand (_16524_, _16523_, _00227_);
  nand (_16525_, _16524_, _16520_);
  nand (_16526_, _16525_, _00561_);
  nand (_16527_, _16526_, _16515_);
  nand (_16528_, _16527_, _00466_);
  nor (_16529_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2]);
  nor (_16530_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2]);
  nor (_16531_, _16530_, _16529_);
  nand (_16532_, _16531_, _00227_);
  nand (_16533_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2]);
  nand (_16534_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2]);
  nand (_16535_, _16534_, _16533_);
  nand (_16536_, _16535_, _01417_);
  nand (_16537_, _16536_, _16532_);
  nand (_16538_, _16537_, _00560_);
  nor (_16539_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2]);
  nor (_16540_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2]);
  nor (_16541_, _16540_, _16539_);
  nand (_16542_, _16541_, _00227_);
  nand (_16543_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2]);
  nand (_16544_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2]);
  nand (_16545_, _16544_, _16543_);
  nand (_16546_, _16545_, _01417_);
  nand (_16547_, _16546_, _16542_);
  nand (_16548_, _16547_, _00561_);
  nand (_16549_, _16548_, _16538_);
  nand (_16551_, _16549_, _00465_);
  nand (_16552_, _16551_, _16528_);
  nand (_16553_, _16552_, _00248_);
  nand (_16554_, _16553_, _16505_);
  nand (_16555_, _16554_, _00320_);
  nand (_16556_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2]);
  nand (_16557_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2]);
  nand (_16558_, _16557_, _16556_);
  nand (_16559_, _16558_, _01417_);
  nand (_16560_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2]);
  nand (_16561_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2]);
  nand (_16562_, _16561_, _16560_);
  nand (_16563_, _16562_, _00227_);
  nand (_16564_, _16563_, _16559_);
  nand (_16565_, _16564_, _00560_);
  nand (_16566_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2]);
  nand (_16567_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2]);
  nand (_16568_, _16567_, _16566_);
  nand (_16569_, _16568_, _01417_);
  nand (_16570_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2]);
  nand (_16571_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2]);
  nand (_16572_, _16571_, _16570_);
  nand (_16573_, _16572_, _00227_);
  nand (_16574_, _16573_, _16569_);
  nand (_16575_, _16574_, _00561_);
  nand (_16576_, _16575_, _16565_);
  nand (_16577_, _16576_, _00466_);
  nor (_16578_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2]);
  nor (_16579_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2]);
  nor (_16580_, _16579_, _16578_);
  nand (_16581_, _16580_, _00227_);
  nand (_16582_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2]);
  nand (_16583_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2]);
  nand (_16584_, _16583_, _16582_);
  nand (_16585_, _16584_, _01417_);
  nand (_16586_, _16585_, _16581_);
  nand (_16587_, _16586_, _00560_);
  nor (_16588_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2]);
  nor (_16589_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2]);
  nor (_16590_, _16589_, _16588_);
  nand (_16591_, _16590_, _00227_);
  nand (_16592_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2]);
  nand (_16593_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2]);
  nand (_16594_, _16593_, _16592_);
  nand (_16595_, _16594_, _01417_);
  nand (_16596_, _16595_, _16591_);
  nand (_16597_, _16596_, _00561_);
  nand (_16598_, _16597_, _16587_);
  nand (_16599_, _16598_, _00465_);
  nand (_16600_, _16599_, _16577_);
  nand (_16602_, _16600_, _00248_);
  nand (_16603_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2]);
  nand (_16604_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2]);
  nand (_16605_, _16604_, _16603_);
  nand (_16606_, _16605_, _01417_);
  nand (_16607_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2]);
  nand (_16608_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2]);
  nand (_16609_, _16608_, _16607_);
  nand (_16610_, _16609_, _00227_);
  nand (_16611_, _16610_, _16606_);
  nand (_16612_, _16611_, _00560_);
  nand (_16613_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2]);
  nand (_16614_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2]);
  nand (_16615_, _16614_, _16613_);
  nand (_16616_, _16615_, _01417_);
  nand (_16617_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2]);
  nand (_16618_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2]);
  nand (_16619_, _16618_, _16617_);
  nand (_16620_, _16619_, _00227_);
  nand (_16621_, _16620_, _16616_);
  nand (_16622_, _16621_, _00561_);
  nand (_16623_, _16622_, _16612_);
  nand (_16624_, _16623_, _00466_);
  nor (_16625_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2]);
  nor (_16626_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2]);
  nor (_16627_, _16626_, _16625_);
  nand (_16628_, _16627_, _01417_);
  nor (_16629_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2]);
  nor (_16630_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2]);
  nor (_16631_, _16630_, _16629_);
  nand (_16632_, _16631_, _00227_);
  nand (_16633_, _16632_, _16628_);
  nand (_16634_, _16633_, _00560_);
  nor (_16635_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2]);
  nor (_16636_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2]);
  nor (_16637_, _16636_, _16635_);
  nand (_16638_, _16637_, _01417_);
  nor (_16639_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2]);
  nor (_16640_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2]);
  nor (_16641_, _16640_, _16639_);
  nand (_16642_, _16641_, _00227_);
  nand (_16643_, _16642_, _16638_);
  nand (_16644_, _16643_, _00561_);
  nand (_16645_, _16644_, _16634_);
  nand (_16646_, _16645_, _00465_);
  nand (_16647_, _16646_, _16624_);
  nand (_16648_, _16647_, _00247_);
  nand (_16649_, _16648_, _16602_);
  nand (_16650_, _16649_, _00319_);
  nand (_16651_, _16650_, _16555_);
  nor (_16652_, _16651_, _00386_);
  nand (_16653_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2]);
  nand (_16654_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2]);
  nand (_16655_, _16654_, _16653_);
  nand (_16656_, _16655_, _01417_);
  nand (_16657_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2]);
  nand (_16658_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2]);
  nand (_16659_, _16658_, _16657_);
  nand (_16660_, _16659_, _00227_);
  nand (_16661_, _16660_, _16656_);
  nand (_16662_, _16661_, _00560_);
  nand (_16663_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2]);
  nand (_16664_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2]);
  nand (_16665_, _16664_, _16663_);
  nand (_16666_, _16665_, _01417_);
  nand (_16667_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2]);
  nand (_16668_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2]);
  nand (_16669_, _16668_, _16667_);
  nand (_16670_, _16669_, _00227_);
  nand (_16671_, _16670_, _16666_);
  nand (_16673_, _16671_, _00561_);
  nand (_16674_, _16673_, _16662_);
  nand (_16675_, _16674_, _00466_);
  nor (_16676_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2]);
  nor (_16677_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2]);
  nor (_16678_, _16677_, _16676_);
  nand (_16679_, _16678_, _00227_);
  nand (_16680_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2]);
  nand (_16681_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2]);
  nand (_16682_, _16681_, _16680_);
  nand (_16683_, _16682_, _01417_);
  nand (_16684_, _16683_, _16679_);
  nand (_16685_, _16684_, _00560_);
  nor (_16686_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2]);
  nor (_16687_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2]);
  nor (_16688_, _16687_, _16686_);
  nand (_16689_, _16688_, _00227_);
  nand (_16690_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2]);
  nand (_16691_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2]);
  nand (_16692_, _16691_, _16690_);
  nand (_16694_, _16692_, _01417_);
  nand (_16695_, _16694_, _16689_);
  nand (_16696_, _16695_, _00561_);
  nand (_16697_, _16696_, _16685_);
  nand (_16698_, _16697_, _00465_);
  nand (_16699_, _16698_, _16675_);
  nand (_16700_, _16699_, _00248_);
  nand (_16701_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2]);
  nand (_16702_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2]);
  nand (_16703_, _16702_, _16701_);
  nand (_16704_, _16703_, _01417_);
  nand (_16705_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2]);
  nand (_16706_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2]);
  nand (_16707_, _16706_, _16705_);
  nand (_16708_, _16707_, _00227_);
  nand (_16709_, _16708_, _16704_);
  nand (_16710_, _16709_, _00560_);
  nand (_16711_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2]);
  nand (_16712_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2]);
  nand (_16713_, _16712_, _16711_);
  nand (_16714_, _16713_, _01417_);
  nand (_16715_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2]);
  nand (_16716_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2]);
  nand (_16717_, _16716_, _16715_);
  nand (_16718_, _16717_, _00227_);
  nand (_16719_, _16718_, _16714_);
  nand (_16720_, _16719_, _00561_);
  nand (_16721_, _16720_, _16710_);
  nand (_16722_, _16721_, _00466_);
  nor (_16723_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2]);
  nor (_16725_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2]);
  nor (_16726_, _16725_, _16723_);
  nand (_16727_, _16726_, _01417_);
  nor (_16728_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2]);
  nor (_16729_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2]);
  nor (_16730_, _16729_, _16728_);
  nand (_16731_, _16730_, _00227_);
  nand (_16732_, _16731_, _16727_);
  nand (_16733_, _16732_, _00560_);
  nor (_16734_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2]);
  nor (_16735_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2]);
  nor (_16736_, _16735_, _16734_);
  nand (_16737_, _16736_, _01417_);
  nor (_16738_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2]);
  nor (_16739_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2]);
  nor (_16740_, _16739_, _16738_);
  nand (_16741_, _16740_, _00227_);
  nand (_16742_, _16741_, _16737_);
  nand (_16743_, _16742_, _00561_);
  nand (_16744_, _16743_, _16733_);
  nand (_16745_, _16744_, _00465_);
  nand (_16746_, _16745_, _16722_);
  nand (_16747_, _16746_, _00247_);
  nand (_16748_, _16747_, _16700_);
  nand (_16749_, _16748_, _00320_);
  nor (_16750_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2]);
  nor (_16751_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2]);
  nor (_16752_, _16751_, _16750_);
  nand (_16753_, _16752_, _01417_);
  nor (_16754_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2]);
  nor (_16755_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2]);
  nor (_16756_, _16755_, _16754_);
  nand (_16757_, _16756_, _00227_);
  nand (_16758_, _16757_, _16753_);
  nand (_16759_, _16758_, _00561_);
  nor (_16760_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2]);
  nor (_16761_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2]);
  nor (_16762_, _16761_, _16760_);
  nand (_16763_, _16762_, _01417_);
  nor (_16764_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2]);
  nor (_16765_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2]);
  nor (_16766_, _16765_, _16764_);
  nand (_16767_, _16766_, _00227_);
  nand (_16768_, _16767_, _16763_);
  nand (_16769_, _16768_, _00560_);
  nand (_16770_, _16769_, _16759_);
  nand (_16771_, _16770_, _00465_);
  nand (_16772_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2]);
  nand (_16773_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2]);
  nand (_16774_, _16773_, _16772_);
  nand (_16775_, _16774_, _01417_);
  nand (_16776_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2]);
  nand (_16777_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2]);
  nand (_16778_, _16777_, _16776_);
  nand (_16779_, _16778_, _00227_);
  nand (_16780_, _16779_, _16775_);
  nand (_16781_, _16780_, _00561_);
  nand (_16782_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2]);
  nand (_16783_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2]);
  nand (_16784_, _16783_, _16782_);
  nand (_16785_, _16784_, _01417_);
  nand (_16786_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2]);
  nand (_16787_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2]);
  nand (_16788_, _16787_, _16786_);
  nand (_16789_, _16788_, _00227_);
  nand (_16790_, _16789_, _16785_);
  nand (_16791_, _16790_, _00560_);
  nand (_16792_, _16791_, _16781_);
  nand (_16793_, _16792_, _00466_);
  nand (_16794_, _16793_, _16771_);
  nand (_16795_, _16794_, _00247_);
  nor (_16796_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2]);
  nor (_16797_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2]);
  nor (_16798_, _16797_, _16796_);
  nand (_16799_, _16798_, _00227_);
  nand (_16800_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2]);
  nand (_16801_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2]);
  nand (_16802_, _16801_, _16800_);
  nand (_16803_, _16802_, _01417_);
  nand (_16804_, _16803_, _16799_);
  nand (_16805_, _16804_, _00561_);
  nor (_16806_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2]);
  nor (_16807_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2]);
  nor (_16808_, _16807_, _16806_);
  nand (_16809_, _16808_, _00227_);
  nand (_16810_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2]);
  nand (_16811_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2]);
  nand (_16812_, _16811_, _16810_);
  nand (_16813_, _16812_, _01417_);
  nand (_16814_, _16813_, _16809_);
  nand (_16815_, _16814_, _00560_);
  nand (_16816_, _16815_, _16805_);
  nand (_16817_, _16816_, _00465_);
  nand (_16818_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2]);
  nand (_16819_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2]);
  nand (_16820_, _16819_, _16818_);
  nand (_16821_, _16820_, _01417_);
  nand (_16822_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2]);
  nand (_16823_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2]);
  nand (_16824_, _16823_, _16822_);
  nand (_16826_, _16824_, _00227_);
  nand (_16827_, _16826_, _16821_);
  nand (_16828_, _16827_, _00561_);
  nand (_16829_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2]);
  nand (_16830_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2]);
  nand (_16831_, _16830_, _16829_);
  nand (_16832_, _16831_, _01417_);
  nand (_16833_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2]);
  nand (_16834_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2]);
  nand (_16835_, _16834_, _16833_);
  nand (_16836_, _16835_, _00227_);
  nand (_16837_, _16836_, _16832_);
  nand (_16838_, _16837_, _00560_);
  nand (_16839_, _16838_, _16828_);
  nand (_16840_, _16839_, _00466_);
  nand (_16841_, _16840_, _16817_);
  nand (_16842_, _16841_, _00248_);
  nand (_16843_, _16842_, _16795_);
  nand (_16844_, _16843_, _00319_);
  nand (_16845_, _16844_, _16749_);
  nor (_16847_, _16845_, _01629_);
  nor (_16848_, _16847_, _16652_);
  nor (_16849_, _16848_, _00156_);
  nand (_16850_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  nand (_16851_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  nand (_16852_, _16851_, _16850_);
  nand (_16853_, _16852_, _01417_);
  nand (_16854_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2]);
  nand (_16855_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2]);
  nand (_16856_, _16855_, _16854_);
  nand (_16857_, _16856_, _00227_);
  nand (_16858_, _16857_, _16853_);
  nand (_16859_, _16858_, _00560_);
  nand (_16860_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2]);
  nand (_16861_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2]);
  nand (_16862_, _16861_, _16860_);
  nand (_16863_, _16862_, _01417_);
  nand (_16864_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  nand (_16865_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2]);
  nand (_16866_, _16865_, _16864_);
  nand (_16868_, _16866_, _00227_);
  nand (_16869_, _16868_, _16863_);
  nand (_16870_, _16869_, _00561_);
  nand (_16871_, _16870_, _16859_);
  nand (_16872_, _16871_, _00466_);
  nor (_16873_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2]);
  nor (_16874_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2]);
  nor (_16875_, _16874_, _16873_);
  nand (_16876_, _16875_, _00227_);
  nand (_16877_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2]);
  nand (_16878_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2]);
  nand (_16879_, _16878_, _16877_);
  nand (_16880_, _16879_, _01417_);
  nand (_16881_, _16880_, _16876_);
  nand (_16882_, _16881_, _00560_);
  nor (_16883_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2]);
  nor (_16884_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2]);
  nor (_16885_, _16884_, _16883_);
  nand (_16886_, _16885_, _00227_);
  nand (_16887_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2]);
  nand (_16888_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2]);
  nand (_16889_, _16888_, _16887_);
  nand (_16890_, _16889_, _01417_);
  nand (_16891_, _16890_, _16886_);
  nand (_16892_, _16891_, _00561_);
  nand (_16893_, _16892_, _16882_);
  nand (_16894_, _16893_, _00465_);
  nand (_16895_, _16894_, _16872_);
  nand (_16896_, _16895_, _00248_);
  nand (_16897_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2]);
  nand (_16898_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2]);
  nand (_16899_, _16898_, _16897_);
  nand (_16900_, _16899_, _01417_);
  nand (_16901_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2]);
  nand (_16902_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2]);
  nand (_16903_, _16902_, _16901_);
  nand (_16904_, _16903_, _00227_);
  nand (_16905_, _16904_, _16900_);
  nand (_16906_, _16905_, _00560_);
  nand (_16907_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2]);
  nand (_16909_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2]);
  nand (_16910_, _16909_, _16907_);
  nand (_16911_, _16910_, _01417_);
  nand (_16912_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2]);
  nand (_16913_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2]);
  nand (_16914_, _16913_, _16912_);
  nand (_16915_, _16914_, _00227_);
  nand (_16916_, _16915_, _16911_);
  nand (_16917_, _16916_, _00561_);
  nand (_16918_, _16917_, _16906_);
  nand (_16919_, _16918_, _00466_);
  nor (_16920_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2]);
  nor (_16921_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2]);
  nor (_16922_, _16921_, _16920_);
  nand (_16923_, _16922_, _01417_);
  nor (_16924_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2]);
  nor (_16925_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2]);
  nor (_16926_, _16925_, _16924_);
  nand (_16927_, _16926_, _00227_);
  nand (_16928_, _16927_, _16923_);
  nand (_16930_, _16928_, _00560_);
  nor (_16931_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2]);
  nor (_16932_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2]);
  nor (_16933_, _16932_, _16931_);
  nand (_16934_, _16933_, _01417_);
  nor (_16935_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2]);
  nor (_16936_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2]);
  nor (_16937_, _16936_, _16935_);
  nand (_16938_, _16937_, _00227_);
  nand (_16939_, _16938_, _16934_);
  nand (_16940_, _16939_, _00561_);
  nand (_16941_, _16940_, _16930_);
  nand (_16942_, _16941_, _00465_);
  nand (_16943_, _16942_, _16919_);
  nand (_16944_, _16943_, _00247_);
  nand (_16945_, _16944_, _16896_);
  nand (_16946_, _16945_, _00319_);
  nand (_16947_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2]);
  nand (_16948_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2]);
  nand (_16949_, _16948_, _16947_);
  nand (_16951_, _16949_, _01417_);
  nand (_16952_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2]);
  nand (_16953_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2]);
  nand (_16954_, _16953_, _16952_);
  nand (_16955_, _16954_, _00227_);
  nand (_16956_, _16955_, _16951_);
  nand (_16957_, _16956_, _00560_);
  nand (_16958_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2]);
  nand (_16959_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2]);
  nand (_16960_, _16959_, _16958_);
  nand (_16961_, _16960_, _01417_);
  nand (_16962_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2]);
  nand (_16963_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2]);
  nand (_16964_, _16963_, _16962_);
  nand (_16965_, _16964_, _00227_);
  nand (_16966_, _16965_, _16961_);
  nand (_16967_, _16966_, _00561_);
  nand (_16968_, _16967_, _16957_);
  nand (_16969_, _16968_, _00466_);
  nor (_16970_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2]);
  nor (_16972_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2]);
  nor (_16973_, _16972_, _16970_);
  nand (_16974_, _16973_, _01417_);
  nor (_16975_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2]);
  nor (_16976_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2]);
  nor (_16977_, _16976_, _16975_);
  nand (_16978_, _16977_, _00227_);
  nand (_16979_, _16978_, _16974_);
  nand (_16980_, _16979_, _00560_);
  nor (_16981_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2]);
  nor (_16982_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2]);
  nor (_16983_, _16982_, _16981_);
  nand (_16984_, _16983_, _01417_);
  nor (_16985_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2]);
  nor (_16986_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2]);
  nor (_16987_, _16986_, _16985_);
  nand (_16988_, _16987_, _00227_);
  nand (_16989_, _16988_, _16984_);
  nand (_16990_, _16989_, _00561_);
  nand (_16991_, _16990_, _16980_);
  nand (_16993_, _16991_, _00465_);
  nand (_16994_, _16993_, _16969_);
  nand (_16995_, _16994_, _00247_);
  nand (_16996_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2]);
  nand (_16997_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2]);
  nand (_16998_, _16997_, _16996_);
  nand (_16999_, _16998_, _01417_);
  nand (_17000_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2]);
  nand (_17001_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2]);
  nand (_17002_, _17001_, _17000_);
  nand (_17003_, _17002_, _00227_);
  nand (_17004_, _17003_, _16999_);
  nand (_17005_, _17004_, _00560_);
  nand (_17006_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2]);
  nand (_17007_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2]);
  nand (_17008_, _17007_, _17006_);
  nand (_17009_, _17008_, _01417_);
  nand (_17010_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2]);
  nand (_17011_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2]);
  nand (_17012_, _17011_, _17010_);
  nand (_17014_, _17012_, _00227_);
  nand (_17015_, _17014_, _17009_);
  nand (_17016_, _17015_, _00561_);
  nand (_17017_, _17016_, _17005_);
  nand (_17018_, _17017_, _00466_);
  nor (_17019_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2]);
  nor (_17020_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2]);
  nor (_17021_, _17020_, _17019_);
  nand (_17022_, _17021_, _00227_);
  nand (_17023_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2]);
  nand (_17024_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2]);
  nand (_17025_, _17024_, _17023_);
  nand (_17026_, _17025_, _01417_);
  nand (_17027_, _17026_, _17022_);
  nand (_17028_, _17027_, _00560_);
  nor (_17029_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2]);
  nor (_17030_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2]);
  nor (_17031_, _17030_, _17029_);
  nand (_17032_, _17031_, _00227_);
  nand (_17033_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2]);
  nand (_17035_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2]);
  nand (_17036_, _17035_, _17033_);
  nand (_17037_, _17036_, _01417_);
  nand (_17038_, _17037_, _17032_);
  nand (_17039_, _17038_, _00561_);
  nand (_17040_, _17039_, _17028_);
  nand (_17041_, _17040_, _00465_);
  nand (_17042_, _17041_, _17018_);
  nand (_17043_, _17042_, _00248_);
  nand (_17044_, _17043_, _16995_);
  nand (_17045_, _17044_, _00320_);
  nand (_17046_, _17045_, _16946_);
  nor (_17047_, _17046_, _00386_);
  nand (_17048_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2]);
  nand (_17049_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2]);
  nand (_17050_, _17049_, _17048_);
  nand (_17051_, _17050_, _00227_);
  nand (_17052_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2]);
  nand (_17053_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2]);
  nand (_17054_, _17053_, _17052_);
  nand (_17055_, _17054_, _01417_);
  nand (_17056_, _17055_, _17051_);
  nand (_17057_, _17056_, _00560_);
  nand (_17058_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2]);
  nand (_17059_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2]);
  nand (_17060_, _17059_, _17058_);
  nand (_17061_, _17060_, _00227_);
  nand (_17062_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2]);
  nand (_17063_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2]);
  nand (_17064_, _17063_, _17062_);
  nand (_17065_, _17064_, _01417_);
  nand (_17066_, _17065_, _17061_);
  nand (_17067_, _17066_, _00561_);
  nand (_17068_, _17067_, _17057_);
  nand (_17069_, _17068_, _00466_);
  nand (_17070_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  nand (_17071_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2]);
  nand (_17072_, _17071_, _17070_);
  nand (_17073_, _17072_, _01417_);
  nor (_17074_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  nor (_17075_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2]);
  nor (_17076_, _17075_, _17074_);
  nand (_17077_, _17076_, _00227_);
  nand (_17078_, _17077_, _17073_);
  nand (_17079_, _17078_, _00560_);
  nand (_17080_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2]);
  nand (_17081_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2]);
  nand (_17082_, _17081_, _17080_);
  nand (_17083_, _17082_, _01417_);
  nor (_17084_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2]);
  nor (_17086_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2]);
  nor (_17087_, _17086_, _17084_);
  nand (_17088_, _17087_, _00227_);
  nand (_17089_, _17088_, _17083_);
  nand (_17090_, _17089_, _00561_);
  nand (_17091_, _17090_, _17079_);
  nand (_17092_, _17091_, _00465_);
  nand (_17093_, _17092_, _17069_);
  nand (_17094_, _17093_, _00248_);
  nand (_17095_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2]);
  nand (_17096_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2]);
  nand (_17097_, _17096_, _17095_);
  nand (_17098_, _17097_, _01417_);
  nand (_17099_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2]);
  nand (_17100_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2]);
  nand (_17101_, _17100_, _17099_);
  nand (_17102_, _17101_, _00227_);
  nand (_17103_, _17102_, _17098_);
  nand (_17104_, _17103_, _00560_);
  nand (_17105_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2]);
  nand (_17107_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2]);
  nand (_17108_, _17107_, _17105_);
  nand (_17109_, _17108_, _01417_);
  nand (_17110_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2]);
  nand (_17111_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2]);
  nand (_17112_, _17111_, _17110_);
  nand (_17113_, _17112_, _00227_);
  nand (_17114_, _17113_, _17109_);
  nand (_17115_, _17114_, _00561_);
  nand (_17116_, _17115_, _17104_);
  nand (_17117_, _17116_, _00466_);
  nor (_17118_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2]);
  nor (_17119_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2]);
  nor (_17120_, _17119_, _17118_);
  nand (_17121_, _17120_, _01417_);
  nor (_17122_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2]);
  nor (_17123_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2]);
  nor (_17124_, _17123_, _17122_);
  nand (_17125_, _17124_, _00227_);
  nand (_17126_, _17125_, _17121_);
  nand (_17127_, _17126_, _00560_);
  nor (_17128_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2]);
  nor (_17129_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2]);
  nor (_17130_, _17129_, _17128_);
  nor (_17131_, _17130_, _00227_);
  nor (_17132_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2]);
  nor (_17133_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2]);
  nor (_17134_, _17133_, _17132_);
  nor (_17135_, _17134_, _01417_);
  nor (_17136_, _17135_, _17131_);
  nand (_17138_, _17136_, _00561_);
  nand (_17139_, _17138_, _17127_);
  nand (_17140_, _17139_, _00465_);
  nand (_17141_, _17140_, _17117_);
  nand (_17142_, _17141_, _00247_);
  nand (_17143_, _17142_, _17094_);
  nand (_17144_, _17143_, _00320_);
  nand (_17145_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2]);
  nand (_17146_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2]);
  nand (_17147_, _17146_, _17145_);
  nand (_17148_, _17147_, _01417_);
  nand (_17149_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2]);
  nand (_17150_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2]);
  nand (_17151_, _17150_, _17149_);
  nand (_17152_, _17151_, _00227_);
  nand (_17153_, _17152_, _17148_);
  nand (_17154_, _17153_, _00560_);
  nand (_17155_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2]);
  nand (_17156_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2]);
  nand (_17157_, _17156_, _17155_);
  nand (_17159_, _17157_, _01417_);
  nand (_17160_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2]);
  nand (_17161_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2]);
  nand (_17162_, _17161_, _17160_);
  nand (_17163_, _17162_, _00227_);
  nand (_17164_, _17163_, _17159_);
  nand (_17165_, _17164_, _00561_);
  nand (_17166_, _17165_, _17154_);
  nand (_17167_, _17166_, _00466_);
  nor (_17168_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2]);
  nor (_17170_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2]);
  nor (_17171_, _17170_, _17168_);
  nand (_17172_, _17171_, _01417_);
  nor (_17173_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2]);
  nor (_17174_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2]);
  nor (_17175_, _17174_, _17173_);
  nand (_17176_, _17175_, _00227_);
  nand (_17177_, _17176_, _17172_);
  nand (_17178_, _17177_, _00560_);
  nor (_17179_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2]);
  nor (_17181_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2]);
  nor (_17182_, _17181_, _17179_);
  nand (_17183_, _17182_, _01417_);
  nor (_17184_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2]);
  nor (_17185_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2]);
  nor (_17186_, _17185_, _17184_);
  nand (_17187_, _17186_, _00227_);
  nand (_17188_, _17187_, _17183_);
  nand (_17189_, _17188_, _00561_);
  nand (_17190_, _17189_, _17178_);
  nand (_17191_, _17190_, _00465_);
  nand (_17192_, _17191_, _17167_);
  nand (_17193_, _17192_, _00247_);
  nand (_17194_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2]);
  nand (_17195_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2]);
  nand (_17196_, _17195_, _17194_);
  nand (_17197_, _17196_, _01417_);
  nand (_17198_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2]);
  nand (_17199_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2]);
  nand (_17200_, _17199_, _17198_);
  nand (_17201_, _17200_, _00227_);
  nand (_17202_, _17201_, _17197_);
  nand (_17203_, _17202_, _00560_);
  nand (_17204_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2]);
  nand (_17205_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2]);
  nand (_17206_, _17205_, _17204_);
  nand (_17207_, _17206_, _01417_);
  nand (_17208_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2]);
  nand (_17209_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2]);
  nand (_17210_, _17209_, _17208_);
  nand (_17212_, _17210_, _00227_);
  nand (_17213_, _17212_, _17207_);
  nand (_17214_, _17213_, _00561_);
  nand (_17215_, _17214_, _17203_);
  nand (_17216_, _17215_, _00466_);
  nor (_17217_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2]);
  nor (_17218_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2]);
  nor (_17219_, _17218_, _17217_);
  nand (_17220_, _17219_, _01417_);
  nor (_17221_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2]);
  nor (_17222_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2]);
  nor (_17223_, _17222_, _17221_);
  nand (_17224_, _17223_, _00227_);
  nand (_17225_, _17224_, _17220_);
  nand (_17226_, _17225_, _00560_);
  nor (_17227_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  nor (_17228_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2]);
  nor (_17229_, _17228_, _17227_);
  nand (_17230_, _17229_, _01417_);
  nor (_17231_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2]);
  nor (_17233_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2]);
  nor (_17234_, _17233_, _17231_);
  nand (_17235_, _17234_, _00227_);
  nand (_17236_, _17235_, _17230_);
  nand (_17237_, _17236_, _00561_);
  nand (_17238_, _17237_, _17226_);
  nand (_17239_, _17238_, _00465_);
  nand (_17240_, _17239_, _17216_);
  nand (_17241_, _17240_, _00248_);
  nand (_17242_, _17241_, _17193_);
  nand (_17243_, _17242_, _00319_);
  nand (_17244_, _17243_, _17144_);
  nor (_17245_, _17244_, _01629_);
  nor (_17246_, _17245_, _17047_);
  nor (_17247_, _17246_, _00556_);
  nor (_17248_, _17247_, _16849_);
  nor (_17249_, _17248_, _01416_);
  not (_17250_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  nand (_17251_, _01416_, _17250_);
  nand (_17252_, _17251_, _23493_);
  nor (_08814_, _17252_, _17249_);
  nor (_17253_, _21733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6]);
  nor (_17254_, _21735_, _21504_);
  nor (_08817_, _17254_, _17253_);
  nor (_25038_[2], _00517_, rst);
  nor (_17255_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7]);
  nor (_17256_, _22448_, _21626_);
  nor (_25092_, _17256_, _17255_);
  nor (_08822_, _00455_, rst);
  nor (_17257_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  nor (_17259_, _22448_, _21414_);
  nor (_08825_, _17259_, _17257_);
  nor (_17260_, _22922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  nor (_17261_, _22924_, _21414_);
  nor (_08827_, _17261_, _17260_);
  nor (_17262_, _21752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2]);
  nor (_17263_, _21754_, _21554_);
  nor (_08829_, _17263_, _17262_);
  nor (_17264_, _09002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6]);
  nor (_17265_, _09004_, _21504_);
  nor (_08831_, _17265_, _17264_);
  nor (_17266_, _12387_, _24170_);
  nor (_17267_, _17266_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_08833_, _17267_, rst);
  nor (_17268_, _22922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2]);
  nor (_17269_, _22924_, _21554_);
  nor (_08836_, _17269_, _17268_);
  not (_17270_, _05289_);
  nor (_17271_, _00225_, _00461_);
  not (_17272_, _17271_);
  nor (_17273_, _17272_, _05222_);
  nand (_17274_, _17273_, _17270_);
  nand (_17275_, _17274_, _11778_);
  nand (_17276_, _05236_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nand (_17277_, _05215_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_17278_, _17277_, _17276_);
  nand (_17279_, _17278_, _00531_);
  not (_17280_, _05236_);
  nor (_17281_, _17280_, _11689_);
  nor (_17282_, _05216_, _11650_);
  nor (_17283_, _17282_, _17281_);
  nor (_17284_, _17283_, _00531_);
  nand (_17285_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand (_17286_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nand (_17287_, _17286_, _17285_);
  nand (_17288_, _17287_, _05303_);
  nand (_17289_, _00671_, _11669_);
  nor (_17290_, _00634_, _00052_);
  not (_17291_, _17290_);
  nor (_17292_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_17293_, _17292_, _17291_);
  nand (_17294_, _17293_, _17289_);
  nand (_17295_, _17294_, _17288_);
  nor (_17296_, _17295_, _17284_);
  nand (_17297_, _17296_, _17279_);
  nand (_17298_, _17297_, _17273_);
  nor (_17299_, _00225_, _00641_);
  not (_17300_, _17299_);
  nor (_17301_, _00318_, _00385_);
  nand (_17302_, _17301_, _00156_);
  nor (_17303_, _17302_, _17300_);
  nand (_17304_, _05236_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nand (_17305_, _05215_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_17306_, _17305_, _17304_);
  nand (_17307_, _17306_, _00671_);
  nor (_17308_, _17280_, _06618_);
  nor (_17309_, _05216_, _01090_);
  nor (_17310_, _17309_, _17308_);
  nor (_17311_, _17310_, _00671_);
  nand (_17312_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_17313_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  nand (_17314_, _17313_, _17312_);
  nand (_17315_, _17314_, _05303_);
  not (_17316_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  nand (_17317_, _00671_, _17316_);
  nor (_17318_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  nor (_17319_, _17318_, _17291_);
  nand (_17320_, _17319_, _17317_);
  nand (_17321_, _17320_, _17315_);
  nor (_17322_, _17321_, _17311_);
  nand (_17323_, _17322_, _17307_);
  nand (_17324_, _17323_, _17303_);
  nand (_17325_, _17324_, _17298_);
  nor (_17326_, _00246_, _00461_);
  not (_17327_, _17326_);
  nor (_17328_, _17327_, _05238_);
  nor (_17329_, _23424_, _23382_);
  nor (_17330_, _14335_, _24761_);
  not (_17331_, _17330_);
  nor (_17332_, _17331_, _17329_);
  nor (_17333_, _23454_, _23326_);
  nor (_17334_, _14340_, _24391_);
  not (_17335_, _17334_);
  nor (_17336_, _17335_, _17333_);
  nor (_17337_, _23436_, _23425_);
  nand (_17338_, _17337_, _17336_);
  nor (_17339_, _14329_, _23469_);
  not (_17340_, _17339_);
  nor (_17341_, _17340_, _17338_);
  nand (_17342_, _17341_, _17332_);
  nor (_17343_, _17342_, _24481_);
  nor (_17344_, _17343_, _24460_);
  not (_17345_, _17344_);
  nor (_17346_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nor (_17347_, _17344_, p1_in[1]);
  nor (_17348_, _17347_, _17346_);
  nand (_17349_, _17348_, _00671_);
  nand (_17350_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  nand (_17351_, _17345_, p1_in[5]);
  nand (_17352_, _17351_, _17350_);
  nand (_17353_, _17352_, _00531_);
  nand (_17354_, _17353_, _17349_);
  nand (_17355_, _17354_, _02437_);
  nor (_17356_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  nor (_17357_, _17344_, p1_in[3]);
  nor (_17358_, _17357_, _17356_);
  nand (_17359_, _17358_, _00671_);
  nand (_17360_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nand (_17361_, _17345_, p1_in[7]);
  nand (_17362_, _17361_, _17360_);
  nand (_17363_, _17362_, _00531_);
  nand (_17364_, _17363_, _17359_);
  nand (_17365_, _17364_, _00052_);
  nand (_17366_, _17365_, _17355_);
  nand (_17367_, _17366_, _00647_);
  nand (_17368_, _17345_, p1_in[4]);
  nand (_17369_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  nand (_17370_, _17369_, _17368_);
  nand (_17371_, _17370_, _00531_);
  nand (_17372_, _17345_, p1_in[0]);
  nand (_17373_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  nand (_17374_, _17373_, _17372_);
  nand (_17375_, _17374_, _00671_);
  nand (_17376_, _17375_, _17371_);
  nand (_17377_, _17376_, _02437_);
  nor (_17378_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  nor (_17379_, _17344_, p1_in[6]);
  nor (_17380_, _17379_, _17378_);
  nand (_17381_, _17380_, _00531_);
  nor (_17382_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  nor (_17383_, _17344_, p1_in[2]);
  nor (_17384_, _17383_, _17382_);
  nand (_17385_, _17384_, _00671_);
  nand (_17386_, _17385_, _17381_);
  nand (_17387_, _17386_, _00052_);
  nand (_17388_, _17387_, _17377_);
  nand (_17389_, _17388_, _00634_);
  nand (_17390_, _17389_, _17367_);
  nand (_17391_, _17390_, _17328_);
  nand (_17392_, _05237_, _00318_);
  nor (_17394_, _17392_, _17300_);
  nand (_17395_, _00531_, _05637_);
  nor (_17396_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  nor (_17397_, _17396_, _00052_);
  nand (_17398_, _17397_, _17395_);
  nor (_17399_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_17400_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nor (_17401_, _17400_, _17399_);
  nand (_17402_, _17401_, _00052_);
  nand (_17403_, _17402_, _17398_);
  nand (_17404_, _17403_, _00647_);
  not (_17405_, _05303_);
  nor (_17406_, _00671_, _14845_);
  nor (_17407_, _00531_, _14952_);
  nor (_17408_, _17407_, _17406_);
  nor (_17409_, _17408_, _17405_);
  nor (_17410_, _00671_, _05645_);
  nor (_17411_, _00531_, _14988_);
  nor (_17412_, _17411_, _17410_);
  nor (_17413_, _17412_, _05216_);
  nor (_17414_, _17413_, _17409_);
  nand (_17415_, _17414_, _17404_);
  nand (_17416_, _17415_, _17394_);
  nand (_17417_, _17416_, _17391_);
  nor (_17418_, _17417_, _17325_);
  not (_17419_, _05283_);
  nand (_17420_, _17419_, \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  not (_17421_, _17302_);
  nand (_17422_, _17326_, _17421_);
  not (_17423_, _17422_);
  nand (_17424_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_17425_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand (_17426_, _17425_, _17424_);
  nand (_17427_, _17426_, _05303_);
  nand (_17428_, _00671_, _24847_);
  nor (_17429_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_17430_, _17429_, _17280_);
  nand (_17431_, _17430_, _17428_);
  nand (_17432_, _00671_, _11504_);
  nor (_17433_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nor (_17434_, _17433_, _17291_);
  nand (_17435_, _17434_, _17432_);
  nand (_17436_, _17435_, _17431_);
  nor (_17437_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_17438_, _11709_, _11697_);
  nand (_17439_, _11709_, _11697_);
  not (_17440_, _17439_);
  nor (_17441_, _17440_, _17438_);
  not (_17442_, _11664_);
  nor (_17443_, _11684_, _17442_);
  nand (_17444_, _11684_, _17442_);
  not (_17445_, _17444_);
  nor (_17446_, _17445_, _17443_);
  nor (_17447_, _17446_, _17441_);
  nand (_17448_, _17446_, _17441_);
  not (_17449_, _17448_);
  nor (_17450_, _17449_, _17447_);
  nor (_17451_, _11724_, _11609_);
  nand (_17452_, _11724_, _11609_);
  not (_17453_, _17452_);
  nor (_17454_, _17453_, _17451_);
  not (_17455_, _11738_);
  nor (_17456_, _11750_, _17455_);
  nor (_17457_, _11751_, _11738_);
  nor (_17458_, _17457_, _17456_);
  not (_17459_, _17458_);
  nor (_17460_, _17459_, _17454_);
  nand (_17461_, _17459_, _17454_);
  not (_17462_, _17461_);
  nor (_17463_, _17462_, _17460_);
  nand (_17465_, _17463_, _17450_);
  not (_17466_, _17450_);
  not (_17467_, _17463_);
  nand (_17468_, _17467_, _17466_);
  nand (_17469_, _17468_, _17465_);
  nand (_17470_, _17469_, _00671_);
  nand (_17471_, _17470_, _05215_);
  nor (_17472_, _17471_, _17437_);
  nor (_17473_, _17472_, _17436_);
  nand (_17474_, _17473_, _17427_);
  nand (_17475_, _17474_, _17423_);
  nand (_17476_, _17475_, _17420_);
  nor (_17477_, _17272_, _05238_);
  nor (_17478_, _17477_, _17273_);
  nand (_17479_, _17478_, _17422_);
  nor (_17480_, _17392_, _00461_);
  not (_17481_, _17480_);
  nor (_17482_, _17327_, _05222_);
  nor (_17483_, _17482_, _17328_);
  nand (_17484_, _17483_, _17481_);
  nor (_17485_, _17484_, _17479_);
  not (_17486_, \oc8051_top_1.oc8051_sfr1.bit_out );
  not (_17487_, _17303_);
  nand (_17488_, _05237_, _00461_);
  nand (_17489_, _17488_, _17487_);
  nor (_17490_, _17489_, _17486_);
  nand (_17491_, _17490_, _17485_);
  nand (_17492_, _00225_, _00461_);
  nor (_17493_, _17492_, _05238_);
  nand (_17494_, _05236_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nand (_17495_, _05215_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_17496_, _17495_, _17494_);
  nand (_17497_, _17496_, _00671_);
  nor (_17498_, _17280_, _14160_);
  nor (_17499_, _05216_, _01060_);
  nor (_17500_, _17499_, _17498_);
  nor (_17501_, _17500_, _00671_);
  nand (_17502_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand (_17503_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nand (_17504_, _17503_, _17502_);
  nand (_17505_, _17504_, _05303_);
  nand (_17506_, _00671_, _16319_);
  nor (_17507_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  nor (_17508_, _17507_, _17291_);
  nand (_17509_, _17508_, _17506_);
  nand (_17510_, _17509_, _17505_);
  nor (_17511_, _17510_, _17501_);
  nand (_17512_, _17511_, _17497_);
  nand (_17513_, _17512_, _17493_);
  nand (_17514_, _17513_, _17491_);
  nor (_17516_, _17514_, _17476_);
  nand (_17517_, _17516_, _17418_);
  nor (_17518_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  nor (_17519_, _17344_, p2_in[1]);
  nor (_17520_, _17519_, _17518_);
  nand (_17521_, _17520_, _00671_);
  nand (_17522_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  nand (_17523_, _17345_, p2_in[5]);
  nand (_17524_, _17523_, _17522_);
  nand (_17525_, _17524_, _00531_);
  nand (_17526_, _17525_, _17521_);
  nand (_17527_, _17526_, _02437_);
  nand (_17528_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nand (_17529_, _17345_, p2_in[7]);
  nand (_17530_, _17529_, _17528_);
  nand (_17531_, _17530_, _00531_);
  nor (_17532_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  nor (_17533_, _17344_, p2_in[3]);
  nor (_17534_, _17533_, _17532_);
  nand (_17535_, _17534_, _00671_);
  nand (_17537_, _17535_, _17531_);
  nand (_17538_, _17537_, _00052_);
  nand (_17539_, _17538_, _17527_);
  nand (_17540_, _17539_, _00647_);
  nand (_17541_, _17345_, p2_in[4]);
  nand (_17542_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  nand (_17543_, _17542_, _17541_);
  nand (_17544_, _17543_, _00531_);
  nand (_17545_, _17345_, p2_in[0]);
  nand (_17546_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  nand (_17547_, _17546_, _17545_);
  nand (_17548_, _17547_, _00671_);
  nand (_17549_, _17548_, _17544_);
  nand (_17550_, _17549_, _02437_);
  nand (_17551_, _17345_, p2_in[2]);
  nand (_17552_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  nand (_17553_, _17552_, _17551_);
  nand (_17554_, _17553_, _00671_);
  nand (_17555_, _17345_, p2_in[6]);
  nand (_17556_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  nand (_17558_, _17556_, _17555_);
  nand (_17559_, _17558_, _00531_);
  nand (_17560_, _17559_, _17554_);
  nand (_17561_, _17560_, _00052_);
  nand (_17562_, _17561_, _17550_);
  nand (_17563_, _17562_, _00634_);
  nand (_17564_, _17563_, _17540_);
  nand (_17565_, _17564_, _00246_);
  nor (_17566_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_17567_, _17344_, p3_in[1]);
  nor (_17568_, _17567_, _17566_);
  nand (_17569_, _17568_, _00671_);
  nand (_17570_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  nand (_17571_, _17345_, p3_in[5]);
  nand (_17572_, _17571_, _17570_);
  nand (_17573_, _17572_, _00531_);
  nand (_17574_, _17573_, _17569_);
  nand (_17575_, _17574_, _02437_);
  nand (_17576_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nand (_17577_, _17345_, p3_in[7]);
  nand (_17579_, _17577_, _17576_);
  nand (_17580_, _17579_, _00531_);
  nor (_17581_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  nor (_17582_, _17344_, p3_in[3]);
  nor (_17583_, _17582_, _17581_);
  nand (_17584_, _17583_, _00671_);
  nand (_17585_, _17584_, _17580_);
  nand (_17586_, _17585_, _00052_);
  nand (_17587_, _17586_, _17575_);
  nand (_17588_, _17587_, _00647_);
  nor (_17589_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  nor (_17590_, _17344_, p3_in[4]);
  nor (_17591_, _17590_, _17589_);
  nand (_17592_, _17591_, _00531_);
  nor (_17593_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  nor (_17594_, _17344_, p3_in[0]);
  nor (_17595_, _17594_, _17593_);
  nand (_17596_, _17595_, _00671_);
  nand (_17597_, _17596_, _17592_);
  nand (_17598_, _17597_, _02437_);
  nor (_17600_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  nor (_17601_, _17344_, p3_in[6]);
  nor (_17602_, _17601_, _17600_);
  nand (_17603_, _17602_, _00531_);
  nor (_17604_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  nor (_17605_, _17344_, p3_in[2]);
  nor (_17606_, _17605_, _17604_);
  nand (_17607_, _17606_, _00671_);
  nand (_17608_, _17607_, _17603_);
  nand (_17609_, _17608_, _00052_);
  nand (_17610_, _17609_, _17598_);
  nand (_17611_, _17610_, _00634_);
  nand (_17612_, _17611_, _17588_);
  nand (_17613_, _17612_, _00225_);
  nand (_17614_, _17613_, _17565_);
  nand (_17615_, _17614_, _17480_);
  nor (_17616_, _05240_, _00641_);
  nand (_17617_, _00531_, _05624_);
  nor (_17618_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nor (_17619_, _17618_, _00052_);
  nand (_17620_, _17619_, _17617_);
  nor (_17621_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nor (_17622_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nor (_17623_, _17622_, _17621_);
  nand (_17624_, _17623_, _00052_);
  nand (_17625_, _17624_, _17620_);
  nand (_17626_, _17625_, _00647_);
  nor (_17627_, _00671_, _02614_);
  nor (_17628_, _00531_, _14665_);
  nor (_17629_, _17628_, _17627_);
  nor (_17630_, _17629_, _17405_);
  nor (_17631_, _00671_, _02678_);
  nor (_17632_, _00531_, _14966_);
  nor (_17633_, _17632_, _17631_);
  nor (_17634_, _17633_, _05216_);
  nor (_17635_, _17634_, _17630_);
  nand (_17636_, _17635_, _17626_);
  nand (_17637_, _17636_, _17616_);
  nor (_17638_, _17492_, _17392_);
  nand (_17639_, _00531_, _05636_);
  nor (_17640_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_17641_, _17640_, _00052_);
  nand (_17642_, _17641_, _17639_);
  nor (_17643_, _00671_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nor (_17644_, _00531_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  nor (_17645_, _17644_, _17643_);
  nand (_17646_, _17645_, _00052_);
  nand (_17647_, _17646_, _17642_);
  nand (_17648_, _17647_, _00647_);
  nor (_17649_, _00671_, _05644_);
  nor (_17651_, _00531_, _05619_);
  nor (_17652_, _17651_, _17649_);
  nor (_17653_, _17652_, _05216_);
  nor (_17654_, _00671_, _14735_);
  nor (_17655_, _00531_, _05629_);
  nor (_17656_, _17655_, _17654_);
  nor (_17657_, _17656_, _17405_);
  nor (_17658_, _17657_, _17653_);
  nand (_17659_, _17658_, _17648_);
  nand (_17660_, _17659_, _17638_);
  nand (_17661_, _17660_, _17637_);
  nor (_17662_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nor (_17663_, _17344_, p0_in[1]);
  nor (_17664_, _17663_, _17662_);
  nand (_17665_, _17664_, _00671_);
  nand (_17666_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  nand (_17667_, _17345_, p0_in[5]);
  nand (_17668_, _17667_, _17666_);
  nand (_17669_, _17668_, _00531_);
  nand (_17670_, _17669_, _17665_);
  nand (_17671_, _17670_, _02437_);
  nand (_17672_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nand (_17673_, _17345_, p0_in[7]);
  nand (_17674_, _17673_, _17672_);
  nand (_17675_, _17674_, _00531_);
  nor (_17676_, _17345_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  nor (_17677_, _17344_, p0_in[3]);
  nor (_17678_, _17677_, _17676_);
  nand (_17679_, _17678_, _00671_);
  nand (_17680_, _17679_, _17675_);
  nand (_17682_, _17680_, _00052_);
  nand (_17683_, _17682_, _17671_);
  nand (_17684_, _17683_, _00647_);
  nand (_17685_, _17345_, p0_in[4]);
  nand (_17686_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  nand (_17687_, _17686_, _17685_);
  nand (_17688_, _17687_, _00531_);
  nand (_17689_, _17345_, p0_in[0]);
  nand (_17690_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  nand (_17691_, _17690_, _17689_);
  nand (_17692_, _17691_, _00671_);
  nand (_17693_, _17692_, _17688_);
  nand (_17694_, _17693_, _02437_);
  nand (_17695_, _17345_, p0_in[2]);
  nand (_17696_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  nand (_17697_, _17696_, _17695_);
  nand (_17698_, _17697_, _00671_);
  nand (_17699_, _17345_, p0_in[6]);
  nand (_17700_, _17344_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  nand (_17701_, _17700_, _17699_);
  nand (_17702_, _17701_, _00531_);
  nand (_17703_, _17702_, _17698_);
  nand (_17704_, _17703_, _00052_);
  nand (_17705_, _17704_, _17694_);
  nand (_17706_, _17705_, _00634_);
  nand (_17707_, _17706_, _17684_);
  nand (_17708_, _17707_, _17477_);
  nand (_17709_, _05215_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nor (_17710_, _17280_, _10825_);
  nor (_17711_, _17710_, _00531_);
  nand (_17712_, _17711_, _17709_);
  nand (_17713_, _05215_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  not (_17714_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor (_17715_, _17280_, _17714_);
  nor (_17716_, _17715_, _00671_);
  nand (_17717_, _17716_, _17713_);
  nand (_17718_, _17717_, _17712_);
  nor (_17719_, _00671_, _10891_);
  nor (_17720_, _00531_, _10840_);
  nor (_17721_, _17720_, _17719_);
  nor (_17722_, _17721_, _17405_);
  nor (_17723_, _00531_, _10811_);
  nor (_17724_, _00671_, _10855_);
  nor (_17725_, _17724_, _17723_);
  nor (_17726_, _17725_, _17291_);
  nor (_17727_, _17726_, _17722_);
  nand (_17728_, _17727_, _17718_);
  nand (_17729_, _17728_, _17482_);
  nand (_17730_, _17729_, _17708_);
  nor (_17731_, _17730_, _17661_);
  nand (_17732_, _17731_, _17615_);
  nor (_17733_, _17732_, _17517_);
  nor (_17734_, _17420_, ABINPUT[0]);
  nor (_17735_, _17734_, _17733_);
  nor (_17736_, _17735_, _17275_);
  nor (_17737_, _00531_, ABINPUT[4]);
  nand (_17738_, _00531_, _00129_);
  nand (_17739_, _17738_, _02437_);
  nor (_17740_, _17739_, _17737_);
  nor (_17741_, _00531_, _24867_);
  nor (_17742_, _00671_, _00106_);
  nor (_17743_, _17742_, _17741_);
  nor (_17744_, _17743_, _02437_);
  nor (_17745_, _17744_, _17740_);
  nor (_17746_, _17745_, _00634_);
  nand (_17747_, _00531_, ABINPUT[7]);
  nand (_17748_, _00671_, ABINPUT[3]);
  nand (_17749_, _17748_, _17747_);
  nand (_17750_, _17749_, _05215_);
  nand (_17751_, _00531_, ABINPUT[9]);
  nand (_17753_, _00671_, ABINPUT[5]);
  nand (_17754_, _17753_, _17751_);
  nand (_17755_, _17754_, _05303_);
  nand (_17756_, _17755_, _17750_);
  nor (_17757_, _17756_, _17746_);
  nand (_17758_, _17757_, _17275_);
  nand (_17759_, _17758_, _23493_);
  nor (_08843_, _17759_, _17736_);
  nand (_17760_, _10411_, _23493_);
  not (_17761_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand (_17762_, _05209_, _17761_);
  not (_17763_, _05209_);
  nand (_17764_, _17763_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand (_17765_, _17764_, _17762_);
  nor (_25455_[3], _17765_, _17760_);
  nor (_17766_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2]);
  nor (_17767_, _22448_, _21554_);
  nor (_25091_, _17767_, _17766_);
  nor (_17768_, _22429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  nor (_17769_, _22431_, _21586_);
  nor (_08851_, _17769_, _17768_);
  nor (_17770_, _22446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3]);
  nor (_17771_, _22448_, _21526_);
  nor (_08853_, _17771_, _17770_);
  nor (_08856_, _00175_, rst);
  nand (_17772_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0]);
  nand (_17773_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0]);
  nand (_17774_, _17773_, _17772_);
  nand (_17775_, _17774_, _01417_);
  nand (_17776_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0]);
  nand (_17778_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0]);
  nand (_17779_, _17778_, _17776_);
  nand (_17780_, _17779_, _00227_);
  nand (_17781_, _17780_, _17775_);
  nand (_17782_, _17781_, _00560_);
  nand (_17783_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0]);
  nand (_17784_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0]);
  nand (_17785_, _17784_, _17783_);
  nand (_17786_, _17785_, _01417_);
  nand (_17787_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0]);
  nand (_17788_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0]);
  nand (_17789_, _17788_, _17787_);
  nand (_17790_, _17789_, _00227_);
  nand (_17791_, _17790_, _17786_);
  nand (_17792_, _17791_, _00561_);
  nand (_17793_, _17792_, _17782_);
  nand (_17794_, _17793_, _00466_);
  nor (_17795_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0]);
  nor (_17796_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0]);
  nor (_17797_, _17796_, _17795_);
  nand (_17799_, _17797_, _01417_);
  nor (_17800_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0]);
  nor (_17801_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0]);
  nor (_17802_, _17801_, _17800_);
  nand (_17803_, _17802_, _00227_);
  nand (_17804_, _17803_, _17799_);
  nand (_17805_, _17804_, _00560_);
  nor (_17806_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0]);
  nor (_17807_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0]);
  nor (_17808_, _17807_, _17806_);
  nand (_17809_, _17808_, _01417_);
  nor (_17810_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0]);
  nor (_17811_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0]);
  nor (_17812_, _17811_, _17810_);
  nand (_17813_, _17812_, _00227_);
  nand (_17814_, _17813_, _17809_);
  nand (_17815_, _17814_, _00561_);
  nand (_17816_, _17815_, _17805_);
  nand (_17817_, _17816_, _00465_);
  nand (_17818_, _17817_, _17794_);
  nand (_17820_, _17818_, _00247_);
  nand (_17821_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0]);
  nand (_17822_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0]);
  nand (_17823_, _17822_, _17821_);
  nand (_17824_, _17823_, _01417_);
  nand (_17825_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0]);
  nand (_17826_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0]);
  nand (_17827_, _17826_, _17825_);
  nand (_17828_, _17827_, _00227_);
  nand (_17829_, _17828_, _17824_);
  nand (_17830_, _17829_, _00560_);
  nand (_17831_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0]);
  nand (_17832_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0]);
  nand (_17833_, _17832_, _17831_);
  nand (_17834_, _17833_, _01417_);
  nand (_17835_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0]);
  nand (_17836_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0]);
  nand (_17837_, _17836_, _17835_);
  nand (_17838_, _17837_, _00227_);
  nand (_17839_, _17838_, _17834_);
  nand (_17841_, _17839_, _00561_);
  nand (_17842_, _17841_, _17830_);
  nand (_17843_, _17842_, _00466_);
  nor (_17844_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0]);
  nor (_17845_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0]);
  nor (_17846_, _17845_, _17844_);
  nand (_17847_, _17846_, _00227_);
  nand (_17848_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0]);
  nand (_17849_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0]);
  nand (_17850_, _17849_, _17848_);
  nand (_17851_, _17850_, _01417_);
  nand (_17852_, _17851_, _17847_);
  nand (_17853_, _17852_, _00560_);
  nor (_17854_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0]);
  nor (_17855_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0]);
  nor (_17856_, _17855_, _17854_);
  nand (_17857_, _17856_, _00227_);
  nand (_17858_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0]);
  nand (_17859_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0]);
  nand (_17860_, _17859_, _17858_);
  nand (_17861_, _17860_, _01417_);
  nand (_17862_, _17861_, _17857_);
  nand (_17863_, _17862_, _00561_);
  nand (_17864_, _17863_, _17853_);
  nand (_17865_, _17864_, _00465_);
  nand (_17866_, _17865_, _17843_);
  nand (_17867_, _17866_, _00248_);
  nand (_17868_, _17867_, _17820_);
  nand (_17869_, _17868_, _00320_);
  nand (_17870_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0]);
  nand (_17872_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0]);
  nand (_17873_, _17872_, _17870_);
  nand (_17874_, _17873_, _01417_);
  nand (_17875_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0]);
  nand (_17876_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0]);
  nand (_17877_, _17876_, _17875_);
  nand (_17878_, _17877_, _00227_);
  nand (_17879_, _17878_, _17874_);
  nand (_17880_, _17879_, _00560_);
  nand (_17881_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0]);
  nand (_17882_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0]);
  nand (_17883_, _17882_, _17881_);
  nand (_17884_, _17883_, _01417_);
  nand (_17885_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0]);
  nand (_17886_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0]);
  nand (_17887_, _17886_, _17885_);
  nand (_17888_, _17887_, _00227_);
  nand (_17889_, _17888_, _17884_);
  nand (_17890_, _17889_, _00561_);
  nand (_17891_, _17890_, _17880_);
  nand (_17893_, _17891_, _00466_);
  nor (_17894_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0]);
  nor (_17895_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0]);
  nor (_17896_, _17895_, _17894_);
  nand (_17897_, _17896_, _00227_);
  nand (_17898_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0]);
  nand (_17899_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0]);
  nand (_17900_, _17899_, _17898_);
  nand (_17901_, _17900_, _01417_);
  nand (_17902_, _17901_, _17897_);
  nand (_17903_, _17902_, _00560_);
  nor (_17904_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0]);
  nor (_17905_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0]);
  nor (_17906_, _17905_, _17904_);
  nand (_17907_, _17906_, _00227_);
  nand (_17908_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0]);
  nand (_17909_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0]);
  nand (_17910_, _17909_, _17908_);
  nand (_17911_, _17910_, _01417_);
  nand (_17912_, _17911_, _17907_);
  nand (_17913_, _17912_, _00561_);
  nand (_17914_, _17913_, _17903_);
  nand (_17915_, _17914_, _00465_);
  nand (_17916_, _17915_, _17893_);
  nand (_17917_, _17916_, _00248_);
  nand (_17918_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0]);
  nand (_17919_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0]);
  nand (_17920_, _17919_, _17918_);
  nand (_17921_, _17920_, _01417_);
  nand (_17922_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0]);
  nand (_17923_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0]);
  nand (_17924_, _17923_, _17922_);
  nand (_17925_, _17924_, _00227_);
  nand (_17926_, _17925_, _17921_);
  nand (_17927_, _17926_, _00560_);
  nand (_17928_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0]);
  nand (_17929_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0]);
  nand (_17930_, _17929_, _17928_);
  nand (_17931_, _17930_, _01417_);
  nand (_17932_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0]);
  nand (_17933_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0]);
  nand (_17934_, _17933_, _17932_);
  nand (_17935_, _17934_, _00227_);
  nand (_17936_, _17935_, _17931_);
  nand (_17937_, _17936_, _00561_);
  nand (_17938_, _17937_, _17927_);
  nand (_17939_, _17938_, _00466_);
  nor (_17940_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0]);
  nor (_17941_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0]);
  nor (_17942_, _17941_, _17940_);
  nand (_17943_, _17942_, _01417_);
  nor (_17944_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0]);
  nor (_17945_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0]);
  nor (_17946_, _17945_, _17944_);
  nand (_17947_, _17946_, _00227_);
  nand (_17948_, _17947_, _17943_);
  nand (_17949_, _17948_, _00560_);
  nor (_17950_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0]);
  nor (_17951_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0]);
  nor (_17952_, _17951_, _17950_);
  nand (_17953_, _17952_, _01417_);
  nor (_17954_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0]);
  nor (_17955_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0]);
  nor (_17956_, _17955_, _17954_);
  nand (_17957_, _17956_, _00227_);
  nand (_17958_, _17957_, _17953_);
  nand (_17959_, _17958_, _00561_);
  nand (_17960_, _17959_, _17949_);
  nand (_17961_, _17960_, _00465_);
  nand (_17962_, _17961_, _17939_);
  nand (_17963_, _17962_, _00247_);
  nand (_17964_, _17963_, _17917_);
  nand (_17965_, _17964_, _00319_);
  nand (_17966_, _17965_, _17869_);
  nor (_17967_, _17966_, _00386_);
  nand (_17968_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0]);
  nand (_17969_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0]);
  nand (_17970_, _17969_, _17968_);
  nand (_17971_, _17970_, _01417_);
  nand (_17972_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0]);
  nand (_17973_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0]);
  nand (_17974_, _17973_, _17972_);
  nand (_17975_, _17974_, _00227_);
  nand (_17976_, _17975_, _17971_);
  nand (_17977_, _17976_, _00560_);
  nand (_17978_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0]);
  nand (_17979_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0]);
  nand (_17980_, _17979_, _17978_);
  nand (_17981_, _17980_, _01417_);
  nand (_17982_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0]);
  nand (_17984_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0]);
  nand (_17985_, _17984_, _17982_);
  nand (_17986_, _17985_, _00227_);
  nand (_17987_, _17986_, _17981_);
  nand (_17988_, _17987_, _00561_);
  nand (_17989_, _17988_, _17977_);
  nand (_17990_, _17989_, _00466_);
  nor (_17991_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0]);
  nor (_17992_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0]);
  nor (_17993_, _17992_, _17991_);
  nand (_17994_, _17993_, _00227_);
  nand (_17995_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0]);
  nand (_17996_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0]);
  nand (_17997_, _17996_, _17995_);
  nand (_17998_, _17997_, _01417_);
  nand (_17999_, _17998_, _17994_);
  nand (_18000_, _17999_, _00560_);
  nor (_18001_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0]);
  nor (_18002_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0]);
  nor (_18003_, _18002_, _18001_);
  nand (_18005_, _18003_, _00227_);
  nand (_18006_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0]);
  nand (_18007_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0]);
  nand (_18008_, _18007_, _18006_);
  nand (_18009_, _18008_, _01417_);
  nand (_18010_, _18009_, _18005_);
  nand (_18011_, _18010_, _00561_);
  nand (_18012_, _18011_, _18000_);
  nand (_18013_, _18012_, _00465_);
  nand (_18014_, _18013_, _17990_);
  nand (_18015_, _18014_, _00248_);
  nand (_18016_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0]);
  nand (_18017_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0]);
  nand (_18018_, _18017_, _18016_);
  nand (_18019_, _18018_, _01417_);
  nand (_18020_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0]);
  nand (_18021_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0]);
  nand (_18022_, _18021_, _18020_);
  nand (_18023_, _18022_, _00227_);
  nand (_18024_, _18023_, _18019_);
  nand (_18026_, _18024_, _00560_);
  nand (_18027_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0]);
  nand (_18028_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0]);
  nand (_18029_, _18028_, _18027_);
  nand (_18030_, _18029_, _01417_);
  nand (_18031_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0]);
  nand (_18032_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0]);
  nand (_18033_, _18032_, _18031_);
  nand (_18034_, _18033_, _00227_);
  nand (_18035_, _18034_, _18030_);
  nand (_18036_, _18035_, _00561_);
  nand (_18037_, _18036_, _18026_);
  nand (_18038_, _18037_, _00466_);
  nor (_18039_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0]);
  nor (_18040_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0]);
  nor (_18041_, _18040_, _18039_);
  nand (_18042_, _18041_, _01417_);
  nor (_18043_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0]);
  nor (_18044_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0]);
  nor (_18045_, _18044_, _18043_);
  nand (_18047_, _18045_, _00227_);
  nand (_18048_, _18047_, _18042_);
  nand (_18049_, _18048_, _00560_);
  nor (_18050_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0]);
  nor (_18051_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0]);
  nor (_18052_, _18051_, _18050_);
  nand (_18053_, _18052_, _01417_);
  nor (_18054_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0]);
  nor (_18055_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0]);
  nor (_18056_, _18055_, _18054_);
  nand (_18057_, _18056_, _00227_);
  nand (_18058_, _18057_, _18053_);
  nand (_18059_, _18058_, _00561_);
  nand (_18060_, _18059_, _18049_);
  nand (_18061_, _18060_, _00465_);
  nand (_18062_, _18061_, _18038_);
  nand (_18063_, _18062_, _00247_);
  nand (_18064_, _18063_, _18015_);
  nand (_18065_, _18064_, _00320_);
  nor (_18066_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0]);
  nor (_18068_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0]);
  nor (_18069_, _18068_, _18066_);
  nand (_18070_, _18069_, _01417_);
  nor (_18071_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0]);
  nor (_18072_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0]);
  nor (_18073_, _18072_, _18071_);
  nand (_18074_, _18073_, _00227_);
  nand (_18075_, _18074_, _18070_);
  nand (_18076_, _18075_, _00561_);
  nor (_18077_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0]);
  nor (_18079_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0]);
  nor (_18080_, _18079_, _18077_);
  nand (_18081_, _18080_, _01417_);
  nor (_18082_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0]);
  nor (_18083_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0]);
  nor (_18084_, _18083_, _18082_);
  nand (_18085_, _18084_, _00227_);
  nand (_18086_, _18085_, _18081_);
  nand (_18087_, _18086_, _00560_);
  nand (_18088_, _18087_, _18076_);
  nand (_18090_, _18088_, _00465_);
  nand (_18091_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0]);
  nand (_18092_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0]);
  nand (_18093_, _18092_, _18091_);
  nand (_18094_, _18093_, _01417_);
  nand (_18095_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0]);
  nand (_18096_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0]);
  nand (_18097_, _18096_, _18095_);
  nand (_18098_, _18097_, _00227_);
  nand (_18099_, _18098_, _18094_);
  nand (_18100_, _18099_, _00561_);
  nand (_18101_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0]);
  nand (_18102_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0]);
  nand (_18103_, _18102_, _18101_);
  nand (_18104_, _18103_, _01417_);
  nand (_18105_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0]);
  nand (_18106_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0]);
  nand (_18107_, _18106_, _18105_);
  nand (_18108_, _18107_, _00227_);
  nand (_18109_, _18108_, _18104_);
  nand (_18111_, _18109_, _00560_);
  nand (_18112_, _18111_, _18100_);
  nand (_18113_, _18112_, _00466_);
  nand (_18114_, _18113_, _18090_);
  nand (_18115_, _18114_, _00247_);
  nor (_18116_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0]);
  nor (_18117_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0]);
  nor (_18118_, _18117_, _18116_);
  nand (_18119_, _18118_, _00227_);
  nand (_18120_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0]);
  nand (_18121_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0]);
  nand (_18122_, _18121_, _18120_);
  nand (_18123_, _18122_, _01417_);
  nand (_18124_, _18123_, _18119_);
  nand (_18125_, _18124_, _00561_);
  nor (_18126_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0]);
  nor (_18127_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0]);
  nor (_18128_, _18127_, _18126_);
  nand (_18129_, _18128_, _00227_);
  nand (_18130_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0]);
  nand (_18132_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0]);
  nand (_18133_, _18132_, _18130_);
  nand (_18134_, _18133_, _01417_);
  nand (_18135_, _18134_, _18129_);
  nand (_18136_, _18135_, _00560_);
  nand (_18137_, _18136_, _18125_);
  nand (_18138_, _18137_, _00465_);
  nand (_18139_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0]);
  nand (_18140_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0]);
  nand (_18141_, _18140_, _18139_);
  nand (_18142_, _18141_, _01417_);
  nand (_18143_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0]);
  nand (_18144_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0]);
  nand (_18145_, _18144_, _18143_);
  nand (_18146_, _18145_, _00227_);
  nand (_18147_, _18146_, _18142_);
  nand (_18148_, _18147_, _00561_);
  nand (_18149_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0]);
  nand (_18150_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0]);
  nand (_18151_, _18150_, _18149_);
  nand (_18153_, _18151_, _01417_);
  nand (_18154_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0]);
  nand (_18155_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0]);
  nand (_18156_, _18155_, _18154_);
  nand (_18157_, _18156_, _00227_);
  nand (_18158_, _18157_, _18153_);
  nand (_18159_, _18158_, _00560_);
  nand (_18160_, _18159_, _18148_);
  nand (_18161_, _18160_, _00466_);
  nand (_18162_, _18161_, _18138_);
  nand (_18163_, _18162_, _00248_);
  nand (_18164_, _18163_, _18115_);
  nand (_18165_, _18164_, _00319_);
  nand (_18166_, _18165_, _18065_);
  nor (_18167_, _18166_, _01629_);
  nor (_18168_, _18167_, _17967_);
  nor (_18169_, _18168_, _00156_);
  nand (_18170_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0]);
  nand (_18171_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0]);
  nand (_18172_, _18171_, _18170_);
  nand (_18173_, _18172_, _00227_);
  nand (_18174_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0]);
  nand (_18175_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0]);
  nand (_18176_, _18175_, _18174_);
  nand (_18177_, _18176_, _01417_);
  nand (_18178_, _18177_, _18173_);
  nand (_18179_, _18178_, _00560_);
  nand (_18180_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0]);
  nand (_18181_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0]);
  nand (_18182_, _18181_, _18180_);
  nand (_18184_, _18182_, _00227_);
  nand (_18185_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0]);
  nand (_18186_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0]);
  nand (_18187_, _18186_, _18185_);
  nand (_18188_, _18187_, _01417_);
  nand (_18189_, _18188_, _18184_);
  nand (_18190_, _18189_, _00561_);
  nand (_18191_, _18190_, _18179_);
  nand (_18192_, _18191_, _00466_);
  nand (_18193_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0]);
  nand (_18194_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0]);
  nand (_18195_, _18194_, _18193_);
  nand (_18196_, _18195_, _01417_);
  nor (_18197_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0]);
  nor (_18198_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0]);
  nor (_18199_, _18198_, _18197_);
  nand (_18200_, _18199_, _00227_);
  nand (_18201_, _18200_, _18196_);
  nand (_18202_, _18201_, _00560_);
  nand (_18203_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0]);
  nand (_18204_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0]);
  nand (_18205_, _18204_, _18203_);
  nand (_18206_, _18205_, _01417_);
  nor (_18207_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0]);
  nor (_18208_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0]);
  nor (_18209_, _18208_, _18207_);
  nand (_18210_, _18209_, _00227_);
  nand (_18211_, _18210_, _18206_);
  nand (_18212_, _18211_, _00561_);
  nand (_18213_, _18212_, _18202_);
  nand (_18214_, _18213_, _00465_);
  nand (_18215_, _18214_, _18192_);
  nand (_18216_, _18215_, _00248_);
  nand (_18217_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0]);
  nand (_18218_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0]);
  nand (_18219_, _18218_, _18217_);
  nand (_18220_, _18219_, _01417_);
  nand (_18221_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0]);
  nand (_18222_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0]);
  nand (_18223_, _18222_, _18221_);
  nand (_18224_, _18223_, _00227_);
  nand (_18225_, _18224_, _18220_);
  nand (_18226_, _18225_, _00560_);
  nand (_18227_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0]);
  nand (_18228_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0]);
  nand (_18229_, _18228_, _18227_);
  nand (_18230_, _18229_, _01417_);
  nand (_18231_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0]);
  nand (_18232_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0]);
  nand (_18233_, _18232_, _18231_);
  nand (_18234_, _18233_, _00227_);
  nand (_18235_, _18234_, _18230_);
  nand (_18236_, _18235_, _00561_);
  nand (_18237_, _18236_, _18226_);
  nand (_18238_, _18237_, _00466_);
  nor (_18239_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0]);
  nor (_18240_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0]);
  nor (_18241_, _18240_, _18239_);
  nand (_18242_, _18241_, _01417_);
  nor (_18243_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0]);
  nor (_18244_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0]);
  nor (_18245_, _18244_, _18243_);
  nand (_18246_, _18245_, _00227_);
  nand (_18247_, _18246_, _18242_);
  nand (_18248_, _18247_, _00560_);
  nor (_18249_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0]);
  nor (_18250_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0]);
  nor (_18251_, _18250_, _18249_);
  nor (_18252_, _18251_, _00227_);
  nor (_18253_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0]);
  nor (_18254_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0]);
  nor (_18255_, _18254_, _18253_);
  nor (_18256_, _18255_, _01417_);
  nor (_18257_, _18256_, _18252_);
  nand (_18258_, _18257_, _00561_);
  nand (_18259_, _18258_, _18248_);
  nand (_18260_, _18259_, _00465_);
  nand (_18261_, _18260_, _18238_);
  nand (_18262_, _18261_, _00247_);
  nand (_18263_, _18262_, _18216_);
  nand (_18265_, _18263_, _00320_);
  nand (_18266_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  nand (_18267_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0]);
  nand (_18268_, _18267_, _18266_);
  nand (_18269_, _18268_, _01417_);
  nand (_18270_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0]);
  nand (_18271_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0]);
  nand (_18272_, _18271_, _18270_);
  nand (_18273_, _18272_, _00227_);
  nand (_18274_, _18273_, _18269_);
  nand (_18275_, _18274_, _00560_);
  nand (_18276_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0]);
  nand (_18277_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0]);
  nand (_18278_, _18277_, _18276_);
  nand (_18279_, _18278_, _01417_);
  nand (_18280_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0]);
  nand (_18281_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0]);
  nand (_18282_, _18281_, _18280_);
  nand (_18283_, _18282_, _00227_);
  nand (_18284_, _18283_, _18279_);
  nand (_18285_, _18284_, _00561_);
  nand (_18286_, _18285_, _18275_);
  nand (_18287_, _18286_, _00466_);
  nor (_18288_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0]);
  nor (_18289_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0]);
  nor (_18290_, _18289_, _18288_);
  nand (_18291_, _18290_, _01417_);
  nor (_18292_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0]);
  nor (_18293_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  nor (_18294_, _18293_, _18292_);
  nand (_18295_, _18294_, _00227_);
  nand (_18296_, _18295_, _18291_);
  nand (_18297_, _18296_, _00560_);
  nor (_18298_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0]);
  nor (_18299_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0]);
  nor (_18300_, _18299_, _18298_);
  nand (_18301_, _18300_, _01417_);
  nor (_18302_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0]);
  nor (_18303_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0]);
  nor (_18304_, _18303_, _18302_);
  nand (_18306_, _18304_, _00227_);
  nand (_18307_, _18306_, _18301_);
  nand (_18308_, _18307_, _00561_);
  nand (_18309_, _18308_, _18297_);
  nand (_18310_, _18309_, _00465_);
  nand (_18311_, _18310_, _18287_);
  nand (_18312_, _18311_, _00248_);
  nand (_18313_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  nand (_18314_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0]);
  nand (_18315_, _18314_, _18313_);
  nand (_18316_, _18315_, _01417_);
  nand (_18317_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0]);
  nand (_18318_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0]);
  nand (_18319_, _18318_, _18317_);
  nand (_18320_, _18319_, _00227_);
  nand (_18321_, _18320_, _18316_);
  nand (_18322_, _18321_, _00560_);
  nand (_18323_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0]);
  nand (_18324_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0]);
  nand (_18325_, _18324_, _18323_);
  nand (_18327_, _18325_, _01417_);
  nand (_18328_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0]);
  nand (_18329_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0]);
  nand (_18330_, _18329_, _18328_);
  nand (_18331_, _18330_, _00227_);
  nand (_18332_, _18331_, _18327_);
  nand (_18333_, _18332_, _00561_);
  nand (_18334_, _18333_, _18322_);
  nand (_18335_, _18334_, _00466_);
  nor (_18336_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0]);
  nor (_18337_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0]);
  nor (_18338_, _18337_, _18336_);
  nand (_18339_, _18338_, _01417_);
  nor (_18340_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0]);
  nor (_18341_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0]);
  nor (_18342_, _18341_, _18340_);
  nand (_18343_, _18342_, _00227_);
  nand (_18344_, _18343_, _18339_);
  nand (_18345_, _18344_, _00560_);
  nor (_18346_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0]);
  nor (_18348_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0]);
  nor (_18349_, _18348_, _18346_);
  nand (_18350_, _18349_, _01417_);
  nor (_18351_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0]);
  nor (_18352_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0]);
  nor (_18353_, _18352_, _18351_);
  nand (_18354_, _18353_, _00227_);
  nand (_18355_, _18354_, _18350_);
  nand (_18356_, _18355_, _00561_);
  nand (_18357_, _18356_, _18345_);
  nand (_18358_, _18357_, _00465_);
  nand (_18359_, _18358_, _18335_);
  nand (_18360_, _18359_, _00247_);
  nand (_18361_, _18360_, _18312_);
  nand (_18362_, _18361_, _00319_);
  nand (_18363_, _18362_, _18265_);
  nor (_18364_, _18363_, _00386_);
  nand (_18365_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0]);
  nand (_18366_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0]);
  nand (_18367_, _18366_, _18365_);
  nand (_18369_, _18367_, _01417_);
  nand (_18370_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0]);
  nand (_18371_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0]);
  nand (_18372_, _18371_, _18370_);
  nand (_18373_, _18372_, _00227_);
  nand (_18374_, _18373_, _18369_);
  nand (_18375_, _18374_, _00560_);
  nand (_18376_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0]);
  nand (_18377_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0]);
  nand (_18378_, _18377_, _18376_);
  nand (_18379_, _18378_, _01417_);
  nand (_18380_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0]);
  nand (_18381_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0]);
  nand (_18382_, _18381_, _18380_);
  nand (_18383_, _18382_, _00227_);
  nand (_18384_, _18383_, _18379_);
  nand (_18385_, _18384_, _00561_);
  nand (_18386_, _18385_, _18375_);
  nand (_18387_, _18386_, _00466_);
  nor (_18388_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  nor (_18389_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  nor (_18390_, _18389_, _18388_);
  nand (_18391_, _18390_, _00227_);
  nand (_18392_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0]);
  nand (_18393_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0]);
  nand (_18394_, _18393_, _18392_);
  nand (_18395_, _18394_, _01417_);
  nand (_18396_, _18395_, _18391_);
  nand (_18397_, _18396_, _00560_);
  nor (_18398_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0]);
  nor (_18399_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0]);
  nor (_18400_, _18399_, _18398_);
  nand (_18401_, _18400_, _00227_);
  nand (_18402_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0]);
  nand (_18403_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0]);
  nand (_18404_, _18403_, _18402_);
  nand (_18405_, _18404_, _01417_);
  nand (_18406_, _18405_, _18401_);
  nand (_18407_, _18406_, _00561_);
  nand (_18408_, _18407_, _18397_);
  nand (_18410_, _18408_, _00465_);
  nand (_18411_, _18410_, _18387_);
  nand (_18412_, _18411_, _00248_);
  nand (_18413_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0]);
  nand (_18414_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0]);
  nand (_18415_, _18414_, _18413_);
  nand (_18416_, _18415_, _01417_);
  nand (_18417_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0]);
  nand (_18418_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0]);
  nand (_18419_, _18418_, _18417_);
  nand (_18420_, _18419_, _00227_);
  nand (_18421_, _18420_, _18416_);
  nand (_18422_, _18421_, _00560_);
  nand (_18423_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0]);
  nand (_18424_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  nand (_18425_, _18424_, _18423_);
  nand (_18426_, _18425_, _01417_);
  nand (_18427_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0]);
  nand (_18428_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0]);
  nand (_18429_, _18428_, _18427_);
  nand (_18431_, _18429_, _00227_);
  nand (_18432_, _18431_, _18426_);
  nand (_18433_, _18432_, _00561_);
  nand (_18434_, _18433_, _18422_);
  nand (_18435_, _18434_, _00466_);
  nor (_18436_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0]);
  nor (_18437_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0]);
  nor (_18438_, _18437_, _18436_);
  nand (_18439_, _18438_, _01417_);
  nor (_18440_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0]);
  nor (_18441_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0]);
  nor (_18442_, _18441_, _18440_);
  nand (_18443_, _18442_, _00227_);
  nand (_18444_, _18443_, _18439_);
  nand (_18445_, _18444_, _00560_);
  nor (_18446_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0]);
  nor (_18447_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0]);
  nor (_18448_, _18447_, _18446_);
  nand (_18449_, _18448_, _01417_);
  nor (_18450_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0]);
  nor (_18451_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0]);
  nor (_18452_, _18451_, _18450_);
  nand (_18453_, _18452_, _00227_);
  nand (_18454_, _18453_, _18449_);
  nand (_18455_, _18454_, _00561_);
  nand (_18456_, _18455_, _18445_);
  nand (_18457_, _18456_, _00465_);
  nand (_18458_, _18457_, _18435_);
  nand (_18459_, _18458_, _00247_);
  nand (_18460_, _18459_, _18412_);
  nand (_18461_, _18460_, _00320_);
  nor (_18462_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0]);
  nor (_18463_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0]);
  nor (_18464_, _18463_, _18462_);
  nand (_18465_, _18464_, _01417_);
  nor (_18466_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0]);
  nor (_18467_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0]);
  nor (_18468_, _18467_, _18466_);
  nand (_18469_, _18468_, _00227_);
  nand (_18470_, _18469_, _18465_);
  nand (_18472_, _18470_, _00561_);
  nor (_18473_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0]);
  nor (_18474_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0]);
  nor (_18475_, _18474_, _18473_);
  nand (_18476_, _18475_, _01417_);
  nor (_18477_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0]);
  nor (_18478_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0]);
  nor (_18479_, _18478_, _18477_);
  nand (_18480_, _18479_, _00227_);
  nand (_18481_, _18480_, _18476_);
  nand (_18482_, _18481_, _00560_);
  nand (_18483_, _18482_, _18472_);
  nand (_18484_, _18483_, _00465_);
  nand (_18485_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0]);
  nand (_18486_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0]);
  nand (_18487_, _18486_, _18485_);
  nand (_18488_, _18487_, _01417_);
  nand (_18489_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0]);
  nand (_18490_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0]);
  nand (_18491_, _18490_, _18489_);
  nand (_18492_, _18491_, _00227_);
  nand (_18493_, _18492_, _18488_);
  nand (_18494_, _18493_, _00561_);
  nand (_18495_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0]);
  nand (_18496_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0]);
  nand (_18497_, _18496_, _18495_);
  nand (_18498_, _18497_, _01417_);
  nand (_18499_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0]);
  nand (_18500_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0]);
  nand (_18501_, _18500_, _18499_);
  nand (_18502_, _18501_, _00227_);
  nand (_18503_, _18502_, _18498_);
  nand (_18504_, _18503_, _00560_);
  nand (_18505_, _18504_, _18494_);
  nand (_18506_, _18505_, _00466_);
  nand (_18507_, _18506_, _18484_);
  nand (_18508_, _18507_, _00247_);
  nor (_18509_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0]);
  nor (_18510_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0]);
  nor (_18511_, _18510_, _18509_);
  nand (_18512_, _18511_, _00227_);
  nand (_18513_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0]);
  nand (_18514_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0]);
  nand (_18515_, _18514_, _18513_);
  nand (_18516_, _18515_, _01417_);
  nand (_18517_, _18516_, _18512_);
  nand (_18518_, _18517_, _00561_);
  nor (_18519_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0]);
  nor (_18520_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0]);
  nor (_18521_, _18520_, _18519_);
  nand (_18523_, _18521_, _00227_);
  nand (_18524_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0]);
  nand (_18525_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0]);
  nand (_18526_, _18525_, _18524_);
  nand (_18527_, _18526_, _01417_);
  nand (_18528_, _18527_, _18523_);
  nand (_18529_, _18528_, _00560_);
  nand (_18530_, _18529_, _18518_);
  nand (_18531_, _18530_, _00465_);
  nand (_18532_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0]);
  nand (_18533_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0]);
  nand (_18534_, _18533_, _18532_);
  nand (_18535_, _18534_, _01417_);
  nand (_18536_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0]);
  nand (_18537_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0]);
  nand (_18538_, _18537_, _18536_);
  nand (_18539_, _18538_, _00227_);
  nand (_18540_, _18539_, _18535_);
  nand (_18541_, _18540_, _00561_);
  nand (_18542_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0]);
  nand (_18543_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0]);
  nand (_18544_, _18543_, _18542_);
  nand (_18545_, _18544_, _01417_);
  nand (_18546_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0]);
  nand (_18547_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0]);
  nand (_18548_, _18547_, _18546_);
  nand (_18549_, _18548_, _00227_);
  nand (_18550_, _18549_, _18545_);
  nand (_18551_, _18550_, _00560_);
  nand (_18552_, _18551_, _18541_);
  nand (_18553_, _18552_, _00466_);
  nand (_18554_, _18553_, _18531_);
  nand (_18555_, _18554_, _00248_);
  nand (_18556_, _18555_, _18508_);
  nand (_18557_, _18556_, _00319_);
  nand (_18558_, _18557_, _18461_);
  nor (_18559_, _18558_, _01629_);
  nor (_18560_, _18559_, _18364_);
  nor (_18561_, _18560_, _00556_);
  nor (_18562_, _18561_, _18169_);
  nor (_18563_, _18562_, _01416_);
  not (_18564_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  nand (_18565_, _01416_, _18564_);
  nand (_18566_, _18565_, _23493_);
  nor (_08862_, _18566_, _18563_);
  nor (_18567_, _21904_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3]);
  nor (_18568_, _21906_, _21526_);
  nor (_08866_, _18568_, _18567_);
  nor (_18569_, _21752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1]);
  nor (_18570_, _21754_, _21474_);
  nor (_08868_, _18570_, _18569_);
  nor (_18571_, _01383_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1]);
  nor (_18572_, _01385_, _21474_);
  nor (_08872_, _18572_, _18571_);
  nor (_08875_, _00301_, rst);
  nand (_18573_, _02393_, _00029_);
  nand (_18574_, _18573_, _23493_);
  not (_18575_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_18576_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _14884_);
  nand (_18577_, _18576_, _01059_);
  nand (_18578_, _18577_, _02485_);
  nand (_18579_, _18578_, _18575_);
  nor (_18580_, _18579_, _02395_);
  nand (_18581_, _24858_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_18582_, _18581_, _10800_);
  nor (_18583_, _18582_, _02390_);
  nor (_18584_, _18583_, _18580_);
  nor (_18585_, _18584_, _02393_);
  nor (_08877_, _18585_, _18574_);
  nor (_18586_, _22922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6]);
  nor (_18588_, _22924_, _21504_);
  nor (_25090_, _18588_, _18586_);
  nor (_18589_, _22429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2]);
  nor (_18590_, _22431_, _21554_);
  nor (_25103_, _18590_, _18589_);
  nor (_18591_, _22450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5]);
  nor (_18592_, _22452_, _21451_);
  nor (_08886_, _18592_, _18591_);
  not (_18593_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nor (_18594_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _18593_);
  nor (_18595_, _01079_, _02448_);
  nor (_18596_, _01066_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  nor (_18597_, _18596_, _14655_);
  nand (_18598_, _01077_, _01058_);
  nor (_18599_, _18598_, _18593_);
  nor (_18600_, _18599_, _18597_);
  nor (_18601_, _18600_, _01071_);
  nor (_18602_, _18601_, _18595_);
  nor (_18603_, _18602_, _01052_);
  nor (_18604_, _18603_, _18594_);
  nor (_08889_, _18604_, rst);
  nor (_18606_, _00880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2]);
  nor (_18607_, _00882_, _21554_);
  nor (_08897_, _18607_, _18606_);
  nor (_18608_, _22408_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0]);
  nor (_18609_, _22410_, _21586_);
  nor (_08910_, _18609_, _18608_);
  nor (_18610_, _23545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5]);
  nor (_18611_, _23547_, _21451_);
  nor (_08914_, _18611_, _18610_);
  nor (_18612_, _23545_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1]);
  nor (_18613_, _23547_, _21474_);
  nor (_08919_, _18613_, _18612_);
  nor (_18614_, _22922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0]);
  nor (_18615_, _22924_, _21586_);
  nor (_08922_, _18615_, _18614_);
  nor (_18616_, _00989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  nor (_18617_, _18616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_18618_, _18617_, _00919_);
  not (_18619_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_18620_, _05052_, _18619_);
  nor (_18621_, _18620_, _05056_);
  nand (_18622_, _18621_, _00930_);
  nand (_18623_, _18622_, _18618_);
  nor (_18624_, _18623_, _00928_);
  nor (_18625_, _00929_, _00114_);
  nor (_18626_, _18625_, _18624_);
  nor (_08928_, _18626_, rst);
  nor (_18627_, _01010_, _00919_);
  nor (_18628_, _18627_, _14692_);
  nand (_18630_, _05018_, _00930_);
  nand (_18631_, _18630_, _00929_);
  nor (_18632_, _18631_, _18628_);
  nand (_18633_, _00928_, _00129_);
  nand (_18634_, _18633_, _23493_);
  nor (_08930_, _18634_, _18632_);
  nor (_18635_, _22450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7]);
  nor (_18636_, _22452_, _21626_);
  nor (_08935_, _18636_, _18635_);
  nor (_18637_, _22450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6]);
  nor (_18638_, _22452_, _21504_);
  nor (_08938_, _18638_, _18637_);
  nor (_18639_, _14304_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2]);
  nor (_18640_, _14306_, _21554_);
  nor (_25284_, _18640_, _18639_);
  nor (_18641_, _21733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5]);
  nor (_18642_, _21735_, _21451_);
  nor (_25244_, _18642_, _18641_);
  nor (_18643_, _12387_, _01330_);
  nor (_18644_, _18643_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  nor (_25036_[5], _18644_, rst);
  nor (_18646_, _05453_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3]);
  nor (_18647_, _05455_, _21526_);
  nor (_08947_, _18647_, _18646_);
  nor (_18648_, _14242_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand (_18649_, _14242_, _14250_);
  nand (_18650_, _18649_, _23493_);
  nor (_08950_, _18650_, _18648_);
  nor (_08952_, _12030_, rst);
  nor (_18651_, _22429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3]);
  nor (_18652_, _22431_, _21526_);
  nor (_08954_, _18652_, _18651_);
  nor (_08956_, _00380_, rst);
  nor (_18653_, _22922_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7]);
  nor (_18654_, _22924_, _21626_);
  nor (_08958_, _18654_, _18653_);
  nand (_18655_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4]);
  nand (_18656_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4]);
  nand (_18657_, _18656_, _18655_);
  nand (_18658_, _18657_, _01417_);
  nand (_18660_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4]);
  nand (_18661_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4]);
  nand (_18662_, _18661_, _18660_);
  nand (_18663_, _18662_, _00227_);
  nand (_18664_, _18663_, _18658_);
  nand (_18665_, _18664_, _00560_);
  nand (_18666_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4]);
  nand (_18667_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4]);
  nand (_18668_, _18667_, _18666_);
  nand (_18669_, _18668_, _01417_);
  nand (_18670_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4]);
  nand (_18671_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4]);
  nand (_18672_, _18671_, _18670_);
  nand (_18673_, _18672_, _00227_);
  nand (_18674_, _18673_, _18669_);
  nand (_18675_, _18674_, _00561_);
  nand (_18676_, _18675_, _18665_);
  nand (_18677_, _18676_, _00466_);
  nor (_18678_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4]);
  nor (_18679_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4]);
  nor (_18680_, _18679_, _18678_);
  nand (_18681_, _18680_, _00227_);
  nand (_18682_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4]);
  nand (_18683_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4]);
  nand (_18684_, _18683_, _18682_);
  nand (_18685_, _18684_, _01417_);
  nand (_18686_, _18685_, _18681_);
  nand (_18687_, _18686_, _00560_);
  nor (_18688_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4]);
  nor (_18689_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4]);
  nor (_18691_, _18689_, _18688_);
  nand (_18692_, _18691_, _00227_);
  nand (_18693_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4]);
  nand (_18694_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4]);
  nand (_18695_, _18694_, _18693_);
  nand (_18696_, _18695_, _01417_);
  nand (_18697_, _18696_, _18692_);
  nand (_18698_, _18697_, _00561_);
  nand (_18699_, _18698_, _18687_);
  nand (_18700_, _18699_, _00465_);
  nand (_18701_, _18700_, _18677_);
  nand (_18702_, _18701_, _00248_);
  nand (_18703_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4]);
  nand (_18704_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4]);
  nand (_18705_, _18704_, _18703_);
  nand (_18706_, _18705_, _01417_);
  nand (_18707_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4]);
  nand (_18708_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4]);
  nand (_18709_, _18708_, _18707_);
  nand (_18710_, _18709_, _00227_);
  nand (_18712_, _18710_, _18706_);
  nand (_18713_, _18712_, _00560_);
  nand (_18714_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4]);
  nand (_18715_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4]);
  nand (_18716_, _18715_, _18714_);
  nand (_18717_, _18716_, _01417_);
  nand (_18718_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4]);
  nand (_18719_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4]);
  nand (_18720_, _18719_, _18718_);
  nand (_18721_, _18720_, _00227_);
  nand (_18722_, _18721_, _18717_);
  nand (_18723_, _18722_, _00561_);
  nand (_18724_, _18723_, _18713_);
  nand (_18725_, _18724_, _00466_);
  nor (_18726_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4]);
  nor (_18727_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4]);
  nor (_18728_, _18727_, _18726_);
  nand (_18729_, _18728_, _01417_);
  nor (_18730_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4]);
  nor (_18731_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4]);
  nor (_18732_, _18731_, _18730_);
  nand (_18733_, _18732_, _00227_);
  nand (_18734_, _18733_, _18729_);
  nand (_18735_, _18734_, _00560_);
  nor (_18736_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4]);
  nor (_18737_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4]);
  nor (_18738_, _18737_, _18736_);
  nand (_18739_, _18738_, _01417_);
  nor (_18740_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4]);
  nor (_18741_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4]);
  nor (_18742_, _18741_, _18740_);
  nand (_18743_, _18742_, _00227_);
  nand (_18744_, _18743_, _18739_);
  nand (_18745_, _18744_, _00561_);
  nand (_18746_, _18745_, _18735_);
  nand (_18747_, _18746_, _00465_);
  nand (_18748_, _18747_, _18725_);
  nand (_18749_, _18748_, _00247_);
  nand (_18750_, _18749_, _18702_);
  nand (_18751_, _18750_, _00319_);
  nand (_18752_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4]);
  nand (_18753_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4]);
  nand (_18754_, _18753_, _18752_);
  nand (_18755_, _18754_, _01417_);
  nand (_18756_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4]);
  nand (_18757_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4]);
  nand (_18758_, _18757_, _18756_);
  nand (_18759_, _18758_, _00227_);
  nand (_18760_, _18759_, _18755_);
  nand (_18761_, _18760_, _00560_);
  nand (_18762_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4]);
  nand (_18763_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4]);
  nand (_18764_, _18763_, _18762_);
  nand (_18765_, _18764_, _01417_);
  nand (_18766_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4]);
  nand (_18767_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4]);
  nand (_18768_, _18767_, _18766_);
  nand (_18769_, _18768_, _00227_);
  nand (_18770_, _18769_, _18765_);
  nand (_18771_, _18770_, _00561_);
  nand (_18772_, _18771_, _18761_);
  nand (_18773_, _18772_, _00466_);
  nor (_18774_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4]);
  nor (_18775_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4]);
  nor (_18776_, _18775_, _18774_);
  nand (_18777_, _18776_, _01417_);
  nor (_18778_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4]);
  nor (_18779_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4]);
  nor (_18780_, _18779_, _18778_);
  nand (_18781_, _18780_, _00227_);
  nand (_18782_, _18781_, _18777_);
  nand (_18783_, _18782_, _00560_);
  nor (_18784_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4]);
  nor (_18785_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4]);
  nor (_18786_, _18785_, _18784_);
  nand (_18787_, _18786_, _01417_);
  nor (_18788_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4]);
  nor (_18789_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4]);
  nor (_18790_, _18789_, _18788_);
  nand (_18791_, _18790_, _00227_);
  nand (_18793_, _18791_, _18787_);
  nand (_18794_, _18793_, _00561_);
  nand (_18795_, _18794_, _18783_);
  nand (_18796_, _18795_, _00465_);
  nand (_18797_, _18796_, _18773_);
  nand (_18798_, _18797_, _00247_);
  nand (_18799_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4]);
  nand (_18800_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4]);
  nand (_18801_, _18800_, _18799_);
  nand (_18802_, _18801_, _01417_);
  nand (_18803_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4]);
  nand (_18804_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4]);
  nand (_18805_, _18804_, _18803_);
  nand (_18806_, _18805_, _00227_);
  nand (_18807_, _18806_, _18802_);
  nand (_18808_, _18807_, _00560_);
  nand (_18809_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4]);
  nand (_18810_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4]);
  nand (_18811_, _18810_, _18809_);
  nand (_18812_, _18811_, _01417_);
  nand (_18813_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4]);
  nand (_18814_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4]);
  nand (_18815_, _18814_, _18813_);
  nand (_18816_, _18815_, _00227_);
  nand (_18817_, _18816_, _18812_);
  nand (_18818_, _18817_, _00561_);
  nand (_18819_, _18818_, _18808_);
  nand (_18820_, _18819_, _00466_);
  nor (_18821_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4]);
  nor (_18822_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4]);
  nor (_18823_, _18822_, _18821_);
  nand (_18824_, _18823_, _00227_);
  nand (_18825_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4]);
  nand (_18826_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4]);
  nand (_18827_, _18826_, _18825_);
  nand (_18828_, _18827_, _01417_);
  nand (_18829_, _18828_, _18824_);
  nand (_18830_, _18829_, _00560_);
  nor (_18831_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4]);
  nor (_18832_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4]);
  nor (_18834_, _18832_, _18831_);
  nand (_18835_, _18834_, _00227_);
  nand (_18836_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4]);
  nand (_18837_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4]);
  nand (_18838_, _18837_, _18836_);
  nand (_18839_, _18838_, _01417_);
  nand (_18840_, _18839_, _18835_);
  nand (_18841_, _18840_, _00561_);
  nand (_18842_, _18841_, _18830_);
  nand (_18843_, _18842_, _00465_);
  nand (_18844_, _18843_, _18820_);
  nand (_18845_, _18844_, _00248_);
  nand (_18846_, _18845_, _18798_);
  nand (_18847_, _18846_, _00320_);
  nand (_18848_, _18847_, _18751_);
  nand (_18849_, _18848_, _01629_);
  nor (_18850_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4]);
  nor (_18851_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4]);
  nor (_18852_, _18851_, _18850_);
  nand (_18853_, _18852_, _01417_);
  nor (_18855_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4]);
  nor (_18856_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4]);
  nor (_18857_, _18856_, _18855_);
  nand (_18858_, _18857_, _00227_);
  nand (_18859_, _18858_, _18853_);
  nand (_18860_, _18859_, _00561_);
  nor (_18861_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4]);
  nor (_18862_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4]);
  nor (_18863_, _18862_, _18861_);
  nand (_18864_, _18863_, _01417_);
  nor (_18865_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4]);
  nor (_18866_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4]);
  nor (_18867_, _18866_, _18865_);
  nand (_18868_, _18867_, _00227_);
  nand (_18869_, _18868_, _18864_);
  nand (_18870_, _18869_, _00560_);
  nand (_18871_, _18870_, _18860_);
  nand (_18872_, _18871_, _00465_);
  nand (_18873_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4]);
  nand (_18874_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4]);
  nand (_18875_, _18874_, _18873_);
  nand (_18876_, _18875_, _01417_);
  nand (_18877_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4]);
  nand (_18878_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4]);
  nand (_18879_, _18878_, _18877_);
  nand (_18880_, _18879_, _00227_);
  nand (_18881_, _18880_, _18876_);
  nand (_18882_, _18881_, _00561_);
  nand (_18883_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4]);
  nand (_18884_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4]);
  nand (_18885_, _18884_, _18883_);
  nand (_18886_, _18885_, _01417_);
  nand (_18887_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4]);
  nand (_18888_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4]);
  nand (_18889_, _18888_, _18887_);
  nand (_18890_, _18889_, _00227_);
  nand (_18891_, _18890_, _18886_);
  nand (_18892_, _18891_, _00560_);
  nand (_18893_, _18892_, _18882_);
  nand (_18894_, _18893_, _00466_);
  nand (_18896_, _18894_, _18872_);
  nand (_18897_, _18896_, _00247_);
  nor (_18898_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4]);
  nor (_18899_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4]);
  nor (_18900_, _18899_, _18898_);
  nand (_18901_, _18900_, _00227_);
  nand (_18902_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4]);
  nand (_18903_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4]);
  nand (_18904_, _18903_, _18902_);
  nand (_18905_, _18904_, _01417_);
  nand (_18906_, _18905_, _18901_);
  nand (_18907_, _18906_, _00561_);
  nor (_18908_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4]);
  nor (_18909_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4]);
  nor (_18910_, _18909_, _18908_);
  nand (_18911_, _18910_, _00227_);
  nand (_18912_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4]);
  nand (_18913_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4]);
  nand (_18914_, _18913_, _18912_);
  nand (_18915_, _18914_, _01417_);
  nand (_18917_, _18915_, _18911_);
  nand (_18918_, _18917_, _00560_);
  nand (_18919_, _18918_, _18907_);
  nand (_18920_, _18919_, _00465_);
  nand (_18921_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4]);
  nand (_18922_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4]);
  nand (_18923_, _18922_, _18921_);
  nand (_18924_, _18923_, _01417_);
  nand (_18925_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4]);
  nand (_18926_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4]);
  nand (_18927_, _18926_, _18925_);
  nand (_18928_, _18927_, _00227_);
  nand (_18929_, _18928_, _18924_);
  nand (_18930_, _18929_, _00561_);
  nand (_18931_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4]);
  nand (_18932_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4]);
  nand (_18933_, _18932_, _18931_);
  nand (_18934_, _18933_, _01417_);
  nand (_18935_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4]);
  nand (_18936_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4]);
  nand (_18938_, _18936_, _18935_);
  nand (_18939_, _18938_, _00227_);
  nand (_18940_, _18939_, _18934_);
  nand (_18941_, _18940_, _00560_);
  nand (_18942_, _18941_, _18930_);
  nand (_18943_, _18942_, _00466_);
  nand (_18944_, _18943_, _18920_);
  nand (_18945_, _18944_, _00248_);
  nand (_18946_, _18945_, _18897_);
  nand (_18947_, _18946_, _00319_);
  nand (_18948_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4]);
  nand (_18949_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4]);
  nand (_18950_, _18949_, _18948_);
  nand (_18951_, _18950_, _01417_);
  nand (_18952_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4]);
  nand (_18953_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4]);
  nand (_18954_, _18953_, _18952_);
  nand (_18955_, _18954_, _00227_);
  nand (_18956_, _18955_, _18951_);
  nand (_18957_, _18956_, _00560_);
  nand (_18959_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4]);
  nand (_18960_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4]);
  nand (_18961_, _18960_, _18959_);
  nand (_18962_, _18961_, _01417_);
  nand (_18963_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4]);
  nand (_18964_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4]);
  nand (_18965_, _18964_, _18963_);
  nand (_18966_, _18965_, _00227_);
  nand (_18967_, _18966_, _18962_);
  nand (_18968_, _18967_, _00561_);
  nand (_18969_, _18968_, _18957_);
  nand (_18970_, _18969_, _00466_);
  nor (_18971_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4]);
  nor (_18972_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4]);
  nor (_18973_, _18972_, _18971_);
  nand (_18974_, _18973_, _00227_);
  nand (_18975_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4]);
  nand (_18976_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4]);
  nand (_18977_, _18976_, _18975_);
  nand (_18978_, _18977_, _01417_);
  nand (_18981_, _18978_, _18974_);
  nand (_18982_, _18981_, _00560_);
  nor (_18983_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4]);
  nor (_18984_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4]);
  nor (_18985_, _18984_, _18983_);
  nand (_18986_, _18985_, _00227_);
  nand (_18987_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4]);
  nand (_18988_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4]);
  nand (_18989_, _18988_, _18987_);
  nand (_18990_, _18989_, _01417_);
  nand (_18991_, _18990_, _18986_);
  nand (_18992_, _18991_, _00561_);
  nand (_18993_, _18992_, _18982_);
  nand (_18994_, _18993_, _00465_);
  nand (_18995_, _18994_, _18970_);
  nand (_18996_, _18995_, _00248_);
  nand (_18997_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4]);
  nand (_18998_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4]);
  nand (_18999_, _18998_, _18997_);
  nand (_19000_, _18999_, _01417_);
  nand (_19001_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4]);
  nand (_19002_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4]);
  nand (_19003_, _19002_, _19001_);
  nand (_19004_, _19003_, _00227_);
  nand (_19005_, _19004_, _19000_);
  nand (_19006_, _19005_, _00560_);
  nand (_19007_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4]);
  nand (_19008_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4]);
  nand (_19009_, _19008_, _19007_);
  nand (_19010_, _19009_, _01417_);
  nand (_19011_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4]);
  nand (_19012_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4]);
  nand (_19013_, _19012_, _19011_);
  nand (_19014_, _19013_, _00227_);
  nand (_19015_, _19014_, _19010_);
  nand (_19016_, _19015_, _00561_);
  nand (_19017_, _19016_, _19006_);
  nand (_19018_, _19017_, _00466_);
  nor (_19019_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4]);
  nor (_19020_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4]);
  nor (_19022_, _19020_, _19019_);
  nand (_19023_, _19022_, _01417_);
  nor (_19024_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4]);
  nor (_19025_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  nor (_19026_, _19025_, _19024_);
  nand (_19027_, _19026_, _00227_);
  nand (_19028_, _19027_, _19023_);
  nand (_19029_, _19028_, _00560_);
  nor (_19030_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4]);
  nor (_19031_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4]);
  nor (_19032_, _19031_, _19030_);
  nand (_19033_, _19032_, _01417_);
  nor (_19034_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4]);
  nor (_19035_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4]);
  nor (_19036_, _19035_, _19034_);
  nand (_19037_, _19036_, _00227_);
  nand (_19038_, _19037_, _19033_);
  nand (_19039_, _19038_, _00561_);
  nand (_19040_, _19039_, _19029_);
  nand (_19041_, _19040_, _00465_);
  nand (_19042_, _19041_, _19018_);
  nand (_19043_, _19042_, _00247_);
  nand (_19044_, _19043_, _18996_);
  nand (_19045_, _19044_, _00320_);
  nand (_19046_, _19045_, _18947_);
  nand (_19047_, _19046_, _00386_);
  nand (_19048_, _19047_, _18849_);
  nor (_19049_, _19048_, _00156_);
  nand (_19050_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4]);
  nand (_19051_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4]);
  nand (_19052_, _19051_, _19050_);
  nand (_19053_, _19052_, _00227_);
  nand (_19054_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4]);
  nand (_19055_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4]);
  nand (_19056_, _19055_, _19054_);
  nand (_19057_, _19056_, _01417_);
  nand (_19058_, _19057_, _19053_);
  nand (_19059_, _19058_, _00560_);
  nand (_19060_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4]);
  nand (_19061_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4]);
  nand (_19062_, _19061_, _19060_);
  nand (_19063_, _19062_, _00227_);
  nand (_19064_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4]);
  nand (_19065_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4]);
  nand (_19066_, _19065_, _19064_);
  nand (_19067_, _19066_, _01417_);
  nand (_19068_, _19067_, _19063_);
  nand (_19069_, _19068_, _00561_);
  nand (_19070_, _19069_, _19059_);
  nand (_19071_, _19070_, _00466_);
  nand (_19073_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4]);
  nand (_19074_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4]);
  nand (_19075_, _19074_, _19073_);
  nand (_19076_, _19075_, _01417_);
  nor (_19077_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  nor (_19078_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4]);
  nor (_19079_, _19078_, _19077_);
  nand (_19080_, _19079_, _00227_);
  nand (_19081_, _19080_, _19076_);
  nand (_19082_, _19081_, _00560_);
  nand (_19083_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4]);
  nand (_19084_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4]);
  nand (_19085_, _19084_, _19083_);
  nand (_19086_, _19085_, _01417_);
  nor (_19087_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4]);
  nor (_19088_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4]);
  nor (_19089_, _19088_, _19087_);
  nand (_19090_, _19089_, _00227_);
  nand (_19091_, _19090_, _19086_);
  nand (_19092_, _19091_, _00561_);
  nand (_19093_, _19092_, _19082_);
  nand (_19094_, _19093_, _00465_);
  nand (_19095_, _19094_, _19071_);
  nand (_19096_, _19095_, _00248_);
  nand (_19097_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4]);
  nand (_19098_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4]);
  nand (_19099_, _19098_, _19097_);
  nand (_19100_, _19099_, _01417_);
  nand (_19101_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4]);
  nand (_19102_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4]);
  nand (_19103_, _19102_, _19101_);
  nand (_19104_, _19103_, _00227_);
  nand (_19105_, _19104_, _19100_);
  nand (_19106_, _19105_, _00560_);
  nand (_19107_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4]);
  nand (_19108_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4]);
  nand (_19109_, _19108_, _19107_);
  nand (_19110_, _19109_, _01417_);
  nand (_19111_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4]);
  nand (_19112_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4]);
  nand (_19113_, _19112_, _19111_);
  nand (_19114_, _19113_, _00227_);
  nand (_19115_, _19114_, _19110_);
  nand (_19116_, _19115_, _00561_);
  nand (_19117_, _19116_, _19106_);
  nand (_19118_, _19117_, _00466_);
  nor (_19119_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4]);
  nor (_19120_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4]);
  nor (_19121_, _19120_, _19119_);
  nand (_19122_, _19121_, _01417_);
  nor (_19123_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4]);
  nor (_19124_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4]);
  nor (_19125_, _19124_, _19123_);
  nand (_19126_, _19125_, _00227_);
  nand (_19127_, _19126_, _19122_);
  nand (_19128_, _19127_, _00560_);
  nor (_19129_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4]);
  nor (_19130_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4]);
  nor (_19131_, _19130_, _19129_);
  nor (_19132_, _19131_, _00227_);
  nor (_19133_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4]);
  nor (_19134_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4]);
  nor (_19135_, _19134_, _19133_);
  nor (_19136_, _19135_, _01417_);
  nor (_19137_, _19136_, _19132_);
  nand (_19138_, _19137_, _00561_);
  nand (_19139_, _19138_, _19128_);
  nand (_19140_, _19139_, _00465_);
  nand (_19141_, _19140_, _19118_);
  nand (_19142_, _19141_, _00247_);
  nand (_19143_, _19142_, _19096_);
  nand (_19144_, _19143_, _00320_);
  nand (_19145_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4]);
  nand (_19146_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4]);
  nand (_19147_, _19146_, _19145_);
  nand (_19148_, _19147_, _01417_);
  nand (_19149_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4]);
  nand (_19150_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4]);
  nand (_19151_, _19150_, _19149_);
  nand (_19152_, _19151_, _00227_);
  nand (_19154_, _19152_, _19148_);
  nand (_19155_, _19154_, _00560_);
  nand (_19156_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4]);
  nand (_19157_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4]);
  nand (_19158_, _19157_, _19156_);
  nand (_19159_, _19158_, _01417_);
  nand (_19160_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4]);
  nand (_19161_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4]);
  nand (_19162_, _19161_, _19160_);
  nand (_19163_, _19162_, _00227_);
  nand (_19164_, _19163_, _19159_);
  nand (_19165_, _19164_, _00561_);
  nand (_19166_, _19165_, _19155_);
  nand (_19167_, _19166_, _00466_);
  nor (_19168_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4]);
  nor (_19169_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4]);
  nor (_19170_, _19169_, _19168_);
  nand (_19171_, _19170_, _01417_);
  nor (_19172_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4]);
  nor (_19173_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4]);
  nor (_19175_, _19173_, _19172_);
  nand (_19176_, _19175_, _00227_);
  nand (_19177_, _19176_, _19171_);
  nand (_19178_, _19177_, _00560_);
  nor (_19179_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4]);
  nor (_19180_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4]);
  nor (_19181_, _19180_, _19179_);
  nand (_19182_, _19181_, _01417_);
  nor (_19183_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4]);
  nor (_19184_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4]);
  nor (_19185_, _19184_, _19183_);
  nand (_19186_, _19185_, _00227_);
  nand (_19187_, _19186_, _19182_);
  nand (_19188_, _19187_, _00561_);
  nand (_19189_, _19188_, _19178_);
  nand (_19190_, _19189_, _00465_);
  nand (_19191_, _19190_, _19167_);
  nand (_19192_, _19191_, _00248_);
  nand (_19193_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4]);
  nand (_19194_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4]);
  nand (_19196_, _19194_, _19193_);
  nand (_19197_, _19196_, _01417_);
  nand (_19198_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4]);
  nand (_19199_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4]);
  nand (_19200_, _19199_, _19198_);
  nand (_19201_, _19200_, _00227_);
  nand (_19202_, _19201_, _19197_);
  nand (_19203_, _19202_, _00560_);
  nand (_19204_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4]);
  nand (_19205_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4]);
  nand (_19206_, _19205_, _19204_);
  nand (_19207_, _19206_, _01417_);
  nand (_19208_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4]);
  nand (_19209_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4]);
  nand (_19210_, _19209_, _19208_);
  nand (_19211_, _19210_, _00227_);
  nand (_19212_, _19211_, _19207_);
  nand (_19213_, _19212_, _00561_);
  nand (_19214_, _19213_, _19203_);
  nand (_19215_, _19214_, _00466_);
  nor (_19217_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4]);
  nor (_19218_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4]);
  nor (_19219_, _19218_, _19217_);
  nand (_19220_, _19219_, _01417_);
  nor (_19221_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4]);
  nor (_19222_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4]);
  nor (_19223_, _19222_, _19221_);
  nand (_19224_, _19223_, _00227_);
  nand (_19225_, _19224_, _19220_);
  nand (_19226_, _19225_, _00560_);
  nor (_19227_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4]);
  nor (_19228_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4]);
  nor (_19229_, _19228_, _19227_);
  nand (_19230_, _19229_, _01417_);
  nor (_19231_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4]);
  nor (_19232_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4]);
  nor (_19233_, _19232_, _19231_);
  nand (_19234_, _19233_, _00227_);
  nand (_19235_, _19234_, _19230_);
  nand (_19236_, _19235_, _00561_);
  nand (_19238_, _19236_, _19226_);
  nand (_19239_, _19238_, _00465_);
  nand (_19240_, _19239_, _19215_);
  nand (_19241_, _19240_, _00247_);
  nand (_19242_, _19241_, _19192_);
  nand (_19243_, _19242_, _00319_);
  nand (_19244_, _19243_, _19144_);
  nand (_19245_, _19244_, _01629_);
  nand (_19246_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4]);
  nand (_19247_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4]);
  nand (_19248_, _19247_, _19246_);
  nand (_19249_, _19248_, _00227_);
  nand (_19250_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4]);
  nand (_19251_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4]);
  nand (_19252_, _19251_, _19250_);
  nand (_19253_, _19252_, _01417_);
  nand (_19254_, _19253_, _19249_);
  nand (_19255_, _19254_, _00560_);
  nand (_19256_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4]);
  nand (_19257_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4]);
  nand (_19259_, _19257_, _19256_);
  nand (_19260_, _19259_, _00227_);
  nand (_19261_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4]);
  nand (_19262_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4]);
  nand (_19263_, _19262_, _19261_);
  nand (_19264_, _19263_, _01417_);
  nand (_19265_, _19264_, _19260_);
  nand (_19266_, _19265_, _00561_);
  nand (_19267_, _19266_, _19255_);
  nand (_19268_, _19267_, _00466_);
  nand (_19269_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4]);
  nand (_19270_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4]);
  nand (_19271_, _19270_, _19269_);
  nand (_19272_, _19271_, _01417_);
  nor (_19273_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4]);
  nor (_19274_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4]);
  nor (_19275_, _19274_, _19273_);
  nand (_19276_, _19275_, _00227_);
  nand (_19277_, _19276_, _19272_);
  nand (_19278_, _19277_, _00560_);
  nand (_19280_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4]);
  nand (_19281_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4]);
  nand (_19282_, _19281_, _19280_);
  nand (_19283_, _19282_, _01417_);
  nor (_19284_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4]);
  nor (_19285_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4]);
  nor (_19286_, _19285_, _19284_);
  nand (_19287_, _19286_, _00227_);
  nand (_19288_, _19287_, _19283_);
  nand (_19289_, _19288_, _00561_);
  nand (_19291_, _19289_, _19278_);
  nand (_19292_, _19291_, _00465_);
  nand (_19293_, _19292_, _19268_);
  nand (_19294_, _19293_, _00248_);
  nand (_19295_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4]);
  nand (_19296_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4]);
  nand (_19297_, _19296_, _19295_);
  nand (_19298_, _19297_, _01417_);
  nand (_19299_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4]);
  nand (_19300_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4]);
  nand (_19302_, _19300_, _19299_);
  nand (_19303_, _19302_, _00227_);
  nand (_19304_, _19303_, _19298_);
  nand (_19305_, _19304_, _00560_);
  nand (_19306_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4]);
  nand (_19307_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4]);
  nand (_19308_, _19307_, _19306_);
  nand (_19309_, _19308_, _01417_);
  nand (_19310_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4]);
  nand (_19311_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4]);
  nand (_19312_, _19311_, _19310_);
  nand (_19313_, _19312_, _00227_);
  nand (_19314_, _19313_, _19309_);
  nand (_19315_, _19314_, _00561_);
  nand (_19316_, _19315_, _19305_);
  nand (_19317_, _19316_, _00466_);
  nor (_19318_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4]);
  nor (_19319_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4]);
  nor (_19320_, _19319_, _19318_);
  nand (_19321_, _19320_, _01417_);
  nor (_19323_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4]);
  nor (_19324_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4]);
  nor (_19325_, _19324_, _19323_);
  nand (_19326_, _19325_, _00227_);
  nand (_19327_, _19326_, _19321_);
  nand (_19328_, _19327_, _00560_);
  nor (_19329_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4]);
  nor (_19330_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4]);
  nor (_19331_, _19330_, _19329_);
  nor (_19332_, _19331_, _00227_);
  nor (_19333_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4]);
  nor (_19334_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4]);
  nor (_19335_, _19334_, _19333_);
  nor (_19336_, _19335_, _01417_);
  nor (_19337_, _19336_, _19332_);
  nand (_19338_, _19337_, _00561_);
  nand (_19339_, _19338_, _19328_);
  nand (_19340_, _19339_, _00465_);
  nand (_19341_, _19340_, _19317_);
  nand (_19342_, _19341_, _00247_);
  nand (_19343_, _19342_, _19294_);
  nand (_19344_, _19343_, _00320_);
  nand (_19345_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  nand (_19346_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4]);
  nand (_19347_, _19346_, _19345_);
  nand (_19348_, _19347_, _01417_);
  nand (_19349_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4]);
  nand (_19350_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4]);
  nand (_19351_, _19350_, _19349_);
  nand (_19352_, _19351_, _00227_);
  nand (_19353_, _19352_, _19348_);
  nand (_19354_, _19353_, _00560_);
  nand (_19355_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4]);
  nand (_19356_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4]);
  nand (_19357_, _19356_, _19355_);
  nand (_19358_, _19357_, _01417_);
  nand (_19359_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4]);
  nand (_19360_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4]);
  nand (_19361_, _19360_, _19359_);
  nand (_19362_, _19361_, _00227_);
  nand (_19363_, _19362_, _19358_);
  nand (_19364_, _19363_, _00561_);
  nand (_19365_, _19364_, _19354_);
  nand (_19366_, _19365_, _00466_);
  nor (_19367_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4]);
  nor (_19368_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4]);
  nor (_19369_, _19368_, _19367_);
  nand (_19370_, _19369_, _01417_);
  nor (_19371_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4]);
  nor (_19372_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4]);
  nor (_19373_, _19372_, _19371_);
  nand (_19374_, _19373_, _00227_);
  nand (_19375_, _19374_, _19370_);
  nand (_19376_, _19375_, _00560_);
  nor (_19377_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4]);
  nor (_19378_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4]);
  nor (_19379_, _19378_, _19377_);
  nand (_19380_, _19379_, _01417_);
  nor (_19381_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4]);
  nor (_19382_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4]);
  nor (_19383_, _19382_, _19381_);
  nand (_19384_, _19383_, _00227_);
  nand (_19385_, _19384_, _19380_);
  nand (_19386_, _19385_, _00561_);
  nand (_19387_, _19386_, _19376_);
  nand (_19388_, _19387_, _00465_);
  nand (_19389_, _19388_, _19366_);
  nand (_19390_, _19389_, _00247_);
  nand (_19391_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4]);
  nand (_19392_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4]);
  nand (_19394_, _19392_, _19391_);
  nand (_19395_, _19394_, _01417_);
  nand (_19396_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4]);
  nand (_19397_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4]);
  nand (_19398_, _19397_, _19396_);
  nand (_19399_, _19398_, _00227_);
  nand (_19400_, _19399_, _19395_);
  nand (_19401_, _19400_, _00560_);
  nand (_19402_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4]);
  nand (_19403_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4]);
  nand (_19404_, _19403_, _19402_);
  nand (_19405_, _19404_, _01417_);
  nand (_19406_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4]);
  nand (_19407_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4]);
  nand (_19408_, _19407_, _19406_);
  nand (_19409_, _19408_, _00227_);
  nand (_19410_, _19409_, _19405_);
  nand (_19411_, _19410_, _00561_);
  nand (_19412_, _19411_, _19401_);
  nand (_19413_, _19412_, _00466_);
  nor (_19414_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4]);
  nor (_19415_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4]);
  nor (_19416_, _19415_, _19414_);
  nand (_19417_, _19416_, _01417_);
  nor (_19418_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4]);
  nor (_19419_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4]);
  nor (_19420_, _19419_, _19418_);
  nand (_19421_, _19420_, _00227_);
  nand (_19422_, _19421_, _19417_);
  nand (_19423_, _19422_, _00560_);
  nor (_19424_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4]);
  nor (_19425_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4]);
  nor (_19426_, _19425_, _19424_);
  nand (_19427_, _19426_, _01417_);
  nor (_19428_, _00643_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  nor (_19429_, _00650_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4]);
  nor (_19430_, _19429_, _19428_);
  nand (_19431_, _19430_, _00227_);
  nand (_19432_, _19431_, _19427_);
  nand (_19433_, _19432_, _00561_);
  nand (_19434_, _19433_, _19423_);
  nand (_19435_, _19434_, _00465_);
  nand (_19436_, _19435_, _19413_);
  nand (_19437_, _19436_, _00248_);
  nand (_19438_, _19437_, _19390_);
  nand (_19439_, _19438_, _00319_);
  nand (_19440_, _19439_, _19344_);
  nand (_19441_, _19440_, _00386_);
  nand (_19442_, _19441_, _19245_);
  nor (_19443_, _19442_, _00556_);
  nor (_19444_, _19443_, _19049_);
  nor (_19445_, _19444_, _01416_);
  not (_19446_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  nand (_19447_, _01416_, _19446_);
  nand (_19448_, _19447_, _23493_);
  nor (_08963_, _19448_, _19445_);
  nor (_19449_, _22429_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1]);
  nor (_19450_, _22431_, _21474_);
  nor (_08965_, _19450_, _19449_);
  nor (_19451_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4]);
  nor (_19453_, _22473_, _21414_);
  nor (_08967_, _19453_, _19451_);
  nor (_19454_, _00919_, _00020_);
  nor (_19455_, _19454_, _17316_);
  nand (_19456_, _05045_, _00930_);
  nand (_19457_, _19456_, _00929_);
  nor (_19458_, _19457_, _19455_);
  nand (_19459_, _00928_, _00006_);
  nand (_19460_, _19459_, _23493_);
  nor (_08969_, _19460_, _19458_);
  nor (_19461_, _06624_, _24858_);
  nor (_19462_, _19461_, _00941_);
  nand (_19463_, _19461_, ABINPUT[0]);
  nand (_19464_, _19463_, _00929_);
  nor (_19465_, _19464_, _19462_);
  nand (_19466_, _00928_, _00029_);
  nand (_19467_, _19466_, _23493_);
  nor (_08971_, _19467_, _19465_);
  nand (_19468_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_19469_, _19468_, _00985_);
  not (_19470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand (_19471_, _00976_, _00954_);
  nand (_19472_, _19471_, _19470_);
  nand (_19473_, _19472_, _01302_);
  nand (_19474_, _19473_, _00996_);
  nor (_19475_, _19474_, _19469_);
  not (_19476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nand (_19477_, _00991_, _19476_);
  nand (_19478_, _19477_, _01006_);
  nor (_19479_, _19478_, _19475_);
  nor (_19480_, _01013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_19481_, _19480_, _01239_);
  nor (_19482_, _19481_, _19479_);
  nand (_19483_, _01013_, _00121_);
  nand (_19484_, _19483_, _23493_);
  nor (_08977_, _19484_, _19482_);
  nand (_19485_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_19486_, _19485_, _00985_);
  not (_19487_, _00975_);
  nand (_19488_, _19487_, _00954_);
  nand (_19489_, _19488_, _00958_);
  nand (_19490_, _19489_, _19471_);
  nand (_19491_, _19490_, _00996_);
  nor (_19492_, _19491_, _19486_);
  not (_19493_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nand (_19494_, _00991_, _19493_);
  nand (_19495_, _19494_, _01006_);
  nor (_19496_, _19495_, _19492_);
  nor (_19497_, _01013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_19498_, _19497_, _01239_);
  nor (_19499_, _19498_, _19496_);
  nand (_19500_, _01013_, _00006_);
  nand (_19501_, _19500_, _23493_);
  nor (_08981_, _19501_, _19499_);
  nor (_19502_, _15182_, _05573_);
  nor (_19503_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_19504_, _19503_, _05622_);
  nand (_19505_, _19504_, _05658_);
  nand (_19506_, _05628_, _05574_);
  nand (_19507_, _19506_, _15320_);
  nor (_19508_, _15166_, _05573_);
  nor (_19509_, _19508_, _15170_);
  nor (_19510_, _15168_, _05574_);
  nor (_19511_, _19510_, _19509_);
  nor (_19512_, _19511_, _05631_);
  nand (_19513_, _19503_, _05631_);
  nand (_19514_, _19513_, _15306_);
  nor (_19515_, _19514_, _19512_);
  nor (_19516_, _19515_, _19507_);
  nor (_19517_, _19516_, _19505_);
  not (_19518_, _19503_);
  nor (_19519_, _19518_, _15329_);
  nor (_19520_, _15146_, _05573_);
  nand (_19521_, _15150_, _15329_);
  nor (_19522_, _19521_, _19520_);
  nor (_19523_, _19522_, _19519_);
  nor (_19524_, _19523_, _05666_);
  nor (_19525_, _05667_, _14122_);
  nor (_19526_, _19525_, _05666_);
  nor (_19527_, _19526_, _05574_);
  nor (_19528_, _19527_, _19524_);
  nor (_19529_, _19528_, _05665_);
  nor (_19530_, _19503_, _14114_);
  nor (_19531_, _19530_, _15336_);
  nor (_19532_, _19531_, _19529_);
  nor (_19533_, _19532_, _19517_);
  nor (_19534_, _19533_, _05606_);
  nor (_19535_, _19534_, _19502_);
  nor (_08983_, _19535_, rst);
  nor (_19536_, _21933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5]);
  nor (_19537_, _21935_, _21451_);
  nor (_08986_, _19537_, _19536_);
  nor (_19538_, _21933_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6]);
  nor (_19539_, _21935_, _21504_);
  nor (_08988_, _19539_, _19538_);
  nor (_19540_, _22198_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5]);
  nor (_19541_, _22200_, _21451_);
  nor (_08990_, _19541_, _19540_);
  nor (_19542_, _12408_, _12404_);
  nor (_19543_, _19542_, _12410_);
  nor (_19544_, _19543_, _23490_);
  nand (_19545_, _23490_, _23056_);
  nand (_19546_, _19545_, _12372_);
  nor (_08992_, _19546_, _19544_);
  not (_19547_, _12326_);
  nand (_19548_, _19547_, _23044_);
  nor (_19549_, _19548_, _23055_);
  nand (_19550_, _19548_, _23055_);
  nand (_19551_, _19550_, _12372_);
  nor (_25037_[0], _19551_, _19549_);
  nor (_19552_, _12387_, _02286_);
  nor (_19553_, _19552_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  nor (_08995_, _19553_, rst);
  nor (_19554_, _07002_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0]);
  nor (_19555_, _07004_, _21586_);
  nor (_09005_, _19555_, _19554_);
  nor (_19556_, _22526_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5]);
  nor (_19557_, _22528_, _21451_);
  nor (_09008_, _19557_, _19556_);
  nand (_19558_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_19559_, _19558_, _00985_);
  not (_19560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_19561_, _00974_, _00954_);
  nand (_19562_, _19561_, _19560_);
  nand (_19563_, _19562_, _19488_);
  nand (_19564_, _19563_, _00996_);
  nor (_19565_, _19564_, _19559_);
  not (_19566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nand (_19567_, _00991_, _19566_);
  nand (_19568_, _19567_, _01006_);
  nor (_19569_, _19568_, _19565_);
  nor (_19570_, _01013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor (_19571_, _19570_, _01239_);
  nor (_19572_, _19571_, _19569_);
  nand (_19573_, _01013_, _00029_);
  nand (_19574_, _19573_, _23493_);
  nor (_09011_, _19574_, _19572_);
  nor (_19575_, _24380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3]);
  nor (_19576_, _24382_, _21526_);
  nor (_09056_, _19576_, _19575_);
  nand (_19579_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_19580_, _19579_, _00985_);
  not (_19581_, _06645_);
  not (_19582_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nand (_19583_, _00980_, _00954_);
  nand (_19584_, _19583_, _19582_);
  nand (_19585_, _19584_, _19581_);
  nand (_19586_, _19585_, _00996_);
  nor (_19587_, _19586_, _19580_);
  not (_19588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nand (_19589_, _00991_, _19588_);
  nand (_19590_, _19589_, _01006_);
  nor (_19591_, _19590_, _19587_);
  nor (_19592_, _01013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_19593_, _19592_, _01239_);
  nor (_19594_, _19593_, _19591_);
  nand (_19595_, _01013_, _00114_);
  nand (_19596_, _19595_, _23493_);
  nor (_09059_, _19596_, _19594_);
  nand (_19597_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nor (_19598_, _19597_, _00985_);
  not (_19599_, _00979_);
  nand (_19600_, _19599_, _00954_);
  nand (_19601_, _19600_, _00956_);
  nand (_19602_, _19601_, _19583_);
  nand (_19603_, _19602_, _00996_);
  nor (_19604_, _19603_, _19598_);
  not (_19605_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nand (_19606_, _00991_, _19605_);
  nand (_19607_, _19606_, _01006_);
  nor (_19608_, _19607_, _19604_);
  nor (_19609_, _01013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_19610_, _19609_, _01239_);
  nor (_19611_, _19610_, _19608_);
  nand (_19612_, _01013_, _00129_);
  nand (_19613_, _19612_, _23493_);
  nor (_09061_, _19613_, _19611_);
  nand (_19614_, _00945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_19615_, _19614_, _00985_);
  not (_19616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nand (_19617_, _00978_, _00954_);
  nand (_19618_, _19617_, _19616_);
  nand (_19619_, _19618_, _19600_);
  nand (_19620_, _19619_, _00996_);
  nor (_19621_, _19620_, _19615_);
  not (_19622_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nand (_19623_, _00991_, _19622_);
  nand (_19624_, _19623_, _01006_);
  nor (_19625_, _19624_, _19621_);
  nor (_19626_, _01013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_19627_, _19626_, _01239_);
  nor (_19628_, _19627_, _19625_);
  nand (_19629_, _01013_, _24900_);
  nand (_19630_, _19629_, _23493_);
  nor (_09064_, _19630_, _19628_);
  nor (_19631_, _00880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0]);
  nor (_19632_, _00882_, _21586_);
  nor (_09077_, _19632_, _19631_);
  nor (_19633_, _10797_, _05559_);
  nor (_19634_, _19633_, _17714_);
  nor (_19635_, _10797_, _06627_);
  nor (_19636_, _19635_, _19634_);
  nor (_19637_, _19636_, _00915_);
  nand (_19638_, _00913_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_19639_, _10798_, _11588_);
  nor (_19640_, _10798_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor (_19641_, _19640_, _00010_);
  nand (_19642_, _19641_, _19639_);
  nand (_19643_, _19642_, _19638_);
  nor (_19644_, _19643_, _19637_);
  nor (_09090_, _19644_, rst);
  nor (_19645_, _21733_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4]);
  nor (_19646_, _21735_, _21414_);
  nor (_09101_, _19646_, _19645_);
  nor (_19647_, _22479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5]);
  nor (_19648_, _22482_, _21451_);
  nor (_09107_, _19648_, _19647_);
  nor (_19649_, _22227_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4]);
  nor (_19650_, _22229_, _21414_);
  nor (_09126_, _19650_, _19649_);
  nor (_19651_, _22479_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7]);
  nor (_19652_, _22482_, _21626_);
  nor (_25069_, _19652_, _19651_);
  nor (_19653_, _22496_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5]);
  nor (_19654_, _22498_, _21451_);
  nor (_25064_, _19654_, _19653_);
  nor (_19655_, _22450_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1]);
  nor (_19656_, _22452_, _21474_);
  nor (_25087_, _19656_, _19655_);
  nor (_19657_, _00880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7]);
  nor (_19658_, _00882_, _21626_);
  nor (_25289_, _19658_, _19657_);
  nand (_19659_, _08687_, first_instr);
  nand (_00000_, _19659_, _23493_);
  nor (_19660_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _15132_);
  nor (_19661_, _15136_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_19662_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_19663_, _19662_, _19661_);
  nand (_19664_, _19663_, _19660_);
  nand (_19665_, _19664_, _15124_);
  nor (_19666_, _15136_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_19667_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_19668_, _19667_, _15132_);
  not (_19669_, _19668_);
  nor (_19670_, _19669_, _19666_);
  nor (_19671_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_19672_, _15136_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_19673_, _19672_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  not (_19674_, _19673_);
  nor (_19675_, _19674_, _19671_);
  nor (_19676_, _19675_, _19670_);
  nor (_19677_, _19676_, _15128_);
  not (_19678_, _19677_);
  nor (_19679_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_19680_, _15136_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_19681_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_19682_, _19681_, _19680_);
  nand (_19683_, _19682_, _19679_);
  nand (_19684_, _19683_, _19678_);
  nor (_19685_, _19684_, _19665_);
  nor (_19686_, _15136_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_19687_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_19688_, _19687_, _19686_);
  nor (_19689_, _19688_, _15132_);
  nor (_19690_, _15136_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_19691_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_19692_, _19691_, _19690_);
  nor (_19693_, _19692_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_19694_, _19693_, _19689_);
  not (_19695_, _19694_);
  nor (_19696_, _19695_, _15128_);
  nor (_19697_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_19698_, _15136_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_19699_, _19698_, _19697_);
  nand (_19700_, _19699_, _19679_);
  not (_19701_, _19700_);
  not (_19702_, _19660_);
  nor (_19703_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_19704_, _15136_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_19705_, _19704_, _19703_);
  not (_19706_, _19705_);
  nor (_19707_, _19706_, _19702_);
  nor (_19708_, _19707_, _19701_);
  not (_19709_, _19708_);
  nor (_19710_, _19709_, _19696_);
  nand (_19711_, _19710_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_19712_, _19711_);
  nor (_19713_, _19712_, _19685_);
  not (_19714_, _19713_);
  nor (_19715_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _15128_);
  not (_19716_, _19715_);
  nor (_19717_, _19716_, _08101_);
  nor (_19718_, _15124_, _15128_);
  not (_19719_, _19718_);
  nor (_19720_, _19719_, _09419_);
  nor (_19721_, _19720_, _19717_);
  nor (_19722_, _15124_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not (_19723_, _19722_);
  nor (_19724_, _19723_, _09413_);
  nor (_19725_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not (_19726_, _19725_);
  nor (_19727_, _19726_, _09415_);
  nor (_19728_, _19727_, _19724_);
  nand (_19729_, _19728_, _19721_);
  nor (_19730_, _19729_, _15132_);
  nor (_19731_, _19716_, _07577_);
  nor (_19732_, _19719_, _07697_);
  nor (_19733_, _19732_, _19731_);
  nor (_19734_, _19723_, _07435_);
  nor (_19735_, _19726_, _07300_);
  nor (_19736_, _19735_, _19734_);
  nand (_19737_, _19736_, _19733_);
  nor (_19738_, _19737_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_19739_, _19738_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_19740_, _19739_);
  nor (_19741_, _19740_, _19730_);
  nor (_19742_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _15136_);
  nor (_19743_, _19719_, _08738_);
  nand (_19744_, _19725_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  not (_19745_, _19744_);
  nor (_19746_, _19745_, _19743_);
  nand (_19747_, _19715_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  not (_19748_, _19747_);
  nor (_19749_, _19723_, _08472_);
  nor (_19750_, _19749_, _19748_);
  nand (_19751_, _19750_, _19746_);
  nand (_19752_, _19751_, _19742_);
  not (_19753_, _19752_);
  nor (_19754_, _15132_, _15136_);
  not (_19755_, _19754_);
  nor (_19756_, _19719_, _09240_);
  not (_19757_, _19756_);
  nand (_19758_, _19715_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand (_19759_, _19758_, _19757_);
  nand (_19760_, _19725_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nand (_19761_, _19722_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand (_19762_, _19761_, _19760_);
  nor (_19763_, _19762_, _19759_);
  nor (_19764_, _19763_, _19755_);
  nor (_19765_, _19764_, _19753_);
  not (_19766_, _19765_);
  nor (_19767_, _19766_, _19741_);
  nor (_19768_, _19767_, _19714_);
  not (_19769_, _19768_);
  nor (_19770_, _19716_, _09469_);
  nor (_19771_, _19719_, _09467_);
  nor (_19772_, _19771_, _19770_);
  nor (_19773_, _19723_, _09462_);
  nor (_19774_, _19726_, _07859_);
  nor (_19775_, _19774_, _19773_);
  nand (_19776_, _19775_, _19772_);
  nor (_19777_, _19776_, _15132_);
  nor (_19778_, _19716_, _07591_);
  nor (_19779_, _19719_, _07711_);
  nor (_19780_, _19779_, _19778_);
  nor (_19781_, _19723_, _07448_);
  nor (_19782_, _19726_, _07316_);
  nor (_19783_, _19782_, _19781_);
  nand (_19784_, _19783_, _19780_);
  nor (_19785_, _19784_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_19786_, _19785_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_19787_, _19786_);
  nor (_19788_, _19787_, _19777_);
  nor (_19789_, _19719_, _08749_);
  nand (_19790_, _19725_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  not (_19791_, _19790_);
  nor (_19792_, _19791_, _19789_);
  nor (_19793_, _19716_, _08615_);
  nor (_19794_, _19723_, _08488_);
  nor (_19795_, _19794_, _19793_);
  nand (_19796_, _19795_, _19792_);
  nand (_19797_, _19796_, _19742_);
  not (_19798_, _19797_);
  nor (_19799_, _19719_, _09252_);
  not (_19800_, _19799_);
  nand (_19801_, _19715_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nand (_19802_, _19801_, _19800_);
  nand (_19803_, _19725_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nand (_19804_, _19722_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nand (_19805_, _19804_, _19803_);
  nor (_19807_, _19805_, _19802_);
  nor (_19808_, _19807_, _19755_);
  nor (_19809_, _19808_, _19798_);
  not (_19810_, _19809_);
  nor (_19811_, _19810_, _19788_);
  nor (_19812_, _19811_, _19714_);
  nand (_19813_, _19715_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  not (_19814_, _19813_);
  nor (_19815_, _19719_, _08182_);
  nor (_19816_, _19815_, _19814_);
  not (_19817_, _19816_);
  nand (_19818_, _19722_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nand (_19819_, _19725_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nand (_19820_, _19819_, _19818_);
  nor (_19821_, _19820_, _19817_);
  nand (_19822_, _19821_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_19823_, _19716_, _07541_);
  nand (_19824_, _19718_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  not (_19825_, _19824_);
  nor (_19826_, _19825_, _19823_);
  nand (_19827_, _19722_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  not (_19828_, _19827_);
  nor (_19829_, _19726_, _07263_);
  nor (_19830_, _19829_, _19828_);
  nand (_19831_, _19830_, _19826_);
  nor (_19832_, _19831_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_19833_, _19832_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nand (_19834_, _19833_, _19822_);
  not (_19835_, _19742_);
  nand (_19836_, _19718_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  nand (_19838_, _19715_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  nand (_19839_, _19838_, _19836_);
  nor (_19840_, _19726_, _08303_);
  not (_19841_, _19840_);
  nand (_19842_, _19722_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nand (_19843_, _19842_, _19841_);
  nor (_19844_, _19843_, _19839_);
  nor (_19845_, _19844_, _19835_);
  nor (_19846_, _19719_, _09214_);
  not (_19847_, _19846_);
  nand (_19848_, _19715_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nand (_19849_, _19848_, _19847_);
  nand (_19850_, _19725_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nand (_19851_, _19722_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nand (_19852_, _19851_, _19850_);
  nor (_19853_, _19852_, _19849_);
  nor (_19854_, _19853_, _19755_);
  nor (_19855_, _19854_, _19845_);
  nand (_19856_, _19855_, _19834_);
  nand (_19857_, _19856_, _19713_);
  not (_19858_, _19857_);
  nor (_19859_, _19858_, _19812_);
  nand (_19860_, _19859_, _19769_);
  nor (_19861_, _19716_, _09370_);
  nor (_19862_, _19719_, _09368_);
  nor (_19863_, _19862_, _19861_);
  nor (_19864_, _19723_, _07965_);
  nor (_19865_, _19726_, _09364_);
  nor (_19866_, _19865_, _19864_);
  nand (_19867_, _19866_, _19863_);
  nor (_19868_, _19867_, _15132_);
  nand (_19869_, _19722_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  not (_19870_, _19869_);
  nor (_19871_, _19870_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_19872_, _19716_, _07562_);
  nand (_19873_, _19718_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nand (_19874_, _19725_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nand (_19875_, _19874_, _19873_);
  nor (_19876_, _19875_, _19872_);
  nand (_19877_, _19876_, _19871_);
  nand (_19878_, _19877_, _15136_);
  nor (_19879_, _19878_, _19868_);
  nand (_19880_, _19718_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  not (_19881_, _19880_);
  nor (_19882_, _19726_, _08320_);
  nor (_19883_, _19882_, _19881_);
  nor (_19884_, _19716_, _08586_);
  nor (_19885_, _19723_, _08457_);
  nor (_19886_, _19885_, _19884_);
  nand (_19887_, _19886_, _19883_);
  nand (_19888_, _19887_, _19742_);
  not (_19889_, _19888_);
  nor (_19890_, _19719_, _09228_);
  not (_19891_, _19890_);
  nand (_19892_, _19715_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nand (_19893_, _19892_, _19891_);
  nand (_19894_, _19725_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nand (_19895_, _19722_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nand (_19896_, _19895_, _19894_);
  nor (_19897_, _19896_, _19893_);
  nor (_19898_, _19897_, _19755_);
  nor (_19899_, _19898_, _19889_);
  not (_19900_, _19899_);
  nor (_19901_, _19900_, _19879_);
  nor (_19902_, _19716_, _09566_);
  nor (_19903_, _19719_, _09564_);
  nor (_19904_, _19903_, _19902_);
  nor (_19905_, _19723_, _08020_);
  nor (_19906_, _19726_, _09560_);
  nor (_19907_, _19906_, _19905_);
  nand (_19908_, _19907_, _19904_);
  nor (_19909_, _19908_, _15132_);
  nor (_19910_, _19716_, _07617_);
  nand (_19911_, _19718_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  not (_19912_, _19911_);
  nor (_19913_, _19912_, _19910_);
  nor (_19914_, _19723_, _07476_);
  nor (_19915_, _19726_, _07347_);
  nor (_19916_, _19915_, _19914_);
  nand (_19917_, _19916_, _19913_);
  nor (_19918_, _19917_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_19919_, _19918_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_19920_, _19919_);
  nor (_19921_, _19920_, _19909_);
  nor (_19922_, _19719_, _08796_);
  nand (_19923_, _19725_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  not (_19924_, _19923_);
  nor (_19925_, _19924_, _19922_);
  nor (_19926_, _19716_, _08642_);
  nor (_19927_, _19723_, _08519_);
  nor (_19928_, _19927_, _19926_);
  nand (_19929_, _19928_, _19925_);
  nand (_19930_, _19929_, _19742_);
  not (_19931_, _19930_);
  nor (_19932_, _19719_, _09276_);
  not (_19933_, _19932_);
  nand (_19934_, _19715_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nand (_19935_, _19934_, _19933_);
  nand (_19936_, _19725_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nand (_19937_, _19722_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nand (_19938_, _19937_, _19936_);
  nor (_19939_, _19938_, _19935_);
  nor (_19940_, _19939_, _19755_);
  nor (_19941_, _19940_, _19931_);
  not (_19942_, _19941_);
  nor (_19943_, _19942_, _19921_);
  nor (_19944_, _19943_, _19714_);
  nor (_19945_, _19716_, _09517_);
  nor (_19946_, _19719_, _09515_);
  nor (_19947_, _19946_, _19945_);
  nor (_19948_, _19723_, _08005_);
  nor (_19949_, _19726_, _07878_);
  nor (_19950_, _19949_, _19948_);
  nand (_19951_, _19950_, _19947_);
  nor (_19952_, _19951_, _15132_);
  nor (_19953_, _19716_, _07604_);
  nor (_19954_, _19719_, _07727_);
  nor (_19955_, _19954_, _19953_);
  nor (_19956_, _19723_, _07463_);
  nor (_19957_, _19726_, _07333_);
  nor (_19958_, _19957_, _19956_);
  nand (_19959_, _19958_, _19955_);
  nor (_19960_, _19959_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_19961_, _19960_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_19962_, _19961_);
  nor (_19963_, _19962_, _19952_);
  nor (_19964_, _19719_, _08769_);
  nor (_19965_, _19726_, _08365_);
  nor (_19966_, _19965_, _19964_);
  nor (_19967_, _19716_, _08629_);
  nand (_19968_, _19722_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  not (_19969_, _19968_);
  nor (_19970_, _19969_, _19967_);
  nand (_19971_, _19970_, _19966_);
  nand (_19972_, _19971_, _19742_);
  not (_19973_, _19972_);
  nor (_19974_, _19719_, _09264_);
  not (_19975_, _19974_);
  nand (_19976_, _19715_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nand (_19977_, _19976_, _19975_);
  nand (_19978_, _19725_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nand (_19979_, _19722_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nand (_19980_, _19979_, _19978_);
  nor (_19981_, _19980_, _19977_);
  nor (_19982_, _19981_, _19755_);
  nor (_19983_, _19982_, _19973_);
  not (_19984_, _19983_);
  nor (_19985_, _19984_, _19963_);
  nor (_19986_, _19985_, _19714_);
  not (_19987_, _19986_);
  nor (_19988_, _19987_, _19944_);
  nand (_19989_, _19988_, _19901_);
  nor (_19990_, _19989_, _19860_);
  not (_19991_, _19944_);
  not (_19992_, _19812_);
  nor (_19993_, _19901_, _19714_);
  nor (_19994_, _19993_, _19769_);
  nand (_19995_, _19994_, _19992_);
  nor (_19996_, _19995_, _19857_);
  nand (_19997_, _19996_, _19991_);
  nor (_19998_, _19997_, _19986_);
  nor (_19999_, _19998_, _19990_);
  nand (_20000_, _19715_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_20001_, _19718_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_20002_, _20001_, _20000_);
  nor (_20003_, _19723_, _06169_);
  nor (_20004_, _19726_, _06171_);
  nor (_20005_, _20004_, _20003_);
  not (_20006_, _20005_);
  nor (_20007_, _20006_, _20002_);
  nand (_20008_, _20007_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_20009_, _19716_, _07641_);
  nor (_20010_, _19719_, _07773_);
  nor (_20011_, _20010_, _20009_);
  nor (_20012_, _19723_, _07503_);
  nor (_20013_, _19726_, _07377_);
  nor (_20014_, _20013_, _20012_);
  nand (_20015_, _20014_, _20011_);
  nor (_20016_, _20015_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_20017_, _20016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nand (_20018_, _20017_, _20008_);
  not (_20019_, _20018_);
  nand (_20020_, _19718_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  not (_20021_, _20020_);
  nor (_20022_, _19726_, _08412_);
  nor (_20023_, _20022_, _20021_);
  nor (_20024_, _19716_, _08672_);
  nor (_20025_, _19723_, _08551_);
  nor (_20026_, _20025_, _20024_);
  nand (_20027_, _20026_, _20023_);
  nand (_20028_, _19742_, _20027_);
  nor (_20029_, _19719_, _06139_);
  nor (_20030_, _19726_, _06135_);
  nor (_20031_, _20030_, _20029_);
  nor (_20032_, _19716_, _06141_);
  nor (_20033_, _19723_, _06131_);
  nor (_20034_, _20033_, _20032_);
  nand (_20035_, _20034_, _20031_);
  nand (_20036_, _20035_, _19754_);
  nand (_20037_, _20036_, _20028_);
  nor (_20038_, _20037_, _20019_);
  nor (_20039_, _20038_, _19714_);
  nor (_20040_, _19716_, _08149_);
  nor (_20041_, _19719_, _09614_);
  nor (_20042_, _20041_, _20040_);
  nor (_20043_, _19723_, _09608_);
  nor (_20044_, _19726_, _09610_);
  nor (_20045_, _20044_, _20043_);
  nand (_20046_, _20045_, _20042_);
  nor (_20047_, _20046_, _15132_);
  nor (_20048_, _19716_, _07629_);
  nand (_20049_, _19718_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  not (_20050_, _20049_);
  nor (_20051_, _20050_, _20048_);
  nand (_20052_, _19722_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  not (_20053_, _20052_);
  nor (_20054_, _19726_, _07362_);
  nor (_20055_, _20054_, _20053_);
  nand (_20056_, _20055_, _20051_);
  nor (_20057_, _20056_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_20058_, _20057_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_20059_, _20058_);
  nor (_20060_, _20059_, _20047_);
  nor (_20061_, _19719_, _08812_);
  nor (_20062_, _19726_, _08398_);
  nor (_20063_, _20062_, _20061_);
  nor (_20064_, _19716_, _08658_);
  nor (_20065_, _19723_, _08535_);
  nor (_20066_, _20065_, _20064_);
  nand (_20067_, _20066_, _20063_);
  nand (_20068_, _20067_, _19742_);
  not (_20069_, _20068_);
  nor (_20070_, _19719_, _09288_);
  not (_20071_, _20070_);
  nand (_20072_, _19715_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nand (_20073_, _20072_, _20071_);
  nand (_20074_, _19725_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nand (_20075_, _19722_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nand (_20076_, _20075_, _20074_);
  nor (_20077_, _20076_, _20073_);
  nor (_20078_, _20077_, _19755_);
  nor (_20079_, _20078_, _20069_);
  not (_20080_, _20079_);
  nor (_20081_, _20080_, _20060_);
  nand (_20082_, _20081_, _20039_);
  nor (_20083_, _20082_, _19999_);
  nor (_20084_, _19987_, _19991_);
  not (_20085_, _19993_);
  nor (_20086_, _20085_, _19857_);
  nand (_20087_, _20086_, _19769_);
  nor (_20088_, _20087_, _19812_);
  nor (_20089_, _20088_, _20084_);
  not (_20090_, _19996_);
  nand (_20091_, _20084_, _20090_);
  not (_20092_, _20038_);
  nor (_20093_, _20081_, _19714_);
  not (_20094_, _20093_);
  nor (_20095_, _20094_, _20092_);
  nand (_20096_, _20095_, _20091_);
  nor (_20097_, _20096_, _20089_);
  nor (_20098_, _20097_, _20083_);
  nor (_20099_, _15264_, _15260_);
  not (_20100_, _20099_);
  nor (_20101_, _20100_, _15274_);
  not (_20102_, _20101_);
  nor (_20103_, _15248_, _15238_);
  nand (_20104_, _20103_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_20105_, _20104_, _15256_);
  not (_20106_, _20105_);
  nor (_20107_, _19725_, _19755_);
  not (_20108_, _20107_);
  nor (_20109_, _20108_, _20106_);
  not (_20110_, _20109_);
  nor (_20111_, _20110_, _20102_);
  not (_20112_, _20111_);
  nor (_20113_, _20112_, _15278_);
  nand (_20114_, _20113_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not (_20115_, _20114_);
  nor (_20116_, _20102_, _15278_);
  not (_20117_, _20116_);
  nor (_20118_, _20110_, _20117_);
  nor (_20119_, _20118_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_20120_, _20119_, _20115_);
  nand (_20121_, _20120_, _15098_);
  nor (_20122_, _20110_, _15260_);
  not (_20123_, _20122_);
  nor (_20124_, _20123_, _15264_);
  nor (_20125_, _20124_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_20126_, _20125_, _20111_);
  nand (_20127_, _20126_, _15089_);
  nand (_20128_, _20127_, _20121_);
  not (_20129_, _20126_);
  nand (_20130_, _20129_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_20131_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_20132_, _15286_, _15102_);
  nor (_20133_, _20132_, _20131_);
  not (_20134_, _20133_);
  nand (_20135_, _20114_, _20134_);
  nand (_20136_, _20115_, _20133_);
  nand (_20137_, _20136_, _20135_);
  nand (_20138_, _20137_, _20130_);
  nor (_20139_, _20138_, _20128_);
  nor (_20140_, _20111_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_20141_, _20140_, _20113_);
  not (_20142_, _20141_);
  nand (_20143_, _20142_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_20144_, _20122_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_20145_, _20144_, _20124_);
  not (_20146_, _20145_);
  nor (_20147_, _20146_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_20148_, _20145_, _15085_);
  nor (_20149_, _20148_, _20147_);
  nand (_20150_, _20149_, _20143_);
  nand (_20151_, _20141_, _15093_);
  nor (_20152_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_20153_, _15248_, _15066_);
  nor (_20154_, _20153_, _20152_);
  nor (_20155_, _20108_, _15238_);
  not (_20156_, _20155_);
  nand (_20157_, _20156_, _20154_);
  nor (_20158_, _19725_, _15132_);
  nor (_20159_, _20158_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_20160_, _20159_, _20107_);
  not (_20161_, _20160_);
  nor (_20162_, _20161_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_20163_, _20156_, _20154_);
  nor (_20164_, _20163_, _20162_);
  nand (_20165_, _20164_, _20157_);
  nor (_20166_, _19715_, _19722_);
  nand (_20167_, _20166_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_20169_, _20166_);
  nand (_20170_, _20169_, _15041_);
  nand (_20171_, _20170_, _20167_);
  nand (_20172_, _19679_, _15124_);
  not (_20173_, _20172_);
  nor (_20174_, _20173_, _20158_);
  nand (_20175_, _20174_, _15048_);
  nand (_20176_, _20175_, _20171_);
  not (_20177_, _20174_);
  nand (_20178_, _20177_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_20179_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_20180_, _15238_, _15056_);
  nor (_20181_, _20180_, _20179_);
  nand (_20182_, _20108_, _20181_);
  nand (_20183_, _20182_, _20178_);
  nor (_20184_, _20183_, _20176_);
  nor (_20185_, _20160_, _15052_);
  nand (_20186_, _15037_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_20187_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], _15124_);
  nand (_20188_, _20187_, _20186_);
  not (_20189_, _20181_);
  nand (_20190_, _20107_, _20189_);
  nand (_20191_, _20190_, _20188_);
  nor (_20192_, _20191_, _20185_);
  nand (_20193_, _20192_, _20184_);
  nor (_20194_, _20193_, _20165_);
  nand (_20195_, _20194_, _20151_);
  nor (_20196_, _20108_, _20104_);
  nor (_20197_, _20156_, _15248_);
  nor (_20198_, _20197_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_20199_, _20198_, _20196_);
  nand (_20200_, _20199_, _15072_);
  not (_20201_, _20199_);
  nand (_20202_, _20201_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_20203_, _20202_, _20200_);
  nor (_20204_, _20203_, _20195_);
  nor (_20205_, _20120_, _15098_);
  nor (_20206_, _20109_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_20207_, _20206_, _20122_);
  nor (_20208_, _20207_, _15081_);
  nor (_20209_, _20196_, _15256_);
  nand (_20210_, _20196_, _15256_);
  not (_20211_, _20210_);
  nor (_20212_, _20211_, _20209_);
  not (_20213_, _20212_);
  nor (_20214_, _20213_, _15077_);
  nor (_20215_, _20214_, _20208_);
  not (_20216_, _20207_);
  nor (_20217_, _20216_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_20218_, _20212_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_20219_, _20218_, _20217_);
  nand (_20220_, _20219_, _20215_);
  nor (_20221_, _20220_, _20205_);
  nand (_20222_, _20221_, _20204_);
  nor (_20223_, _20222_, _20150_);
  nand (_20224_, _20223_, _20139_);
  nand (_20225_, _20118_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_20226_, _20225_, _15286_);
  not (_20227_, _20226_);
  nor (_20228_, _20227_, _15290_);
  not (_20229_, _20228_);
  nand (_20230_, _20229_, _08696_);
  nand (_20231_, _20228_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nand (_20232_, _20231_, _20230_);
  nand (_20233_, _20232_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_20234_, _20232_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_20235_, _20226_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_20236_, _20235_, _20228_);
  not (_20237_, _20236_);
  nor (_20238_, _20237_, _15106_);
  nor (_20239_, _20236_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_20240_, _20239_, _20238_);
  nor (_20241_, _20240_, _20234_);
  nand (_20242_, _20241_, _20233_);
  nor (_20243_, _20242_, _20224_);
  nor (_20244_, _20243_, _20098_);
  nor (_20245_, _19755_, _15128_);
  not (_20246_, _20245_);
  nor (_20247_, _20246_, _20106_);
  not (_20248_, _20247_);
  nor (_20249_, _20248_, _20100_);
  not (_20250_, _20249_);
  nor (_20251_, _20250_, _15274_);
  not (_20252_, _20251_);
  nor (_20253_, _20252_, _15278_);
  nand (_20254_, _20253_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_20255_, _20254_, _15286_);
  not (_20256_, _20255_);
  nor (_20257_, _20256_, _15290_);
  not (_20258_, _20257_);
  nor (_20259_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_20260_, _08696_, _08690_);
  nor (_20261_, _20260_, _20259_);
  not (_20262_, _20261_);
  nor (_20263_, _20255_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not (_20264_, _20263_);
  nand (_20265_, _20264_, _15106_);
  nand (_20266_, _20265_, _20262_);
  nand (_20267_, _20266_, _20258_);
  nor (_20268_, _20263_, _20257_);
  nor (_20269_, _20268_, _15106_);
  not (_20270_, _20254_);
  nand (_20271_, _20134_, _20270_);
  nor (_20272_, _15128_, _15132_);
  nand (_20273_, _20272_, _15136_);
  not (_20274_, _20272_);
  nand (_20275_, _20274_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nand (_20276_, _20275_, _20273_);
  nand (_20277_, _20276_, _15052_);
  nor (_20278_, _20276_, _15052_);
  nand (_20279_, _20189_, _20245_);
  nor (_20280_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _15128_);
  nor (_20281_, _15041_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_20282_, _20281_, _20280_);
  nor (_20283_, _20188_, _20282_);
  nand (_20284_, _20283_, _20279_);
  nor (_20285_, _20284_, _20278_);
  nand (_20286_, _20285_, _20277_);
  nor (_20287_, _20246_, _15238_);
  nand (_20288_, _20154_, _20287_);
  not (_20289_, _20287_);
  not (_20290_, _20154_);
  nand (_20291_, _20290_, _20289_);
  nand (_20292_, _20291_, _20288_);
  nor (_20293_, _15128_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  not (_20294_, _20293_);
  nand (_20295_, _20294_, _19702_);
  nor (_20296_, _20295_, _15048_);
  nand (_20297_, _20295_, _15048_);
  nand (_20298_, _20181_, _20246_);
  nand (_20299_, _20298_, _20297_);
  nor (_20300_, _20299_, _20296_);
  nand (_20301_, _20300_, _20292_);
  nor (_20302_, _20301_, _20286_);
  nor (_20303_, _20248_, _15260_);
  nor (_20304_, _20247_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_20305_, _20304_, _20303_);
  not (_20306_, _20305_);
  nor (_20307_, _20306_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_20308_, _20305_, _15081_);
  nor (_20309_, _20308_, _20307_);
  nand (_20310_, _20309_, _20302_);
  nor (_20311_, _20102_, _20248_);
  nor (_20312_, _20249_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_20313_, _20312_, _20311_);
  nand (_20314_, _20313_, _15089_);
  nor (_20315_, _20246_, _20104_);
  nor (_20316_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_20317_, _15256_, _15077_);
  nor (_20318_, _20317_, _20316_);
  not (_20319_, _20318_);
  nand (_20320_, _20319_, _20315_);
  not (_20321_, _20315_);
  nand (_20322_, _20318_, _20321_);
  nand (_20323_, _20322_, _20320_);
  nor (_20324_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nor (_20325_, _15264_, _15085_);
  nor (_20326_, _20325_, _20324_);
  not (_20327_, _20326_);
  nand (_20328_, _20327_, _20303_);
  not (_20329_, _20303_);
  nand (_20330_, _20326_, _20329_);
  nand (_20331_, _20330_, _20328_);
  nor (_20332_, _20331_, _20323_);
  nand (_20333_, _20332_, _20314_);
  nor (_20334_, _20333_, _20310_);
  nand (_20335_, _20334_, _20271_);
  not (_20336_, _20311_);
  nor (_20337_, _20336_, _15278_);
  nor (_20338_, _20337_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_20339_, _20338_, _20270_);
  not (_20340_, _20339_);
  nand (_20341_, _20340_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_20342_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_20343_, _15278_, _15093_);
  nor (_20344_, _20343_, _20342_);
  not (_20345_, _20344_);
  nand (_20346_, _20345_, _20311_);
  nand (_20347_, _20344_, _20336_);
  nand (_20348_, _20347_, _20346_);
  not (_20349_, _20313_);
  nand (_20350_, _20349_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_20351_, _20289_, _15248_);
  nor (_20352_, _20351_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_20353_, _20352_, _20315_);
  nand (_20354_, _20353_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  not (_20355_, _20353_);
  nand (_20356_, _20355_, _15072_);
  nand (_20357_, _20356_, _20354_);
  nand (_20358_, _20357_, _20350_);
  nor (_20359_, _20358_, _20348_);
  nand (_20360_, _20359_, _20341_);
  nor (_20361_, _20360_, _20335_);
  nor (_20362_, _20338_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_20363_, _20362_, _20133_);
  nor (_20364_, _20363_, _20270_);
  nor (_20365_, _20261_, _20258_);
  nor (_20366_, _20365_, _20364_);
  nand (_20367_, _20366_, _20361_);
  nor (_20368_, _20367_, _20269_);
  nand (_20370_, _20368_, _20267_);
  not (_20371_, _19988_);
  nor (_20372_, _19995_, _20371_);
  not (_20373_, _19860_);
  nand (_20374_, _20373_, _19944_);
  nor (_20375_, _20085_, _19769_);
  nor (_20376_, _20375_, _19812_);
  not (_20377_, _20376_);
  nand (_20378_, _20377_, _19985_);
  nand (_20379_, _20378_, _20374_);
  nor (_20380_, _20379_, _20372_);
  nand (_20381_, _20380_, _20094_);
  nor (_20382_, _20090_, _19986_);
  nor (_20383_, _20382_, _20094_);
  nand (_20384_, _20090_, _19944_);
  nand (_20385_, _19860_, _19991_);
  nand (_20386_, _20385_, _20384_);
  nand (_20387_, _20386_, _20383_);
  nand (_20388_, _20387_, _20381_);
  nor (_20389_, _20085_, _19860_);
  nand (_20390_, _20389_, _19991_);
  nand (_20391_, _20390_, _20388_);
  nand (_20392_, _20391_, _20039_);
  not (_20393_, _20039_);
  not (_20394_, _19995_);
  nand (_20395_, _20394_, _19944_);
  nand (_20396_, _20395_, _20094_);
  nand (_20397_, _20394_, _19857_);
  nand (_20398_, _20084_, _19812_);
  nand (_20399_, _20398_, _20397_);
  not (_20400_, _20389_);
  nand (_20401_, _19986_, _20375_);
  not (_20402_, _20401_);
  nand (_20403_, _20402_, _19944_);
  nand (_20404_, _20403_, _20400_);
  nor (_20405_, _20404_, _20399_);
  nand (_20406_, _20405_, _20383_);
  nand (_20407_, _20406_, _20396_);
  nand (_20408_, _20407_, _19997_);
  nand (_20409_, _20408_, _20393_);
  nand (_20410_, _20409_, _20392_);
  nand (_20411_, _20410_, _20370_);
  nand (_20412_, _19812_, _19991_);
  nand (_20413_, _19857_, _19768_);
  nor (_20414_, _19993_, _19858_);
  nand (_20415_, _20414_, _19987_);
  nand (_20416_, _20415_, _20413_);
  nand (_20417_, _20416_, _19991_);
  nand (_20418_, _20417_, _20376_);
  nand (_20419_, _20418_, _20094_);
  nand (_20420_, _20419_, _20412_);
  nand (_20421_, _20420_, _20393_);
  nand (_20422_, _19858_, _19811_);
  nor (_20423_, _20422_, _19901_);
  nor (_20424_, _20413_, _19812_);
  nor (_20425_, _20424_, _20423_);
  nor (_20426_, _20425_, _20393_);
  nor (_20427_, _19991_, _20393_);
  nand (_20428_, _20422_, _20427_);
  nand (_20429_, _20428_, _20378_);
  nor (_20430_, _20429_, _20426_);
  nor (_20431_, _20430_, _20094_);
  nor (_20432_, _19812_, _19944_);
  nand (_20433_, _20432_, _20402_);
  nor (_20434_, _19995_, _19986_);
  not (_20435_, _20427_);
  nand (_20436_, _19857_, _19991_);
  nand (_20437_, _20436_, _20435_);
  nand (_20438_, _20437_, _20434_);
  nor (_20439_, _20371_, _19992_);
  nor (_20440_, _20439_, _20088_);
  nand (_20441_, _20440_, _20438_);
  nand (_20442_, _20441_, _20094_);
  nand (_20443_, _20442_, _20433_);
  nor (_20444_, _20443_, _20431_);
  nand (_20445_, _20444_, _20421_);
  nor (_20446_, _20258_, _15124_);
  not (_20447_, _20446_);
  nand (_20448_, _20255_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_20449_, _20448_, _15290_);
  nand (_20450_, _20449_, _15106_);
  nand (_20451_, _20450_, _20262_);
  nand (_20452_, _20451_, _20447_);
  nor (_20453_, _19719_, _19755_);
  not (_20454_, _20453_);
  nor (_20455_, _20454_, _20106_);
  not (_20456_, _20455_);
  nor (_20457_, _20456_, _20117_);
  not (_20458_, _20457_);
  nor (_20459_, _20458_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_20460_, _20457_, _15282_);
  nor (_20461_, _20460_, _20459_);
  nand (_20462_, _20461_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_20463_, _20461_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nor (_20464_, _20456_, _15260_);
  nor (_20465_, _20455_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_20466_, _20465_, _20464_);
  nand (_20467_, _20466_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  not (_20468_, _20466_);
  nand (_20469_, _20468_, _15081_);
  nand (_20471_, _20469_, _20467_);
  nor (_20472_, _20454_, _20104_);
  nor (_20473_, _20472_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_20474_, _20473_, _20455_);
  not (_20475_, _20474_);
  nor (_20476_, _20475_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_20477_, _20474_, _15077_);
  nor (_20478_, _20477_, _20476_);
  nand (_20479_, _20478_, _20471_);
  nor (_20480_, _20479_, _20463_);
  nand (_20481_, _20480_, _20462_);
  nand (_20482_, _20261_, _15106_);
  nand (_20483_, _20482_, _20446_);
  nor (_20484_, _20449_, _15106_);
  nor (_20485_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20486_, _20456_, _20102_);
  nor (_20487_, _20486_, _20485_);
  not (_20488_, _20487_);
  nor (_20489_, _20488_, _20312_);
  nor (_20490_, _20489_, _15089_);
  not (_20491_, _20489_);
  nor (_20492_, _20491_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_20493_, _20492_, _20490_);
  nand (_20494_, _20453_, _20103_);
  nand (_20495_, _20494_, _15252_);
  not (_20496_, _20495_);
  nor (_20497_, _20496_, _20472_);
  not (_20498_, _20497_);
  nor (_20499_, _20498_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_20500_, _20497_, _15072_);
  nor (_20501_, _20500_, _20499_);
  nand (_20502_, _20501_, _20493_);
  nand (_20503_, _20464_, _20327_);
  not (_20504_, _20464_);
  nand (_20505_, _20504_, _20326_);
  nand (_20506_, _20505_, _20503_);
  nor (_20507_, _20273_, _15124_);
  nor (_20508_, _19719_, _15132_);
  nor (_20509_, _20508_, _15136_);
  nor (_20510_, _20509_, _20507_);
  not (_20511_, _20510_);
  nor (_20512_, _20511_, _15052_);
  nand (_20513_, _20511_, _15052_);
  nor (_20514_, _20453_, _20189_);
  nand (_20515_, _20453_, _20189_);
  nand (_20516_, _20515_, _20188_);
  nor (_20517_, _20516_, _20514_);
  nand (_20518_, _20517_, _20513_);
  nor (_20519_, _20518_, _20512_);
  nor (_20520_, _20454_, _15238_);
  nor (_20521_, _20520_, _20154_);
  nor (_20522_, _20288_, _15124_);
  nor (_20523_, _20522_, _20521_);
  nor (_20524_, _19718_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_20525_, _20524_, _20508_);
  not (_20526_, _20525_);
  nand (_20527_, _20526_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_20528_, _20526_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_20529_, _20528_, _20171_);
  nand (_20530_, _20529_, _20527_);
  nor (_20531_, _20530_, _20523_);
  nand (_20532_, _20531_, _20519_);
  nor (_20533_, _20532_, _20506_);
  nor (_20534_, _20486_, _15278_);
  not (_20535_, _20534_);
  nand (_20536_, _20486_, _15278_);
  nand (_20537_, _20536_, _20535_);
  nor (_20538_, _20537_, _15093_);
  not (_20539_, _20537_);
  nor (_20540_, _20539_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_20541_, _20540_, _20538_);
  nand (_20542_, _20541_, _20533_);
  nor (_20543_, _20542_, _20502_);
  nor (_20544_, _20254_, _15124_);
  nor (_20545_, _20544_, _20134_);
  nor (_20546_, _20271_, _15124_);
  nor (_20547_, _20546_, _20545_);
  nand (_20548_, _20547_, _20543_);
  nor (_20549_, _20548_, _20484_);
  nand (_20550_, _20549_, _20483_);
  nor (_20551_, _20550_, _20481_);
  nand (_20552_, _20551_, _20452_);
  nand (_20553_, _20552_, _20445_);
  nand (_20554_, _20553_, _20411_);
  nor (_20555_, _20554_, _20244_);
  nor (_20556_, _15048_, _15041_);
  not (_20557_, _20556_);
  nor (_20558_, _20557_, _15037_);
  nor (_20559_, _20558_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_20560_, _20558_);
  nor (_20561_, _20560_, _15052_);
  nor (_20562_, _20561_, _20559_);
  nor (_20563_, _20562_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_20564_, _15041_, _15037_);
  nor (_20565_, _20564_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_20566_, _20565_, _20558_);
  nand (_20567_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _06097_);
  nand (_20568_, _20567_, _20566_);
  nor (_20569_, _20568_, _20563_);
  nor (_20570_, _20562_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_20571_, _20566_);
  nand (_20572_, _20562_, _06101_);
  nand (_20573_, _20572_, _20571_);
  nor (_20574_, _20573_, _20570_);
  nor (_20575_, _20574_, _20569_);
  nand (_20576_, _20575_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_20577_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _06226_);
  nor (_20578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_20579_, _20578_, _20557_);
  nand (_20580_, _20579_, _20577_);
  nor (_20581_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _06395_);
  not (_20582_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_20583_, _15052_, _20582_);
  nor (_20584_, _20583_, _20581_);
  not (_20585_, _20584_);
  nor (_20586_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2], _15041_);
  nand (_20587_, _20586_, _20585_);
  nand (_20588_, _20587_, _20580_);
  nor (_20589_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_20590_, _20589_, _15048_);
  nor (_20591_, _20590_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_20592_, _20590_);
  nor (_20593_, _20592_, _15052_);
  nor (_20594_, _20593_, _20591_);
  nand (_20595_, _20594_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand (_20596_, _20589_, _15048_);
  nand (_20597_, _20596_, _20592_);
  nor (_20598_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _06103_);
  nor (_20599_, _20598_, _20597_);
  nand (_20600_, _20599_, _20595_);
  nand (_20601_, _20600_, _15041_);
  not (_20602_, _20594_);
  nor (_20603_, _20602_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_20604_, _20594_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_20605_, _20604_, _20603_);
  not (_20606_, _20597_);
  nor (_20607_, _20606_, _20605_);
  nor (_20608_, _20607_, _20601_);
  nor (_20609_, _20608_, _20588_);
  nand (_20610_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_20611_, _15052_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nand (_20612_, _20611_, _20610_);
  nand (_20613_, _20612_, _15048_);
  nor (_20614_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _06747_);
  not (_20615_, _20614_);
  nand (_20616_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  nand (_20617_, _20616_, _20615_);
  nand (_20618_, _20617_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_20619_, _20618_, _20613_);
  nand (_20620_, _20619_, _15041_);
  nor (_20621_, _15052_, _07201_);
  nor (_20622_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _06245_);
  nor (_20623_, _20622_, _15048_);
  not (_20624_, _20623_);
  nor (_20625_, _20624_, _20621_);
  nor (_20626_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_20627_, _15052_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_20628_, _20627_, _20626_);
  nor (_20629_, _20628_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_20630_, _20629_, _20625_);
  nand (_20631_, _20630_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_20632_, _20631_, _20620_);
  nand (_20633_, _20632_, _15037_);
  nand (_20634_, _20617_, _20586_);
  nand (_20635_, _15052_, _06065_);
  nor (_20636_, _15052_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_20637_, _20636_, _20557_);
  nand (_20638_, _20637_, _20635_);
  nand (_20639_, _20638_, _20634_);
  not (_20640_, _20630_);
  nor (_20641_, _20640_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_20642_, _20641_, _20639_);
  nor (_20643_, _20642_, _20633_);
  nor (_20644_, _20562_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nand (_20645_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _20582_);
  nand (_20646_, _20566_, _20645_);
  nor (_20647_, _20646_, _20644_);
  nor (_20648_, _20562_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand (_20649_, _20562_, _06045_);
  nand (_20650_, _20649_, _20571_);
  nor (_20651_, _20650_, _20648_);
  nor (_20652_, _20651_, _20647_);
  nand (_20653_, _20652_, _15041_);
  nand (_20654_, _20653_, _20643_);
  nor (_20655_, _20654_, _20609_);
  nand (_20656_, _20655_, _20576_);
  nor (_20657_, _20594_, _06056_);
  nor (_20658_, _20602_, _06065_);
  nor (_20659_, _20658_, _20657_);
  nand (_20660_, _20659_, _20597_);
  nand (_20661_, _20594_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nand (_20662_, _20661_, _20606_);
  nor (_20663_, _20662_, _20614_);
  nor (_20664_, _20663_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_20665_, _20664_, _20660_);
  nand (_20666_, _20594_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_20667_, _20622_, _20597_);
  nand (_20668_, _20667_, _20666_);
  nand (_20669_, _20602_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_20670_, _20594_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand (_20671_, _20670_, _20669_);
  nor (_20672_, _20671_, _20606_);
  nor (_20673_, _20672_, _15041_);
  nand (_20674_, _20673_, _20668_);
  nand (_20675_, _20674_, _20665_);
  nor (_20676_, _20562_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_20677_, _15052_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_20678_, _20677_, _20676_);
  nor (_20679_, _20678_, _20571_);
  not (_20680_, _20562_);
  nor (_20681_, _20680_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_20682_, _20562_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_20683_, _20682_, _20681_);
  nor (_20684_, _20683_, _20566_);
  nor (_20685_, _20684_, _20679_);
  nor (_20686_, _20685_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_20687_, _20562_, _06065_);
  nor (_20688_, _20562_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_20689_, _20688_, _20566_);
  nand (_20690_, _20689_, _20687_);
  nor (_20691_, _20562_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nand (_20692_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _07043_);
  nand (_20693_, _20692_, _20566_);
  nor (_20694_, _20693_, _20691_);
  nor (_20695_, _20694_, _15041_);
  nand (_20696_, _20695_, _20690_);
  not (_20697_, _20564_);
  nand (_20698_, _15052_, _06103_);
  nand (_20699_, _20698_, _20567_);
  nand (_20700_, _20699_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_20701_, _15052_, _06095_);
  nand (_20702_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _06101_);
  nand (_20703_, _20702_, _20701_);
  nand (_20704_, _20703_, _15048_);
  nand (_20705_, _20704_, _20700_);
  nor (_20706_, _20705_, _20697_);
  nand (_20707_, _15041_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nand (_20708_, _20584_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_20709_, _15052_, _06226_);
  nand (_20710_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _06045_);
  nand (_20711_, _20710_, _20709_);
  nand (_20712_, _20711_, _15048_);
  nand (_20713_, _20712_, _20708_);
  nor (_20714_, _20713_, _20707_);
  nor (_20715_, _20714_, _20706_);
  nor (_20716_, _20705_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_20717_, _20716_, _20588_);
  nor (_20718_, _20717_, _20715_);
  nand (_20719_, _20718_, _20696_);
  nor (_20720_, _20719_, _20686_);
  nand (_20721_, _20720_, _20675_);
  nand (_20722_, _20721_, _20656_);
  nand (_20723_, _20510_, _06395_);
  nor (_20724_, _20510_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_20725_, _20724_, _20526_);
  nand (_20726_, _20725_, _20723_);
  nand (_20727_, _20510_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand (_20728_, _20511_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nand (_20729_, _20728_, _20727_);
  nand (_20730_, _20729_, _20526_);
  nand (_20731_, _20730_, _20726_);
  nand (_20732_, _20731_, _19725_);
  nand (_20733_, _20510_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nand (_20734_, _20511_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nand (_20735_, _20734_, _20733_);
  nand (_20736_, _20735_, _20525_);
  nand (_20737_, _20510_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_20738_, _20511_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand (_20739_, _20738_, _20737_);
  nand (_20740_, _20739_, _20526_);
  nand (_20741_, _20740_, _20736_);
  nand (_20742_, _20741_, _19722_);
  nand (_20743_, _20742_, _20732_);
  nand (_20744_, _20510_, _06747_);
  nor (_20745_, _20510_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_20746_, _20745_, _20526_);
  nand (_20747_, _20746_, _20744_);
  nand (_20748_, _20510_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nand (_20749_, _20511_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_20750_, _20749_, _20748_);
  nand (_20751_, _20750_, _20526_);
  nand (_20752_, _20751_, _20747_);
  nand (_20753_, _20752_, _19718_);
  nand (_20754_, _20510_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand (_20755_, _20511_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand (_20756_, _20755_, _20754_);
  nand (_20757_, _20756_, _20525_);
  nand (_20758_, _20510_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand (_20759_, _20511_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nand (_20760_, _20759_, _20758_);
  nand (_20761_, _20760_, _20526_);
  nand (_20762_, _20761_, _20757_);
  nand (_20763_, _20762_, _19715_);
  nand (_20764_, _20763_, _20753_);
  nor (_20765_, _20764_, _20743_);
  nor (_20766_, _20161_, _06045_);
  nor (_20767_, _20160_, _06226_);
  nor (_20768_, _20767_, _20766_);
  nor (_20769_, _20768_, _19716_);
  nor (_20770_, _20769_, _20174_);
  nor (_20771_, _20161_, _06082_);
  nor (_20772_, _20160_, _06084_);
  nor (_20773_, _20772_, _20771_);
  nor (_20774_, _20773_, _19719_);
  nand (_20775_, _20160_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nand (_20776_, _20161_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand (_20777_, _20776_, _20775_);
  nand (_20778_, _20777_, _19725_);
  nand (_20779_, _20160_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_20780_, _20161_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nand (_20781_, _20780_, _20779_);
  nand (_20782_, _20781_, _19722_);
  nand (_20783_, _20782_, _20778_);
  nor (_20784_, _20783_, _20774_);
  nand (_20785_, _20784_, _20770_);
  nand (_20786_, _20160_, _20582_);
  nor (_20787_, _19716_, _19703_);
  nand (_20788_, _20787_, _20786_);
  nand (_20789_, _20788_, _20174_);
  nand (_20790_, _20160_, _07201_);
  nor (_20791_, _19719_, _19667_);
  nand (_20792_, _20791_, _20790_);
  nor (_20793_, _20160_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_20794_, _19686_);
  nand (_20795_, _19725_, _20794_);
  nor (_20796_, _20795_, _20793_);
  nor (_20797_, _20160_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not (_20798_, _19661_);
  nand (_20799_, _19722_, _20798_);
  nor (_20800_, _20799_, _20797_);
  nor (_20801_, _20800_, _20796_);
  nand (_20802_, _20801_, _20792_);
  nor (_20803_, _20802_, _20789_);
  nand (_20804_, _20245_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_20805_, _20273_, _06045_);
  nor (_20806_, _19706_, _20294_);
  nor (_20807_, _20806_, _20805_);
  nand (_20808_, _20807_, _20804_);
  nand (_20809_, _20808_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_20810_, _19726_, _19676_);
  nand (_20811_, _19722_, _19694_);
  nand (_20812_, _19715_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nand (_20813_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _06056_);
  nand (_20814_, _15136_, _06065_);
  nand (_20815_, _20814_, _20813_);
  nor (_20816_, _20815_, _20812_);
  not (_20817_, _19663_);
  nand (_20818_, _20293_, _15124_);
  nor (_20819_, _20818_, _20817_);
  nor (_20820_, _20819_, _20816_);
  nand (_20821_, _20820_, _20811_);
  nor (_20822_, _20821_, _20810_);
  nand (_20823_, _20822_, _20809_);
  not (_20824_, first_instr);
  nand (_20825_, _08692_, _20824_);
  nor (_20826_, _20825_, _19714_);
  nand (_20827_, _20826_, _20823_);
  nor (_20828_, _20827_, _20803_);
  nand (_20829_, _20828_, _20785_);
  nor (_20830_, _20829_, _20765_);
  nand (_20831_, _20830_, _20722_);
  nor (property_invalid, _20831_, _20555_);
  nor (_20832_, _24380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1]);
  nor (_20833_, _24382_, _21474_);
  nor (_25291_, _20833_, _20832_);
  nor (_20834_, _22838_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5]);
  nor (_20835_, _22840_, _21451_);
  nor (_25067_, _20835_, _20834_);
  nor (_20836_, _22561_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1]);
  nor (_20837_, _22563_, _21474_);
  nor (_25075_, _20837_, _20836_);
  nor (_20838_, _23025_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0]);
  nor (_20839_, _23027_, _21586_);
  nor (_25117_, _20839_, _20838_);
  nor (_20840_, _24380_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0]);
  nor (_20841_, _24382_, _21586_);
  nor (_25290_, _20841_, _20840_);
  nor (_20842_, _21752_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6]);
  nor (_20843_, _21754_, _21504_);
  nor (_25237_, _20843_, _20842_);
  nor (_20844_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand (_20845_, _23553_, _00599_);
  nand (_20846_, _20845_, _23493_);
  nor (_25042_[0], _20846_, _20844_);
  nor (_20847_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand (_20848_, _23553_, _23257_);
  nand (_20849_, _20848_, _23493_);
  nor (_25042_[1], _20849_, _20847_);
  nor (_20850_, _21741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4]);
  nor (_20851_, _21744_, _21414_);
  nor (_25241_, _20851_, _20850_);
  nor (_20852_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand (_20853_, _23553_, _23215_);
  nand (_20854_, _20853_, _23493_);
  nor (_25042_[2], _20854_, _20852_);
  nor (_20855_, _00880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3]);
  nor (_20856_, _00882_, _21526_);
  nor (_25287_, _20856_, _20855_);
  nor (_20857_, _23553_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand (_20858_, _23553_, _23188_);
  nand (_20859_, _20858_, _23493_);
  nor (_25042_[3], _20859_, _20857_);
  nor (_20860_, _22470_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1]);
  nor (_20861_, _22473_, _21474_);
  nor (_25079_, _20861_, _20860_);
  nor (_20862_, _21741_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5]);
  nor (_20863_, _21744_, _21451_);
  nor (_25242_, _20863_, _20862_);
  nor (_09412_, rst, _05924_);
  nor (_20864_, _00880_, \oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5]);
  nor (_20865_, _00882_, _21451_);
  nor (_25288_, _20865_, _20864_);
  dff (first_instr, _00000_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _25011_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _25011_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _25011_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _25011_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _25011_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _25011_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _25011_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _25011_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _24989_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _24990_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _24991_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _24992_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _24993_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _24994_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _24995_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _24996_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _25009_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _25009_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _25009_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _25009_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _25009_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _25009_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _25009_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _25009_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _24997_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _24998_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _24999_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _25000_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _25001_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _25002_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _25003_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _25004_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _25010_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _25010_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _25010_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _25010_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _25010_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _25010_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _25010_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _25010_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _25005_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _25005_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _25005_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _25005_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _25005_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _25005_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _25005_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _25005_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _24973_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _24974_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _24975_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _24976_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _24977_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _24978_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _24979_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _24980_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _24965_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _24966_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _24967_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _24968_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _24969_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _24970_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _24971_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _24972_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _25015_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _25015_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _25015_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _25015_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _25015_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _25015_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _25015_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _25015_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _25014_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _25014_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _25014_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _25014_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _25014_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _25014_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _25014_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _25014_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _24964_[0]);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _24964_[1]);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _24964_[2]);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _24964_[3]);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _24964_[4]);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _24964_[5]);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _24964_[6]);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _24964_[7]);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _24964_[8]);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _24964_[9]);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _24964_[10]);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _24964_[11]);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _24964_[12]);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _24964_[13]);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _24964_[14]);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _24964_[15]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _25006_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _25006_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _25006_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _25006_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _25006_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _25006_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _25006_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _25006_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _25007_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _25007_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _25007_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _25007_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _25007_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _25007_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _25007_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _25007_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _25008_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _25008_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _25008_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _25008_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _25008_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _25008_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _25008_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _25008_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _24981_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _24982_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _24983_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _24984_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _24985_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _24986_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _24987_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _24988_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _25013_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _25013_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _25013_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _25013_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _25013_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _25013_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _25013_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _25013_[7]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _25012_[0]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _25012_[1]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _25012_[2]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _25012_[3]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _25012_[4]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _25012_[5]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _25012_[6]);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _25012_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _25016_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _25016_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _25016_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _25017_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _25017_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _25017_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _25018_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _25018_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _25019_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _25019_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _25019_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _25019_[3]);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _25019_[4]);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _25019_[5]);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _25019_[6]);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _25019_[7]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _25020_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _25020_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _25021_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _25021_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _25021_[2]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _25022_[0]);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _25022_[1]);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _25023_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _03778_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _03782_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _03789_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _03791_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _03797_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _03800_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _03801_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _23357_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _03813_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _03816_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _03818_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _03820_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _25024_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _25024_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _25024_[6]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _23361_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _03859_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _03861_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _03863_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _03865_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _25025_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _25025_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _03873_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _23363_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _25026_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _03892_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _03901_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _03904_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _03906_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _03908_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _03911_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _23380_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _03928_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _03930_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _25027_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _03936_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _03938_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _03941_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _03943_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _23390_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _25028_[0]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _25028_[1]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _03962_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _03964_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _03967_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _03969_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _03971_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _25028_[7]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _04008_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _04013_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _04016_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _04019_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _04021_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _25029_[5]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _04031_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _23395_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _04054_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _04056_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _25030_[2]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _04059_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _25030_[4]);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _04068_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _04077_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _23401_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _07730_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _07757_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _07781_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _07783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _05527_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _08345_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _25031_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _08356_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _08358_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _08360_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _25031_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _25031_[6]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _08377_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _08379_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _08381_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _08384_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _08386_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _08388_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _25031_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _25031_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _00735_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08440_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _08443_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _08445_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08447_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _25032_[4]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _08514_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _08516_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _08518_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _08520_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _08522_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _08537_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _08550_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _25032_[12]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _25032_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _25032_[14]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _00758_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _25042_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _25042_[1]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _25042_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _25042_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _23916_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _22400_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _21062_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _05685_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _05022_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _04276_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _10326_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _25042_[11]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _21170_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _25042_[13]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _18004_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _19174_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _21099_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _21211_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _21387_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _21765_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _21896_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _21908_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _21916_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _22177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _25042_[24]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _22247_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _22518_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _25042_[27]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _25042_[28]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _25042_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _25042_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _25042_[31]);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _05495_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _08151_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _08206_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _08268_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _08274_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _08348_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _25033_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _08464_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _05538_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _08717_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _08808_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [2], _25038_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _08822_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _08856_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _08875_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _08956_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [7], _05552_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], _08952_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _22589_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _25039_[2]);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _02018_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _18025_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _21087_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], _21124_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _05576_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _05689_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _06432_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _06435_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _06441_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _06453_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _06456_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _06459_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _06463_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _25034_[7]);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _06467_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _06470_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _06472_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _06475_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _06478_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _06484_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _06488_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _05750_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _06518_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _06521_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _06523_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _06525_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _06528_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _06532_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _06537_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _06542_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _06545_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _06548_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _06550_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _06552_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _06554_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _06559_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _06560_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _05752_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _05757_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _05759_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _25035_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _06580_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _06584_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _06586_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _08689_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _08833_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _25036_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _08995_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _05761_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _25037_[0]);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _08992_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _05769_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], _05570_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _05780_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _06402_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _06389_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _06386_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _25040_[3]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _06380_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _25040_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _06374_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _05782_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _05783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _25041_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _06357_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _06354_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _06350_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _05833_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _06288_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _06285_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _06282_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _06279_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _06276_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _25043_[5]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _06266_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _06251_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _06248_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _06242_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _06239_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _06236_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _06233_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _06224_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _06221_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _25043_[15]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _06208_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _06205_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _06201_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _06198_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _06179_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _25043_[21]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _06174_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _25043_[23]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _06161_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _06158_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _06152_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _06146_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _06132_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _25043_[29]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _25043_[30]);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _05867_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _05880_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _05882_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _05884_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _05973_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _05969_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _05965_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _05963_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _05888_);
  dff (\oc8051_top_1.oc8051_ram_top1.rd_en_r , _20959_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [0], _25044_[0]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [1], _21143_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [2], _21144_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [3], _21149_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [4], _25044_[4]);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [5], _21153_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [6], _21154_);
  dff (\oc8051_top_1.oc8051_ram_top1.wr_data_r [7], _20960_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_addr_r , _20961_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [0], _21159_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [1], _21161_);
  dff (\oc8051_top_1.oc8051_ram_top1.bit_select [2], _20963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [0], _23291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [1], _23252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [2], _02282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [3], _08947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [4], _22788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [5], _25336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [6], _22774_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[255] [7], _02277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [0], _23314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [1], _23336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [2], _23344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [3], _23340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [4], _21065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [5], _23089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [6], _23053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[254] [7], _02285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [0], _23446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [1], _23437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [2], _25334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [3], _25335_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [4], _23533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [5], _23526_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [6], _04011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[253] [7], _23311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [0], _21069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [1], _03699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [2], _23550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [3], _23548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [4], _04028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [5], _23724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [6], _23703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[252] [7], _04025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [0], _24001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [1], _23988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [2], _04039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [3], _25332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [4], _25333_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [5], _04036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [6], _23765_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[251] [7], _23762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [0], _24037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [1], _04047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [2], _25329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [3], _25330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [4], _04050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [5], _21140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [6], _23787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[250] [7], _25331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [0], _21167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [1], _24124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [2], _24116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [3], _24114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [4], _24139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [5], _24141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [6], _21075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[249] [7], _24056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [0], _24237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [1], _04074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [2], _24262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [3], _04071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [4], _25324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [5], _24182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [6], _25325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[248] [7], _25326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [0], _25320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [1], _24285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [2], _24281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [3], _24321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [4], _25321_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [5], _24311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [6], _25322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[247] [7], _25323_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [0], _03707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [1], _24354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [2], _25319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [3], _24341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [4], _24371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [5], _24377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [6], _24374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[246] [7], _21070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [0], _09005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [1], _25315_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [2], _24418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [3], _24415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [4], _25316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [5], _25317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [6], _25318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[245] [7], _04093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [0], _25309_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [1], _25310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [2], _21151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [3], _25311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [4], _04100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [5], _25312_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [6], _25313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[244] [7], _25314_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [0], _24639_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [1], _24334_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [2], _25303_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [3], _25304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [4], _25305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [5], _25306_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [6], _25307_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[243] [7], _25308_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [0], _24658_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [1], _00289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [2], _00065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [3], _05695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [4], _25300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [5], _25301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [6], _24388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[242] [7], _25302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [0], _00679_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [1], _00614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [2], _25299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [3], _01512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [4], _01440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [5], _05697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [6], _24656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[241] [7], _24660_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [0], _05893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [1], _01903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [2], _02425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [3], _25298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [4], _03637_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [5], _03501_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [6], _08831_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[240] [7], _00846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [0], _21828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [1], _05207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [2], _05196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [3], _25296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [4], _03713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [5], _04227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [6], _04144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[239] [7], _25297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [0], _02273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [1], _24806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [2], _05621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [3], _25295_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [4], _05776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [5], _05692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [6], _23071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[238] [7], _04984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [0], _03274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [1], _06799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [2], _06795_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [3], _06788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [4], _05877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [5], _06602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [6], _06190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[237] [7], _06665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [0], _21043_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [1], _08919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [2], _01332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [3], _22345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [4], _25294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [5], _08914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [6], _06749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[236] [7], _06744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [0], _25290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [1], _25291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [2], _25292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [3], _09056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [4], _06722_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [5], _25293_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [6], _21023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[235] [7], _20882_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [0], _09077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [1], _05139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [2], _08897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [3], _25287_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [4], _21025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [5], _25288_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [6], _23605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[234] [7], _25289_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [0], _07060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [1], _07050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [2], _06828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [3], _25285_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [4], _03360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [5], _06953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [6], _06944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[233] [7], _25286_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [0], _07078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [1], _07080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [2], _25284_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [3], _07137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [4], _07152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [5], _06987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [6], _07007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[232] [7], _06989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [0], _07360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [1], _08217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [2], _07186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [3], _25282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [4], _07196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [5], _25283_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [6], _07269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[231] [7], _07242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [0], _08367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [1], _21145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [2], _07394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [3], _07933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [4], _07434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [5], _08089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [6], _25281_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[230] [7], _07317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [0], _21103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [1], _25278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [2], _07538_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [3], _07625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [4], _08585_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [5], _07456_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [6], _07453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[229] [7], _07989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [0], _22720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [1], _07837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [2], _07828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [3], _06496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [4], _07895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [5], _21162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [6], _07702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[228] [7], _23024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [0], _25276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [1], _08220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [2], _05268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [3], _07986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [4], _07930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [5], _07967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [6], _25277_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[227] [7], _08030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [0], _25273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [1], _25274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [2], _23820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [3], _08512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [4], _08482_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [5], _25275_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [6], _08570_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[226] [7], _22575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [0], _25271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [1], _08872_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [2], _07818_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [3], _22985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [4], _25272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [5], _23780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [6], _08799_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[225] [7], _23483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [0], _06997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [1], _02853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [2], _03119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [3], _03183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [4], _03465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [5], _08242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [6], _03545_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[224] [7], _00635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [0], _25269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [1], _07190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [2], _01008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [3], _00012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [4], _01019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [5], _25270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [6], _01567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[223] [7], _02629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [0], _25264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [1], _23494_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [2], _07486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [3], _25265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [4], _00215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [5], _25266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [6], _25267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[222] [7], _25268_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [0], _24338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [1], _24339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [2], _02301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [3], _10116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [4], _25261_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [5], _25262_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [6], _06677_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[221] [7], _25263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [0], _25260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [1], _03003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [2], _23712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [3], _02651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [4], _24047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [5], _22384_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [6], _24228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[220] [7], _02483_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [0], _22580_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [1], _22597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [2], _03577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [3], _25259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [4], _22643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [5], _22888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [6], _10367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[219] [7], _22906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [0], _10576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [1], _25255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [2], _22375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [3], _25256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [4], _25257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [5], _21018_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [6], _22472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[218] [7], _25258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [0], _21457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [1], _06469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [2], _09726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [3], _21460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [4], _21463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [5], _21471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [6], _21489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[217] [7], _24106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [0], _22129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [1], _04410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [2], _22157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [3], _22254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [4], _21091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [5], _08929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [6], _11258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[216] [7], _25254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [0], _22154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [1], _21886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [2], _04956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [3], _21898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [4], _21909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [5], _21415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [6], _09148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[215] [7], _21941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [0], _09528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [1], _21522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [2], _21527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [3], _21539_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [4], _22554_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [5], _21543_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [6], _25253_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[214] [7], _10441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [0], _02342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [1], _25251_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [2], _21492_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [3], _21509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [4], _23633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [5], _21516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [6], _23451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[213] [7], _25252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [0], _21408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [1], _21399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [2], _03690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [3], _04141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [4], _03846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [5], _21053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [6], _25249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[212] [7], _25250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [0], _06779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [1], _22079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [2], _20962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [3], _05890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [4], _05214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [5], _25247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [6], _06623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[211] [7], _25248_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [0], _07652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [1], _25246_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [2], _07598_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [3], _22057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [4], _06737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [5], _06728_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [6], _06717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[210] [7], _06867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [0], _07714_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [1], _07712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [2], _07922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [3], _07916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [4], _13311_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [5], _21031_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [6], _07504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[209] [7], _07205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [0], _13642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [1], _25243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [2], _08301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [3], _08236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [4], _09101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [5], _25244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [6], _08817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[208] [7], _22001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [0], _24664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [1], _25240_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [2], _00102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [3], _13930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [4], _25241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [5], _25242_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [6], _21171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[207] [7], _20877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [0], _21924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [1], _25239_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [2], _06656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [3], _21901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [4], _20964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [5], _22522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [6], _22185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[206] [7], _22163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [0], _07863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [1], _07790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [2], _21879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [3], _08473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [4], _25238_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [5], _14445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [6], _04753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[205] [7], _04697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [0], _25235_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [1], _08868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [2], _08829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [3], _21840_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [4], _25236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [5], _00396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [6], _25237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[204] [7], _14712_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [0], _06438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [1], _21751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [2], _20979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [3], _22218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [4], _21936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [5], _21204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [6], _00082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[203] [7], _02270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [0], _06480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [1], _06515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [2], _06503_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [3], _06500_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [4], _15202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [5], _19279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [6], _18089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[202] [7], _25234_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [0], _06540_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [1], _06530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [2], _25232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [3], _06567_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [4], _25233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [5], _21696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [6], _20987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[201] [7], _06486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [0], _21033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [1], _21068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [2], _06588_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [3], _06582_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [4], _21680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [5], _08986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [6], _08988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[200] [7], _21665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [0], _06360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [1], _06369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [2], _15777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [3], _06697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [4], _25227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [5], _06422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [6], _06713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[199] [7], _21624_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [0], _06340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [1], _21575_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [2], _06331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [3], _25225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [4], _06318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [5], _21556_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [6], _25226_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[198] [7], _06408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [0], _21036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [1], _06305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [2], _06296_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [3], _06299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [4], _06273_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [5], _06263_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [6], _06269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[197] [7], _21535_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [0], _21470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [1], _06216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [2], _06210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [3], _06213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [4], _06154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [5], _06134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [6], _06149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[196] [7], _21513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [0], _06030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [1], _06032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [2], _21416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [3], _20992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [4], _06113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [5], _06107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [6], _06110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[195] [7], _06088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [0], _05984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [1], _05986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [2], _21369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [3], _06058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [4], _06049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [5], _25223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [6], _25224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[194] [7], _06025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [0], _05941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [1], _05948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [2], _21317_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [3], _21001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [4], _21064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [5], _06012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [6], _25222_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[193] [7], _06004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [0], _05902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [1], _25220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [2], _05906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [3], _17169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [4], _05972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [5], _25221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [6], _05967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[192] [7], _05939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [0], _01349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [1], _01343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [2], _21265_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [3], _01225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [4], _25219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [5], _01221_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [6], _17464_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[191] [7], _05919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [0], _25217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [1], _18078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [2], _21040_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [3], _22469_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [4], _22480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [5], _25218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [6], _22391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[190] [7], _21182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [0], _21054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [1], _21060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [2], _21180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [3], _21035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [4], _21037_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [5], _25214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [6], _21120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[189] [7], _21181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [0], _15614_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [1], _25212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [2], _18979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [3], _21024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [4], _21026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [5], _20974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [6], _20978_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[188] [7], _25213_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [0], _21097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [1], _05399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [2], _25211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [3], _21098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [4], _21027_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [5], _21066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [6], _20892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[187] [7], _21177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [0], _03219_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [1], _21092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [2], _25210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [3], _03505_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [4], _03533_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [5], _21095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [6], _21094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[186] [7], _21029_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [0], _21088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [1], _25209_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [2], _02605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [3], _20947_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [4], _03110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [5], _02832_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [6], _21090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[185] [7], _21030_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [0], _14320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [1], _21173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [2], _23778_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [3], _23814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [4], _19290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [5], _02460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [6], _02504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[184] [7], _02643_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [0], _23576_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [1], _23463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [2], _23559_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [3], _22746_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [4], _22445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [5], _25207_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [6], _19578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[183] [7], _25208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [0], _21082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [1], _21079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [2], _25160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [3], _21055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [4], _25161_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [5], _25162_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [6], _25163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[165] [7], _00792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [0], _01785_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [1], _01772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [2], _25164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [3], _25165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [4], _00001_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [5], _01730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [6], _25166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[166] [7], _25167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [0], _01579_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [1], _25168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [2], _01569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [3], _00457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [4], _00823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [5], _20928_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [6], _25169_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[167] [7], _20906_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [0], _20893_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [1], _25170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [2], _20889_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [3], _00278_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [4], _20872_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [5], _25171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [6], _20871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[168] [7], _00257_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [0], _25172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [1], _25173_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [2], _00236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [3], _00776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [4], _25174_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [5], _18522_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [6], _25175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[169] [7], _18264_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [0], _18131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [1], _25176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [2], _25177_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [3], _07695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [4], _09126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [5], _25178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [6], _25179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[170] [7], _25180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [0], _25181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [1], _00571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [2], _00854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [3], _05613_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [4], _21113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [5], _25182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [6], _03478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[171] [7], _25183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [0], _25184_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [1], _25185_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [2], _20972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [3], _08454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [4], _25186_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [5], _11410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [6], _25187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[172] [7], _25188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [0], _00530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [1], _22171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [2], _25189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [3], _25190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [4], _00087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [5], _05937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [6], _06090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[173] [7], _25191_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [0], _06416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [1], _25192_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [2], _25193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [3], _25194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [4], _06707_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [5], _08990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [6], _25195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[174] [7], _00509_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [0], _25196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [1], _21781_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [2], _22112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [3], _05421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [4], _05423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [5], _20923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [6], _25197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[175] [7], _22814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [0], _00061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [1], _00166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [2], _25198_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [3], _04693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [4], _20909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [5], _21114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [6], _21117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[176] [7], _25199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [0], _20898_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [1], _06070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [2], _06044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [3], _21118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [4], _25200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [5], _20894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [6], _05943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[177] [7], _06023_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [0], _05993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [1], _21119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [2], _21022_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [3], _21128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [4], _08010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [5], _04467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [6], _20879_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[178] [7], _08194_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [0], _08021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [1], _25201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [2], _21021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [3], _08866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [4], _21133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [5], _25202_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [6], _21132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[179] [7], _21107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [0], _21137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [1], _21115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [2], _23267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [3], _20866_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [4], _25204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [5], _21139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [6], _21110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[180] [7], _21138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [0], _22755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [1], _04541_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [2], _22729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [3], _25205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [4], _20470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [5], _03467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [6], _21096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[181] [7], _02243_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [0], _02279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [1], _05426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [2], _20168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [3], _20953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [4], _21032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [5], _04932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [6], _20973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[182] [7], _25206_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [0], _10779_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [1], _21157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [2], _01474_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [3], _25153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [4], _01472_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [5], _00436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [6], _23886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[162] [7], _23706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [0], _00414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [1], _25154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [2], _25155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [3], _23656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [4], _00392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [5], _23649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [6], _22944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[163] [7], _25156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [0], _00807_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [1], _21158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [2], _21105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [3], _25157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [4], _21093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [5], _25158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [6], _25159_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[164] [7], _00330_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [0], _10666_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [1], _11157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [2], _23417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [3], _10590_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [4], _06399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [5], _07664_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [6], _00787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[161] [7], _10757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [0], _08656_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [1], _08790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [2], _04397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [3], _25152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [4], _11041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [5], _10894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [6], _10912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[160] [7], _24772_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [0], _03448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [1], _08407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [2], _03422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [3], _08455_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [4], _04422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [5], _08549_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [6], _25149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[159] [7], _25150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [0], _07999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [1], _03578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [2], _08057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [3], _08144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [4], _03520_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [5], _08188_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [6], _25148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[158] [7], _03487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [0], _03671_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [1], _07717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [2], _03645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [3], _07760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [4], _25146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [5], _07848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [6], _25147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[157] [7], _03612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [0], _25143_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [1], _25144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [2], _04569_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [3], _07444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [4], _03725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [5], _07487_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [6], _04548_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[156] [7], _25145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [0], _03877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [1], _07017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [2], _25141_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [3], _07055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [4], _07150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [5], _03815_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [6], _07199_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[155] [7], _25142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [0], _03987_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [1], _06565_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [2], _04689_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [3], _06649_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [4], _06801_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [5], _03949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [6], _06899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[154] [7], _03920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [0], _25138_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [1], _04341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [2], _25139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [3], _04871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [4], _05410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [5], _05466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [6], _04298_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[153] [7], _25140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [0], _25136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [1], _04024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [2], _25137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [3], _05249_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [4], _04376_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [5], _05271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [6], _04890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[152] [7], _05200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [0], _06105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [1], _04130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [2], _06157_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [3], _04747_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [4], _06259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [5], _04083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [6], _06301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[151] [7], _04725_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [0], _04816_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [1], _25133_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [2], _05916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [3], _25134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [4], _25135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [5], _05980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [6], _04164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[150] [7], _05999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [0], _25129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [1], _04837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [2], _25130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [3], _05705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [4], _04244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [5], _05039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [6], _05739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[149] [7], _25131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [0], _25126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [1], _25127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [2], _25128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [3], _04090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [4], _21625_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [5], _10652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [6], _11142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[148] [7], _05504_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [0], _21038_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [1], _21019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [2], _25123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [3], _21156_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [4], _11228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [5], _25124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [6], _10631_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[147] [7], _25125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [0], _01788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [1], _11057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [2], _21061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [3], _20896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [4], _19577_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [5], _10849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [6], _20914_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[146] [7], _25122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [0], _25120_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [1], _03210_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [2], _01751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [3], _11010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [4], _09923_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [5], _25121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [6], _10974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[145] [7], _07732_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [0], _25117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [1], _25118_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [2], _25119_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [3], _02050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [4], _08820_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [5], _07302_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [6], _08486_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[144] [7], _08758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [0], _07460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [1], _06764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [2], _06790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [3], _06917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [4], _00951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [5], _04993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [6], _22530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[143] [7], _24787_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [0], _02355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [1], _05089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [2], _05149_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [3], _25116_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [4], _00419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [5], _00630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [6], _08527_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[142] [7], _07155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [0], _21179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [1], _01024_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [2], _22610_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [3], _23406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [4], _24270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [5], _08490_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [6], _25114_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[141] [7], _25115_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [0], _08702_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [1], _08015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [2], _25113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [3], _08344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [4], _02378_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [5], _03130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [6], _08427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[140] [7], _21447_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [0], _25111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [1], _04845_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [2], _08292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [3], _05106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [4], _08276_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [5], _08247_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [6], _07096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[139] [7], _25112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [0], _08910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [1], _08507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [2], _08212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [3], _25110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [4], _07853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [5], _07743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [6], _01082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[138] [7], _02842_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [0], _02417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [1], _08052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [2], _08068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [3], _08168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [4], _08147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [5], _08272_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [6], _08086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[137] [7], _01109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [0], _08528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [1], _08498_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [2], _01155_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [3], _08175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [4], _08233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [5], _08215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [6], _25108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[136] [7], _25109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [0], _08652_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [1], _25106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [2], _01180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [3], _25107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [4], _08410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [5], _08394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [6], _08337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[135] [7], _08471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [0], _08851_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [1], _08965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [2], _25103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [3], _08954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [4], _25104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [5], _25105_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [6], _08609_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[134] [7], _07956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [0], _25101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [1], _08034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [2], _08007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [3], _07822_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [4], _25102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [5], _07959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [6], _01232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[133] [7], _08756_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [0], _25099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [1], _03091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [2], _08438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [3], _25100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [4], _08197_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [5], _07739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [6], _08450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[132] [7], _08324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [0], _08566_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [1], _08668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [2], _25096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [3], _08484_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [4], _25097_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [5], _08373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [6], _25098_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[131] [7], _08607_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [0], _07423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [1], _08665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [2], _08620_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [3], _07557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [4], _25094_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [5], _07506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [6], _25095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[130] [7], _08705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [0], _01368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [1], _02894_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [2], _25091_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [3], _08853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [4], _08825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [5], _07466_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [6], _08761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[129] [7], _25092_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [0], _08922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [1], _25089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [2], _08836_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [3], _08748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [4], _08827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [5], _07391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [6], _25090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[128] [7], _08958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [0], _24093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [1], _25087_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [2], _22687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [3], _25088_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [4], _01399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [5], _08886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [6], _08938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[127] [7], _08935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [0], _25085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [1], _21017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [2], _25086_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [3], _22405_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [4], _01339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [5], _21121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [6], _01421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[126] [7], _06813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [0], _06053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [1], _21888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [2], _21890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [3], _22244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [4], _07070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [5], _25083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [6], _03113_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[125] [7], _25084_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [0], _02571_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [1], _21228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [2], _21108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [3], _21299_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [4], _07036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [5], _24259_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [6], _06998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[124] [7], _06127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [0], _22715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [1], _01511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [2], _23453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [3], _04371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [4], _25080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [5], _25081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [6], _25082_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[123] [7], _22777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [0], _22742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [1], _25079_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [2], _01544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [3], _02916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [4], _08967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [5], _01744_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [6], _08650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[122] [7], _21405_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [0], _02592_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [1], _25075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [2], _06726_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [3], _06594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [4], _25076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [5], _06672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [6], _25077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[121] [7], _25078_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [0], _25074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [1], _21705_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [2], _06511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [3], _20943_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [4], _21676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [5], _06632_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [6], _23325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[120] [7], _21650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [0], _25072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [1], _02123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [2], _21063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [3], _05480_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [4], _05451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [5], _02742_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [6], _03187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[119] [7], _21755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [0], _05359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [1], _25070_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [2], _05327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [3], _21034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [4], _25071_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [5], _14465_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [6], _05392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[118] [7], _02764_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [0], _03310_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [1], _05292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [2], _02791_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [3], _05036_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [4], _04979_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [5], _09008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [6], _21076_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[117] [7], _02266_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [0], _01695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [1], _06383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [2], _02608_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [3], _03140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [4], _03212_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [5], _04537_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [6], _04291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[116] [7], _02233_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [0], _21127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [1], _05414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [2], _23136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [3], _01684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [4], _22880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [5], _09107_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [6], _25068_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[115] [7], _25069_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [0], _05956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [1], _06046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [2], _06324_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [3], _02970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [4], _20977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [5], _01717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [6], _05444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[114] [7], _06121_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [0], _23033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [1], _01763_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [2], _04681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [3], _12953_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [4], _07014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [5], _21172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [6], _04771_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[113] [7], _06232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [0], _23260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [1], _21122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [2], _25066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [3], _21089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [4], _23699_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [5], _25067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [6], _06182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[112] [7], _23158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [0], _25065_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [1], _08657_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [2], _05959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [3], _23322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [4], _22419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [5], _21131_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [6], _21630_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[111] [7], _01827_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [0], _05491_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [1], _05896_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [2], _05875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [3], _08680_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [4], _05936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [5], _25064_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [6], _01870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[110] [7], _08599_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [0], _05792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [1], _22618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [2], _25059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [3], _08331_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [4], _04865_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [5], _25060_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [6], _24347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[109] [7], _01935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [0], _05618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [1], _25057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [2], _05720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [3], _02452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [4], _05683_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [5], _02695_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [6], _25058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[108] [7], _24099_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [0], _25056_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [1], _22753_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [2], _23530_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [3], _05578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [4], _02721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [5], _07642_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [6], _05662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[107] [7], _10241_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [0], _01968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [1], _02089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [2], _11290_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [3], _12623_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [4], _12932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [5], _20369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [6], _05542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[106] [7], _23962_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [0], _25052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [1], _01478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [2], _01600_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [3], _25053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [4], _12644_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [5], _25054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [6], _01849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[105] [7], _25055_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [0], _11446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [1], _01126_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [2], _11432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [3], _01270_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [4], _12269_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [5], _12828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [6], _01313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[104] [7], _01443_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [0], _00729_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [1], _11515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [2], _00761_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [3], _11497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [4], _00838_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [5], _25051_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [6], _00972_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[103] [7], _11460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [0], _00488_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [1], _11602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [2], _00612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [3], _11583_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [4], _00636_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [5], _12340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [6], _25050_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[102] [7], _00700_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [0], _00140_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [1], _00172_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [2], _11665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [3], _00193_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [4], _25049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [5], _00214_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [6], _12378_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[101] [7], _00351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [0], _25045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [1], _11740_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [2], _25046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [3], _12450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [4], _25047_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [5], _00109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [6], _25048_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[100] [7], _12717_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [0], _12911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [1], _25448_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [2], _11797_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [3], _25449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [4], _12470_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [5], _25450_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [6], _25451_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[99] [7], _11757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [0], _12168_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [1], _21595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [2], _12117_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [3], _21713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [4], _12581_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [5], _21730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [6], _21862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[98] [7], _12075_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [0], _11828_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [1], _25446_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [2], _12485_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [3], _12869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [4], _21436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [5], _12147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [6], _25447_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[97] [7], _12602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [0], _23665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [1], _11909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [2], _25443_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [3], _12513_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [4], _25444_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [5], _11869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [6], _25445_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[96] [7], _12499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [0], _11971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [1], _22662_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [2], _25441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [3], _22704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [4], _25442_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [5], _12890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [6], _22913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[95] [7], _23254_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [0], _22017_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [1], _12033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [2], _22033_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [3], _12012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [4], _22095_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [5], _12557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [6], _25439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[94] [7], _25440_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [0], _25436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [1], _20873_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [2], _25437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [3], _02260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [4], _02267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [5], _20880_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [6], _02255_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[93] [7], _25438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [0], _20875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [1], _25434_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [2], _02220_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [3], _02077_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [4], _02083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [5], _20867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [6], _25435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[92] [7], _02227_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [0], _14546_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [1], _20887_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [2], _20891_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [3], _20885_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [4], _20869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [5], _25432_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [6], _25433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[91] [7], _20876_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [0], _19216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [1], _14627_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [2], _19237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [3], _15292_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [4], _19301_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [5], _25430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [6], _19452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[90] [7], _25431_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [0], _18854_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [1], _14720_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [2], _18916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [3], _14704_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [4], _18958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [5], _15337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [6], _19072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[89] [7], _25429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [0], _15400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [1], _18471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [2], _18605_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [3], _25427_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [4], _18629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [5], _18711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [6], _14739_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[88] [7], _25428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [0], _18152_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [1], _14819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [2], _15736_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [3], _18183_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [4], _18326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [5], _14800_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [6], _18347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[87] [7], _18430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [0], _17840_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [1], _14883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [2], _17871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [3], _15481_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [4], _25426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [5], _18067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [6], _14844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[86] [7], _18110_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [0], _17515_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [1], _17599_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [2], _25424_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [3], _17650_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [4], _25425_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [5], _14909_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [6], _17777_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[85] [7], _17819_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [0], _16011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [1], _25423_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [2], _16154_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [3], _16224_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [4], _15165_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [5], _16291_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [6], _15144_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[84] [7], _16318_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [0], _15573_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [1], _17180_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [2], _17232_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [3], _17258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [4], _25421_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [5], _25422_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [6], _16074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[83] [7], _16135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [0], _15042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [1], _16867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [2], _15788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [3], _16908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [4], _17013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [5], _15020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [6], _17085_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[82] [7], _15003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [0], _16443_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [1], _25420_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [2], _16519_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [3], _16601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [4], _16693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [5], _15074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [6], _16724_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[81] [7], _15635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [0], _02297_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [1], _02294_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [2], _02339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [3], _02336_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [4], _02329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [5], _25418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [6], _25419_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[80] [7], _16384_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [0], _25415_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [1], _25416_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [2], _25417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [3], _02364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [4], _02409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [5], _02406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [6], _02401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[79] [7], _20878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [0], _02052_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [1], _02044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [2], _20870_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [3], _02109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [4], _02103_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [5], _02090_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [6], _02074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[78] [7], _02428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [0], _20884_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [1], _02147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [2], _02145_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [3], _02139_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [4], _02179_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [5], _02170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [6], _02166_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[77] [7], _20868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [0], _02477_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [1], _02463_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [2], _02457_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [3], _20890_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [4], _25413_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [5], _02566_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [6], _25414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[76] [7], _02593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [0], _13878_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [1], _02506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [2], _20888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [3], _02531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [4], _02528_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [5], _20886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [6], _02441_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[75] [7], _02438_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [0], _04792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [1], _04635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [2], _13005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [3], _21146_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [4], _25411_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [5], _25412_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [6], _02396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[74] [7], _02200_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [0], _05218_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [1], _19393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [2], _05640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [3], _05524_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [4], _25410_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [5], _02949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [6], _03163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[73] [7], _03016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [0], _07780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [1], _13057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [2], _06204_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [3], _25408_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [4], _06035_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [5], _25409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [6], _06776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[72] [7], _19322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [0], _08905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [1], _09578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [2], _19195_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [3], _07371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [4], _07237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [5], _07223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [6], _07181_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[71] [7], _07913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [0], _11073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [1], _11025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [2], _10995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [3], _19153_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [4], _11366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [5], _11417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [6], _08383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[70] [7], _25407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [0], _18980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [1], _13949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [2], _12096_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [3], _12054_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [4], _11930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [5], _12696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [6], _12665_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[69] [7], _12529_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [0], _14868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [1], _18895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [2], _13108_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [3], _13026_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [4], _12974_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [5], _19021_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [6], _13622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[68] [7], _25404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [0], _16053_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [1], _15959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [2], _18833_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [3], _13976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [4], _14252_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [5], _14124_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [6], _18937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[67] [7], _25403_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [0], _16404_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [1], _18792_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [2], _16971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [3], _16950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [4], _25401_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [5], _13189_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [6], _15502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[66] [7], _25402_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [0], _17557_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [1], _17393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [2], _25399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [3], _17983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [4], _17892_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [5], _18690_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [6], _25400_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[65] [7], _16478_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [0], _20874_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [1], _18587_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [2], _18368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [3], _18305_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [4], _18659_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [5], _19258_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [6], _25398_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[64] [7], _18645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [0], _20883_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [1], _20881_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [2], _25396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [3], _20903_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [4], _20895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [5], _25397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [6], _19837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[63] [7], _19806_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [0], _20965_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [1], _13250_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [2], _20925_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [3], _25393_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [4], _25394_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [5], _25395_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [6], _18409_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[62] [7], _14341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [0], _21002_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [1], _25390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [2], _21015_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [3], _25391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [4], _25392_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [5], _20955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [6], _20952_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[61] [7], _20950_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [0], _21041_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [1], _21039_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [2], _21028_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [3], _21020_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [4], _21049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [5], _25388_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [6], _21044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[60] [7], _25389_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [0], _13353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [1], _21059_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [2], _21058_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [3], _21057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [4], _25387_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [5], _21073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [6], _21067_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[59] [7], _13332_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [0], _18046_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [1], _14074_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [2], _21083_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [3], _21081_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [4], _21080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [5], _21102_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [6], _21101_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[58] [7], _21100_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [0], _21135_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [1], _21134_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [2], _25386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [3], _21104_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [4], _21106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [5], _21109_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [6], _21112_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[57] [7], _21111_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [0], _21163_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [1], _21160_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [2], _13391_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [3], _21130_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [4], _21129_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [5], _21125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [6], _21123_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[56] [7], _21136_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [0], _21178_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [1], _21176_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [2], _21225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [3], _21201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [4], _13414_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [5], _21148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [6], _21147_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[55] [7], _21164_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [0], _25385_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [1], _21402_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [2], _21326_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [3], _21633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [4], _21628_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [5], _21594_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [6], _13437_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[54] [7], _21175_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [0], _22089_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [1], _13467_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [2], _21721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [3], _21710_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [4], _25383_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [5], _17798_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [6], _21770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[53] [7], _25384_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [0], _22237_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [1], _25380_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [2], _25381_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [3], _22267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [4], _17681_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [5], _25382_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [6], _21921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[52] [7], _17752_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [0], _17536_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [1], _22552_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [2], _25379_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [3], _22350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [4], _22340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [5], _22436_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [6], _22433_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[51] [7], _17578_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [0], _01735_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [1], _16271_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [2], _25377_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [3], _01673_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [4], _25378_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [5], _13760_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [6], _14428_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[50] [7], _22460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [0], _01877_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [1], _01908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [2], _01886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [3], _13810_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [4], _16244_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [5], _25375_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [6], _01835_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[49] [7], _13790_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [0], _01938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [1], _01955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [2], _25373_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [3], _02012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [4], _25374_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [5], _16032_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [6], _02025_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[48] [7], _15990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [0], _22691_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [1], _25371_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [2], _22809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [3], _22748_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [4], _22737_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [5], _13516_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [6], _01977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[47] [7], _25372_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [0], _22964_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [1], _13555_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [2], _22859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [3], _22850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [4], _22868_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [5], _22875_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [6], _22871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[46] [7], _22711_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [0], _25369_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [1], _25370_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [2], _23093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [3], _17211_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [4], _22916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [5], _22935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [6], _22926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[45] [7], _22959_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [0], _23171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [1], _23142_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [2], _17158_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [3], _23196_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [4], _23205_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [5], _17137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [6], _14171_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[44] [7], _23019_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [0], _17034_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [1], _25368_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [2], _16992_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [3], _14190_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [4], _23274_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [5], _17106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [6], _23399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[43] [7], _13602_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [0], _23635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [1], _13653_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [2], _14386_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [3], _23506_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [4], _23511_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [5], _25367_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [6], _16929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[42] [7], _23439_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [0], _23715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [1], _25366_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [2], _14225_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [3], _23645_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [4], _16846_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [5], _16825_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [6], _23621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[41] [7], _23618_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [0], _23823_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [1], _23773_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [2], _23804_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [3], _25364_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [4], _23869_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [5], _16672_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [6], _25365_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[40] [7], _23688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [0], _01454_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [1], _25359_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [2], _01507_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [3], _01497_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [4], _16550_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [5], _25360_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [6], _25361_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[39] [7], _25362_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [0], _02435_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [1], _01595_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [2], _01648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [3], _01621_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [4], _13730_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [5], _01542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [6], _01572_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[38] [7], _25358_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [0], _20900_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [1], _20935_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [2], _02872_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [3], _02886_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [4], _20899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [5], _02888_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [6], _02911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[37] [7], _20897_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [0], _02857_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [1], _20930_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [2], _25357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [3], _02859_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [4], _02863_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [5], _20902_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [6], _02867_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[36] [7], _20901_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [0], _20905_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [1], _25355_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [2], _25356_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [3], _02844_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [4], _20904_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [5], _02847_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [6], _20931_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[35] [7], _02850_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [0], _02829_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [1], _02834_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [2], _20908_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [3], _20936_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [4], _25354_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [5], _20907_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [6], _02837_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[34] [7], _20932_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [0], _20911_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [1], _25352_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [2], _02809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [3], _25353_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [4], _20937_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [5], _02812_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [6], _02817_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[33] [7], _20910_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [0], _20915_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [1], _02793_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [2], _25350_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [3], _02796_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [4], _25351_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [5], _20913_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [6], _02802_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[32] [7], _20912_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [0], _02661_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [1], _20942_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [2], _02776_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [3], _02783_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [4], _20917_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [5], _02786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [6], _20916_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[31] [7], _02788_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [0], _20938_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [1], _02668_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [2], _20929_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [3], _25348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [4], _20934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [5], _25349_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [6], _02676_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[30] [7], _20933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [0], _20920_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [1], _20939_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [2], _02755_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [3], _25346_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [4], _20919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [5], _02767_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [6], _20918_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[29] [7], _02770_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [0], _02716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [1], _20922_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [2], _20940_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [3], _25343_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [4], _02733_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [5], _20921_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [6], _25344_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[28] [7], _25345_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [0], _02692_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [1], _02697_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [2], _20926_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [3], _20941_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [4], _02703_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [5], _02706_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [6], _20924_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[27] [7], _02713_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [0], _05429_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [1], _25338_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [2], _25339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [3], _25340_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [4], _25341_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [5], _25342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [6], _02688_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[26] [7], _20927_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [0], _03014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [1], _03005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [2], _21016_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [3], _02622_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [4], _02617_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [5], _02934_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [6], _25337_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[25] [7], _02919_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [0], _03049_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [1], _03045_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [2], _25327_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [3], _25328_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [4], _03072_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [5], _20944_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [6], _02977_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[24] [7], _02971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [0], _03201_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [1], _20945_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [2], _03127_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [3], _03122_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [4], _03150_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [5], _03148_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [6], _03137_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[23] [7], _03057_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [0], _03267_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [1], _03260_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [2], _03256_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [3], _20946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [4], _25279_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [5], _03167_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [6], _25280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[22] [7], _03208_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [0], _03282_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [1], _03329_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [2], _03325_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [3], _03320_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [4], _21014_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [5], _20966_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [6], _03223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[21] [7], _03231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [0], _25245_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [1], _03356_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [2], _03397_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [3], _03390_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [4], _03387_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [5], _21013_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [6], _03304_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[20] [7], _03300_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [0], _20949_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [1], _03426_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [2], _03418_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [3], _03460_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [4], _25228_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [5], _03473_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [6], _20948_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[19] [7], _20975_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [0], _21012_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [1], _20967_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [2], _03547_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [3], _03542_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [4], _03531_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [5], _03561_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [6], _25215_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[18] [7], _25216_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [0], _03663_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [1], _25203_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [2], _21011_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [3], _03597_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [4], _03606_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [5], _03601_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [6], _03640_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[17] [7], _03634_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [0], _03684_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [1], _21010_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [2], _03696_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [3], _03693_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [4], _20951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [5], _20976_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [6], _03651_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[16] [7], _03647_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [0], _21008_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [1], _20968_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [2], _03716_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [3], _03715_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [4], _25151_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [5], _03762_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [6], _03757_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[15] [7], _03749_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [0], _03853_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [1], _03848_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [2], _21007_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [3], _03871_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [4], _25132_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [5], _03786_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [6], _03780_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[14] [7], _21009_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [0], _03973_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [1], _21004_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [2], _03895_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [3], _03899_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [4], _21006_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [5], _03933_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [6], _21005_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[13] [7], _20969_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [0], _04044_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [1], _04042_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [2], _20954_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [3], _03957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [4], _03955_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [5], _03951_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [6], _03946_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[12] [7], _25093_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [0], _04066_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [1], _04128_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [2], _04125_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [3], _04106_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [4], _21003_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [5], _03983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [6], _03991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[11] [7], _25073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [0], _25061_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [1], _04170_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [2], _04187_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [3], _04182_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [4], _25062_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [5], _20956_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [6], _25063_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[10] [7], _04080_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [0], _04217_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [1], _04236_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [2], _04223_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [3], _21000_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [4], _25452_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [5], _25453_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [6], _04280_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[9] [7], _20999_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [0], _04430_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [1], _20997_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [2], _04322_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [3], _04313_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [4], _20998_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [5], _04342_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [6], _04357_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[8] [7], _04348_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [0], _04449_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [1], _04443_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [2], _04489_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [3], _04471_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [4], _04462_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [5], _20957_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [6], _04399_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[7] [7], _04407_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [0], _20995_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [1], _20970_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [2], _04496_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [3], _04502_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [4], _04499_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [5], _25405_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [6], _04512_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[6] [7], _25406_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [0], _04593_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [1], _20994_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [2], _04616_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [3], _04612_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [4], _20993_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [5], _04544_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [6], _04534_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[5] [7], _20996_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [0], _04701_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [1], _20990_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [2], _04633_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [3], _04629_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [4], _20991_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [5], _04648_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [6], _25376_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[4] [7], _20958_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [0], _04731_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [1], _04721_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [2], _04719_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [3], _04758_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [4], _25363_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [5], _04751_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [6], _20989_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[3] [7], _04687_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [0], _20982_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [1], _05417_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [2], _20981_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [3], _20980_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [4], _04794_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [5], _25347_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [6], _04809_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[2] [7], _04813_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [0], _25229_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [1], _20985_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [2], _05339_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [3], _25230_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [4], _20986_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [5], _05319_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [6], _05316_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[1] [7], _25231_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [0], _04849_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [1], _20988_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [2], _20971_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [3], _05396_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [4], _20984_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [5], _05402_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [6], _20983_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.buff[0] [7], _05352_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0], _08862_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1], _25454_[1]);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2], _08814_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3], _08635_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4], _08963_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5], _21743_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6], _06073_);
  dff (\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7], _21116_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _22304_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _01701_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _01761_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _25455_[2]);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _25455_[3]);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _08843_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _22309_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _05494_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _05510_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _05515_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _05514_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _05518_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _05525_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _05523_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _05354_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _03430_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _03438_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _03444_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _03441_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _03457_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _03453_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _03470_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _09090_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _09412_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _08691_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _08734_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _08662_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _08730_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _08699_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _08614_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _08678_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _22979_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _08534_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _23281_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _06724_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _08589_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _08476_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _06730_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _08983_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _08452_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _06732_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _08363_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _08425_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _07550_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _07517_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _07560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _23270_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _08203_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _08155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _08285_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _06921_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _08244_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _08279_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _08163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _08146_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _08266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _08050_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _07948_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _06930_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _07844_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _07961_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _08100_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _07840_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _07849_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _07876_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _07823_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _06965_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _22097_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _07420_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _07412_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _07415_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _22093_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _21927_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _21953_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _07886_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _21925_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _07282_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _07279_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _22104_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _07325_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _07321_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _07315_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _07865_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _07214_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _22110_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _07253_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _07250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _07247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _07245_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _22107_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _07851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _21918_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _21950_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _07094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _07092_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _07084_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _22120_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _07123_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _07835_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _05155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _05157_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _05167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _05163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _05165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _05172_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _04416_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _03875_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _03878_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _03880_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _03884_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _03882_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _03888_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _03887_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _03658_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _03655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _23674_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _23573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _21815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _21854_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _08754_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _08751_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _21813_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _08765_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _08763_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _23566_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _21809_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _21851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _08771_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _08768_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _21807_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _08775_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _08773_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _21746_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _23734_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _23731_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _21848_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _08782_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _08780_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _21803_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _08786_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _08784_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _21802_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _23720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _21845_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _08791_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _08789_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _21800_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _08795_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _08793_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _21797_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _21740_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _21715_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _21795_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _21841_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _08801_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _21793_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _08806_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _08804_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _23538_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _24323_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _24392_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _24358_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _24356_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _21072_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _05778_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _05763_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _21071_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _21046_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _21051_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _06681_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _21174_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _21047_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _21052_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _05141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _21074_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _05433_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _05416_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _05325_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _24040_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _24024_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _04198_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _04136_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _21078_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _21077_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _21045_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _03164_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _03114_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _24009_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _09011_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _08981_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _08977_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _21084_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _09064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _09061_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _09059_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _24007_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _23995_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _08971_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _08969_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _21085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _21042_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _21050_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _08930_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _08928_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _23986_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _21086_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _21126_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _22694_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _21166_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _05643_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _00044_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _08601_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _21048_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _08889_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _21165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _21833_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _06857_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _07521_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _07579_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _07574_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _07534_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _06863_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _06872_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _08950_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _06870_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _24846_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _24825_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _21155_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _06866_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _06855_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _06852_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _06832_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _06843_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _21142_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _21150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _01458_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _06840_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _21141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _04193_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _23866_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _23503_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _06662_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _21168_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _21912_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _21056_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _22727_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _22722_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _06837_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _06835_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _08877_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _08778_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _21169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _21152_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _08043_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _08032_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _08036_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _06808_);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.desOv , ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_sfr1.desAc , ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_sfr1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [0], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [0]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [1], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [1]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [2], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [2]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [3], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [3]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [4], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [4]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [5], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [5]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [6], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [6]);
  buf(\oc8051_top_1.oc8051_ram_top1.rd_data_m [7], \oc8051_top_1.oc8051_ram_top1.oc8051_idata.rd_data [7]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_ram_top1.wr_data [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_ram_top1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.bit_data_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_ram_top1.clk , clk);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_comp1.des [0], ABINPUT[27]);
  buf(\oc8051_top_1.oc8051_comp1.des [1], ABINPUT[28]);
  buf(\oc8051_top_1.oc8051_comp1.des [2], ABINPUT[29]);
  buf(\oc8051_top_1.oc8051_comp1.des [3], ABINPUT[30]);
  buf(\oc8051_top_1.oc8051_comp1.des [4], ABINPUT[31]);
  buf(\oc8051_top_1.oc8051_comp1.des [5], ABINPUT[32]);
  buf(\oc8051_top_1.oc8051_comp1.des [6], ABINPUT[33]);
  buf(\oc8051_top_1.oc8051_comp1.des [7], ABINPUT[34]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], \oc8051_top_1.oc8051_sfr1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [8], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [9], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [10], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [11], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [12], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [13], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [14], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.alu [15], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_memory_interface1.imm2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_memory_interface1.imm2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_memory_interface1.imm_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_memory_interface1.imm_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_memory_interface1.op3_buff [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.wr_dat [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_indi_addr1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.rst , rst);
  buf(\oc8051_top_1.oc8051_ram_top1.oc8051_idata.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data2_in [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.ov_in , ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.ac_in , ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.cy_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data2_in [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.sub_result [0], ABINPUT[27]);
  buf(\oc8051_top_1.sub_result [1], ABINPUT[28]);
  buf(\oc8051_top_1.sub_result [2], ABINPUT[29]);
  buf(\oc8051_top_1.sub_result [3], ABINPUT[30]);
  buf(\oc8051_top_1.sub_result [4], ABINPUT[31]);
  buf(\oc8051_top_1.sub_result [5], ABINPUT[32]);
  buf(\oc8051_top_1.sub_result [6], ABINPUT[33]);
  buf(\oc8051_top_1.sub_result [7], ABINPUT[34]);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.ABINPUT [9], ABINPUT[9]);
  buf(\oc8051_top_1.ABINPUT [10], ABINPUT[10]);
  buf(\oc8051_top_1.ABINPUT [11], ABINPUT[11]);
  buf(\oc8051_top_1.ABINPUT [12], ABINPUT[12]);
  buf(\oc8051_top_1.ABINPUT [13], ABINPUT[13]);
  buf(\oc8051_top_1.ABINPUT [14], ABINPUT[14]);
  buf(\oc8051_top_1.ABINPUT [15], ABINPUT[15]);
  buf(\oc8051_top_1.ABINPUT [16], ABINPUT[16]);
  buf(\oc8051_top_1.ABINPUT [17], ABINPUT[17]);
  buf(\oc8051_top_1.ABINPUT [18], ABINPUT[18]);
  buf(\oc8051_top_1.ABINPUT [19], ABINPUT[19]);
  buf(\oc8051_top_1.ABINPUT [20], ABINPUT[20]);
  buf(\oc8051_top_1.ABINPUT [21], ABINPUT[21]);
  buf(\oc8051_top_1.ABINPUT [22], ABINPUT[22]);
  buf(\oc8051_top_1.ABINPUT [23], ABINPUT[23]);
  buf(\oc8051_top_1.ABINPUT [24], ABINPUT[24]);
  buf(\oc8051_top_1.ABINPUT [25], ABINPUT[25]);
  buf(\oc8051_top_1.ABINPUT [26], ABINPUT[26]);
  buf(\oc8051_top_1.ABINPUT [27], ABINPUT[27]);
  buf(\oc8051_top_1.ABINPUT [28], ABINPUT[28]);
  buf(\oc8051_top_1.ABINPUT [29], ABINPUT[29]);
  buf(\oc8051_top_1.ABINPUT [30], ABINPUT[30]);
  buf(\oc8051_top_1.ABINPUT [31], ABINPUT[31]);
  buf(\oc8051_top_1.ABINPUT [32], ABINPUT[32]);
  buf(\oc8051_top_1.ABINPUT [33], ABINPUT[33]);
  buf(\oc8051_top_1.ABINPUT [34], ABINPUT[34]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.desOv , ABINPUT[2]);
  buf(\oc8051_top_1.desAc , ABINPUT[1]);
  buf(\oc8051_top_1.desCy , ABINPUT[0]);
  buf(\oc8051_top_1.des2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.des2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.des2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.des2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.des2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.des2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.des2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.des2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.des1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.des1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.des1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.des1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.des1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.des1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.des1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.des1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.des_acc [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.wr_dat [0], ABINPUT[3]);
  buf(\oc8051_top_1.wr_dat [1], ABINPUT[4]);
  buf(\oc8051_top_1.wr_dat [2], ABINPUT[5]);
  buf(\oc8051_top_1.wr_dat [3], ABINPUT[6]);
  buf(\oc8051_top_1.wr_dat [4], ABINPUT[7]);
  buf(\oc8051_top_1.wr_dat [5], ABINPUT[8]);
  buf(\oc8051_top_1.wr_dat [6], ABINPUT[9]);
  buf(\oc8051_top_1.wr_dat [7], ABINPUT[10]);
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], \oc8051_top_1.oc8051_sfr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], \oc8051_top_1.oc8051_sfr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], \oc8051_top_1.oc8051_sfr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], \oc8051_top_1.oc8051_sfr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], \oc8051_top_1.oc8051_sfr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], \oc8051_top_1.oc8051_sfr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], \oc8051_top_1.oc8051_sfr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.intr , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.data_in [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.wr_bit_r , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [0], ABINPUT[11]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [1], ABINPUT[12]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [2], ABINPUT[13]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [3], ABINPUT[14]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [4], ABINPUT[15]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [5], ABINPUT[16]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [6], ABINPUT[17]);
  buf(\oc8051_top_1.oc8051_sfr1.dat2 [7], ABINPUT[18]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [0], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [1], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [2], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [3], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [4], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [5], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [6], ABINPUT[9]);
  buf(\oc8051_top_1.oc8051_sfr1.dat1 [7], ABINPUT[10]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.des_acc [7], ABINPUT[26]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [0], ABINPUT[19]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [1], ABINPUT[20]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [2], ABINPUT[21]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [3], ABINPUT[22]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [4], ABINPUT[23]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [5], ABINPUT[24]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [6], ABINPUT[25]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_in [7], ABINPUT[26]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_ram_top1.bit_addr_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
