
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pcp1, property_invalid_pcp2, property_invalid_pcp3, property_invalid_sjmp, property_invalid_ljmp, property_invalid_ajmp, ABINPUT);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  input [8:0] ABINPUT;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid_ajmp;
  output property_invalid_ljmp;
  output property_invalid_pcp1;
  output property_invalid_pcp2;
  output property_invalid_pcp3;
  output property_invalid_sjmp;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  or (_06399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_06400_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_06401_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_06402_, _06401_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_06403_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_06404_, _06403_);
  not (_06405_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_06406_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06407_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _06406_);
  and (_06408_, _06407_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_06409_, _06408_, _06405_);
  not (_06410_, _06409_);
  nor (_06411_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_06412_, _06411_, _06410_);
  and (_06413_, _06412_, _06404_);
  not (_06414_, _06413_);
  not (_06415_, _06407_);
  and (_06416_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _06406_);
  and (_06417_, _06416_, _06415_);
  and (_06418_, _06417_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_06419_, _06418_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  and (_06420_, _06408_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_06421_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _06406_);
  nor (_06422_, _06421_, _06416_);
  and (_06423_, _06422_, _06407_);
  and (_06424_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  or (_06425_, _06424_, _06420_);
  nor (_06426_, _06425_, _06419_);
  and (_06427_, _06417_, _06405_);
  and (_06428_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nand (_06429_, _06422_, _06415_);
  not (_06430_, _06429_);
  and (_06431_, _06430_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_06432_, _06431_, _06428_);
  and (_06433_, _06432_, _06426_);
  and (_06434_, _06433_, _06414_);
  not (_06435_, _06402_);
  nor (_06436_, _06401_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_06437_, _06436_, _06410_);
  and (_06438_, _06437_, _06435_);
  not (_06439_, _06438_);
  and (_06440_, _06430_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and (_06441_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor (_06442_, _06441_, _06440_);
  and (_06443_, _06418_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_06444_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_06445_, _06444_, _06443_);
  and (_06446_, _06445_, _06442_);
  and (_06447_, _06446_, _06439_);
  not (_06448_, _06447_);
  and (_06449_, _06448_, _06434_);
  and (_06450_, _06403_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_06451_, _06450_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_06452_, _06451_);
  nor (_06453_, _06450_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_06454_, _06453_, _06410_);
  and (_06455_, _06454_, _06452_);
  not (_06456_, _06455_);
  and (_06457_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_06458_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  and (_06459_, _06418_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or (_06460_, _06459_, _06458_);
  or (_06461_, _06460_, _06420_);
  nor (_06462_, _06461_, _06457_);
  and (_06463_, _06462_, _06456_);
  not (_06464_, _06450_);
  nor (_06465_, _06403_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_06466_, _06465_, _06410_);
  and (_06467_, _06466_, _06464_);
  not (_06468_, _06467_);
  and (_06469_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  not (_06470_, _06469_);
  and (_06471_, _06418_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  not (_06472_, _06471_);
  and (_06473_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  nor (_06474_, _06473_, _06420_);
  and (_06475_, _06474_, _06472_);
  and (_06476_, _06475_, _06470_);
  and (_06477_, _06476_, _06468_);
  not (_06478_, _06477_);
  nor (_06479_, _06478_, _06463_);
  and (_06480_, _06479_, _06449_);
  and (_06481_, \oc8051_top_1.oc8051_decoder1.wr , _06406_);
  not (_06482_, _06481_);
  and (_06483_, _06407_, _06405_);
  nor (_06484_, _06483_, _06482_);
  and (_06485_, _06484_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not (_06486_, _06485_);
  not (_06487_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_06488_, _06451_, _06487_);
  and (_06489_, _06451_, _06487_);
  nor (_06490_, _06489_, _06488_);
  nor (_06491_, _06490_, _06410_);
  not (_06492_, _06491_);
  and (_06493_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and (_06494_, _06427_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_06495_, _06418_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  or (_06496_, _06495_, _06494_);
  or (_06497_, _06496_, _06420_);
  nor (_06498_, _06497_, _06493_);
  and (_06499_, _06498_, _06492_);
  nor (_06500_, _06499_, _06486_);
  and (_06501_, _06500_, _06480_);
  or (_06502_, _06501_, _06399_);
  and (_06503_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_06504_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_06505_, _06504_, _06503_);
  and (_06506_, _06418_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  not (_06507_, _06506_);
  not (_06508_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_06509_, _06409_, _06508_);
  and (_06510_, _06430_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_06511_, _06510_, _06509_);
  and (_06512_, _06511_, _06507_);
  and (_06513_, _06512_, _06505_);
  not (_06514_, _06513_);
  nor (_06515_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_06516_, _06515_, _06401_);
  and (_06517_, _06516_, _06409_);
  and (_06518_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_06519_, _06518_, _06517_);
  and (_06520_, _06418_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_06521_, _06427_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and (_06522_, _06430_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_06523_, _06522_, _06521_);
  nor (_06524_, _06523_, _06520_);
  and (_06525_, _06524_, _06519_);
  nor (_06526_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_06527_, _06526_, _06400_);
  and (_06528_, _06527_, _06409_);
  and (_06529_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_06530_, _06529_, _06528_);
  and (_06531_, _06418_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_06532_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_06533_, _06430_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_06534_, _06533_, _06532_);
  nor (_06535_, _06534_, _06531_);
  and (_06537_, _06535_, _06530_);
  nor (_06538_, _06537_, _06525_);
  and (_06539_, _06538_, _06514_);
  not (_06540_, _06539_);
  not (_06541_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_06543_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _06406_);
  and (_06544_, _06543_, _06541_);
  and (_06545_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _06406_);
  and (_06546_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _06406_);
  nor (_06547_, _06546_, _06545_);
  and (_06548_, _06547_, _06544_);
  not (_06549_, _06548_);
  not (_06550_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not (_06551_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_06552_, _06551_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_06553_, _06552_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_06554_, _06553_, _06550_);
  nor (_06555_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_06556_, _06555_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand (_06557_, _06556_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_06558_, _06557_, _06554_);
  not (_06559_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or (_06560_, _06552_, _06559_);
  not (_06561_, _06560_);
  nand (_06562_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_06563_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_06564_, _06563_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_06565_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_06566_, _06565_, _06562_);
  and (_06567_, _06566_, _06558_);
  and (_06568_, _06555_, _06551_);
  not (_06569_, _06568_);
  not (_06570_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_06572_, _06570_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or (_06573_, _06572_, ABINPUT[8]);
  nand (_06574_, _06570_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or (_06575_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_06576_, _06575_, _06573_);
  or (_06577_, _06576_, _06569_);
  and (_06578_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_06579_, _06578_, _06559_);
  nand (_06581_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_06582_, _06578_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_06583_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and (_06584_, _06583_, _06581_);
  and (_06585_, _06584_, _06577_);
  and (_06586_, _06585_, _06567_);
  nor (_06587_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not (_06588_, _06587_);
  or (_06589_, _06588_, _06576_);
  nand (_06590_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_06591_, _06590_, _06550_);
  not (_06592_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not (_06593_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_06594_, _06593_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_06595_, _06594_, _06592_);
  and (_06596_, _06595_, _06591_);
  and (_06597_, _06596_, _06589_);
  nor (_06598_, _06597_, _06586_);
  not (_06599_, _06598_);
  not (_06600_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  or (_06601_, _06553_, _06600_);
  nand (_06602_, _06556_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  and (_06603_, _06602_, _06601_);
  nand (_06604_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand (_06605_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_06606_, _06605_, _06604_);
  and (_06607_, _06606_, _06603_);
  or (_06608_, _06572_, ABINPUT[6]);
  or (_06609_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_06610_, _06609_, _06608_);
  or (_06611_, _06610_, _06569_);
  nand (_06612_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  nand (_06613_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_06614_, _06613_, _06612_);
  and (_06615_, _06614_, _06611_);
  nand (_06616_, _06615_, _06607_);
  or (_06617_, _06610_, _06588_);
  or (_06618_, _06590_, _06600_);
  not (_06619_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_06620_, _06594_, _06619_);
  and (_06621_, _06620_, _06618_);
  and (_06622_, _06621_, _06617_);
  not (_06623_, _06622_);
  and (_06624_, _06623_, _06616_);
  nor (_06625_, _06623_, _06616_);
  nor (_06627_, _06625_, _06624_);
  not (_06628_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  or (_06629_, _06553_, _06628_);
  nand (_06630_, _06556_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  and (_06631_, _06630_, _06629_);
  nand (_06632_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand (_06633_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_06634_, _06633_, _06632_);
  and (_06635_, _06634_, _06631_);
  or (_06636_, _06572_, ABINPUT[5]);
  or (_06637_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_06639_, _06637_, _06636_);
  or (_06640_, _06639_, _06569_);
  nand (_06642_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_06643_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and (_06644_, _06643_, _06642_);
  and (_06645_, _06644_, _06640_);
  and (_06646_, _06645_, _06635_);
  or (_06647_, _06639_, _06588_);
  or (_06648_, _06590_, _06628_);
  not (_06649_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_06650_, _06594_, _06649_);
  and (_06651_, _06650_, _06648_);
  and (_06652_, _06651_, _06647_);
  nor (_06653_, _06652_, _06646_);
  and (_06654_, _06652_, _06646_);
  nor (_06655_, _06654_, _06653_);
  nand (_06656_, _06556_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  not (_06657_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  or (_06658_, _06553_, _06657_);
  and (_06659_, _06658_, _06656_);
  nand (_06660_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand (_06661_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_06662_, _06661_, _06660_);
  and (_06663_, _06662_, _06659_);
  or (_06664_, _06572_, ABINPUT[4]);
  or (_06665_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_06666_, _06665_, _06664_);
  or (_06667_, _06666_, _06569_);
  nand (_06668_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand (_06669_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and (_06670_, _06669_, _06668_);
  and (_06672_, _06670_, _06667_);
  and (_06673_, _06672_, _06663_);
  or (_06675_, _06666_, _06588_);
  or (_06676_, _06590_, _06657_);
  not (_06677_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_06678_, _06594_, _06677_);
  and (_06679_, _06678_, _06676_);
  and (_06680_, _06679_, _06675_);
  nor (_06681_, _06680_, _06673_);
  and (_06682_, _06680_, _06673_);
  nor (_06683_, _06682_, _06681_);
  nand (_06684_, _06556_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  not (_06685_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_06686_, _06553_, _06685_);
  and (_06687_, _06686_, _06684_);
  nand (_06688_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nand (_06689_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_06690_, _06689_, _06688_);
  and (_06691_, _06690_, _06687_);
  nand (_06692_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_06693_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_06694_, _06693_, _06692_);
  or (_06695_, _06572_, ABINPUT[3]);
  or (_06696_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_06697_, _06696_, _06695_);
  or (_06698_, _06697_, _06569_);
  and (_06699_, _06698_, _06694_);
  nand (_06700_, _06699_, _06691_);
  or (_06701_, _06697_, _06588_);
  or (_06702_, _06590_, _06685_);
  not (_06703_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_06704_, _06594_, _06703_);
  and (_06705_, _06704_, _06702_);
  nand (_06706_, _06705_, _06701_);
  and (_06707_, _06706_, _06700_);
  nor (_06708_, _06706_, _06700_);
  nor (_06709_, _06708_, _06707_);
  not (_06710_, _06709_);
  nand (_06711_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  nand (_06712_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_06713_, _06712_, _06711_);
  not (_06714_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_06715_, _06560_, _06714_);
  not (_06716_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or (_06717_, _06553_, _06716_);
  and (_06718_, _06717_, _06715_);
  and (_06719_, _06718_, _06713_);
  or (_06720_, _06572_, ABINPUT[2]);
  or (_06721_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_06722_, _06721_, _06720_);
  or (_06723_, _06722_, _06569_);
  nand (_06724_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_06725_, _06556_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_06726_, _06725_, _06724_);
  and (_06727_, _06726_, _06723_);
  and (_06728_, _06727_, _06719_);
  or (_06729_, _06722_, _06588_);
  or (_06730_, _06590_, _06716_);
  not (_06731_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_06732_, _06594_, _06731_);
  and (_06733_, _06732_, _06730_);
  nand (_06734_, _06733_, _06729_);
  not (_06735_, _06734_);
  nor (_06736_, _06735_, _06728_);
  not (_06737_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_06738_, _06553_, _06737_);
  and (_06739_, _06556_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor (_06740_, _06739_, _06738_);
  and (_06741_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_06742_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_06743_, _06742_, _06741_);
  and (_06744_, _06743_, _06740_);
  or (_06745_, _06572_, ABINPUT[1]);
  or (_06746_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_06747_, _06746_, _06745_);
  and (_06748_, _06747_, _06568_);
  not (_06749_, _06748_);
  and (_06750_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_06751_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor (_06752_, _06751_, _06750_);
  and (_06753_, _06752_, _06749_);
  and (_06754_, _06753_, _06744_);
  nand (_06755_, _06747_, _06587_);
  or (_06756_, _06590_, _06737_);
  not (_06757_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_06758_, _06594_, _06757_);
  and (_06759_, _06758_, _06756_);
  nand (_06760_, _06759_, _06755_);
  not (_06761_, _06760_);
  nor (_06762_, _06761_, _06754_);
  and (_06763_, _06735_, _06728_);
  nor (_06764_, _06763_, _06736_);
  and (_06765_, _06764_, _06762_);
  nor (_06766_, _06765_, _06736_);
  nor (_06767_, _06766_, _06710_);
  nor (_06768_, _06767_, _06707_);
  nor (_06769_, _06768_, _06683_);
  and (_06770_, _06768_, _06683_);
  nor (_06771_, _06770_, _06769_);
  and (_06772_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_06773_, _06772_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nor (_06774_, _06572_, ABINPUT[0]);
  nor (_06775_, _06574_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_06776_, _06775_, _06774_);
  nor (_06777_, _06776_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_06778_, _06777_, _06773_);
  and (_06779_, _06761_, _06754_);
  nor (_06780_, _06779_, _06762_);
  and (_06781_, _06780_, _06778_);
  and (_06782_, _06781_, _06764_);
  and (_06783_, _06766_, _06710_);
  nor (_06784_, _06783_, _06767_);
  and (_06785_, _06784_, _06782_);
  not (_06786_, _06785_);
  nor (_06787_, _06786_, _06771_);
  nor (_06788_, _06768_, _06682_);
  or (_06789_, _06788_, _06681_);
  or (_06790_, _06789_, _06787_);
  and (_06791_, _06790_, _06655_);
  and (_06792_, _06791_, _06627_);
  nand (_06793_, _06556_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_06794_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  or (_06795_, _06553_, _06794_);
  and (_06796_, _06795_, _06793_);
  nand (_06797_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_06798_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_06799_, _06560_, _06798_);
  and (_06800_, _06799_, _06797_);
  and (_06801_, _06800_, _06796_);
  or (_06802_, _06572_, ABINPUT[7]);
  or (_06803_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_06804_, _06803_, _06802_);
  or (_06805_, _06804_, _06569_);
  nand (_06806_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand (_06807_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_06808_, _06807_, _06806_);
  and (_06809_, _06808_, _06805_);
  and (_06810_, _06809_, _06801_);
  or (_06811_, _06804_, _06588_);
  or (_06812_, _06590_, _06794_);
  not (_06813_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_06814_, _06594_, _06813_);
  and (_06815_, _06814_, _06812_);
  and (_06816_, _06815_, _06811_);
  nor (_06817_, _06816_, _06810_);
  and (_06818_, _06816_, _06810_);
  nor (_06819_, _06818_, _06817_);
  not (_06820_, _06819_);
  and (_06821_, _06653_, _06627_);
  nor (_06822_, _06821_, _06624_);
  nor (_06823_, _06822_, _06820_);
  and (_06824_, _06822_, _06820_);
  nor (_06826_, _06824_, _06823_);
  and (_06828_, _06826_, _06792_);
  nor (_06830_, _06823_, _06817_);
  not (_06832_, _06830_);
  nor (_06834_, _06832_, _06828_);
  and (_06835_, _06597_, _06586_);
  or (_06837_, _06835_, _06834_);
  and (_06839_, _06837_, _06599_);
  nor (_06840_, _06839_, _06549_);
  not (_06841_, _06840_);
  not (_06842_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_06843_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _06406_);
  and (_06844_, _06843_, _06842_);
  and (_06845_, _06844_, _06547_);
  not (_06846_, _06845_);
  not (_06847_, _06597_);
  and (_06848_, _06847_, _06586_);
  nor (_06849_, _06835_, _06598_);
  not (_06850_, _06816_);
  nor (_06851_, _06850_, _06810_);
  and (_06852_, _06622_, _06616_);
  nand (_06853_, _06651_, _06647_);
  and (_06854_, _06853_, _06646_);
  nor (_06855_, _06854_, _06627_);
  nor (_06856_, _06855_, _06852_);
  nor (_06857_, _06856_, _06819_);
  nor (_06858_, _06857_, _06851_);
  and (_06859_, _06856_, _06819_);
  nor (_06860_, _06859_, _06857_);
  not (_06861_, _06860_);
  and (_06862_, _06854_, _06627_);
  nor (_06863_, _06862_, _06855_);
  not (_06864_, _06863_);
  not (_06865_, _06655_);
  and (_06866_, _06760_, _06754_);
  nor (_06867_, _06866_, _06764_);
  nor (_06868_, _06734_, _06728_);
  nor (_06869_, _06868_, _06867_);
  nor (_06870_, _06869_, _06709_);
  and (_06871_, _06705_, _06701_);
  and (_06872_, _06871_, _06700_);
  nor (_06873_, _06872_, _06870_);
  nor (_06874_, _06873_, _06683_);
  and (_06875_, _06873_, _06683_);
  nor (_06876_, _06875_, _06874_);
  and (_06877_, _06869_, _06709_);
  nor (_06878_, _06877_, _06870_);
  not (_06879_, _06878_);
  and (_06880_, _06866_, _06764_);
  nor (_06881_, _06880_, _06867_);
  not (_06882_, _06881_);
  not (_06883_, _06778_);
  nor (_06884_, _06780_, _06883_);
  and (_06885_, _06884_, _06882_);
  and (_06886_, _06885_, _06879_);
  not (_06887_, _06886_);
  nor (_06888_, _06887_, _06876_);
  not (_06889_, _06680_);
  or (_06890_, _06889_, _06673_);
  and (_06891_, _06889_, _06673_);
  or (_06892_, _06873_, _06891_);
  and (_06893_, _06892_, _06890_);
  or (_06894_, _06893_, _06888_);
  and (_06895_, _06894_, _06865_);
  and (_06896_, _06895_, _06864_);
  and (_06897_, _06896_, _06861_);
  nor (_06898_, _06897_, _06858_);
  nor (_06899_, _06898_, _06849_);
  nor (_06900_, _06899_, _06848_);
  nor (_06901_, _06900_, _06846_);
  not (_06902_, _06810_);
  nor (_06903_, _06902_, _06616_);
  not (_06904_, _06903_);
  not (_06905_, _06646_);
  not (_06906_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_06907_, _06545_, _06906_);
  and (_06908_, _06907_, _06544_);
  not (_06909_, _06728_);
  nor (_06910_, _06909_, _06700_);
  nor (_06911_, _06910_, _06673_);
  and (_06912_, _06911_, _06908_);
  and (_06913_, _06912_, _06905_);
  nor (_06914_, _06913_, _06904_);
  nor (_06915_, _06914_, _06586_);
  nor (_06916_, _06915_, _06778_);
  not (_06917_, _06916_);
  not (_06918_, _06908_);
  nor (_06919_, _06883_, _06586_);
  not (_06920_, _06919_);
  nor (_06921_, _06920_, _06914_);
  nor (_06922_, _06921_, _06918_);
  and (_06923_, _06922_, _06917_);
  not (_06924_, _06754_);
  and (_06925_, _06546_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_06926_, _06925_, _06544_);
  and (_06927_, _06926_, _06924_);
  and (_06928_, _06776_, _06773_);
  not (_06929_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_06930_, _06546_, _06929_);
  and (_06931_, _06930_, _06844_);
  and (_06932_, _06843_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_06933_, _06932_, _06907_);
  and (_06934_, _06933_, _06776_);
  nor (_06935_, _06934_, _06931_);
  nor (_06936_, _06935_, _06928_);
  nor (_06937_, _06936_, _06927_);
  not (_06938_, _06912_);
  nor (_06939_, _06778_, _06776_);
  and (_06940_, _06930_, _06544_);
  nor (_06941_, _06843_, _06543_);
  and (_06942_, _06930_, _06941_);
  not (_06943_, _06942_);
  not (_06944_, _06776_);
  nor (_06945_, _06944_, _06773_);
  nor (_06946_, _06945_, _06943_);
  nor (_06947_, _06946_, _06940_);
  nor (_06948_, _06947_, _06939_);
  and (_06949_, _06941_, _06925_);
  and (_06950_, _06949_, _06944_);
  and (_06951_, _06941_, _06547_);
  nor (_06952_, _06951_, _06950_);
  and (_06953_, _06952_, _06778_);
  and (_06954_, _06907_, _06844_);
  nor (_06955_, _06954_, _06778_);
  nor (_06956_, _06955_, _06953_);
  not (_06957_, _06586_);
  and (_06958_, _06930_, _06932_);
  and (_06959_, _06958_, _06957_);
  or (_06960_, _06959_, _06956_);
  nor (_06961_, _06960_, _06948_);
  and (_06962_, _06961_, _06938_);
  and (_06963_, _06962_, _06937_);
  not (_06964_, _06963_);
  nor (_06965_, _06964_, _06923_);
  not (_06966_, _06965_);
  nor (_06967_, _06966_, _06901_);
  and (_06968_, _06967_, _06841_);
  nor (_06969_, _06968_, _06540_);
  not (_06970_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_06971_, _06539_, _06970_);
  nand (_06972_, _06971_, _06501_);
  or (_06973_, _06972_, _06969_);
  and (_06974_, _06973_, _06502_);
  and (_06975_, _06477_, _06434_);
  nor (_06976_, _06499_, _06463_);
  and (_06977_, _06976_, _06975_);
  and (_06978_, _06537_, _06513_);
  and (_06979_, _06978_, _06525_);
  not (_06980_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_06981_, _06481_, _06980_);
  not (_06982_, _06981_);
  nor (_06983_, _06982_, _06483_);
  not (_06984_, _06983_);
  nor (_06985_, _06984_, _06447_);
  and (_06986_, _06985_, _06979_);
  and (_06987_, _06986_, _06977_);
  or (_06988_, _06987_, _06974_);
  not (_06989_, rst);
  and (_06990_, _06883_, _06586_);
  and (_06991_, _06932_, _06925_);
  not (_06992_, _06991_);
  and (_06993_, _06778_, _06597_);
  nor (_06994_, _06993_, _06992_);
  not (_06995_, _06994_);
  nor (_06996_, _06995_, _06990_);
  and (_06997_, _06925_, _06844_);
  and (_06998_, _06910_, _06754_);
  and (_06999_, _06998_, _06673_);
  and (_07000_, _06999_, _06646_);
  and (_07001_, _07000_, _06903_);
  nor (_07002_, _07001_, _06883_);
  not (_07003_, _06673_);
  nor (_07004_, _06754_, _06728_);
  and (_07005_, _07004_, _06700_);
  and (_07006_, _07005_, _07003_);
  and (_07007_, _07006_, _06905_);
  and (_07008_, _07007_, _06616_);
  and (_07009_, _07008_, _06902_);
  nor (_07010_, _07009_, _06778_);
  or (_07011_, _07010_, _07002_);
  and (_07012_, _07011_, _06586_);
  nor (_07013_, _07011_, _06586_);
  nor (_07014_, _07013_, _07012_);
  and (_07015_, _07014_, _06997_);
  nor (_07016_, _07015_, _06996_);
  not (_07017_, _06940_);
  nor (_07018_, _07017_, _06835_);
  and (_07019_, _06942_, _06849_);
  nor (_07020_, _07019_, _07018_);
  and (_07021_, _06933_, _06598_);
  and (_07022_, _06954_, _06586_);
  nor (_07023_, _07022_, _07021_);
  and (_07024_, _06941_, _06907_);
  not (_07025_, _07024_);
  and (_07026_, _06544_, _06906_);
  and (_07027_, _06932_, _06547_);
  nor (_07028_, _07027_, _07026_);
  and (_07029_, _07028_, _07025_);
  and (_07030_, _06925_, _06541_);
  not (_07031_, _07030_);
  and (_07032_, _06930_, _06843_);
  nor (_07033_, _07032_, _06951_);
  and (_07034_, _07033_, _07031_);
  and (_07035_, _07034_, _07029_);
  nor (_07036_, _07035_, _06586_);
  not (_07037_, _07036_);
  and (_07038_, _07037_, _07023_);
  and (_07039_, _07038_, _07020_);
  and (_07040_, _07039_, _07016_);
  nand (_07041_, _07040_, _06987_);
  and (_07042_, _07041_, _06989_);
  and (_11486_, _07042_, _06988_);
  not (_07043_, _06525_);
  and (_07044_, _06978_, _07043_);
  and (_07045_, _06985_, _07044_);
  and (_07046_, _07045_, _06977_);
  and (_07047_, _06537_, _06514_);
  and (_07048_, _07047_, _07043_);
  and (_07049_, _06985_, _07048_);
  and (_07050_, _07049_, _06977_);
  nor (_07051_, _07050_, _07046_);
  and (_07052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_07053_, _07052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_07054_, _07053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_07055_, _07054_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_07056_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_07057_, _07056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_07058_, _07057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_07059_, _07058_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_07060_, _07059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_07061_, _07060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_07062_, _07061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_07063_, _07062_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_07064_, _07063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_07065_, _07064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_07066_, _07065_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_07067_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not (_07068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_07069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _07068_);
  and (_07070_, _07069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_07071_, _07070_, _07067_);
  nor (_07072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not (_07073_, _07072_);
  not (_07074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_07075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_07076_, _07075_, _07072_);
  and (_07077_, _07076_, _07074_);
  nor (_07078_, _07077_, _07073_);
  and (_07079_, _07078_, _07071_);
  nand (_07080_, _07079_, _07066_);
  nand (_07081_, _07080_, _07051_);
  or (_07082_, _07051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_07083_, _07082_, _06989_);
  and (_13884_, _07083_, _07081_);
  not (_07084_, _06434_);
  and (_07085_, _06477_, _07084_);
  and (_07086_, _06499_, _06463_);
  and (_07087_, _07086_, _07085_);
  and (_07088_, _06537_, _06525_);
  and (_07089_, _07088_, _06514_);
  and (_07090_, _07089_, _06448_);
  and (_07091_, _07090_, _07087_);
  and (_07092_, _06778_, _06623_);
  and (_07093_, _06883_, _06616_);
  or (_07094_, _07093_, _07092_);
  and (_07095_, _07094_, _06991_);
  not (_07096_, _06616_);
  and (_07097_, _07007_, _06883_);
  and (_07098_, _07000_, _06778_);
  nor (_07099_, _07098_, _07097_);
  and (_07100_, _07099_, _07096_);
  not (_07101_, _06997_);
  nor (_07102_, _07099_, _07096_);
  or (_07103_, _07102_, _07101_);
  nor (_07104_, _07103_, _07100_);
  nor (_07105_, _07104_, _07095_);
  not (_07106_, _07035_);
  and (_07107_, _07106_, _06616_);
  not (_07108_, _07107_);
  and (_07109_, _06942_, _06627_);
  nor (_07110_, _07017_, _06625_);
  not (_07111_, _07110_);
  and (_07112_, _06933_, _06624_);
  and (_07113_, _06954_, _07096_);
  nor (_07114_, _07113_, _07112_);
  nand (_07115_, _07114_, _07111_);
  nor (_07116_, _07115_, _07109_);
  and (_07117_, _07116_, _07108_);
  and (_07118_, _07117_, _07105_);
  not (_07119_, _07118_);
  and (_07120_, _07119_, _07091_);
  not (_07121_, _07087_);
  nand (_07122_, _07089_, _06447_);
  nor (_07123_, _07122_, _07121_);
  and (_07124_, _06525_, _06447_);
  and (_07125_, _07124_, _06978_);
  and (_07126_, _07125_, _07087_);
  nor (_07127_, _07126_, _07123_);
  and (_07128_, _06979_, _06448_);
  and (_07129_, _07087_, _07128_);
  not (_07130_, _07129_);
  and (_07131_, _07130_, _07127_);
  not (_07132_, _07131_);
  and (_07133_, _06981_, _07088_);
  nand (_07134_, _07133_, _07087_);
  or (_07135_, _07134_, _07132_);
  and (_07136_, _07135_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  or (_07137_, _07136_, _07120_);
  or (_07138_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_07139_, _07138_, _06989_);
  and (_06571_, _07139_, _07137_);
  and (_07140_, _07071_, _07064_);
  and (_07141_, _07140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_07142_, _07141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_07143_, _07141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_07144_, _07143_, _07142_);
  and (_07145_, _07072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not (_07146_, _07145_);
  and (_07147_, _07146_, _07071_);
  and (_07148_, _07147_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_07149_, _07148_, _07066_);
  or (_07150_, _07149_, _07077_);
  or (_07151_, _07150_, _07144_);
  not (_07152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_07153_, _07077_, _07152_);
  nor (_07154_, _07153_, _07046_);
  and (_07155_, _07154_, _07151_);
  and (_07156_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_07157_, _07156_, _07050_);
  or (_07158_, _07157_, _07155_);
  nand (_07159_, _07050_, _07040_);
  and (_07160_, _07159_, _06989_);
  and (_10680_, _07160_, _07158_);
  and (_07161_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_07162_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_12565_, _07162_, _07161_);
  not (_07164_, _07161_);
  not (_07165_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_07167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _07166_);
  and (_07168_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_07169_, _07168_, _07167_);
  and (_07170_, _07169_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_07171_, _07170_, _07165_);
  not (_07172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_07173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_07174_, _07173_, _07172_);
  and (_07175_, _07174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_07176_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_07177_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor (_07178_, _07177_, _07176_);
  and (_07179_, _07178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nor (_07180_, _07179_, _07175_);
  and (_07181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_07182_, _07181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_07183_, _07182_);
  and (_07184_, _07183_, _07180_);
  and (_07185_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_07186_, _07185_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_07187_, _07186_);
  and (_07188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_07189_, _07188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_07190_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_07191_, _07190_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_07193_, _07191_, _07189_);
  and (_07194_, _07193_, _07187_);
  and (_07195_, _07194_, _07184_);
  nor (_07196_, _07195_, _07171_);
  not (_07197_, _07196_);
  and (_07198_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _07165_);
  not (_07199_, _07198_);
  not (_07200_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_07201_, _07185_, _07200_);
  not (_07202_, _07201_);
  not (_07203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_07204_, _07188_, _07203_);
  not (_07205_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_07206_, _07190_, _07205_);
  nor (_07207_, _07206_, _07204_);
  and (_07208_, _07207_, _07202_);
  nor (_07209_, _07208_, _07199_);
  not (_07210_, _07209_);
  not (_07211_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_07212_, _07174_, _07211_);
  not (_07213_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_07215_, _07178_, _07213_);
  nor (_07216_, _07215_, _07212_);
  not (_07217_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_07218_, _07181_, _07217_);
  not (_07219_, _07218_);
  and (_07220_, _07219_, _07216_);
  or (_07221_, _07220_, _07199_);
  and (_07222_, _07221_, _07210_);
  and (_07223_, _07222_, _07197_);
  and (_07224_, _07223_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_07225_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_07226_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_07227_, _07226_, _07225_);
  nor (_07228_, _07227_, _07197_);
  or (_07229_, _07228_, _07224_);
  and (_07230_, _07229_, _07164_);
  and (_07231_, _07227_, _07161_);
  or (_07232_, _07231_, _07230_);
  and (_12832_, _07232_, _06989_);
  and (_07233_, _07195_, _07165_);
  nand (_07234_, _07233_, _07222_);
  nand (_07235_, _07225_, _07161_);
  and (_07236_, _07235_, _06989_);
  and (_12851_, _07236_, _07234_);
  nor (_07237_, _06778_, _06646_);
  and (_07238_, _06778_, _06853_);
  or (_07239_, _07238_, _07237_);
  and (_07240_, _07239_, _06991_);
  nor (_07242_, _07006_, _06778_);
  nor (_07243_, _06999_, _06883_);
  nor (_07244_, _07243_, _07242_);
  nor (_07245_, _07244_, _06905_);
  and (_07246_, _07244_, _06905_);
  nor (_07247_, _07246_, _07245_);
  and (_07248_, _07247_, _06997_);
  nor (_07249_, _07248_, _07240_);
  and (_07250_, _06942_, _06655_);
  and (_07251_, _06933_, _06653_);
  nor (_07252_, _07017_, _06654_);
  and (_07253_, _06954_, _06646_);
  or (_07254_, _07253_, _07252_);
  or (_07255_, _07254_, _07251_);
  nor (_07256_, _07255_, _07250_);
  nor (_07257_, _07035_, _06646_);
  not (_07258_, _07257_);
  and (_07259_, _07258_, _07256_);
  and (_07260_, _07259_, _07249_);
  and (_07261_, _07129_, _06981_);
  not (_07262_, _07261_);
  nor (_07263_, _07262_, _07260_);
  and (_07264_, _07262_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  or (_07265_, _07264_, _07263_);
  and (_13225_, _07265_, _06989_);
  and (_07266_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not (_07267_, _07184_);
  or (_07268_, _07194_, _07171_);
  or (_07269_, _07268_, _07267_);
  and (_07270_, _07269_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_07271_, _07221_, _07197_);
  and (_07272_, _07271_, _07270_);
  or (_07273_, _07272_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor (_07274_, _07222_, _07196_);
  nor (_07275_, _07208_, _07166_);
  nand (_07276_, _07275_, _07274_);
  nor (_07277_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_07278_, _07268_, _07164_);
  or (_07279_, _07278_, _07277_);
  and (_07281_, _07279_, _07276_);
  and (_07282_, _07281_, _07273_);
  or (_07283_, _07282_, _07266_);
  and (_13415_, _07283_, _06989_);
  and (_07284_, _07125_, _06983_);
  and (_07285_, _07284_, _06976_);
  and (_07286_, _06434_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_07287_, _07085_, _06976_);
  and (_07288_, _07287_, _07284_);
  not (_07289_, _07288_);
  and (_07290_, _07289_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_07291_, _07285_, _07085_);
  not (_07292_, _07291_);
  nor (_07293_, _07292_, _07260_);
  nor (_07294_, _07293_, _07290_);
  and (_07295_, _07294_, _07084_);
  nor (_07296_, _07295_, _07286_);
  and (_07297_, _07289_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_07298_, _06998_, _06883_);
  nor (_07299_, _07005_, _06778_);
  nor (_07300_, _07299_, _07298_);
  nor (_07301_, _07300_, _07003_);
  not (_07302_, _07301_);
  and (_07303_, _07300_, _07003_);
  nor (_07304_, _07303_, _07101_);
  and (_07305_, _07304_, _07302_);
  nor (_07306_, _06992_, _06680_);
  nor (_07307_, _07306_, _07305_);
  and (_07308_, _06933_, _06681_);
  and (_07309_, _06954_, _06673_);
  nor (_07310_, _07309_, _07308_);
  nor (_07311_, _07035_, _06673_);
  and (_07312_, _06942_, _06683_);
  nor (_07313_, _07017_, _06682_);
  or (_07314_, _07313_, _07312_);
  nor (_07315_, _07314_, _07311_);
  and (_07316_, _07315_, _07310_);
  and (_07317_, _07316_, _07307_);
  nor (_07318_, _07317_, _07292_);
  nor (_07319_, _07318_, _07297_);
  and (_07320_, _07319_, _06448_);
  not (_07321_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor (_07322_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_07323_, _07322_, _07321_);
  nor (_07324_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_07325_, _07324_, _06406_);
  and (_07326_, _07325_, _07323_);
  not (_07327_, _07326_);
  not (_07328_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_07330_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_07331_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_07332_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_07333_, _07332_, _07331_);
  and (_07334_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not (_07335_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_07337_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _07335_);
  and (_07338_, _07337_, _07331_);
  and (_07339_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_07340_, _07339_, _07334_);
  nor (_07341_, _07332_, _07331_);
  nand (_07342_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_07343_, _07332_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_07344_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_07345_, _07344_, _07342_);
  and (_07346_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_07347_, _07346_, _07331_);
  nand (_07348_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  not (_07349_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_07350_, _07349_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_07351_, _07350_, _07331_);
  nand (_07352_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_07353_, _07352_, _07348_);
  and (_07354_, _07353_, _07345_);
  nand (_07355_, _07354_, _07340_);
  nand (_07356_, _07355_, _07330_);
  nand (_07357_, _07356_, _07328_);
  nor (_07358_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _07328_);
  not (_07359_, _07358_);
  and (_07360_, _07359_, _07357_);
  or (_07361_, _07360_, _07327_);
  not (_07362_, _07323_);
  nor (_07363_, _07325_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_07364_, _07363_, _07362_);
  and (_07365_, _07364_, _07361_);
  nor (_07366_, _07365_, _06513_);
  not (_07367_, _07366_);
  nand (_07368_, _07367_, _07086_);
  nor (_07369_, _07368_, _07320_);
  nor (_07370_, _07319_, _06448_);
  and (_07371_, _07365_, _06513_);
  nand (_07372_, _06981_, _06525_);
  nand (_07373_, _06537_, _06477_);
  or (_07374_, _07373_, _07372_);
  or (_07375_, _07374_, _07371_);
  nor (_07376_, _07375_, _07370_);
  and (_07377_, _07376_, _07369_);
  and (_07378_, _07377_, _07296_);
  nor (_07379_, _07365_, _07319_);
  and (_07380_, _07379_, _07294_);
  and (_07381_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  not (_07382_, _07294_);
  not (_07383_, _07365_);
  nor (_07384_, _07383_, _07319_);
  and (_07385_, _07384_, _07382_);
  and (_07386_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_07387_, _07386_, _07381_);
  and (_07389_, _07379_, _07382_);
  and (_07390_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_07391_, _07383_, _07319_);
  and (_07392_, _07391_, _07382_);
  and (_07393_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_07394_, _07393_, _07390_);
  and (_07395_, _07394_, _07387_);
  and (_07396_, _07391_, _07294_);
  and (_07397_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_07398_, _07384_, _07294_);
  and (_07399_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_07400_, _07399_, _07397_);
  and (_07401_, _07365_, _07319_);
  and (_07402_, _07401_, _07382_);
  and (_07403_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and (_07404_, _07401_, _07294_);
  and (_07405_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_07406_, _07405_, _07403_);
  and (_07407_, _07406_, _07400_);
  and (_07408_, _07407_, _07395_);
  nor (_07409_, _07408_, _07378_);
  not (_07410_, _07317_);
  and (_07411_, _07378_, _07410_);
  nor (_07412_, _07411_, _07409_);
  nor (_14142_, _07412_, rst);
  and (_07413_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_07414_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor (_07415_, _07414_, _07413_);
  and (_07416_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_07417_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_07418_, _07417_, _07416_);
  and (_07419_, _07418_, _07415_);
  and (_07420_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_07421_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_07422_, _07421_, _07420_);
  and (_07423_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_07424_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_07425_, _07424_, _07423_);
  and (_07426_, _07425_, _07422_);
  and (_07427_, _07426_, _07419_);
  nor (_07428_, _07427_, _07378_);
  not (_07429_, _07260_);
  and (_07430_, _07378_, _07429_);
  nor (_07431_, _07430_, _07428_);
  nor (_14393_, _07431_, rst);
  and (_07432_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_07433_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_07434_, _07433_, _07432_);
  and (_07435_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_07436_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_07437_, _07436_, _07435_);
  and (_07438_, _07437_, _07434_);
  and (_07439_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_07440_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor (_07441_, _07440_, _07439_);
  and (_07442_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_07443_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor (_07444_, _07443_, _07442_);
  and (_07445_, _07444_, _07441_);
  and (_07446_, _07445_, _07438_);
  nor (_07447_, _07446_, _07378_);
  and (_07449_, _07378_, _07119_);
  nor (_07450_, _07449_, _07447_);
  nor (_01178_, _07450_, rst);
  not (_07452_, _06463_);
  nor (_07453_, _06499_, _07452_);
  and (_07454_, _07453_, _06975_);
  nor (_07455_, _06486_, _06447_);
  and (_07456_, _07455_, _06539_);
  and (_07457_, _07456_, _07454_);
  nand (_07458_, _07457_, _06968_);
  and (_07459_, _07454_, _06986_);
  not (_07460_, _07459_);
  nor (_07461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_07462_, _07461_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  not (_07463_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and (_07464_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_07465_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor (_07466_, _07465_, _07464_);
  nor (_07467_, _07466_, _07165_);
  or (_07468_, _07467_, _07463_);
  nor (_07469_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_07470_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_07471_, _07470_, _07165_);
  nor (_07472_, _07471_, _07469_);
  and (_07473_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_07474_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor (_07475_, _07474_, _07473_);
  nand (_07476_, _07475_, _07472_);
  or (_07477_, _07476_, _07468_);
  and (_07478_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_07479_, _07478_, _07462_);
  or (_07480_, _07479_, _07457_);
  and (_07481_, _07480_, _07460_);
  and (_07482_, _07481_, _07458_);
  nor (_07483_, _07460_, _07040_);
  or (_07484_, _07483_, _07482_);
  and (_01362_, _07484_, _06989_);
  and (_07485_, _07126_, _06981_);
  not (_07486_, _07485_);
  nor (_07487_, _07486_, _07317_);
  and (_07488_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or (_07489_, _07488_, _07487_);
  and (_01526_, _07489_, _06989_);
  not (_07490_, _07325_);
  nor (_07491_, _07346_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_07492_, _07491_, _07490_);
  nor (_07493_, _07492_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_07494_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  not (_07495_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor (_07496_, _07493_, _07495_);
  or (_07497_, _07496_, _07494_);
  and (_03985_, _07497_, _06989_);
  and (_07498_, _06951_, _06734_);
  and (_07499_, _06958_, _06616_);
  and (_07500_, _07001_, _06586_);
  and (_07501_, _07500_, _06761_);
  and (_07502_, _07501_, _06778_);
  nor (_07504_, _06761_, _06586_);
  and (_07505_, _07504_, _07009_);
  and (_07506_, _07505_, _06883_);
  nor (_07507_, _07506_, _07502_);
  nor (_07508_, _07507_, _06734_);
  and (_07509_, _07507_, _06734_);
  nor (_07510_, _07509_, _07508_);
  nor (_07511_, _07510_, _07101_);
  nor (_07512_, _06992_, _06728_);
  or (_07513_, _07512_, _07511_);
  or (_07514_, _07513_, _07499_);
  nor (_07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07516_, _07515_, _06586_);
  nor (_07517_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_07518_, _07517_);
  and (_07519_, _07518_, _07516_);
  not (_07520_, _07519_);
  or (_07521_, _06760_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not (_07522_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07523_, _06706_, _07522_);
  and (_07524_, _07523_, _07521_);
  or (_07525_, _07524_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07526_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07527_, _06853_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07528_, _06816_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_07529_, _07528_, _07527_);
  or (_07530_, _07529_, _07526_);
  and (_07531_, _07530_, _07525_);
  or (_07532_, _07531_, _07520_);
  not (_07533_, _07531_);
  or (_07534_, _07533_, _07519_);
  not (_07535_, _07534_);
  nand (_07536_, _07515_, _06810_);
  nor (_07537_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_07538_, _07537_);
  and (_07539_, _07538_, _07536_);
  not (_07540_, _07539_);
  and (_07541_, _06734_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07542_, _07541_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07543_, _06680_, _07522_);
  nand (_07544_, _06622_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_07545_, _07544_, _07543_);
  or (_07546_, _07545_, _07526_);
  and (_07547_, _07546_, _07542_);
  or (_07548_, _07547_, _07540_);
  or (_07549_, _07548_, _07535_);
  and (_07550_, _07549_, _07532_);
  and (_07551_, _07534_, _07532_);
  nand (_07552_, _07547_, _07540_);
  and (_07553_, _07552_, _07548_);
  and (_07554_, _07553_, _07551_);
  not (_07555_, _07515_);
  or (_07556_, _07555_, _06616_);
  nor (_07557_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_07558_, _07557_);
  nand (_07559_, _07558_, _07556_);
  and (_07560_, _06760_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07561_, _07560_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or (_07562_, _06706_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07563_, _06853_, _07522_);
  and (_07564_, _07563_, _07562_);
  or (_07565_, _07564_, _07526_);
  and (_07566_, _07565_, _07561_);
  nor (_07567_, _07566_, _07559_);
  or (_07568_, _06734_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07569_, _06680_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_07570_, _07569_, _07568_);
  and (_07571_, _07570_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07572_, _07571_);
  nand (_07573_, _07515_, _06646_);
  nor (_07574_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_07575_, _07574_);
  and (_07576_, _07575_, _07573_);
  and (_07577_, _07576_, _07572_);
  and (_07579_, _07566_, _07559_);
  or (_07580_, _07579_, _07567_);
  not (_07582_, _07580_);
  and (_07583_, _07582_, _07577_);
  or (_07585_, _07583_, _07567_);
  nand (_07586_, _07585_, _07554_);
  and (_07587_, _07586_, _07550_);
  and (_07588_, _07524_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07589_, _07588_);
  nand (_07590_, _07515_, _06673_);
  nor (_07591_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_07593_, _07591_);
  and (_07594_, _07593_, _07590_);
  nand (_07595_, _07594_, _07589_);
  or (_07596_, _07594_, _07589_);
  nand (_07597_, _07596_, _07595_);
  and (_07598_, _07541_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07600_, _07598_);
  or (_07601_, _07555_, _06700_);
  nor (_07602_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_07603_, _07602_);
  and (_07604_, _07603_, _07601_);
  nand (_07605_, _07604_, _07600_);
  and (_07606_, _07560_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07607_, _07606_);
  nand (_07608_, _07515_, _06728_);
  nor (_07609_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_07610_, _07609_);
  and (_07611_, _07610_, _07608_);
  nor (_07612_, _07611_, _07607_);
  or (_07613_, _07604_, _07600_);
  nand (_07614_, _07613_, _07605_);
  or (_07615_, _07614_, _07612_);
  and (_07617_, _07615_, _07605_);
  or (_07618_, _07617_, _07597_);
  nand (_07619_, _07618_, _07595_);
  nor (_07621_, _07576_, _07572_);
  nor (_07622_, _07621_, _07577_);
  and (_07623_, _07582_, _07622_);
  and (_07624_, _07623_, _07554_);
  nand (_07625_, _07624_, _07619_);
  nand (_07626_, _07625_, _07587_);
  nor (_07627_, _07570_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_07628_, _06622_, _07522_);
  and (_07629_, _06597_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_07630_, _07629_, _07628_);
  nor (_07631_, _07630_, _07526_);
  nor (_07632_, _07631_, _07627_);
  not (_07633_, _07632_);
  and (_07634_, _06816_, _06597_);
  nor (_07636_, _07634_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_07637_, _07545_, _07529_);
  nor (_07638_, _07630_, _07564_);
  and (_07639_, _07638_, _07637_);
  nor (_07640_, _07639_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_07641_, _07640_, _07636_);
  and (_07642_, _07641_, _07633_);
  and (_07643_, _07642_, _07626_);
  and (_07644_, _07643_, _07024_);
  nor (_07645_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_07646_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_07647_, _07646_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07648_, _07647_, _07645_);
  not (_07649_, _07648_);
  nor (_07650_, _07649_, _06839_);
  nor (_07651_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_07652_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_07653_, _07652_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07654_, _07653_, _07651_);
  nor (_07655_, _07654_, _07650_);
  not (_07656_, _07655_);
  and (_07657_, _07654_, _07650_);
  nor (_07658_, _07657_, _06549_);
  and (_07659_, _07658_, _07656_);
  nor (_07660_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  nand (_07661_, _07660_, _06597_);
  not (_07662_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  or (_07663_, _07662_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  or (_07664_, _07663_, _06622_);
  not (_07665_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  or (_07666_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _07665_);
  or (_07667_, _07666_, _06680_);
  and (_07668_, _07667_, _07664_);
  and (_07669_, _07666_, _07663_);
  or (_07670_, _06734_, _07665_);
  nand (_07671_, _07670_, _07669_);
  nand (_07672_, _07671_, _07668_);
  and (_07674_, _07672_, _07661_);
  and (_07675_, _07674_, _06909_);
  nand (_07676_, _07660_, _06816_);
  or (_07677_, _07663_, _06652_);
  or (_07678_, _07666_, _06871_);
  and (_07679_, _07678_, _07677_);
  or (_07680_, _06760_, _07665_);
  nand (_07681_, _07680_, _07669_);
  nand (_07682_, _07681_, _07679_);
  and (_07683_, _07682_, _07676_);
  and (_07684_, _07683_, _06924_);
  and (_07685_, _07684_, _07675_);
  and (_07686_, _07674_, _06924_);
  not (_07687_, _07686_);
  nand (_07688_, _07682_, _07676_);
  or (_07689_, _07688_, _06728_);
  and (_07690_, _07689_, _07687_);
  nor (_07691_, _07690_, _07685_);
  and (_07692_, _07691_, _07027_);
  or (_07693_, _07692_, _07659_);
  or (_07694_, _07693_, _07644_);
  or (_07695_, _07694_, _07514_);
  nor (_07696_, _07695_, _07498_);
  not (_07697_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_07698_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _06406_);
  and (_07699_, _07698_, _07697_);
  not (_07700_, _07699_);
  nor (_07701_, _07700_, _07696_);
  not (_07702_, _07701_);
  not (_07703_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_07704_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _06406_);
  and (_07705_, _07704_, _07703_);
  nor (_07706_, _06477_, _07084_);
  and (_07707_, _07706_, _06976_);
  and (_07708_, _07707_, _07125_);
  and (_07709_, _07708_, _06983_);
  nor (_07710_, _07709_, _07705_);
  nand (_07711_, _07642_, _07626_);
  not (_07712_, _07553_);
  and (_07713_, _07622_, _07619_);
  nor (_07714_, _07713_, _07577_);
  nor (_07715_, _07714_, _07579_);
  nor (_07716_, _07715_, _07567_);
  nor (_07717_, _07716_, _07712_);
  and (_07718_, _07716_, _07712_);
  nor (_07719_, _07718_, _07717_);
  nor (_07720_, _07719_, _07711_);
  and (_07721_, _07711_, _07540_);
  nor (_07722_, _07721_, _07720_);
  and (_07723_, _07722_, _07533_);
  nor (_07724_, _07722_, _07533_);
  nor (_07725_, _07724_, _07723_);
  not (_07726_, _07547_);
  and (_07727_, _07580_, _07714_);
  nor (_07728_, _07580_, _07714_);
  nor (_07729_, _07728_, _07727_);
  nor (_07730_, _07729_, _07711_);
  and (_07731_, _07711_, _07559_);
  nor (_07732_, _07731_, _07730_);
  and (_07733_, _07732_, _07726_);
  nand (_07734_, _07565_, _07561_);
  nor (_07735_, _07622_, _07619_);
  or (_07736_, _07735_, _07713_);
  and (_07737_, _07736_, _07643_);
  nor (_07738_, _07643_, _07576_);
  nor (_07739_, _07738_, _07737_);
  and (_07740_, _07739_, _07734_);
  not (_07741_, _07740_);
  nor (_07742_, _07732_, _07726_);
  or (_07743_, _07733_, _07742_);
  nor (_07744_, _07743_, _07741_);
  nor (_07745_, _07744_, _07733_);
  not (_07746_, _07745_);
  and (_07747_, _07617_, _07597_);
  not (_07748_, _07747_);
  and (_07749_, _07748_, _07618_);
  nor (_07750_, _07749_, _07711_);
  nor (_07751_, _07643_, _07594_);
  nor (_07752_, _07751_, _07750_);
  nor (_07753_, _07752_, _07572_);
  not (_07754_, _07753_);
  not (_07755_, _07611_);
  or (_07756_, _07711_, _07607_);
  nand (_07757_, _07756_, _07755_);
  or (_07758_, _07756_, _07755_);
  and (_07759_, _07758_, _07757_);
  nand (_07760_, _07759_, _07600_);
  or (_07761_, _07759_, _07600_);
  and (_07762_, _07761_, _07760_);
  and (_07763_, _07515_, _06754_);
  nor (_07765_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor (_07766_, _07765_, _07763_);
  nor (_07768_, _07766_, _07607_);
  not (_07769_, _07768_);
  nand (_07770_, _07769_, _07762_);
  and (_07771_, _07770_, _07760_);
  and (_07772_, _07614_, _07612_);
  not (_07774_, _07772_);
  and (_07775_, _07774_, _07615_);
  or (_07776_, _07775_, _07711_);
  or (_07777_, _07643_, _07604_);
  and (_07778_, _07777_, _07776_);
  and (_07779_, _07778_, _07589_);
  nor (_07780_, _07778_, _07589_);
  or (_07781_, _07780_, _07779_);
  or (_07782_, _07781_, _07771_);
  and (_07783_, _07752_, _07572_);
  nor (_07784_, _07783_, _07779_);
  nand (_07786_, _07784_, _07782_);
  and (_07787_, _07786_, _07754_);
  nor (_07788_, _07739_, _07734_);
  nor (_07789_, _07788_, _07740_);
  not (_07790_, _07743_);
  and (_07791_, _07790_, _07789_);
  and (_07792_, _07791_, _07787_);
  or (_07793_, _07792_, _07746_);
  and (_07794_, _07793_, _07725_);
  and (_07795_, _07711_, _07519_);
  not (_07796_, _07717_);
  and (_07797_, _07796_, _07548_);
  and (_07798_, _07797_, _07551_);
  nor (_07799_, _07797_, _07551_);
  or (_07800_, _07799_, _07798_);
  and (_07801_, _07800_, _07643_);
  or (_07802_, _07801_, _07795_);
  and (_07803_, _07802_, _07633_);
  or (_07804_, _07803_, _07723_);
  or (_07805_, _07804_, _07794_);
  not (_07807_, _07641_);
  nor (_07808_, _07802_, _07633_);
  nor (_07809_, _07808_, _07807_);
  nand (_07810_, _07809_, _07805_);
  or (_07811_, _07769_, _07762_);
  and (_07812_, _07811_, _07770_);
  or (_07813_, _07812_, _07810_);
  and (_07814_, _07809_, _07805_);
  or (_07815_, _07814_, _07759_);
  and (_07816_, _07815_, _07813_);
  nand (_07817_, _07816_, _07024_);
  not (_07818_, _07660_);
  and (_07819_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_07821_, _07674_, _06905_);
  and (_07822_, _07683_, _07003_);
  and (_07823_, _07822_, _07821_);
  and (_07824_, _07683_, _06905_);
  and (_07825_, _07674_, _06616_);
  nand (_07826_, _07825_, _07824_);
  and (_07827_, _07683_, _06616_);
  or (_07828_, _07827_, _07821_);
  and (_07830_, _07828_, _07826_);
  and (_07831_, _07830_, _07823_);
  or (_07832_, _07826_, _06810_);
  and (_07833_, _07683_, _06902_);
  not (_07835_, _07833_);
  nand (_07836_, _07835_, _07826_);
  and (_07837_, _07836_, _07832_);
  nand (_07838_, _07837_, _07825_);
  or (_07839_, _07833_, _07825_);
  and (_07840_, _07839_, _07838_);
  nand (_07841_, _07840_, _07831_);
  not (_07842_, _07841_);
  not (_07843_, _07832_);
  or (_07844_, _07688_, _06586_);
  nand (_07845_, _07672_, _07661_);
  or (_07846_, _07845_, _06810_);
  or (_07847_, _07846_, _07844_);
  nand (_07848_, _07846_, _07844_);
  and (_07849_, _07848_, _07847_);
  and (_07850_, _07849_, _07843_);
  not (_07851_, _07850_);
  and (_07852_, _07837_, _07825_);
  nand (_07853_, _07849_, _07852_);
  or (_07854_, _07849_, _07852_);
  nand (_07855_, _07854_, _07853_);
  nand (_07856_, _07855_, _07832_);
  and (_07857_, _07856_, _07851_);
  nand (_07858_, _07857_, _07842_);
  or (_07859_, _07857_, _07842_);
  nand (_07860_, _07859_, _07858_);
  not (_07861_, _07860_);
  and (_07862_, _07683_, _06700_);
  nand (_07863_, _07862_, _07675_);
  and (_07864_, _07674_, _06700_);
  and (_07865_, _07864_, _07689_);
  nand (_07866_, _07865_, _07822_);
  nand (_07867_, _07866_, _07863_);
  not (_07868_, _07823_);
  and (_07870_, _07674_, _07003_);
  or (_07871_, _07870_, _07824_);
  and (_07872_, _07871_, _07868_);
  nand (_07873_, _07872_, _07867_);
  not (_07874_, _07873_);
  not (_07875_, _07831_);
  or (_07876_, _07830_, _07823_);
  and (_07877_, _07876_, _07875_);
  and (_07878_, _07877_, _07874_);
  or (_07879_, _07840_, _07831_);
  and (_07880_, _07879_, _07841_);
  nand (_07881_, _07880_, _07878_);
  or (_07882_, _07862_, _07675_);
  and (_07883_, _07882_, _07863_);
  and (_07884_, _07883_, _07685_);
  or (_07885_, _07865_, _07822_);
  and (_07886_, _07885_, _07866_);
  nand (_07887_, _07886_, _07884_);
  not (_07888_, _07887_);
  or (_07889_, _07872_, _07867_);
  and (_07890_, _07889_, _07873_);
  nand (_07891_, _07890_, _07888_);
  not (_07892_, _07891_);
  nand (_07893_, _07877_, _07874_);
  or (_07894_, _07877_, _07874_);
  and (_07895_, _07894_, _07893_);
  nand (_07896_, _07895_, _07892_);
  not (_07897_, _07896_);
  or (_07898_, _07880_, _07878_);
  and (_07899_, _07898_, _07881_);
  nand (_07900_, _07899_, _07897_);
  nand (_07901_, _07900_, _07881_);
  nand (_07902_, _07901_, _07861_);
  nand (_07903_, _07902_, _07858_);
  and (_07904_, _07674_, _06957_);
  and (_07905_, _07904_, _07835_);
  not (_07906_, _07905_);
  and (_07907_, _07851_, _07853_);
  nor (_07908_, _07907_, _07906_);
  and (_07909_, _07907_, _07906_);
  nor (_07910_, _07909_, _07908_);
  nand (_07911_, _07910_, _07903_);
  or (_07912_, _07910_, _07903_);
  and (_07913_, _07912_, _07911_);
  nand (_07914_, _07913_, _07819_);
  and (_07915_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  or (_07916_, _07901_, _07861_);
  and (_07917_, _07916_, _07902_);
  nand (_07918_, _07917_, _07915_);
  or (_07919_, _07917_, _07915_);
  nand (_07920_, _07919_, _07918_);
  and (_07921_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or (_07922_, _07899_, _07897_);
  and (_07923_, _07922_, _07900_);
  nand (_07924_, _07923_, _07921_);
  or (_07925_, _07923_, _07921_);
  nand (_07926_, _07925_, _07924_);
  and (_07927_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  or (_07928_, _07895_, _07892_);
  and (_07929_, _07928_, _07896_);
  nand (_07930_, _07929_, _07927_);
  or (_07931_, _07929_, _07927_);
  nand (_07932_, _07931_, _07930_);
  and (_07934_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or (_07935_, _07890_, _07888_);
  and (_07936_, _07935_, _07891_);
  nand (_07937_, _07936_, _07934_);
  and (_07938_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or (_07939_, _07886_, _07884_);
  and (_07940_, _07939_, _07887_);
  nand (_07941_, _07940_, _07938_);
  and (_07942_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  not (_07943_, _07942_);
  nor (_07944_, _07883_, _07685_);
  or (_07945_, _07944_, _07884_);
  or (_07946_, _07945_, _07943_);
  or (_07947_, _07940_, _07938_);
  nand (_07948_, _07947_, _07941_);
  or (_07949_, _07948_, _07946_);
  and (_07950_, _07949_, _07941_);
  or (_07951_, _07936_, _07934_);
  nand (_07952_, _07951_, _07937_);
  or (_07953_, _07952_, _07950_);
  and (_07954_, _07953_, _07937_);
  or (_07955_, _07954_, _07932_);
  and (_07956_, _07955_, _07930_);
  or (_07957_, _07956_, _07926_);
  and (_07958_, _07957_, _07924_);
  or (_07960_, _07958_, _07920_);
  and (_07961_, _07960_, _07918_);
  or (_07962_, _07913_, _07819_);
  nand (_07963_, _07962_, _07914_);
  or (_07964_, _07963_, _07961_);
  and (_07965_, _07964_, _07914_);
  and (_07966_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not (_07967_, _07908_);
  and (_07968_, _07967_, _07847_);
  nand (_07970_, _07968_, _07911_);
  nand (_07971_, _07970_, _07966_);
  or (_07972_, _07970_, _07966_);
  nand (_07974_, _07972_, _07971_);
  or (_07975_, _07974_, _07965_);
  nand (_07977_, _07974_, _07965_);
  and (_07978_, _07977_, _07975_);
  nand (_07979_, _07978_, _07027_);
  nor (_07981_, _06884_, _06882_);
  nor (_07982_, _07981_, _06885_);
  nor (_07983_, _07982_, _06846_);
  not (_07984_, _07983_);
  nor (_07985_, _06911_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_07986_, _07985_, _06909_);
  nor (_07987_, _07985_, _06909_);
  nor (_07988_, _07987_, _07986_);
  nor (_07990_, _07988_, _06918_);
  and (_07991_, _06942_, _06764_);
  nor (_07993_, _07017_, _06763_);
  not (_07994_, _07993_);
  and (_07995_, _06933_, _06736_);
  and (_07996_, _06954_, _06728_);
  nor (_07998_, _07996_, _07995_);
  nand (_07999_, _07998_, _07994_);
  nor (_08000_, _07999_, _07991_);
  not (_08001_, _07032_);
  nor (_08002_, _08001_, _06754_);
  not (_08003_, _08002_);
  and (_08004_, _06951_, _06909_);
  and (_08005_, _07030_, _06700_);
  nor (_08006_, _08005_, _08004_);
  and (_08007_, _08006_, _08003_);
  and (_08008_, _08007_, _08000_);
  not (_08009_, _08008_);
  nor (_08010_, _08009_, _07990_);
  and (_08011_, _06991_, _06734_);
  and (_08012_, _06754_, _06728_);
  nor (_08013_, _08012_, _07004_);
  nor (_08014_, _08013_, _06778_);
  and (_08015_, _08013_, _06778_);
  nor (_08016_, _08015_, _08014_);
  and (_08017_, _08016_, _06997_);
  nor (_08018_, _08017_, _08011_);
  not (_08019_, _08018_);
  nor (_08020_, _06764_, _06762_);
  or (_08021_, _08020_, _06765_);
  and (_08022_, _08021_, _06781_);
  nor (_08023_, _08021_, _06781_);
  or (_08024_, _08023_, _08022_);
  and (_08025_, _08024_, _06548_);
  nor (_08026_, _08025_, _08019_);
  and (_08027_, _08026_, _08010_);
  and (_08028_, _08027_, _07984_);
  and (_08029_, _08028_, _07979_);
  nand (_08030_, _08029_, _07817_);
  or (_08031_, _08030_, _07710_);
  not (_08032_, _07089_);
  nor (_08033_, _06968_, _08032_);
  nor (_08034_, _07089_, _06731_);
  nor (_08035_, _08034_, _08033_);
  nor (_08036_, _06499_, _06448_);
  and (_08037_, _08036_, _06434_);
  nor (_08038_, _06477_, _06463_);
  and (_08039_, _08038_, _06485_);
  and (_08040_, _08039_, _08037_);
  and (_08041_, _07710_, _07700_);
  and (_08042_, _08041_, _08040_);
  not (_08043_, _08042_);
  nor (_08044_, _08043_, _08035_);
  not (_08045_, _07710_);
  nor (_08046_, _08040_, _06731_);
  nor (_08047_, _08046_, _08045_);
  not (_08048_, _08047_);
  nor (_08049_, _08048_, _08044_);
  nor (_08050_, _08049_, _07699_);
  nand (_08051_, _08050_, _08031_);
  nand (_08052_, _08051_, _07702_);
  and (_06536_, _08052_, _06989_);
  and (_08053_, _06951_, _06760_);
  and (_08055_, _06958_, _06905_);
  nor (_08056_, _06990_, _06919_);
  not (_08057_, _08056_);
  nor (_08058_, _08057_, _07011_);
  nor (_08059_, _08058_, _06760_);
  and (_08060_, _08058_, _06760_);
  nor (_08061_, _08060_, _08059_);
  and (_08062_, _08061_, _06997_);
  nor (_08063_, _06992_, _06754_);
  or (_08064_, _08063_, _08062_);
  or (_08065_, _08064_, _08055_);
  and (_08066_, _07814_, _07024_);
  and (_08067_, _07649_, _06839_);
  nor (_08068_, _08067_, _07650_);
  and (_08069_, _08068_, _06548_);
  and (_08070_, _07684_, _07027_);
  or (_08071_, _08070_, _08069_);
  or (_08072_, _08071_, _08066_);
  or (_08074_, _08072_, _08065_);
  or (_08075_, _08074_, _08053_);
  nand (_08076_, _08075_, _07699_);
  nand (_08077_, _07814_, _07606_);
  and (_08078_, _08077_, _07766_);
  nor (_08079_, _08077_, _07766_);
  or (_08080_, _08079_, _08078_);
  nand (_08082_, _08080_, _07024_);
  not (_08083_, _07964_);
  and (_08084_, _07963_, _07961_);
  nor (_08085_, _08084_, _08083_);
  and (_08086_, _08085_, _07027_);
  nor (_08087_, _06780_, _06778_);
  nor (_08089_, _08087_, _06781_);
  nor (_08090_, _06845_, _06548_);
  not (_08091_, _08090_);
  and (_08092_, _08091_, _08089_);
  not (_08093_, _08092_);
  nor (_08095_, _06943_, _06762_);
  nor (_08096_, _08095_, _06940_);
  or (_08098_, _08096_, _06779_);
  and (_08099_, _06997_, _06754_);
  and (_08101_, _06991_, _06760_);
  nor (_08102_, _08101_, _08099_);
  and (_08103_, _06933_, _06762_);
  and (_08104_, _06954_, _06754_);
  nor (_08106_, _08104_, _08103_);
  and (_08107_, _08106_, _08102_);
  and (_08109_, _06958_, _06778_);
  nor (_08110_, _06951_, _06908_);
  nor (_08112_, _08110_, _06754_);
  nor (_08113_, _08112_, _08109_);
  and (_08114_, _06931_, _06957_);
  nor (_08115_, _07031_, _06728_);
  nor (_08116_, _08115_, _08114_);
  and (_08117_, _08116_, _08113_);
  and (_08118_, _08117_, _08107_);
  and (_08119_, _08118_, _08098_);
  and (_08120_, _08119_, _08093_);
  not (_08121_, _08120_);
  nor (_08122_, _08121_, _08086_);
  nand (_08123_, _08122_, _08082_);
  or (_08124_, _08123_, _07710_);
  not (_08125_, _08040_);
  not (_08126_, _06968_);
  and (_08127_, _08126_, _06979_);
  nor (_08128_, _06979_, _06757_);
  nor (_08129_, _08128_, _08127_);
  nor (_08130_, _08129_, _08125_);
  nor (_08131_, _08040_, _06757_);
  nor (_08132_, _08131_, _08045_);
  not (_08133_, _08132_);
  nor (_08134_, _08133_, _08130_);
  nor (_08136_, _08134_, _07699_);
  nand (_08137_, _08136_, _08124_);
  nand (_08138_, _08137_, _08076_);
  and (_06542_, _08138_, _06989_);
  and (_08139_, _07326_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_08140_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not (_08141_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_08142_, _08139_, _08141_);
  or (_08143_, _08142_, _08140_);
  and (_06580_, _08143_, _06989_);
  and (_08144_, _06951_, _06623_);
  and (_08145_, _06958_, _06909_);
  and (_08146_, _07505_, _06734_);
  and (_08147_, _08146_, _06706_);
  and (_08148_, _08147_, _06889_);
  nor (_08149_, _08148_, _06778_);
  nor (_08150_, _06760_, _06734_);
  and (_08151_, _06871_, _06680_);
  and (_08152_, _08151_, _08150_);
  and (_08153_, _08152_, _07500_);
  and (_08154_, _08153_, _06652_);
  nor (_08155_, _08154_, _06883_);
  nor (_08156_, _06778_, _06853_);
  or (_08157_, _08156_, _08155_);
  nor (_08158_, _08157_, _08149_);
  and (_08159_, _08158_, _06622_);
  nor (_08160_, _08158_, _06622_);
  nor (_08161_, _08160_, _08159_);
  nor (_08162_, _08161_, _07101_);
  nor (_08163_, _06778_, _06622_);
  and (_08164_, _06778_, _06616_);
  or (_08165_, _08164_, _08163_);
  and (_08166_, _08165_, _06991_);
  or (_08167_, _08166_, _08162_);
  or (_08168_, _08167_, _08145_);
  and (_08169_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_08170_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_08171_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_08172_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08171_);
  nor (_08173_, _08172_, _08170_);
  nor (_08174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_08175_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_08176_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08175_);
  nor (_08177_, _08176_, _08174_);
  and (_08178_, _08177_, _07657_);
  and (_08179_, _08178_, _08173_);
  nor (_08180_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_08182_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_08183_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08182_);
  nor (_08184_, _08183_, _08180_);
  and (_08185_, _08184_, _08179_);
  nor (_08186_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_08187_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_08188_, _08187_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_08189_, _08188_, _08186_);
  nor (_08190_, _08189_, _08185_);
  and (_08191_, _08189_, _08185_);
  nor (_08192_, _08191_, _08190_);
  and (_08193_, _08192_, _06548_);
  and (_08195_, _07954_, _07932_);
  not (_08196_, _08195_);
  and (_08197_, _08196_, _07955_);
  and (_08198_, _08197_, _07027_);
  or (_08199_, _08198_, _08193_);
  or (_08200_, _08199_, _08169_);
  or (_08201_, _08200_, _08168_);
  nor (_08202_, _08201_, _08144_);
  nor (_08203_, _08202_, _07700_);
  not (_08204_, _08203_);
  nand (_08205_, _07810_, _07732_);
  nand (_08206_, _07789_, _07787_);
  and (_08207_, _08206_, _07741_);
  nand (_08208_, _08207_, _07790_);
  or (_08209_, _08207_, _07790_);
  nand (_08210_, _08209_, _08208_);
  nand (_08211_, _08210_, _07814_);
  nand (_08212_, _08211_, _08205_);
  nand (_08213_, _08212_, _07024_);
  or (_08214_, _07974_, _07914_);
  nand (_08215_, _08214_, _07971_);
  and (_08216_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_08218_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_08219_, _08218_, _08216_);
  and (_08220_, _08219_, _08215_);
  nor (_08221_, _07974_, _07963_);
  nand (_08222_, _08219_, _08221_);
  nor (_08223_, _08222_, _07961_);
  or (_08224_, _08223_, _08220_);
  and (_08225_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_08226_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_08227_, _08226_, _08225_);
  nand (_08228_, _08227_, _08224_);
  and (_08229_, _08224_, _08225_);
  or (_08230_, _08226_, _08229_);
  and (_08231_, _08230_, _08228_);
  nand (_08232_, _08231_, _07027_);
  nor (_08233_, _06895_, _06864_);
  nor (_08234_, _08233_, _06896_);
  nor (_08235_, _08234_, _06846_);
  not (_08236_, _08235_);
  nor (_08237_, _06653_, _06627_);
  nor (_08238_, _08237_, _06821_);
  nor (_08239_, _08238_, _06791_);
  not (_08240_, _08239_);
  nor (_08241_, _06792_, _06549_);
  and (_08242_, _08241_, _08240_);
  nor (_08243_, _06903_, _06586_);
  nor (_08244_, _08243_, _06778_);
  and (_08245_, _08244_, _06938_);
  nor (_08246_, _08245_, _06913_);
  and (_08247_, _08246_, _07096_);
  nor (_08248_, _08246_, _07096_);
  nor (_08249_, _08248_, _08247_);
  nor (_08251_, _08249_, _06918_);
  nor (_08252_, _07031_, _06810_);
  not (_08253_, _08252_);
  and (_08254_, _06951_, _06616_);
  not (_08255_, _08254_);
  or (_08256_, _08001_, _06646_);
  and (_08257_, _08256_, _08255_);
  and (_08258_, _08257_, _08253_);
  and (_08259_, _08258_, _07116_);
  not (_08260_, _08259_);
  nor (_08261_, _08260_, _08251_);
  and (_08262_, _08261_, _07105_);
  not (_08263_, _08262_);
  nor (_08264_, _08263_, _08242_);
  and (_08265_, _08264_, _08236_);
  and (_08267_, _08265_, _08232_);
  nand (_08268_, _08267_, _08213_);
  or (_08269_, _08268_, _07710_);
  nor (_08270_, _08040_, _06619_);
  nor (_08271_, _08270_, _08045_);
  and (_08272_, _06968_, _07048_);
  or (_08273_, _07048_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_08274_, _08273_, _08040_);
  or (_08275_, _08274_, _08272_);
  and (_08276_, _08275_, _08271_);
  nor (_08277_, _08276_, _07699_);
  nand (_08278_, _08277_, _08269_);
  nand (_08279_, _08278_, _08204_);
  and (_06626_, _08279_, _06989_);
  and (_08280_, _06951_, _06853_);
  and (_08281_, _06958_, _06924_);
  nor (_08282_, _08153_, _06883_);
  nor (_08283_, _08282_, _08149_);
  nor (_08284_, _08283_, _06853_);
  and (_08285_, _08283_, _06853_);
  nor (_08286_, _08285_, _08284_);
  and (_08287_, _08286_, _06997_);
  and (_08288_, _06778_, _06646_);
  nor (_08289_, _08156_, _06992_);
  not (_08290_, _08289_);
  nor (_08291_, _08290_, _08288_);
  or (_08292_, _08291_, _08287_);
  or (_08293_, _08292_, _08281_);
  and (_08294_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor (_08295_, _08184_, _08179_);
  not (_08296_, _08295_);
  nor (_08298_, _08185_, _06549_);
  and (_08299_, _08298_, _08296_);
  and (_08300_, _07952_, _07950_);
  not (_08301_, _08300_);
  and (_08302_, _08301_, _07953_);
  and (_08303_, _08302_, _07027_);
  or (_08304_, _08303_, _08299_);
  or (_08305_, _08304_, _08294_);
  or (_08306_, _08305_, _08293_);
  nor (_08307_, _08306_, _08280_);
  nor (_08308_, _08307_, _07700_);
  not (_08309_, _08308_);
  or (_08310_, _07789_, _07787_);
  and (_08311_, _08310_, _08206_);
  and (_08312_, _08311_, _07814_);
  and (_08313_, _07810_, _07739_);
  or (_08314_, _08313_, _08312_);
  nand (_08315_, _08314_, _07024_);
  nor (_08316_, _08224_, _08225_);
  nor (_08317_, _08316_, _08229_);
  nand (_08318_, _08317_, _07027_);
  nor (_08319_, _06894_, _06655_);
  and (_08320_, _06894_, _06655_);
  nor (_08322_, _08320_, _08319_);
  and (_08323_, _08322_, _06845_);
  not (_08324_, _08323_);
  nor (_08325_, _06790_, _06655_);
  nor (_08326_, _08325_, _06791_);
  and (_08327_, _08326_, _06548_);
  nor (_08328_, _06912_, _06905_);
  or (_08329_, _08328_, _06918_);
  nor (_08331_, _08329_, _06913_);
  not (_08332_, _08331_);
  or (_08333_, _08001_, _06673_);
  nand (_08334_, _07030_, _06616_);
  not (_08335_, _08334_);
  and (_08336_, _06951_, _06905_);
  nor (_08337_, _08336_, _08335_);
  and (_08338_, _08337_, _08333_);
  and (_08339_, _08338_, _07256_);
  and (_08340_, _08339_, _08332_);
  and (_08341_, _08340_, _07249_);
  not (_08342_, _08341_);
  nor (_08343_, _08342_, _08327_);
  and (_08344_, _08343_, _08324_);
  and (_08345_, _08344_, _08318_);
  nand (_08346_, _08345_, _08315_);
  or (_08348_, _08346_, _07710_);
  and (_08349_, _08126_, _07044_);
  nor (_08350_, _07044_, _06649_);
  nor (_08351_, _08350_, _08349_);
  nor (_08352_, _08351_, _08043_);
  nor (_08353_, _08040_, _06649_);
  nor (_08354_, _08353_, _08045_);
  not (_08355_, _08354_);
  nor (_08356_, _08355_, _08352_);
  nor (_08357_, _08356_, _07699_);
  nand (_08358_, _08357_, _08348_);
  nand (_08359_, _08358_, _08309_);
  and (_06638_, _08359_, _06989_);
  and (_08360_, _06951_, _06889_);
  and (_08361_, _08150_, _07500_);
  and (_08362_, _08361_, _06871_);
  nor (_08363_, _08362_, _06883_);
  nor (_08364_, _08147_, _06778_);
  nor (_08365_, _08364_, _08363_);
  and (_08366_, _08365_, _06889_);
  not (_08367_, _08366_);
  nor (_08368_, _08365_, _06889_);
  nor (_08369_, _08368_, _07101_);
  and (_08370_, _08369_, _08367_);
  nor (_08371_, _06992_, _06673_);
  or (_08372_, _08371_, _08370_);
  or (_08373_, _08372_, _06959_);
  and (_08374_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor (_08375_, _08178_, _08173_);
  nor (_08376_, _08375_, _08179_);
  and (_08377_, _08376_, _06548_);
  and (_08378_, _07948_, _07946_);
  not (_08379_, _08378_);
  and (_08380_, _08379_, _07949_);
  and (_08381_, _08380_, _07027_);
  or (_08382_, _08381_, _08377_);
  or (_08383_, _08382_, _08374_);
  or (_08384_, _08383_, _08373_);
  nor (_08385_, _08384_, _08360_);
  nor (_08386_, _08385_, _07700_);
  not (_08387_, _08386_);
  nand (_08388_, _07810_, _07752_);
  or (_08389_, _07783_, _07753_);
  not (_08390_, _07779_);
  and (_08391_, _07782_, _08390_);
  and (_08392_, _08391_, _08389_);
  nor (_08393_, _08391_, _08389_);
  or (_08394_, _08393_, _08392_);
  or (_08395_, _08394_, _07810_);
  nand (_08396_, _08395_, _08388_);
  nand (_08397_, _08396_, _07024_);
  nand (_08398_, _07975_, _07971_);
  nand (_08399_, _08398_, _08216_);
  not (_08400_, _08218_);
  and (_08401_, _08400_, _08399_);
  nor (_08402_, _08401_, _08224_);
  nand (_08403_, _08402_, _07027_);
  and (_08404_, _06887_, _06876_);
  nor (_08405_, _08404_, _06888_);
  nor (_08406_, _08405_, _06846_);
  not (_08407_, _08406_);
  and (_08408_, _06786_, _06771_);
  or (_08409_, _08408_, _06549_);
  nor (_08410_, _08409_, _06787_);
  not (_08411_, _08410_);
  not (_08412_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_08413_, _06910_, _08412_);
  nor (_08414_, _08413_, _07003_);
  not (_08415_, _08414_);
  nor (_08416_, _06911_, _06918_);
  and (_08417_, _08416_, _08415_);
  not (_08418_, _08417_);
  and (_08419_, _06951_, _07003_);
  not (_08420_, _08419_);
  and (_08421_, _08420_, _07310_);
  or (_08422_, _07031_, _06646_);
  and (_08423_, _07032_, _06700_);
  not (_08424_, _08423_);
  nand (_08425_, _08424_, _08422_);
  nor (_08426_, _08425_, _07314_);
  and (_08427_, _08426_, _08421_);
  and (_08428_, _08427_, _07307_);
  and (_08429_, _08428_, _08418_);
  and (_08430_, _08429_, _08411_);
  and (_08431_, _08430_, _08407_);
  and (_08432_, _08431_, _08403_);
  nand (_08433_, _08432_, _08397_);
  or (_08434_, _08433_, _07710_);
  nor (_08435_, _06537_, _06513_);
  and (_08436_, _08435_, _06525_);
  and (_08437_, _08126_, _08436_);
  nor (_08438_, _08436_, _06677_);
  nor (_08439_, _08438_, _08437_);
  nor (_08440_, _08439_, _08125_);
  nor (_08441_, _08040_, _06677_);
  nor (_08442_, _08441_, _08045_);
  not (_08443_, _08442_);
  nor (_08444_, _08443_, _08440_);
  nor (_08445_, _08444_, _07699_);
  nand (_08446_, _08445_, _08434_);
  nand (_08447_, _08446_, _08387_);
  and (_06641_, _08447_, _06989_);
  nand (_08448_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nand (_08449_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_08450_, _08449_, _08448_);
  nand (_08451_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_08452_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_08453_, _08452_, _08451_);
  nand (_08454_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_08455_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_08456_, _08455_, _08454_);
  and (_08457_, _08456_, _08453_);
  nand (_08458_, _08457_, _08450_);
  nand (_08459_, _08458_, _07330_);
  nand (_08460_, _08459_, _07328_);
  nor (_08461_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _07328_);
  not (_08462_, _08461_);
  and (_08463_, _08462_, _08460_);
  and (_06671_, _08463_, _06989_);
  nor (_08464_, _07325_, _06550_);
  and (_08465_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_08466_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_08467_, _08466_, _08465_);
  and (_08468_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_08469_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_08470_, _08469_, _08468_);
  and (_08471_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_08472_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_08473_, _08472_, _08471_);
  and (_08474_, _08473_, _08470_);
  and (_08475_, _08474_, _08467_);
  and (_08476_, _07325_, _07330_);
  not (_08477_, _08476_);
  nor (_08478_, _08477_, _08475_);
  nor (_08479_, _08478_, _08464_);
  nor (_06674_, _08479_, rst);
  and (_06825_, _07360_, _06989_);
  and (_08480_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_08481_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_08482_, _08481_, _08480_);
  nand (_08483_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_08484_, _08483_, _07330_);
  and (_08485_, _08484_, _08482_);
  and (_08486_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not (_08487_, _08486_);
  and (_08488_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_08489_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_08490_, _08489_, _08488_);
  and (_08491_, _08490_, _08487_);
  nand (_08492_, _08491_, _08485_);
  or (_08493_, _08492_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_08494_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _07328_);
  not (_08495_, _08494_);
  and (_08496_, _08495_, _08493_);
  and (_06827_, _08496_, _06989_);
  and (_08497_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_08498_, _08497_);
  nand (_08499_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand (_08500_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_08501_, _08500_, _08499_);
  nand (_08502_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nand (_08503_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and (_08504_, _08503_, _08502_);
  and (_08505_, _08504_, _08501_);
  and (_08506_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_08507_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_08508_, _08507_, _08506_);
  and (_08509_, _08508_, _08505_);
  or (_08510_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_08511_, _08510_, _08509_);
  and (_08512_, _08511_, _08498_);
  nor (_06829_, _08512_, rst);
  nand (_08513_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nand (_08514_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_08515_, _08514_, _08513_);
  nand (_08516_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_08517_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_08518_, _08517_, _08516_);
  nand (_08519_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_08520_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_08522_, _08520_, _08519_);
  and (_08523_, _08522_, _08518_);
  nand (_08524_, _08523_, _08515_);
  nand (_08525_, _08524_, _07330_);
  nand (_08526_, _08525_, _07328_);
  nor (_08527_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _07328_);
  not (_08528_, _08527_);
  and (_08529_, _08528_, _08526_);
  and (_06831_, _08529_, _06989_);
  and (_08530_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_08531_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_08532_, _08531_, _08530_);
  and (_08533_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  not (_08534_, _08533_);
  and (_08535_, _08534_, _08532_);
  and (_08536_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_08537_, _08536_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_08538_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_08539_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_08540_, _08539_, _08538_);
  and (_08541_, _08540_, _08537_);
  and (_08542_, _08541_, _08535_);
  and (_08543_, _08542_, _07328_);
  nor (_08544_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _07328_);
  nor (_08545_, _08544_, _08543_);
  and (_06833_, _08545_, _06989_);
  nand (_08546_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nand (_08547_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_08548_, _08547_, _08546_);
  nand (_08549_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_08550_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_08551_, _08550_, _08549_);
  nand (_08552_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand (_08553_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and (_08554_, _08553_, _08552_);
  and (_08555_, _08554_, _08551_);
  nand (_08556_, _08555_, _08548_);
  and (_08557_, _08556_, _07330_);
  or (_08558_, _08557_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_08559_, _07328_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  not (_08560_, _08559_);
  and (_08561_, _08560_, _08558_);
  and (_06836_, _08561_, _06989_);
  nand (_08562_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nand (_08563_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_08564_, _08563_, _08562_);
  nand (_08565_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_08566_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_08567_, _08566_, _08565_);
  nand (_08568_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand (_08569_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_08570_, _08569_, _08568_);
  and (_08571_, _08570_, _08567_);
  and (_08572_, _08571_, _08564_);
  or (_08573_, _08572_, _08510_);
  and (_08574_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_08575_, _08574_);
  and (_08576_, _08575_, _08573_);
  nor (_06838_, _08576_, rst);
  nor (_08577_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_08578_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08579_, _08578_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor (_08580_, _08579_, _08577_);
  nor (_08581_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_08582_, _08578_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nor (_08583_, _08582_, _08581_);
  not (_08584_, _08583_);
  not (_08585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_08586_, _07493_, _08585_);
  and (_08587_, _07493_, _08585_);
  nor (_08588_, _08587_, _08586_);
  nor (_08589_, _08588_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08590_, _08578_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor (_08591_, _08590_, _08589_);
  and (_08592_, _08591_, _08584_);
  not (_08593_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor (_08594_, _08586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_08595_, _08586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_08596_, _08595_, _08594_);
  nor (_08597_, _08596_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08598_, _08578_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor (_08599_, _08598_, _08597_);
  and (_08600_, _08599_, _08593_);
  nor (_08601_, _08599_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08602_, _08601_, _08600_);
  not (_08603_, _08602_);
  nand (_08604_, _08603_, _08592_);
  and (_08605_, _08604_, _08580_);
  nor (_08606_, _08591_, _08584_);
  not (_08607_, _08606_);
  not (_08608_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_08609_, _08599_, _08608_);
  and (_08610_, _08599_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08611_, _08610_, _08609_);
  nor (_08612_, _08611_, _08607_);
  and (_08613_, _08591_, _08583_);
  not (_08614_, _08613_);
  not (_08615_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_08616_, _08599_, _08615_);
  and (_08617_, _08599_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_08618_, _08617_, _08616_);
  nor (_08619_, _08618_, _08614_);
  nor (_08620_, _08619_, _08612_);
  not (_08621_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08622_, _08599_, _08621_);
  nor (_08623_, _08591_, _08583_);
  nor (_08624_, _08599_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_08625_, _08624_);
  nand (_08626_, _08625_, _08623_);
  or (_08627_, _08626_, _08622_);
  and (_08628_, _08627_, _08620_);
  and (_08629_, _08628_, _08605_);
  and (_08630_, _08599_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08631_, _08630_, _08606_);
  not (_08632_, _08599_);
  and (_08633_, _08606_, _08632_);
  and (_08634_, _08633_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08635_, _08634_, _08580_);
  or (_08636_, _08635_, _08631_);
  not (_08637_, _08623_);
  and (_08638_, _08599_, \oc8051_symbolic_cxrom1.regvalid [8]);
  not (_08639_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_08640_, _08599_, _08639_);
  nor (_08641_, _08640_, _08638_);
  nor (_08642_, _08641_, _08637_);
  and (_08643_, _08632_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08644_, _08599_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_08645_, _08644_, _08643_);
  nor (_08646_, _08645_, _08614_);
  not (_08647_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_08648_, _08599_, _08647_);
  nor (_08649_, _08599_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_08650_, _08649_, _08648_);
  not (_08651_, _08650_);
  and (_08652_, _08651_, _08592_);
  or (_08653_, _08652_, _08646_);
  or (_08654_, _08653_, _08642_);
  nor (_08655_, _08654_, _08636_);
  nor (_08656_, _08655_, _08629_);
  not (_08657_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_08658_, _08580_, _08657_);
  or (_08659_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_08661_, _08659_, _08658_);
  and (_08662_, _08661_, _08613_);
  not (_08663_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_08664_, _08580_, _08663_);
  or (_08665_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_08666_, _08665_, _08664_);
  and (_08667_, _08666_, _08606_);
  or (_08668_, _08667_, _08662_);
  not (_08669_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_08670_, _08580_, _08669_);
  or (_08671_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_08672_, _08671_, _08670_);
  and (_08673_, _08672_, _08592_);
  not (_08674_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_08675_, _08580_, _08674_);
  or (_08676_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_08677_, _08676_, _08675_);
  and (_08678_, _08677_, _08623_);
  or (_08679_, _08678_, _08673_);
  or (_08680_, _08679_, _08668_);
  and (_08681_, _08680_, _08599_);
  not (_08682_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_08683_, _08580_, _08682_);
  or (_08684_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_08685_, _08684_, _08683_);
  and (_08686_, _08685_, _08606_);
  not (_08687_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_08688_, _08580_, _08687_);
  or (_08689_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_08690_, _08689_, _08688_);
  and (_08691_, _08690_, _08613_);
  or (_08692_, _08691_, _08686_);
  not (_08693_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_08694_, _08580_, _08693_);
  or (_08695_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_08696_, _08695_, _08694_);
  and (_08697_, _08696_, _08592_);
  not (_08698_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_08699_, _08580_, _08698_);
  or (_08700_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_08701_, _08700_, _08699_);
  and (_08702_, _08701_, _08623_);
  or (_08703_, _08702_, _08697_);
  or (_08704_, _08703_, _08692_);
  and (_08705_, _08704_, _08632_);
  or (_08706_, _08705_, _08681_);
  and (_08707_, _08706_, _08656_);
  not (_08708_, _08656_);
  and (_08709_, _08708_, word_in[7]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _08709_, _08707_);
  not (_08710_, _08580_);
  and (_08711_, _08583_, _08710_);
  not (_08712_, _08711_);
  and (_08713_, _08583_, _08580_);
  and (_08714_, _08713_, _08591_);
  nor (_08715_, _08713_, _08591_);
  nor (_08716_, _08715_, _08714_);
  not (_08717_, _08716_);
  nor (_08718_, _08717_, _08618_);
  nor (_08719_, _08714_, _08632_);
  not (_08720_, _08591_);
  nor (_08721_, _08599_, _08720_);
  and (_08722_, _08713_, _08721_);
  nor (_08723_, _08722_, _08719_);
  and (_08724_, _08723_, _08717_);
  and (_08725_, _08724_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_08726_, _08723_, _08716_);
  and (_08727_, _08726_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08728_, _08727_, _08725_);
  nor (_08729_, _08728_, _08718_);
  nor (_08730_, _08729_, _08712_);
  nor (_08731_, _08583_, _08580_);
  not (_08732_, _08731_);
  nor (_08733_, _08717_, _08602_);
  and (_08734_, _08724_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_08735_, _08726_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_08736_, _08735_, _08734_);
  nor (_08737_, _08736_, _08733_);
  nor (_08738_, _08737_, _08732_);
  nor (_08739_, _08738_, _08730_);
  and (_08740_, _08584_, _08580_);
  not (_08741_, _08740_);
  nor (_08742_, _08717_, _08645_);
  and (_08743_, _08724_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_08744_, _08726_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08745_, _08744_, _08743_);
  nor (_08746_, _08745_, _08742_);
  nor (_08747_, _08746_, _08741_);
  not (_08748_, _08713_);
  nor (_08750_, _08717_, _08650_);
  and (_08751_, _08724_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_08752_, _08726_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_08753_, _08752_, _08751_);
  nor (_08754_, _08753_, _08750_);
  nor (_08755_, _08754_, _08748_);
  nor (_08756_, _08755_, _08747_);
  and (_08757_, _08756_, _08739_);
  or (_08758_, _08713_, _08731_);
  not (_08759_, _08758_);
  not (_08760_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_08761_, _08580_, _08760_);
  or (_08762_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_08763_, _08762_, _08761_);
  and (_08764_, _08763_, _08759_);
  not (_08765_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_08766_, _08580_, _08765_);
  or (_08767_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_08768_, _08767_, _08766_);
  and (_08769_, _08768_, _08758_);
  or (_08770_, _08769_, _08764_);
  and (_08771_, _08770_, _08726_);
  not (_08772_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_08773_, _08580_, _08772_);
  or (_08774_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_08775_, _08774_, _08773_);
  and (_08776_, _08775_, _08759_);
  not (_08777_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_08778_, _08580_, _08777_);
  or (_08779_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_08780_, _08779_, _08778_);
  and (_08781_, _08780_, _08758_);
  or (_08782_, _08781_, _08776_);
  and (_08783_, _08782_, _08724_);
  and (_08784_, _08716_, _08632_);
  not (_08785_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_08786_, _08580_, _08785_);
  or (_08787_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_08788_, _08787_, _08786_);
  and (_08789_, _08788_, _08759_);
  not (_08790_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_08791_, _08580_, _08790_);
  or (_08792_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_08793_, _08792_, _08791_);
  and (_08794_, _08793_, _08758_);
  or (_08795_, _08794_, _08789_);
  and (_08796_, _08795_, _08784_);
  and (_08797_, _08716_, _08599_);
  not (_08798_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_08799_, _08580_, _08798_);
  or (_08800_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_08801_, _08800_, _08799_);
  and (_08802_, _08801_, _08759_);
  not (_08803_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_08804_, _08580_, _08803_);
  or (_08805_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_08806_, _08805_, _08804_);
  and (_08807_, _08806_, _08758_);
  or (_08808_, _08807_, _08802_);
  and (_08810_, _08808_, _08797_);
  or (_08811_, _08810_, _08796_);
  or (_08812_, _08811_, _08783_);
  nor (_08813_, _08812_, _08771_);
  nor (_08814_, _08813_, _08757_);
  and (_08815_, _08757_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _08815_, _08814_);
  nor (_08816_, _08613_, _08623_);
  not (_08817_, _08816_);
  nor (_08818_, _08817_, _08602_);
  and (_08819_, _08613_, _08599_);
  nor (_08820_, _08613_, _08599_);
  nor (_08821_, _08820_, _08819_);
  and (_08822_, _08821_, _08817_);
  and (_08823_, _08822_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_08824_, _08821_, _08816_);
  and (_08825_, _08824_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08826_, _08825_, _08823_);
  nor (_08827_, _08826_, _08818_);
  nor (_08828_, _08827_, _08748_);
  nor (_08829_, _08817_, _08618_);
  and (_08830_, _08824_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_08831_, _08822_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_08832_, _08831_, _08830_);
  nor (_08833_, _08832_, _08829_);
  nor (_08834_, _08833_, _08741_);
  nor (_08835_, _08834_, _08828_);
  nor (_08836_, _08817_, _08645_);
  and (_08837_, _08824_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_08838_, _08822_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_08839_, _08838_, _08837_);
  nor (_08841_, _08839_, _08836_);
  nor (_08842_, _08841_, _08732_);
  nor (_08843_, _08817_, _08650_);
  and (_08844_, _08822_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08845_, _08824_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_08846_, _08845_, _08844_);
  nor (_08847_, _08846_, _08843_);
  nor (_08848_, _08847_, _08712_);
  nor (_08849_, _08848_, _08842_);
  and (_08850_, _08849_, _08835_);
  and (_08851_, _08850_, word_in[23]);
  and (_08852_, _08696_, _08606_);
  and (_08853_, _08685_, _08623_);
  or (_08854_, _08853_, _08852_);
  and (_08855_, _08690_, _08592_);
  and (_08856_, _08701_, _08613_);
  or (_08857_, _08856_, _08855_);
  or (_08858_, _08857_, _08854_);
  or (_08859_, _08858_, _08821_);
  not (_08860_, _08821_);
  and (_08861_, _08672_, _08606_);
  and (_08862_, _08677_, _08632_);
  or (_08863_, _08862_, _08861_);
  and (_08864_, _08661_, _08592_);
  and (_08865_, _08666_, _08623_);
  or (_08866_, _08865_, _08864_);
  or (_08867_, _08866_, _08863_);
  or (_08868_, _08867_, _08860_);
  nand (_08869_, _08868_, _08859_);
  nor (_08870_, _08869_, _08850_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _08870_, _08851_);
  nand (_08871_, _08732_, _08591_);
  nor (_08872_, _08732_, _08591_);
  not (_08873_, _08872_);
  and (_08874_, _08873_, _08871_);
  not (_08875_, _08874_);
  nor (_08876_, _08875_, _08618_);
  nor (_08877_, _08871_, _08599_);
  and (_08878_, _08871_, _08599_);
  nor (_08879_, _08878_, _08877_);
  nor (_08880_, _08879_, _08874_);
  and (_08881_, _08880_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08882_, _08881_, _08876_);
  nor (_08883_, _08882_, _08732_);
  nor (_08884_, _08650_, _08875_);
  and (_08885_, _08879_, _08875_);
  and (_08886_, _08885_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_08887_, _08886_, _08884_);
  and (_08888_, _08887_, _08740_);
  and (_08889_, _08872_, _08609_);
  and (_08890_, _08740_, _08721_);
  and (_08891_, _08890_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_08892_, _08891_, _08889_);
  or (_08893_, _08892_, _08888_);
  or (_08894_, _08893_, _08883_);
  nor (_08895_, _08645_, _08875_);
  and (_08896_, _08880_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08897_, _08885_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08898_, _08897_, _08896_);
  nor (_08899_, _08898_, _08895_);
  nor (_08900_, _08899_, _08748_);
  nor (_08901_, _08875_, _08602_);
  and (_08902_, _08885_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_08903_, _08880_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_08904_, _08903_, _08902_);
  nor (_08905_, _08904_, _08901_);
  nor (_08906_, _08905_, _08712_);
  or (_08907_, _08906_, _08900_);
  nor (_08908_, _08907_, _08894_);
  and (_08909_, _08768_, _08759_);
  and (_08910_, _08763_, _08758_);
  or (_08911_, _08910_, _08909_);
  and (_08912_, _08911_, _08880_);
  and (_08913_, _08780_, _08759_);
  and (_08914_, _08775_, _08758_);
  or (_08915_, _08914_, _08913_);
  and (_08916_, _08915_, _08885_);
  and (_08917_, _08874_, _08632_);
  and (_08918_, _08793_, _08759_);
  and (_08919_, _08788_, _08758_);
  or (_08920_, _08919_, _08918_);
  and (_08921_, _08920_, _08917_);
  and (_08922_, _08806_, _08759_);
  and (_08923_, _08801_, _08758_);
  or (_08924_, _08923_, _08922_);
  and (_08925_, _08878_, _08873_);
  and (_08926_, _08925_, _08924_);
  or (_08927_, _08926_, _08921_);
  or (_08928_, _08927_, _08916_);
  nor (_08929_, _08928_, _08912_);
  nor (_08930_, _08929_, _08908_);
  and (_08931_, _08908_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08931_, _08930_);
  and (_08932_, _08599_, _08591_);
  or (_08933_, _08932_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_07163_, _08933_, _06989_);
  and (_08934_, _08932_, _08731_);
  and (_08935_, _08908_, _06989_);
  and (_08936_, _08935_, _08934_);
  and (_08937_, _08850_, _06989_);
  and (_08938_, _08937_, _08816_);
  and (_08939_, _08938_, _08821_);
  and (_08940_, _08939_, _08740_);
  not (_08941_, _08940_);
  and (_08942_, _08937_, word_in[23]);
  or (_08943_, _08942_, _08941_);
  and (_08944_, _08757_, _06989_);
  and (_08945_, _08944_, _08711_);
  and (_08946_, _08945_, _08797_);
  and (_08947_, _08629_, _06989_);
  and (_08948_, _08947_, _08583_);
  nor (_08949_, _08656_, rst);
  and (_08950_, _08949_, _08932_);
  and (_08951_, _08950_, _08948_);
  nor (_08952_, _08951_, _08657_);
  and (_08953_, _08949_, word_in[7]);
  and (_08954_, _08953_, _08951_);
  or (_08955_, _08954_, _08952_);
  or (_08956_, _08955_, _08946_);
  not (_08957_, _08946_);
  or (_08958_, _08957_, word_in[15]);
  and (_08959_, _08958_, _08956_);
  or (_08960_, _08959_, _08940_);
  and (_08961_, _08960_, _08943_);
  or (_08963_, _08961_, _08936_);
  not (_08964_, _08936_);
  or (_08965_, _08964_, word_in[31]);
  and (_07192_, _08965_, _08963_);
  or (_08966_, _08885_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_07214_, _08966_, _06989_);
  not (_08967_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand (_08968_, _08623_, _08632_);
  nand (_08969_, _08968_, _08967_);
  or (_08970_, _08969_, _08819_);
  and (_07241_, _08970_, _06989_);
  and (_08971_, _08714_, _08599_);
  not (_08972_, _08971_);
  and (_08973_, _08968_, _08972_);
  not (_08974_, _08973_);
  and (_08975_, _08740_, _08917_);
  and (_08976_, _08711_, _08917_);
  nor (_08977_, _08976_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_08978_, _08977_, _08975_);
  or (_08979_, _08978_, _08974_);
  and (_07280_, _08979_, _06989_);
  not (_08980_, _08724_);
  and (_08981_, _08713_, _08917_);
  or (_08982_, _08981_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_08983_, _08982_, _08980_);
  and (_08984_, _08609_, _08623_);
  or (_08985_, _08984_, _08976_);
  or (_08986_, _08985_, _08983_);
  and (_08987_, _08986_, _08973_);
  not (_08988_, _08968_);
  and (_08989_, _08982_, _08971_);
  or (_08990_, _08989_, _08988_);
  or (_08991_, _08990_, _08987_);
  and (_07329_, _08991_, _06989_);
  not (_08992_, _07090_);
  nand (_08993_, _07086_, _06975_);
  nor (_08994_, _08993_, _08992_);
  not (_08995_, _07128_);
  nor (_08996_, _08993_, _08995_);
  nor (_08997_, _08996_, _08994_);
  and (_08998_, _08997_, _07127_);
  or (_08999_, _08998_, _06982_);
  and (_09000_, _08999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  not (_09001_, _07126_);
  nand (_09002_, _08997_, _09001_);
  and (_09003_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_09004_, _09003_, _09002_);
  nor (_09005_, _07035_, _06728_);
  not (_09006_, _09005_);
  and (_09007_, _09006_, _08000_);
  and (_09008_, _09007_, _08018_);
  not (_09009_, _09008_);
  and (_09010_, _07123_, _06981_);
  and (_09011_, _09010_, _09009_);
  or (_09012_, _09011_, _09004_);
  or (_09013_, _09012_, _09000_);
  and (_07336_, _09013_, _06989_);
  or (_09014_, _08975_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_09015_, _09014_, _08974_);
  and (_09016_, _08721_, _08731_);
  or (_09017_, _09016_, _08981_);
  or (_09018_, _09017_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_09019_, _09018_, _08980_);
  or (_09020_, _09019_, _09015_);
  or (_09021_, _09020_, _08976_);
  and (_07388_, _09021_, _06989_);
  and (_09022_, _06478_, _06463_);
  and (_09023_, _09022_, _08037_);
  and (_09024_, _09023_, _06539_);
  nand (_09025_, _09024_, _06968_);
  or (_09026_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_09027_, _09026_, _06485_);
  and (_09028_, _09027_, _09025_);
  and (_09029_, _07706_, _07453_);
  and (_09030_, _09029_, _07125_);
  not (_09031_, _09030_);
  nor (_09032_, _09031_, _07040_);
  not (_09033_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor (_09034_, _09030_, _09033_);
  or (_09035_, _09034_, _09032_);
  and (_09036_, _09035_, _06983_);
  nor (_09037_, _06484_, _09033_);
  or (_09038_, _09037_, rst);
  or (_09039_, _09038_, _09036_);
  or (_07448_, _09039_, _09028_);
  and (_09040_, _08872_, _08632_);
  nor (_09041_, _09040_, _08917_);
  not (_09042_, _08820_);
  or (_09043_, _09042_, _09017_);
  and (_09044_, _09043_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_09045_, _08976_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_09046_, _09045_, _08890_);
  or (_09048_, _09046_, _09044_);
  and (_09049_, _09048_, _09041_);
  and (_09050_, _08988_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_09051_, _09050_, _08976_);
  or (_09052_, _09051_, _09016_);
  or (_09053_, _09052_, _08981_);
  or (_09054_, _09053_, _09049_);
  and (_07451_, _09054_, _06989_);
  or (_09055_, _08719_, _08877_);
  and (_09056_, _08932_, _08711_);
  or (_09057_, _08821_, _09056_);
  and (_09058_, _08711_, _08721_);
  or (_09059_, _09058_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_09060_, _09059_, _09057_);
  and (_09061_, _09017_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_09062_, _09061_, _08890_);
  or (_09063_, _09062_, _09060_);
  and (_09064_, _09063_, _09055_);
  and (_09065_, _09059_, _08971_);
  and (_09066_, _08715_, _08643_);
  or (_09067_, _09066_, _08981_);
  or (_09068_, _09067_, _09016_);
  or (_09069_, _09068_, _09065_);
  or (_09070_, _09069_, _09064_);
  and (_07503_, _09070_, _06989_);
  and (_09071_, _07704_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_09072_, _06983_, _06447_);
  nor (_09073_, _06537_, _06514_);
  and (_09074_, _09073_, _06525_);
  and (_09075_, _07454_, _09074_);
  and (_09076_, _09075_, _09072_);
  nor (_09077_, _09076_, _09071_);
  or (_09078_, _09077_, _08123_);
  not (_09079_, _09077_);
  or (_09080_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_09081_, _09080_, _06989_);
  and (_07578_, _09081_, _09078_);
  nor (_09082_, _07793_, _07725_);
  or (_09083_, _09082_, _07794_);
  nand (_09084_, _09083_, _07814_);
  or (_09085_, _07814_, _07722_);
  and (_09086_, _09085_, _09084_);
  nand (_09087_, _09086_, _07024_);
  and (_09088_, _08227_, _08224_);
  and (_09089_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  nand (_09090_, _09089_, _09088_);
  or (_09091_, _09089_, _09088_);
  and (_09092_, _09091_, _09090_);
  nand (_09093_, _09092_, _07027_);
  nor (_09094_, _06826_, _06792_);
  not (_09095_, _09094_);
  nor (_09096_, _06828_, _06549_);
  and (_09097_, _09096_, _09095_);
  not (_09098_, _09097_);
  nor (_09099_, _06896_, _06861_);
  nor (_09100_, _09099_, _06897_);
  nor (_09101_, _09100_, _06846_);
  and (_09102_, _06810_, _06883_);
  not (_09103_, _09102_);
  and (_09104_, _06816_, _06778_);
  nor (_09105_, _09104_, _06992_);
  and (_09106_, _09105_, _09103_);
  or (_09107_, _07008_, _06902_);
  and (_09108_, _09107_, _07010_);
  and (_09109_, _07000_, _07096_);
  nor (_09110_, _09109_, _06810_);
  or (_09111_, _09110_, _07001_);
  and (_09112_, _09111_, _06778_);
  or (_09113_, _09112_, _09108_);
  and (_09114_, _09113_, _06997_);
  nor (_09115_, _09114_, _09106_);
  nor (_09116_, _08247_, _06810_);
  and (_09117_, _08247_, _06810_);
  nor (_09118_, _09117_, _09116_);
  nor (_09119_, _09118_, _06918_);
  and (_09120_, _06951_, _06902_);
  not (_09121_, _09120_);
  or (_09123_, _07031_, _06586_);
  nand (_09124_, _07032_, _06616_);
  and (_09125_, _09124_, _09123_);
  and (_09126_, _09125_, _09121_);
  and (_09127_, _06942_, _06819_);
  and (_09128_, _06933_, _06817_);
  nor (_09129_, _07017_, _06818_);
  and (_09130_, _06954_, _06810_);
  or (_09131_, _09130_, _09129_);
  or (_09132_, _09131_, _09128_);
  nor (_09133_, _09132_, _09127_);
  and (_09134_, _09133_, _09126_);
  not (_09136_, _09134_);
  nor (_09138_, _09136_, _09119_);
  and (_09139_, _09138_, _09115_);
  not (_09140_, _09139_);
  nor (_09142_, _09140_, _09101_);
  and (_09143_, _09142_, _09098_);
  and (_09144_, _09143_, _09093_);
  and (_09145_, _09144_, _09087_);
  nand (_09146_, _09145_, _09079_);
  or (_09147_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_09148_, _09147_, _06989_);
  and (_07581_, _09148_, _09146_);
  or (_09149_, _09077_, _08268_);
  or (_09150_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_09151_, _09150_, _06989_);
  and (_07584_, _09151_, _09149_);
  or (_09153_, _09077_, _08346_);
  or (_09155_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_09156_, _09155_, _06989_);
  and (_07592_, _09156_, _09153_);
  or (_09157_, _08714_, _08599_);
  nor (_09158_, _08599_, _08710_);
  or (_09159_, _09158_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_09160_, _09159_, _09042_);
  and (_09161_, _08616_, _08614_);
  or (_09162_, _09161_, _09160_);
  and (_09163_, _09162_, _09157_);
  and (_09164_, _08874_, _08616_);
  and (_09165_, _09040_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_09166_, _09165_, _09016_);
  or (_09167_, _09166_, _09164_);
  or (_09168_, _09167_, _08890_);
  or (_09169_, _09168_, _09058_);
  or (_09170_, _09169_, _09163_);
  and (_07599_, _09170_, _06989_);
  or (_09171_, _09077_, _08433_);
  or (_09172_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_09173_, _09172_, _06989_);
  and (_07616_, _09173_, _09171_);
  and (_09174_, _07781_, _07771_);
  not (_09175_, _09174_);
  and (_09176_, _09175_, _07782_);
  or (_09177_, _09176_, _07810_);
  or (_09178_, _07814_, _07778_);
  and (_09179_, _09178_, _09177_);
  nand (_09180_, _09179_, _07024_);
  or (_09181_, _08398_, _08216_);
  and (_09182_, _09181_, _08399_);
  nand (_09183_, _09182_, _07027_);
  nor (_09184_, _06784_, _06782_);
  not (_09185_, _09184_);
  nor (_09186_, _06785_, _06549_);
  and (_09187_, _09186_, _09185_);
  not (_09188_, _09187_);
  nor (_09189_, _06885_, _06879_);
  nor (_09190_, _09189_, _06886_);
  nor (_09191_, _09190_, _06846_);
  not (_09192_, _09191_);
  and (_09193_, _06991_, _06706_);
  nor (_09194_, _07004_, _06778_);
  nor (_09195_, _08012_, _06883_);
  nor (_09196_, _09195_, _09194_);
  and (_09197_, _09196_, _06700_);
  not (_09198_, _09197_);
  nor (_09199_, _09196_, _06700_);
  nor (_09200_, _09199_, _07101_);
  and (_09201_, _09200_, _09198_);
  nor (_09202_, _09201_, _09193_);
  and (_09203_, _06910_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  not (_09204_, _06700_);
  nor (_09205_, _07987_, _09204_);
  nor (_09206_, _09205_, _09203_);
  nor (_09207_, _09206_, _06918_);
  nor (_09208_, _07017_, _06708_);
  and (_09209_, _06942_, _06709_);
  nor (_09210_, _09209_, _09208_);
  and (_09211_, _06933_, _06707_);
  and (_09212_, _06954_, _09204_);
  nor (_09213_, _09212_, _09211_);
  or (_09214_, _07031_, _06673_);
  nor (_09215_, _08001_, _06728_);
  and (_09216_, _06951_, _06700_);
  nor (_09217_, _09216_, _09215_);
  and (_09218_, _09217_, _09214_);
  and (_09219_, _09218_, _09213_);
  and (_09220_, _09219_, _09210_);
  not (_09221_, _09220_);
  nor (_09222_, _09221_, _09207_);
  and (_09223_, _09222_, _09202_);
  and (_09224_, _09223_, _09192_);
  and (_09225_, _09224_, _09188_);
  and (_09226_, _09225_, _09183_);
  and (_09227_, _09226_, _09180_);
  nand (_09228_, _09227_, _09079_);
  or (_09229_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_09230_, _09229_, _06989_);
  and (_07620_, _09230_, _09228_);
  or (_09231_, _09077_, _08030_);
  or (_09232_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_09233_, _09232_, _06989_);
  and (_07635_, _09233_, _09231_);
  not (_09234_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_09236_, _08877_, _09234_);
  or (_09237_, _09236_, _08880_);
  and (_07673_, _09237_, _06989_);
  and (_09239_, _07454_, _09072_);
  nand (_09240_, _09239_, _08436_);
  nor (_09241_, _09240_, _09145_);
  and (_09242_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_09244_, _09242_, _09071_);
  or (_09245_, _09244_, _09241_);
  and (_09246_, _06951_, _06850_);
  and (_09248_, _06958_, _06700_);
  and (_09249_, _08148_, _06853_);
  and (_09250_, _09249_, _06623_);
  or (_09252_, _09250_, _06778_);
  and (_09253_, _08154_, _06622_);
  or (_09255_, _09253_, _06883_);
  and (_09256_, _09255_, _09252_);
  and (_09258_, _09256_, _06816_);
  nor (_09259_, _09256_, _06816_);
  or (_09260_, _09259_, _09258_);
  and (_09261_, _09260_, _06997_);
  nor (_09262_, _06816_, _06778_);
  nor (_09263_, _06810_, _06883_);
  or (_09264_, _09263_, _09262_);
  and (_09265_, _09264_, _06991_);
  or (_09266_, _09265_, _09261_);
  or (_09267_, _09266_, _09248_);
  and (_09268_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_09269_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_09270_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_09271_, _09270_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_09272_, _09271_, _09269_);
  nor (_09273_, _09272_, _08191_);
  not (_09274_, _09273_);
  and (_09275_, _09272_, _08191_);
  nor (_09276_, _09275_, _06549_);
  and (_09277_, _09276_, _09274_);
  and (_09278_, _07956_, _07926_);
  not (_09279_, _09278_);
  and (_09280_, _09279_, _07957_);
  and (_09281_, _09280_, _07027_);
  or (_09282_, _09281_, _09277_);
  or (_09283_, _09282_, _09268_);
  or (_09284_, _09283_, _09267_);
  nor (_09285_, _09284_, _09246_);
  nand (_09286_, _09285_, _09071_);
  and (_09287_, _09286_, _06989_);
  and (_07764_, _09287_, _09245_);
  and (_09288_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_09289_, _07124_, _08435_);
  and (_09290_, _09289_, _07454_);
  and (_09291_, _09290_, _06484_);
  and (_09292_, _09291_, _06980_);
  and (_09293_, _09292_, _08268_);
  or (_09294_, _09293_, _09288_);
  or (_09295_, _09294_, _09071_);
  nand (_09296_, _09071_, _08202_);
  and (_09297_, _09296_, _06989_);
  and (_07767_, _09297_, _09295_);
  and (_09298_, _08820_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_09299_, _08872_, _08599_);
  and (_09300_, _08719_, _08873_);
  and (_09301_, _08925_, _08740_);
  nor (_09302_, _08820_, _08621_);
  or (_09303_, _09302_, _09301_);
  and (_09304_, _09303_, _09300_);
  or (_09306_, _09304_, _09299_);
  and (_09307_, _09303_, _08971_);
  or (_09308_, _09307_, _09058_);
  or (_09309_, _09308_, _08722_);
  or (_09310_, _09309_, _09306_);
  or (_09311_, _09310_, _09298_);
  and (_07773_, _09311_, _06989_);
  and (_09312_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_09313_, _09292_, _08346_);
  or (_09314_, _09313_, _09312_);
  or (_09315_, _09314_, _09071_);
  nand (_09316_, _09071_, _08307_);
  and (_09317_, _09316_, _06989_);
  and (_07785_, _09317_, _09315_);
  and (_09318_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and (_09319_, _09292_, _08433_);
  or (_09320_, _09319_, _09318_);
  or (_09321_, _09320_, _09071_);
  nand (_09322_, _09071_, _08385_);
  and (_09323_, _09322_, _06989_);
  and (_07806_, _09323_, _09321_);
  nor (_09324_, _09240_, _09227_);
  and (_09325_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_09326_, _09325_, _09071_);
  or (_09327_, _09326_, _09324_);
  and (_09329_, _06951_, _06706_);
  and (_09330_, _06958_, _06902_);
  nor (_09331_, _08146_, _06778_);
  nor (_09332_, _08361_, _06883_);
  nor (_09333_, _09332_, _09331_);
  nor (_09334_, _09333_, _06706_);
  and (_09336_, _09333_, _06706_);
  nor (_09337_, _09336_, _09334_);
  and (_09338_, _09337_, _06997_);
  and (_09339_, _06991_, _06700_);
  or (_09340_, _09339_, _09338_);
  or (_09341_, _09340_, _09330_);
  and (_09342_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_09343_, _08177_, _07657_);
  nor (_09344_, _09343_, _08178_);
  and (_09345_, _09344_, _06548_);
  and (_09347_, _07945_, _07943_);
  not (_09348_, _09347_);
  and (_09349_, _09348_, _07946_);
  and (_09350_, _09349_, _07027_);
  or (_09352_, _09350_, _09345_);
  or (_09353_, _09352_, _09342_);
  or (_09355_, _09353_, _09341_);
  nor (_09356_, _09355_, _09329_);
  nand (_09357_, _09356_, _09071_);
  and (_09358_, _09357_, _06989_);
  and (_07820_, _09358_, _09327_);
  and (_09359_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and (_09360_, _09292_, _08030_);
  or (_09361_, _09360_, _09359_);
  or (_09362_, _09361_, _09071_);
  nand (_09363_, _09071_, _07696_);
  and (_09364_, _09363_, _06989_);
  and (_07829_, _09364_, _09362_);
  and (_09365_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_09366_, _09292_, _08123_);
  or (_09367_, _09366_, _09365_);
  or (_09368_, _09367_, _09071_);
  not (_09369_, _09071_);
  or (_09370_, _09369_, _08075_);
  and (_09371_, _09370_, _06989_);
  and (_07834_, _09371_, _09368_);
  and (_09372_, _08711_, _08878_);
  not (_09373_, _08715_);
  and (_09374_, _09373_, _08630_);
  or (_09375_, _09374_, _09372_);
  or (_09376_, _09058_, _08988_);
  and (_09377_, _09376_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_09378_, _08816_, _08632_);
  and (_09379_, _09378_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_09380_, _09379_, _08722_);
  or (_09381_, _09380_, _09377_);
  or (_09382_, _09381_, _09301_);
  or (_09383_, _09382_, _09299_);
  or (_09384_, _09383_, _09375_);
  and (_07869_, _09384_, _06989_);
  nand (_09385_, _08512_, _07326_);
  nor (_09386_, _07325_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_09387_, _09386_, _07362_);
  and (_09388_, _09387_, _09385_);
  and (_07933_, _09388_, _06989_);
  not (_09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_09390_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_09391_, _09390_, _06989_);
  nor (_09392_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_09393_, _09392_);
  and (_09394_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_09395_, _09394_, _09393_);
  not (_09396_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_09397_, _09396_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not (_09398_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_09399_, _09398_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_09400_, _09399_, _09397_);
  not (_09401_, _09400_);
  and (_09402_, _09401_, _09395_);
  and (_09403_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_09404_, _09403_, _09393_);
  not (_09405_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_09406_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _09405_);
  not (_09407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_09408_, _09392_, _09407_);
  and (_09409_, _09408_, _09406_);
  nor (_09410_, _09409_, _09395_);
  not (_09411_, _09410_);
  nor (_09412_, _09411_, _09404_);
  nor (_09413_, _09412_, _09402_);
  and (_09414_, _09392_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_09415_, _09414_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or (_09416_, _09415_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_09417_, _09416_, _09413_);
  and (_09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _06989_);
  and (_09419_, _09400_, _09395_);
  nor (_09420_, _09419_, _09415_);
  or (_09421_, _09420_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_09422_, _09421_, _09418_);
  and (_09423_, _09422_, _09417_);
  or (_07959_, _09423_, _09391_);
  not (_09424_, _09420_);
  nor (_09425_, _09409_, _09404_);
  nor (_09426_, _09425_, _09395_);
  nor (_09427_, _09426_, _09424_);
  nor (_09428_, _09427_, _09389_);
  or (_09429_, _09428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_09430_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_09431_, _09430_, _09420_);
  and (_09432_, _09431_, _06989_);
  and (_07969_, _09432_, _09429_);
  and (_09433_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_09434_, _09433_, _06989_);
  or (_09435_, _09426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_09436_, _09435_, _09424_);
  or (_09437_, _09420_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_09438_, _09437_, _09418_);
  and (_09439_, _09438_, _09436_);
  or (_07973_, _09439_, _09434_);
  and (_09440_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_09441_, _09440_, _06989_);
  or (_09442_, _09426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_09443_, _09442_, _09420_);
  and (_09444_, _09424_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_09445_, _09444_, _09443_);
  and (_09446_, _09445_, _09418_);
  or (_07976_, _09446_, _09441_);
  and (_09447_, _08713_, _08878_);
  and (_09448_, _08932_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_09449_, _09448_, _09447_);
  or (_09450_, _08599_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_09451_, _09450_, _08872_);
  or (_09452_, _09451_, _09301_);
  or (_09453_, _09452_, _09449_);
  nor (_09454_, _08872_, _08599_);
  and (_09455_, _09454_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_09456_, _09455_, _09372_);
  or (_09457_, _09456_, _09453_);
  and (_07980_, _09457_, _06989_);
  and (_09458_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_09459_, _09458_, _06989_);
  or (_09460_, _09426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_09461_, _09460_, _09420_);
  and (_09462_, _09424_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_09463_, _09462_, _09461_);
  and (_09464_, _09463_, _09418_);
  or (_07989_, _09464_, _09459_);
  and (_09465_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_09466_, _09465_, _06989_);
  or (_09467_, _09426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_09468_, _09467_, _09420_);
  and (_09469_, _09424_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_09470_, _09469_, _09468_);
  and (_09471_, _09470_, _09418_);
  or (_07992_, _09471_, _09466_);
  or (_09472_, _09428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_09473_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_09474_, _09473_, _09420_);
  and (_09475_, _09474_, _06989_);
  and (_07997_, _09475_, _09472_);
  and (_09476_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_09477_, _09476_, _06989_);
  and (_09478_, _09424_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_09479_, _09402_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_09480_, _09479_, _09410_);
  not (_09481_, _09415_);
  or (_09482_, _09404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_09483_, _09482_, _09481_);
  and (_09484_, _09483_, _09480_);
  or (_09485_, _09484_, _09478_);
  and (_09486_, _09485_, _09418_);
  or (_08054_, _09486_, _09477_);
  and (_09487_, _07135_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_09488_, _07091_, _06981_);
  not (_09489_, _09488_);
  nor (_09490_, _09489_, _07260_);
  or (_09491_, _09490_, _09487_);
  and (_08073_, _09491_, _06989_);
  and (_09492_, _08932_, _08732_);
  and (_09493_, _09492_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_09494_, _08721_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_09495_, _08633_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_09496_, _09495_, _08925_);
  or (_09497_, _08975_, _08872_);
  and (_09498_, _09497_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_09499_, _09498_, _09496_);
  or (_09500_, _09499_, _09494_);
  or (_09501_, _09500_, _09493_);
  and (_08081_, _09501_, _06989_);
  nor (_08088_, _07319_, rst);
  or (_09502_, _09428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_09503_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_09504_, _09503_, _09420_);
  and (_09505_, _09504_, _06989_);
  and (_08094_, _09505_, _09502_);
  and (_09506_, _09400_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_09507_, _09506_, _09425_);
  or (_09508_, _09507_, _09427_);
  and (_09509_, _09508_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_09510_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nand (_09511_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_09512_, _09511_, _09420_);
  or (_09513_, _09512_, _09510_);
  or (_09514_, _09513_, _09509_);
  and (_08097_, _09514_, _06989_);
  not (_09515_, _09428_);
  and (_09516_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_09517_, _09516_, _09515_);
  and (_09518_, _09400_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nand (_09519_, _09518_, _09425_);
  nand (_09520_, _09519_, _09420_);
  and (_09521_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_09523_, _09521_, _09520_);
  or (_08100_, _09523_, _09517_);
  and (_09524_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  not (_09525_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor (_09527_, _07493_, _09525_);
  or (_09528_, _09527_, _09524_);
  and (_08105_, _09528_, _06989_);
  and (_09529_, _08436_, _06448_);
  and (_09530_, _09529_, _06983_);
  and (_09531_, _09530_, _06977_);
  nand (_09532_, _09531_, _07040_);
  and (_09533_, _07145_, _07075_);
  not (_09534_, _09533_);
  and (_09535_, _06985_, _09074_);
  and (_09536_, _09535_, _06977_);
  nor (_09537_, _09536_, _09534_);
  nor (_09538_, _09537_, _07152_);
  and (_09539_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_09541_, _09539_, _09538_);
  or (_09542_, _09531_, _09541_);
  and (_09543_, _09542_, _06989_);
  and (_08108_, _09543_, _09532_);
  or (_09544_, _08496_, _07327_);
  nor (_09545_, _07325_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_09546_, _09545_, _07362_);
  and (_09547_, _09546_, _09544_);
  and (_08111_, _09547_, _06989_);
  and (_09548_, _07958_, _07920_);
  not (_09549_, _09548_);
  and (_09550_, _09549_, _07960_);
  and (_08135_, _09550_, _06989_);
  nand (_09551_, _09536_, _07040_);
  not (_09552_, _09531_);
  not (_09553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor (_09554_, _09533_, _09553_);
  and (_09555_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_09556_, _09555_, _09554_);
  or (_09557_, _09556_, _09536_);
  and (_09558_, _09557_, _09552_);
  and (_09559_, _09558_, _09551_);
  and (_09560_, _06985_, _08436_);
  and (_09561_, _09560_, _06977_);
  and (_09562_, _09561_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_09563_, _09562_, _09559_);
  and (_08181_, _09563_, _06989_);
  and (_08194_, _07365_, _06989_);
  and (_09564_, _08821_, _08816_);
  or (_09565_, _09564_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_08217_, _09565_, _06989_);
  nor (_09566_, t2_i, rst);
  and (_08250_, _09566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  not (_09567_, _07066_);
  and (_09568_, _07073_, _07071_);
  and (_09569_, _09568_, _07051_);
  nand (_09570_, _09569_, _09567_);
  or (_09571_, _09569_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_09572_, _09571_, _06989_);
  and (_08266_, _09572_, _09570_);
  nand (_09573_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _06989_);
  nor (_08297_, _09573_, t2ex_i);
  and (_08321_, t2ex_i, _06989_);
  not (_09574_, _07077_);
  and (_09575_, _07071_, _07057_);
  or (_09576_, _09575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_09577_, _07071_, _07058_);
  and (_09578_, _09577_, _09576_);
  nor (_09579_, _07145_, _09553_);
  and (_09580_, _07071_, _07066_);
  and (_09581_, _09580_, _09579_);
  or (_09582_, _09581_, _09578_);
  and (_09583_, _09582_, _09574_);
  and (_09584_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_09585_, _09584_, _07046_);
  or (_09586_, _09585_, _09583_);
  nand (_09587_, _07046_, _07040_);
  and (_09588_, _09587_, _09586_);
  or (_09589_, _09588_, _07050_);
  not (_09590_, _07050_);
  or (_09591_, _09590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_09592_, _09591_, _06989_);
  and (_08330_, _09592_, _09589_);
  or (_09593_, _08797_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_08347_, _09593_, _06989_);
  nor (_09594_, _07035_, _06754_);
  not (_09595_, _09594_);
  and (_09597_, _09595_, _08107_);
  and (_09598_, _09597_, _08098_);
  not (_09599_, _09598_);
  and (_09600_, _09599_, _07485_);
  and (_09601_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  or (_09602_, _09601_, _09600_);
  and (_08521_, _09602_, _06989_);
  not (_09603_, _07125_);
  nor (_09604_, _08993_, _09603_);
  nor (_09605_, _08993_, _07122_);
  nor (_09606_, _09604_, _09605_);
  and (_09607_, _09606_, _08997_);
  and (_09608_, _09607_, _09001_);
  or (_09609_, _09608_, _06982_);
  or (_09610_, _09609_, _09604_);
  and (_09611_, _09610_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_09613_, _09009_, _07485_);
  not (_09614_, _09605_);
  nand (_09615_, _09614_, _08997_);
  and (_09616_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_09618_, _09616_, _09615_);
  or (_09619_, _09618_, _09613_);
  or (_09621_, _09619_, _09611_);
  and (_08660_, _09621_, _06989_);
  and (_09623_, _08944_, _08971_);
  not (_09625_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_09626_, _08949_, _08583_);
  nor (_09627_, _09626_, _08947_);
  and (_09629_, _08949_, _08591_);
  and (_09630_, _08949_, _08599_);
  nor (_09631_, _09630_, _09629_);
  and (_09632_, _09631_, _08949_);
  and (_09633_, _09632_, _09627_);
  nor (_09634_, _09633_, _09625_);
  and (_09636_, _08949_, word_in[0]);
  and (_09637_, _09636_, _09633_);
  or (_09638_, _09637_, _09634_);
  or (_09639_, _09638_, _09623_);
  and (_09640_, _08937_, _09056_);
  not (_09641_, _09640_);
  not (_09642_, _09623_);
  or (_09643_, _09642_, word_in[8]);
  and (_09644_, _09643_, _09641_);
  and (_09645_, _09644_, _09639_);
  and (_09646_, _08740_, _08932_);
  and (_09647_, _08935_, _09646_);
  and (_09648_, _08937_, word_in[16]);
  and (_09649_, _09648_, _09056_);
  or (_09650_, _09649_, _09647_);
  or (_09652_, _09650_, _09645_);
  not (_09653_, _09647_);
  or (_09654_, _09653_, word_in[24]);
  and (_14642_, _09654_, _09652_);
  and (_09656_, _08935_, word_in[25]);
  and (_09657_, _09656_, _09647_);
  not (_09658_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_09659_, _09633_, _09658_);
  and (_09660_, _08949_, word_in[1]);
  and (_09661_, _09660_, _09633_);
  or (_09663_, _09661_, _09659_);
  or (_09664_, _09663_, _09623_);
  or (_09665_, _09642_, word_in[9]);
  and (_09666_, _09665_, _09664_);
  or (_09667_, _09666_, _09640_);
  nor (_09668_, _09641_, word_in[17]);
  nor (_09670_, _09668_, _09647_);
  and (_09671_, _09670_, _09667_);
  or (_14643_, _09671_, _09657_);
  not (_09672_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_09673_, _09633_, _09672_);
  and (_09674_, _08949_, word_in[2]);
  and (_09675_, _09674_, _09633_);
  or (_09676_, _09675_, _09673_);
  and (_09678_, _09676_, _09642_);
  and (_09679_, _09623_, word_in[10]);
  or (_09680_, _09679_, _09678_);
  or (_09681_, _09680_, _09640_);
  or (_09682_, _09641_, word_in[18]);
  and (_09683_, _09682_, _09653_);
  and (_09684_, _09683_, _09681_);
  and (_09685_, _08935_, word_in[26]);
  and (_09686_, _09685_, _09647_);
  or (_14644_, _09686_, _09684_);
  not (_09688_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_09689_, _09633_, _09688_);
  and (_09690_, _08949_, word_in[3]);
  and (_09692_, _09690_, _09633_);
  or (_09693_, _09692_, _09689_);
  or (_09694_, _09693_, _09623_);
  or (_09695_, _09642_, word_in[11]);
  and (_09696_, _09695_, _09694_);
  or (_09697_, _09696_, _09640_);
  or (_09698_, _09641_, word_in[19]);
  and (_09699_, _09698_, _09653_);
  and (_09700_, _09699_, _09697_);
  and (_09701_, _08935_, word_in[27]);
  and (_09702_, _09701_, _09647_);
  or (_14645_, _09702_, _09700_);
  and (_09703_, _08935_, word_in[28]);
  and (_09704_, _09703_, _09647_);
  not (_09705_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_09706_, _09633_, _09705_);
  and (_09707_, _08949_, word_in[4]);
  and (_09708_, _09707_, _09633_);
  or (_09709_, _09708_, _09706_);
  and (_09710_, _09709_, _09642_);
  and (_09712_, _09623_, word_in[12]);
  or (_09713_, _09712_, _09710_);
  or (_09714_, _09713_, _09640_);
  nor (_09715_, _09641_, word_in[20]);
  nor (_09716_, _09715_, _09647_);
  and (_09717_, _09716_, _09714_);
  or (_08749_, _09717_, _09704_);
  and (_09718_, _08935_, word_in[29]);
  and (_09719_, _09718_, _09647_);
  not (_09720_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_09721_, _09633_, _09720_);
  and (_09722_, _08949_, word_in[5]);
  and (_09723_, _09722_, _09633_);
  or (_09724_, _09723_, _09721_);
  or (_09725_, _09724_, _09623_);
  or (_09726_, _09642_, word_in[13]);
  and (_09727_, _09726_, _09725_);
  or (_09728_, _09727_, _09640_);
  nor (_09729_, _09641_, word_in[21]);
  nor (_09730_, _09729_, _09647_);
  and (_09731_, _09730_, _09728_);
  or (_14646_, _09731_, _09719_);
  not (_09732_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_09734_, _09633_, _09732_);
  and (_09735_, _08949_, word_in[6]);
  and (_09736_, _09735_, _09633_);
  or (_09737_, _09736_, _09734_);
  or (_09738_, _09737_, _09623_);
  or (_09739_, _09642_, word_in[14]);
  and (_09740_, _09739_, _09738_);
  or (_09741_, _09740_, _09640_);
  nor (_09742_, _09641_, word_in[22]);
  nor (_09743_, _09742_, _09647_);
  and (_09744_, _09743_, _09741_);
  and (_09745_, _08935_, word_in[30]);
  and (_09746_, _09745_, _09647_);
  or (_14647_, _09746_, _09744_);
  nor (_09748_, _09633_, _08777_);
  and (_09749_, _09633_, _08953_);
  or (_09750_, _09749_, _09748_);
  and (_09751_, _09750_, _09642_);
  and (_09752_, _09623_, word_in[15]);
  or (_09753_, _09752_, _09751_);
  or (_09754_, _09753_, _09640_);
  or (_09755_, _09641_, word_in[23]);
  and (_09756_, _09755_, _09653_);
  and (_09757_, _09756_, _09754_);
  and (_09758_, _09647_, word_in[31]);
  or (_14648_, _09758_, _09757_);
  nor (_09759_, _09404_, _09395_);
  or (_09760_, _09759_, _09389_);
  and (_09761_, _09760_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_09762_, _09395_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_09763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_09764_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_09765_, _09764_, _09763_);
  and (_09766_, _09765_, _09762_);
  or (_09767_, _09766_, _09761_);
  and (_08809_, _09767_, _06989_);
  and (_09768_, _08944_, _08731_);
  and (_09769_, _09768_, _08724_);
  not (_09770_, _09769_);
  not (_09771_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_09772_, _08947_, _08584_);
  and (_09773_, _09772_, _09631_);
  nor (_09774_, _09773_, _09771_);
  and (_09775_, _09773_, _09636_);
  or (_09776_, _09775_, _09774_);
  and (_09777_, _09776_, _09770_);
  and (_09778_, _08937_, _08713_);
  and (_09780_, _09778_, _08824_);
  and (_09781_, _09769_, word_in[8]);
  or (_09782_, _09781_, _09780_);
  or (_09783_, _09782_, _09777_);
  and (_09784_, _08935_, _09056_);
  not (_09785_, _09784_);
  not (_09786_, _09780_);
  or (_09787_, _09786_, _09648_);
  and (_09788_, _09787_, _09785_);
  and (_09789_, _09788_, _09783_);
  and (_09790_, _09784_, word_in[24]);
  or (_08840_, _09790_, _09789_);
  not (_09792_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_09793_, _09773_, _09792_);
  and (_09794_, _09773_, _09660_);
  or (_09796_, _09794_, _09793_);
  and (_09797_, _09796_, _09770_);
  and (_09798_, _09769_, word_in[9]);
  or (_09799_, _09798_, _09780_);
  or (_09800_, _09799_, _09797_);
  and (_09801_, _08937_, word_in[17]);
  or (_09802_, _09786_, _09801_);
  and (_09803_, _09802_, _09785_);
  and (_09805_, _09803_, _09800_);
  and (_09806_, _09784_, word_in[25]);
  or (_14666_, _09806_, _09805_);
  not (_09807_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_09808_, _09773_, _09807_);
  and (_09809_, _09773_, _09674_);
  or (_09810_, _09809_, _09808_);
  and (_09811_, _09810_, _09770_);
  and (_09813_, _09769_, word_in[10]);
  or (_09814_, _09813_, _09780_);
  or (_09815_, _09814_, _09811_);
  and (_09816_, _08937_, word_in[18]);
  or (_09817_, _09786_, _09816_);
  and (_09818_, _09817_, _09785_);
  and (_09819_, _09818_, _09815_);
  and (_09820_, _09784_, word_in[26]);
  or (_14667_, _09820_, _09819_);
  not (_09821_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_09822_, _09773_, _09821_);
  and (_09823_, _09773_, _09690_);
  or (_09824_, _09823_, _09822_);
  and (_09825_, _09824_, _09770_);
  and (_09826_, _09769_, word_in[11]);
  or (_09827_, _09826_, _09780_);
  or (_09828_, _09827_, _09825_);
  and (_09829_, _08937_, word_in[19]);
  or (_09830_, _09786_, _09829_);
  and (_09831_, _09830_, _09785_);
  and (_09832_, _09831_, _09828_);
  and (_09833_, _09784_, word_in[27]);
  or (_14668_, _09833_, _09832_);
  not (_09834_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_09835_, _09773_, _09834_);
  and (_09836_, _09773_, _09707_);
  or (_09837_, _09836_, _09835_);
  and (_09838_, _09837_, _09770_);
  and (_09839_, _09769_, word_in[12]);
  or (_09840_, _09839_, _09780_);
  or (_09841_, _09840_, _09838_);
  and (_09842_, _08937_, word_in[20]);
  or (_09843_, _09786_, _09842_);
  and (_09844_, _09843_, _09785_);
  and (_09845_, _09844_, _09841_);
  and (_09846_, _09784_, word_in[28]);
  or (_14669_, _09846_, _09845_);
  not (_09847_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_09848_, _09773_, _09847_);
  and (_09849_, _09773_, _09722_);
  or (_09850_, _09849_, _09848_);
  and (_09851_, _09850_, _09770_);
  and (_09852_, _09769_, word_in[13]);
  or (_09853_, _09852_, _09780_);
  or (_09854_, _09853_, _09851_);
  and (_09855_, _08937_, word_in[21]);
  or (_09856_, _09786_, _09855_);
  and (_09857_, _09856_, _09785_);
  and (_09858_, _09857_, _09854_);
  and (_09859_, _09784_, word_in[29]);
  or (_14670_, _09859_, _09858_);
  not (_09860_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_09861_, _09773_, _09860_);
  and (_09862_, _09773_, _09735_);
  or (_09863_, _09862_, _09861_);
  and (_09865_, _09863_, _09770_);
  and (_09866_, _09769_, word_in[14]);
  or (_09868_, _09866_, _09780_);
  or (_09870_, _09868_, _09865_);
  and (_09871_, _08937_, word_in[22]);
  or (_09872_, _09786_, _09871_);
  and (_09873_, _09872_, _09785_);
  and (_09875_, _09873_, _09870_);
  and (_09876_, _09784_, word_in[30]);
  or (_14671_, _09876_, _09875_);
  nor (_09878_, _09773_, _08698_);
  and (_09879_, _09773_, _08953_);
  or (_09881_, _09879_, _09878_);
  and (_09882_, _09881_, _09770_);
  and (_09883_, _09769_, word_in[15]);
  or (_09884_, _09883_, _09780_);
  or (_09886_, _09884_, _09882_);
  or (_09887_, _09786_, _08942_);
  and (_09888_, _09887_, _09785_);
  and (_09889_, _09888_, _09886_);
  and (_09890_, _09784_, word_in[31]);
  or (_14672_, _09890_, _09889_);
  and (_09891_, _08935_, _08713_);
  and (_09892_, _09891_, _08885_);
  and (_09893_, _08937_, _08731_);
  and (_09894_, _09893_, _08824_);
  not (_09895_, _09894_);
  or (_09896_, _09895_, _09648_);
  and (_09897_, _08944_, _08740_);
  and (_09898_, _09897_, _08724_);
  not (_09899_, _09898_);
  not (_09900_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  not (_09901_, _08947_);
  and (_09902_, _09626_, _09901_);
  and (_09903_, _09902_, _09631_);
  nor (_09904_, _09903_, _09900_);
  and (_09905_, _09903_, _09636_);
  or (_09906_, _09905_, _09904_);
  and (_09907_, _09906_, _09899_);
  and (_09908_, _09898_, word_in[8]);
  or (_09909_, _09908_, _09894_);
  or (_09910_, _09909_, _09907_);
  and (_09911_, _09910_, _09896_);
  or (_09912_, _09911_, _09892_);
  not (_09913_, _09892_);
  or (_09914_, _09913_, word_in[24]);
  and (_14673_, _09914_, _09912_);
  or (_09915_, _09895_, _09801_);
  not (_09916_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_09917_, _09903_, _09916_);
  and (_09918_, _09903_, _09660_);
  or (_09920_, _09918_, _09917_);
  and (_09921_, _09920_, _09899_);
  and (_09923_, _09898_, word_in[9]);
  or (_09924_, _09923_, _09894_);
  or (_09925_, _09924_, _09921_);
  and (_09926_, _09925_, _09915_);
  or (_09927_, _09926_, _09892_);
  or (_09928_, _09913_, word_in[25]);
  and (_14674_, _09928_, _09927_);
  or (_09930_, _09895_, _09816_);
  not (_09931_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_09932_, _09903_, _09931_);
  and (_09933_, _09903_, _09674_);
  or (_09934_, _09933_, _09932_);
  and (_09935_, _09934_, _09899_);
  and (_09937_, _09898_, word_in[10]);
  or (_09938_, _09937_, _09894_);
  or (_09939_, _09938_, _09935_);
  and (_09940_, _09939_, _09930_);
  or (_09941_, _09940_, _09892_);
  or (_09942_, _09913_, word_in[26]);
  and (_14675_, _09942_, _09941_);
  or (_09943_, _09895_, _09829_);
  not (_09944_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_09945_, _09903_, _09944_);
  and (_09946_, _09903_, _09690_);
  or (_09947_, _09946_, _09945_);
  and (_09948_, _09947_, _09899_);
  and (_09949_, _09898_, word_in[11]);
  or (_09950_, _09949_, _09894_);
  or (_09951_, _09950_, _09948_);
  and (_09952_, _09951_, _09943_);
  or (_09953_, _09952_, _09892_);
  or (_09954_, _09913_, word_in[27]);
  and (_14676_, _09954_, _09953_);
  or (_09955_, _09895_, _09842_);
  not (_09957_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_09958_, _09903_, _09957_);
  and (_09959_, _09903_, _09707_);
  or (_09960_, _09959_, _09958_);
  and (_09962_, _09960_, _09899_);
  and (_09964_, _09898_, word_in[12]);
  or (_09965_, _09964_, _09894_);
  or (_09966_, _09965_, _09962_);
  and (_09968_, _09966_, _09955_);
  or (_09969_, _09968_, _09892_);
  or (_09970_, _09913_, word_in[28]);
  and (_14677_, _09970_, _09969_);
  or (_09972_, _09895_, _09855_);
  not (_09974_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_09975_, _09903_, _09974_);
  and (_09977_, _09903_, _09722_);
  or (_09979_, _09977_, _09975_);
  and (_09980_, _09979_, _09899_);
  and (_09981_, _09898_, word_in[13]);
  or (_09982_, _09981_, _09894_);
  or (_09983_, _09982_, _09980_);
  and (_09984_, _09983_, _09972_);
  and (_09985_, _09984_, _09913_);
  and (_09986_, _09892_, word_in[29]);
  or (_08962_, _09986_, _09985_);
  or (_09987_, _09895_, _09871_);
  not (_09988_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_09989_, _09903_, _09988_);
  and (_09990_, _09903_, _09735_);
  or (_09991_, _09990_, _09989_);
  and (_09992_, _09991_, _09899_);
  and (_09993_, _09898_, word_in[14]);
  or (_09994_, _09993_, _09894_);
  or (_09995_, _09994_, _09992_);
  and (_09996_, _09995_, _09987_);
  and (_09997_, _09996_, _09913_);
  and (_09998_, _09892_, word_in[30]);
  or (_14678_, _09998_, _09997_);
  or (_10000_, _09895_, _08942_);
  nor (_10001_, _09903_, _08772_);
  and (_10002_, _09903_, _08953_);
  or (_10003_, _10002_, _10001_);
  and (_10004_, _10003_, _09899_);
  and (_10005_, _09898_, word_in[15]);
  or (_10006_, _10005_, _09894_);
  or (_10007_, _10006_, _10004_);
  and (_10008_, _10007_, _10000_);
  and (_10009_, _10008_, _09913_);
  and (_10010_, _09892_, word_in[31]);
  or (_14679_, _10010_, _10009_);
  and (_10011_, _08935_, _08731_);
  and (_10012_, _10011_, _08885_);
  not (_10013_, _10012_);
  and (_10014_, _08945_, _08724_);
  not (_10015_, _10014_);
  not (_10016_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_10017_, _09631_, _08948_);
  nor (_10018_, _10017_, _10016_);
  and (_10019_, _10017_, _09636_);
  or (_10021_, _10019_, _10018_);
  and (_10022_, _10021_, _10015_);
  and (_10023_, _08937_, _08740_);
  and (_10024_, _10023_, _08824_);
  and (_10026_, _10014_, word_in[8]);
  or (_10027_, _10026_, _10024_);
  or (_10028_, _10027_, _10022_);
  not (_10030_, _10024_);
  or (_10031_, _10030_, _09648_);
  and (_10032_, _10031_, _10028_);
  and (_10034_, _10032_, _10013_);
  and (_10035_, _10012_, word_in[24]);
  or (_14680_, _10035_, _10034_);
  not (_10037_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_10038_, _10017_, _10037_);
  and (_10039_, _10017_, _09660_);
  or (_10040_, _10039_, _10038_);
  and (_10041_, _10040_, _10015_);
  and (_10043_, _10014_, word_in[9]);
  or (_10044_, _10043_, _10024_);
  or (_10046_, _10044_, _10041_);
  or (_10048_, _10030_, _09801_);
  and (_10050_, _10048_, _10046_);
  or (_10052_, _10050_, _10012_);
  or (_10054_, _10013_, word_in[25]);
  and (_14681_, _10054_, _10052_);
  not (_10057_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_10059_, _10017_, _10057_);
  and (_10060_, _10017_, _09674_);
  or (_10061_, _10060_, _10059_);
  and (_10063_, _10061_, _10015_);
  and (_10064_, _10014_, word_in[10]);
  or (_10065_, _10064_, _10024_);
  or (_10066_, _10065_, _10063_);
  or (_10067_, _10030_, _09816_);
  and (_10068_, _10067_, _10066_);
  or (_10069_, _10068_, _10012_);
  or (_10070_, _10013_, word_in[26]);
  and (_14682_, _10070_, _10069_);
  and (_10071_, _10017_, _09690_);
  not (_10072_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_10073_, _10017_, _10072_);
  or (_10075_, _10073_, _10071_);
  and (_10076_, _10075_, _10015_);
  and (_10077_, _10014_, word_in[11]);
  or (_10078_, _10077_, _10024_);
  or (_10080_, _10078_, _10076_);
  or (_10081_, _10030_, _09829_);
  and (_10082_, _10081_, _10080_);
  and (_10083_, _10082_, _10013_);
  and (_10084_, _10012_, word_in[27]);
  or (_14683_, _10084_, _10083_);
  and (_10085_, _10017_, _09707_);
  not (_10086_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_10087_, _10017_, _10086_);
  or (_10088_, _10087_, _10085_);
  and (_10089_, _10088_, _10015_);
  and (_10090_, _10014_, word_in[12]);
  or (_10091_, _10090_, _10024_);
  or (_10093_, _10091_, _10089_);
  or (_10094_, _10030_, _09842_);
  and (_10095_, _10094_, _10093_);
  and (_10096_, _10095_, _10013_);
  and (_10097_, _10012_, word_in[28]);
  or (_14684_, _10097_, _10096_);
  or (_10099_, _10030_, _09855_);
  not (_10100_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_10102_, _10017_, _10100_);
  and (_10103_, _10017_, _09722_);
  or (_10104_, _10103_, _10102_);
  and (_10105_, _10104_, _10015_);
  and (_10106_, _10014_, word_in[13]);
  or (_10107_, _10106_, _10024_);
  or (_10108_, _10107_, _10105_);
  and (_10109_, _10108_, _10099_);
  or (_10110_, _10109_, _10012_);
  or (_10111_, _10013_, word_in[29]);
  and (_14685_, _10111_, _10110_);
  not (_10113_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_10115_, _10017_, _10113_);
  and (_10116_, _10017_, _09735_);
  or (_10117_, _10116_, _10115_);
  and (_10118_, _10117_, _10015_);
  and (_10119_, _10014_, word_in[14]);
  or (_10120_, _10119_, _10024_);
  or (_10121_, _10120_, _10118_);
  or (_10122_, _10030_, _09871_);
  and (_10123_, _10122_, _10121_);
  and (_10124_, _10123_, _10013_);
  and (_10125_, _10012_, word_in[30]);
  or (_14686_, _10125_, _10124_);
  and (_10127_, _10017_, _08953_);
  nor (_10128_, _10017_, _08682_);
  or (_10130_, _10128_, _10127_);
  and (_10132_, _10130_, _10015_);
  and (_10134_, _10014_, word_in[15]);
  or (_10136_, _10134_, _10024_);
  or (_10138_, _10136_, _10132_);
  or (_10140_, _10030_, _08942_);
  and (_10141_, _10140_, _10138_);
  and (_10143_, _10141_, _10013_);
  and (_10145_, _10012_, word_in[31]);
  or (_09047_, _10145_, _10143_);
  and (_10146_, _09604_, _06981_);
  nand (_10147_, _10146_, _07118_);
  or (_10148_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_10149_, _10148_, _06989_);
  and (_09122_, _10149_, _10147_);
  and (_10150_, _08935_, _08874_);
  and (_10151_, _10150_, _08879_);
  and (_10152_, _10151_, _08740_);
  and (_10153_, _08938_, _08860_);
  and (_10154_, _10153_, _08711_);
  not (_10155_, _10154_);
  or (_10156_, _10155_, _09648_);
  and (_10157_, _08944_, _08981_);
  not (_10158_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_10159_, _08949_, _08721_);
  and (_10160_, _10159_, _09627_);
  nor (_10161_, _10160_, _10158_);
  and (_10162_, _10160_, _09636_);
  or (_10163_, _10162_, _10161_);
  or (_10164_, _10163_, _10157_);
  not (_10165_, _10157_);
  or (_10166_, _10165_, word_in[8]);
  and (_10167_, _10166_, _10164_);
  or (_10168_, _10167_, _10154_);
  and (_10169_, _10168_, _10156_);
  or (_10170_, _10169_, _10152_);
  and (_10171_, _08935_, word_in[24]);
  not (_10172_, _10152_);
  or (_10173_, _10172_, _10171_);
  and (_09135_, _10173_, _10170_);
  or (_10174_, _10155_, _09801_);
  not (_10175_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_10176_, _10160_, _10175_);
  and (_10177_, _10160_, _09660_);
  or (_10178_, _10177_, _10176_);
  or (_10179_, _10178_, _10157_);
  or (_10180_, _10165_, word_in[9]);
  and (_10181_, _10180_, _10179_);
  or (_10182_, _10181_, _10154_);
  and (_10183_, _10182_, _10174_);
  or (_10184_, _10183_, _10152_);
  or (_10185_, _10172_, _09656_);
  and (_09137_, _10185_, _10184_);
  or (_10186_, _10155_, _09816_);
  not (_10187_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_10188_, _10160_, _10187_);
  and (_10189_, _10160_, _09674_);
  or (_10190_, _10189_, _10188_);
  or (_10191_, _10190_, _10157_);
  or (_10192_, _10165_, word_in[10]);
  and (_10193_, _10192_, _10191_);
  or (_10194_, _10193_, _10154_);
  and (_10195_, _10194_, _10186_);
  or (_10196_, _10195_, _10152_);
  or (_10197_, _10172_, _09685_);
  and (_09141_, _10197_, _10196_);
  or (_10198_, _10155_, _09829_);
  not (_10199_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_10200_, _10160_, _10199_);
  and (_10201_, _10160_, _09690_);
  or (_10202_, _10201_, _10200_);
  or (_10203_, _10202_, _10157_);
  or (_10204_, _10165_, word_in[11]);
  and (_10205_, _10204_, _10203_);
  or (_10206_, _10205_, _10154_);
  and (_10207_, _10206_, _10198_);
  or (_10208_, _10207_, _10152_);
  or (_10209_, _10172_, _09701_);
  and (_14687_, _10209_, _10208_);
  and (_10210_, _10154_, _09842_);
  and (_10211_, _10160_, word_in[4]);
  not (_10212_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_10213_, _10160_, _10212_);
  or (_10214_, _10213_, _10211_);
  and (_10215_, _10214_, _10165_);
  and (_10216_, _10157_, word_in[12]);
  or (_10217_, _10216_, _10215_);
  and (_10218_, _10217_, _10155_);
  or (_10219_, _10218_, _10210_);
  and (_10220_, _10219_, _10172_);
  and (_10221_, _10152_, _09703_);
  or (_14688_, _10221_, _10220_);
  or (_10222_, _10155_, _09855_);
  not (_10223_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_10224_, _10160_, _10223_);
  and (_10225_, _10160_, _09722_);
  or (_10226_, _10225_, _10224_);
  or (_10227_, _10226_, _10157_);
  or (_10228_, _10165_, word_in[13]);
  and (_10229_, _10228_, _10227_);
  or (_10230_, _10229_, _10154_);
  and (_10231_, _10230_, _10222_);
  or (_10232_, _10231_, _10152_);
  or (_10233_, _10172_, _09718_);
  and (_14689_, _10233_, _10232_);
  and (_10234_, _10160_, word_in[6]);
  not (_10235_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_10236_, _10160_, _10235_);
  or (_10237_, _10236_, _10234_);
  or (_10238_, _10237_, _10157_);
  or (_10239_, _10165_, word_in[14]);
  and (_10240_, _10239_, _10155_);
  and (_10241_, _10240_, _10238_);
  and (_10242_, _10154_, _09871_);
  or (_10243_, _10242_, _10152_);
  or (_10244_, _10243_, _10241_);
  or (_10245_, _10172_, _09745_);
  and (_09152_, _10245_, _10244_);
  and (_10246_, _10154_, _08942_);
  and (_10247_, _10160_, word_in[7]);
  nor (_10248_, _10160_, _08790_);
  or (_10249_, _10248_, _10247_);
  and (_10250_, _10249_, _10165_);
  and (_10251_, _10157_, word_in[15]);
  or (_10252_, _10251_, _10250_);
  and (_10253_, _10252_, _10155_);
  or (_10254_, _10253_, _10246_);
  and (_10255_, _10254_, _10172_);
  and (_10256_, _08935_, word_in[31]);
  and (_10257_, _10152_, _10256_);
  or (_09154_, _10257_, _10255_);
  and (_10258_, _10153_, _08713_);
  not (_10259_, _10258_);
  and (_10260_, _09768_, _08784_);
  and (_10261_, _10159_, _09772_);
  and (_10262_, _10261_, _09636_);
  not (_10263_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_10264_, _10261_, _10263_);
  nor (_10265_, _10264_, _10262_);
  nor (_10266_, _10265_, _10260_);
  and (_10267_, _10260_, word_in[8]);
  or (_10268_, _10267_, _10266_);
  and (_10269_, _10268_, _10259_);
  and (_10270_, _10151_, _08711_);
  and (_10271_, _10258_, _09648_);
  or (_10272_, _10271_, _10270_);
  or (_10273_, _10272_, _10269_);
  not (_10274_, _10270_);
  or (_10275_, _10274_, word_in[24]);
  and (_09235_, _10275_, _10273_);
  not (_10276_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_10277_, _10261_, _10276_);
  and (_10278_, _10261_, _09660_);
  nor (_10279_, _10278_, _10277_);
  nor (_10280_, _10279_, _10260_);
  and (_10281_, _10260_, word_in[9]);
  or (_10282_, _10281_, _10280_);
  and (_10283_, _10282_, _10259_);
  and (_10284_, _10258_, _09801_);
  or (_10285_, _10284_, _10270_);
  or (_10286_, _10285_, _10283_);
  or (_10287_, _10274_, word_in[25]);
  and (_09238_, _10287_, _10286_);
  not (_10288_, _10260_);
  or (_10289_, _10288_, word_in[10]);
  not (_10290_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_10291_, _10261_, _10290_);
  and (_10292_, _10261_, _09674_);
  or (_10293_, _10292_, _10291_);
  or (_10294_, _10293_, _10260_);
  and (_10295_, _10294_, _10259_);
  and (_10296_, _10295_, _10289_);
  and (_10297_, _10258_, _09816_);
  or (_10298_, _10297_, _10270_);
  or (_10299_, _10298_, _10296_);
  or (_10300_, _10274_, word_in[26]);
  and (_14690_, _10300_, _10299_);
  not (_10301_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_10302_, _10261_, _10301_);
  and (_10303_, _10261_, _09690_);
  or (_10304_, _10303_, _10302_);
  or (_10305_, _10304_, _10260_);
  or (_10306_, _10288_, word_in[11]);
  and (_10307_, _10306_, _10305_);
  or (_10308_, _10307_, _10258_);
  or (_10309_, _10259_, _09829_);
  and (_10310_, _10309_, _10308_);
  or (_10311_, _10310_, _10270_);
  or (_10312_, _10274_, word_in[27]);
  and (_09243_, _10312_, _10311_);
  and (_10313_, _10258_, _09842_);
  and (_10314_, _10261_, _09707_);
  not (_10315_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_10316_, _10261_, _10315_);
  nor (_10317_, _10316_, _10314_);
  nor (_10318_, _10317_, _10260_);
  and (_10319_, _10260_, word_in[12]);
  or (_10320_, _10319_, _10318_);
  and (_10321_, _10320_, _10259_);
  or (_10322_, _10321_, _10313_);
  and (_10323_, _10322_, _10274_);
  and (_10324_, _10270_, word_in[28]);
  or (_09247_, _10324_, _10323_);
  not (_10325_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_10326_, _10261_, _10325_);
  and (_10327_, _10261_, _09722_);
  or (_10328_, _10327_, _10326_);
  or (_10329_, _10328_, _10260_);
  or (_10330_, _10288_, word_in[13]);
  and (_10331_, _10330_, _10329_);
  or (_10332_, _10331_, _10258_);
  or (_10333_, _10259_, _09855_);
  and (_10334_, _10333_, _10332_);
  or (_10335_, _10334_, _10270_);
  or (_10336_, _10274_, word_in[29]);
  and (_09251_, _10336_, _10335_);
  or (_10337_, _10288_, word_in[14]);
  not (_10338_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_10339_, _10261_, _10338_);
  and (_10340_, _10261_, _09735_);
  or (_10341_, _10340_, _10339_);
  or (_10342_, _10341_, _10260_);
  and (_10343_, _10342_, _10259_);
  and (_10344_, _10343_, _10337_);
  and (_10345_, _10258_, _09871_);
  or (_10346_, _10345_, _10270_);
  or (_10347_, _10346_, _10344_);
  or (_10348_, _10274_, word_in[30]);
  and (_09254_, _10348_, _10347_);
  nor (_10349_, _10261_, _08693_);
  and (_10350_, _10261_, _08953_);
  or (_10351_, _10350_, _10349_);
  or (_10352_, _10351_, _10260_);
  or (_10353_, _10288_, word_in[15]);
  and (_10354_, _10353_, _10352_);
  or (_10355_, _10354_, _10258_);
  or (_10356_, _10259_, _08942_);
  and (_10357_, _10356_, _10355_);
  or (_10358_, _10357_, _10270_);
  or (_10359_, _10274_, word_in[31]);
  and (_09257_, _10359_, _10358_);
  nand (_10360_, _10146_, _07317_);
  or (_10361_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_10362_, _10361_, _06989_);
  and (_09305_, _10362_, _10360_);
  and (_10363_, _10151_, _08713_);
  and (_10364_, _10153_, _08731_);
  not (_10365_, _10364_);
  or (_10366_, _10365_, _09648_);
  and (_10367_, _09897_, _08784_);
  not (_10368_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_10369_, _09902_, _08721_);
  nor (_10370_, _10369_, _10368_);
  and (_10371_, _10369_, _09636_);
  or (_10372_, _10371_, _10370_);
  or (_10373_, _10372_, _10367_);
  not (_10374_, _10367_);
  or (_10375_, _10374_, word_in[8]);
  and (_10376_, _10375_, _10373_);
  or (_10377_, _10376_, _10364_);
  and (_10378_, _10377_, _10366_);
  or (_10379_, _10378_, _10363_);
  not (_10380_, _10363_);
  or (_10381_, _10380_, word_in[24]);
  and (_09328_, _10381_, _10379_);
  not (_10382_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_10383_, _10369_, _10382_);
  and (_10384_, _10369_, _09660_);
  or (_10385_, _10384_, _10383_);
  and (_10386_, _10385_, _10374_);
  and (_10387_, _10367_, word_in[9]);
  or (_10388_, _10387_, _10364_);
  or (_10389_, _10388_, _10386_);
  or (_10390_, _10365_, _09801_);
  and (_10391_, _10390_, _10389_);
  or (_10392_, _10391_, _10363_);
  or (_10393_, _10380_, word_in[25]);
  and (_14691_, _10393_, _10392_);
  or (_10394_, _10365_, _09816_);
  not (_10395_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_10396_, _10369_, _10395_);
  and (_10397_, _10369_, _09674_);
  or (_10398_, _10397_, _10396_);
  and (_10399_, _10398_, _10374_);
  and (_10401_, _10367_, word_in[10]);
  or (_10402_, _10401_, _10364_);
  or (_10403_, _10402_, _10399_);
  and (_10404_, _10403_, _10394_);
  or (_10405_, _10404_, _10363_);
  or (_10406_, _10380_, word_in[26]);
  and (_09335_, _10406_, _10405_);
  not (_10407_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_10408_, _10369_, _10407_);
  and (_10409_, _10369_, _09690_);
  or (_10410_, _10409_, _10408_);
  or (_10411_, _10410_, _10367_);
  or (_10412_, _10374_, word_in[11]);
  and (_10413_, _10412_, _10411_);
  or (_10414_, _10413_, _10364_);
  or (_10415_, _10365_, _09829_);
  and (_10416_, _10415_, _10414_);
  and (_10417_, _10416_, _10380_);
  and (_10418_, _10363_, word_in[27]);
  or (_14692_, _10418_, _10417_);
  or (_10419_, _10365_, _09842_);
  not (_10420_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_10421_, _10369_, _10420_);
  and (_10422_, _10369_, _09707_);
  or (_10423_, _10422_, _10421_);
  and (_10424_, _10423_, _10374_);
  and (_10425_, _10367_, word_in[12]);
  or (_10426_, _10425_, _10364_);
  or (_10427_, _10426_, _10424_);
  and (_10428_, _10427_, _10419_);
  or (_10429_, _10428_, _10363_);
  or (_10430_, _10380_, word_in[28]);
  and (_14693_, _10430_, _10429_);
  not (_10431_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_10432_, _10369_, _10431_);
  and (_10433_, _10369_, _09722_);
  or (_10434_, _10433_, _10432_);
  or (_10435_, _10434_, _10367_);
  or (_10436_, _10374_, word_in[13]);
  and (_10437_, _10436_, _10435_);
  or (_10438_, _10437_, _10364_);
  or (_10439_, _10365_, _09855_);
  and (_10440_, _10439_, _10438_);
  and (_10441_, _10440_, _10380_);
  and (_10442_, _10363_, word_in[29]);
  or (_09346_, _10442_, _10441_);
  or (_10443_, _10365_, _09871_);
  not (_10444_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_10445_, _10369_, _10444_);
  and (_10447_, _10369_, _09735_);
  or (_10448_, _10447_, _10445_);
  and (_10450_, _10448_, _10374_);
  and (_10451_, _10367_, word_in[14]);
  or (_10453_, _10451_, _10364_);
  or (_10454_, _10453_, _10450_);
  and (_10455_, _10454_, _10443_);
  or (_10456_, _10455_, _10363_);
  or (_10457_, _10380_, word_in[30]);
  and (_09351_, _10457_, _10456_);
  or (_10458_, _10365_, _08942_);
  nor (_10459_, _10369_, _08785_);
  and (_10460_, _10369_, _08953_);
  or (_10461_, _10460_, _10459_);
  and (_10462_, _10461_, _10374_);
  and (_10463_, _10367_, word_in[15]);
  or (_10464_, _10463_, _10364_);
  or (_10465_, _10464_, _10462_);
  and (_10466_, _10465_, _10458_);
  or (_10467_, _10466_, _10363_);
  or (_10468_, _10380_, word_in[31]);
  and (_09354_, _10468_, _10467_);
  and (_10469_, _08935_, _09016_);
  and (_10470_, _10153_, _08740_);
  not (_10471_, _10470_);
  or (_10472_, _10471_, _09648_);
  and (_10473_, _08945_, _08784_);
  not (_10474_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_10475_, _10159_, _08948_);
  nor (_10476_, _10475_, _10474_);
  and (_10477_, _10475_, _09636_);
  or (_10478_, _10477_, _10476_);
  or (_10479_, _10478_, _10473_);
  not (_10480_, _10473_);
  or (_10481_, _10480_, word_in[8]);
  and (_10482_, _10481_, _10479_);
  or (_10483_, _10482_, _10470_);
  and (_10484_, _10483_, _10472_);
  or (_10485_, _10484_, _10469_);
  not (_10486_, _10469_);
  or (_10487_, _10486_, word_in[24]);
  and (_14694_, _10487_, _10485_);
  or (_10488_, _10480_, word_in[9]);
  not (_10489_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_10490_, _10475_, _10489_);
  and (_10491_, _10475_, _09660_);
  or (_10492_, _10491_, _10490_);
  or (_10493_, _10492_, _10473_);
  and (_10494_, _10493_, _10471_);
  and (_10495_, _10494_, _10488_);
  and (_10496_, _10470_, _09801_);
  or (_10497_, _10496_, _10469_);
  or (_10498_, _10497_, _10495_);
  or (_10499_, _10486_, word_in[25]);
  and (_14695_, _10499_, _10498_);
  or (_10500_, _10471_, _09816_);
  not (_10501_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_10502_, _10475_, _10501_);
  and (_10503_, _10475_, _09674_);
  or (_10504_, _10503_, _10502_);
  or (_10505_, _10504_, _10473_);
  or (_10506_, _10480_, word_in[10]);
  and (_10507_, _10506_, _10505_);
  or (_10508_, _10507_, _10470_);
  and (_10509_, _10508_, _10500_);
  and (_10510_, _10509_, _10486_);
  and (_10511_, _10469_, word_in[26]);
  or (_14696_, _10511_, _10510_);
  not (_10512_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_10513_, _10475_, _10512_);
  and (_10514_, _10475_, _09690_);
  nor (_10515_, _10514_, _10513_);
  nor (_10516_, _10515_, _10473_);
  and (_10517_, _10473_, word_in[11]);
  or (_10518_, _10517_, _10516_);
  and (_10519_, _10518_, _10471_);
  and (_10520_, _10470_, _09829_);
  or (_10521_, _10520_, _10469_);
  or (_10522_, _10521_, _10519_);
  or (_10523_, _10486_, word_in[27]);
  and (_14697_, _10523_, _10522_);
  or (_10524_, _10480_, word_in[12]);
  not (_10525_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_10526_, _10475_, _10525_);
  and (_10527_, _10475_, _09707_);
  or (_10528_, _10527_, _10526_);
  or (_10529_, _10528_, _10473_);
  and (_10530_, _10529_, _10471_);
  and (_10531_, _10530_, _10524_);
  and (_10532_, _10470_, _09842_);
  or (_10533_, _10532_, _10469_);
  or (_10534_, _10533_, _10531_);
  or (_10535_, _10486_, word_in[28]);
  and (_14698_, _10535_, _10534_);
  or (_10536_, _10471_, _09855_);
  not (_10537_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_10538_, _10475_, _10537_);
  and (_10539_, _10475_, _09722_);
  or (_10540_, _10539_, _10538_);
  or (_10541_, _10540_, _10473_);
  or (_10542_, _10480_, word_in[13]);
  and (_10543_, _10542_, _10541_);
  or (_10544_, _10543_, _10470_);
  and (_10545_, _10544_, _10536_);
  or (_10546_, _10545_, _10469_);
  or (_10547_, _10486_, word_in[29]);
  and (_14699_, _10547_, _10546_);
  not (_10548_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_10549_, _10475_, _10548_);
  and (_10550_, _10475_, _09735_);
  nor (_10551_, _10550_, _10549_);
  nor (_10552_, _10551_, _10473_);
  and (_10553_, _10473_, word_in[14]);
  or (_10554_, _10553_, _10552_);
  and (_10555_, _10554_, _10471_);
  and (_10556_, _10470_, _09871_);
  or (_10557_, _10556_, _10469_);
  or (_10558_, _10557_, _10555_);
  or (_10559_, _10486_, word_in[30]);
  and (_14700_, _10559_, _10558_);
  or (_10560_, _10471_, _08942_);
  nor (_10561_, _10475_, _08687_);
  and (_10562_, _10475_, _08953_);
  or (_10563_, _10562_, _10561_);
  or (_10564_, _10563_, _10473_);
  or (_10565_, _10480_, word_in[15]);
  and (_10566_, _10565_, _10564_);
  or (_10567_, _10566_, _10470_);
  and (_10568_, _10567_, _10560_);
  or (_10569_, _10568_, _10469_);
  or (_10570_, _10486_, word_in[31]);
  and (_14701_, _10570_, _10569_);
  and (_10571_, _08937_, _09058_);
  and (_10572_, _08944_, _08722_);
  not (_10573_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_10574_, _09630_, _08720_);
  and (_10575_, _10574_, _09627_);
  nor (_10576_, _10575_, _10573_);
  and (_10577_, _10575_, _09636_);
  or (_10578_, _10577_, _10576_);
  or (_10579_, _10578_, _10572_);
  not (_10580_, _10572_);
  or (_10581_, _10580_, word_in[8]);
  and (_10582_, _10581_, _10579_);
  or (_10583_, _10582_, _10571_);
  and (_10584_, _08935_, _08890_);
  not (_10585_, _10584_);
  not (_10586_, _10571_);
  or (_10587_, _10586_, word_in[16]);
  and (_10588_, _10587_, _10585_);
  and (_10589_, _10588_, _10583_);
  and (_10590_, _10584_, word_in[24]);
  or (_09522_, _10590_, _10589_);
  not (_10591_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_10592_, _10575_, _10591_);
  and (_10593_, _10575_, _09660_);
  or (_10594_, _10593_, _10592_);
  or (_10595_, _10594_, _10572_);
  or (_10596_, _10580_, word_in[9]);
  and (_10597_, _10596_, _10595_);
  or (_10598_, _10597_, _10571_);
  or (_10599_, _10586_, word_in[17]);
  and (_10600_, _10599_, _10585_);
  and (_10601_, _10600_, _10598_);
  and (_10602_, _10584_, word_in[25]);
  or (_14702_, _10602_, _10601_);
  not (_10603_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_10604_, _10575_, _10603_);
  and (_10605_, _10575_, _09674_);
  or (_10606_, _10605_, _10604_);
  or (_10607_, _10606_, _10572_);
  or (_10608_, _10580_, word_in[10]);
  and (_10609_, _10608_, _10607_);
  or (_10610_, _10609_, _10571_);
  or (_10611_, _10586_, word_in[18]);
  and (_10612_, _10611_, _10585_);
  and (_10613_, _10612_, _10610_);
  and (_10614_, _10584_, word_in[26]);
  or (_09526_, _10614_, _10613_);
  not (_10615_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_10616_, _10575_, _10615_);
  and (_10617_, _10575_, _09690_);
  or (_10618_, _10617_, _10616_);
  or (_10619_, _10618_, _10572_);
  or (_10620_, _10580_, word_in[11]);
  and (_10621_, _10620_, _10619_);
  or (_10622_, _10621_, _10571_);
  or (_10623_, _10586_, word_in[19]);
  and (_10624_, _10623_, _10585_);
  and (_10625_, _10624_, _10622_);
  and (_10626_, _10584_, word_in[27]);
  or (_14703_, _10626_, _10625_);
  not (_10627_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_10628_, _10575_, _10627_);
  and (_10629_, _10575_, _09707_);
  or (_10630_, _10629_, _10628_);
  or (_10631_, _10630_, _10572_);
  or (_10632_, _10580_, word_in[12]);
  and (_10633_, _10632_, _10631_);
  or (_10634_, _10633_, _10571_);
  or (_10635_, _10586_, word_in[20]);
  and (_10636_, _10635_, _10585_);
  and (_10637_, _10636_, _10634_);
  and (_10638_, _10584_, word_in[28]);
  or (_14704_, _10638_, _10637_);
  not (_10639_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_10640_, _10575_, _10639_);
  and (_10641_, _10575_, _09722_);
  or (_10642_, _10641_, _10640_);
  or (_10643_, _10642_, _10572_);
  or (_10644_, _10580_, word_in[13]);
  and (_10645_, _10644_, _10643_);
  or (_10646_, _10645_, _10571_);
  or (_10647_, _10586_, word_in[21]);
  and (_10648_, _10647_, _10585_);
  and (_10649_, _10648_, _10646_);
  and (_10650_, _10584_, word_in[29]);
  or (_14705_, _10650_, _10649_);
  and (_10651_, _10584_, word_in[30]);
  not (_10652_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_10653_, _10575_, _10652_);
  and (_10654_, _10575_, _09735_);
  or (_10655_, _10654_, _10653_);
  and (_10656_, _10655_, _10580_);
  and (_10657_, _10572_, word_in[14]);
  or (_10658_, _10657_, _10656_);
  or (_10659_, _10658_, _10571_);
  nor (_10660_, _10586_, word_in[22]);
  nor (_10661_, _10660_, _10584_);
  and (_10662_, _10661_, _10659_);
  or (_09540_, _10662_, _10651_);
  nor (_10663_, _10575_, _08765_);
  and (_10664_, _10575_, _08953_);
  or (_10665_, _10664_, _10663_);
  or (_10666_, _10665_, _10572_);
  or (_10667_, _10580_, word_in[15]);
  and (_10668_, _10667_, _10666_);
  or (_10669_, _10668_, _10571_);
  or (_10670_, _10586_, word_in[23]);
  and (_10671_, _10670_, _10585_);
  and (_10672_, _10671_, _10669_);
  and (_10673_, _10584_, word_in[31]);
  or (_14706_, _10673_, _10672_);
  and (_10674_, _07262_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor (_10675_, _07317_, _07262_);
  or (_10676_, _10675_, _10674_);
  and (_09596_, _10676_, _06989_);
  and (_10677_, _08935_, _08711_);
  and (_10678_, _10677_, _08880_);
  and (_10679_, _09778_, _08822_);
  not (_10681_, _10679_);
  or (_10682_, _10681_, _09648_);
  and (_10683_, _09768_, _08726_);
  not (_10684_, _10683_);
  not (_10685_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_10686_, _10574_, _09772_);
  nor (_10687_, _10686_, _10685_);
  and (_10688_, _10686_, _09636_);
  or (_10689_, _10688_, _10687_);
  and (_10690_, _10689_, _10684_);
  and (_10691_, _10683_, word_in[8]);
  or (_10692_, _10691_, _10679_);
  or (_10693_, _10692_, _10690_);
  and (_10694_, _10693_, _10682_);
  or (_10695_, _10694_, _10678_);
  not (_10696_, _10678_);
  or (_10697_, _10696_, word_in[24]);
  and (_14707_, _10697_, _10695_);
  or (_10698_, _10681_, _09801_);
  not (_10699_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_10700_, _10686_, _10699_);
  and (_10701_, _10686_, _09660_);
  or (_10702_, _10701_, _10700_);
  and (_10703_, _10702_, _10684_);
  and (_10704_, _10683_, word_in[9]);
  or (_10705_, _10704_, _10679_);
  or (_10706_, _10705_, _10703_);
  and (_10707_, _10706_, _10698_);
  or (_10708_, _10707_, _10678_);
  or (_10709_, _10696_, word_in[25]);
  and (_09612_, _10709_, _10708_);
  not (_10710_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_10711_, _10686_, _10710_);
  and (_10712_, _10686_, _09674_);
  or (_10713_, _10712_, _10711_);
  and (_10714_, _10713_, _10684_);
  and (_10715_, _10683_, word_in[10]);
  or (_10716_, _10715_, _10679_);
  or (_10717_, _10716_, _10714_);
  or (_10718_, _10681_, _09816_);
  and (_10719_, _10718_, _10717_);
  or (_10720_, _10719_, _10678_);
  or (_10721_, _10696_, word_in[26]);
  and (_09617_, _10721_, _10720_);
  and (_10722_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  not (_10723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor (_10724_, _07493_, _10723_);
  or (_10725_, _10724_, _10722_);
  and (_09620_, _10725_, _06989_);
  or (_10726_, _10681_, _09829_);
  not (_10727_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_10728_, _10686_, _10727_);
  and (_10729_, _10686_, _09690_);
  or (_10730_, _10729_, _10728_);
  and (_10731_, _10730_, _10684_);
  and (_10732_, _10683_, word_in[11]);
  or (_10733_, _10732_, _10679_);
  or (_10734_, _10733_, _10731_);
  and (_10735_, _10734_, _10726_);
  or (_10736_, _10735_, _10678_);
  or (_10737_, _10696_, word_in[27]);
  and (_09622_, _10737_, _10736_);
  and (_10738_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  not (_10739_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor (_10740_, _07493_, _10739_);
  or (_10741_, _10740_, _10738_);
  and (_09624_, _10741_, _06989_);
  or (_10742_, _10681_, _09842_);
  not (_10743_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_10744_, _10686_, _10743_);
  and (_10745_, _10686_, _09707_);
  or (_10746_, _10745_, _10744_);
  and (_10747_, _10746_, _10684_);
  and (_10748_, _10683_, word_in[12]);
  or (_10749_, _10748_, _10679_);
  or (_10750_, _10749_, _10747_);
  and (_10751_, _10750_, _10742_);
  or (_10752_, _10751_, _10678_);
  or (_10753_, _10696_, word_in[28]);
  and (_14708_, _10753_, _10752_);
  and (_10754_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not (_10755_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_10756_, _07493_, _10755_);
  or (_10757_, _10756_, _10754_);
  and (_09628_, _10757_, _06989_);
  or (_10758_, _10681_, _09855_);
  not (_10759_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_10760_, _10686_, _10759_);
  and (_10761_, _10686_, _09722_);
  or (_10762_, _10761_, _10760_);
  and (_10763_, _10762_, _10684_);
  and (_10764_, _10683_, word_in[13]);
  or (_10765_, _10764_, _10679_);
  or (_10766_, _10765_, _10763_);
  and (_10767_, _10766_, _10758_);
  or (_10768_, _10767_, _10678_);
  or (_10769_, _10696_, word_in[29]);
  and (_14709_, _10769_, _10768_);
  or (_10770_, _10681_, _09871_);
  not (_10771_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_10772_, _10686_, _10771_);
  and (_10773_, _10686_, _09735_);
  or (_10774_, _10773_, _10772_);
  and (_10775_, _10774_, _10684_);
  and (_10776_, _10683_, word_in[14]);
  or (_10777_, _10776_, _10679_);
  or (_10778_, _10777_, _10775_);
  and (_10779_, _10778_, _10770_);
  or (_10780_, _10779_, _10678_);
  or (_10781_, _10696_, word_in[30]);
  and (_14710_, _10781_, _10780_);
  or (_10782_, _10681_, _08942_);
  nor (_10783_, _10686_, _08674_);
  and (_10784_, _10686_, _08953_);
  or (_10785_, _10784_, _10783_);
  and (_10786_, _10785_, _10684_);
  and (_10787_, _10683_, word_in[15]);
  or (_10788_, _10787_, _10679_);
  or (_10789_, _10788_, _10786_);
  and (_10790_, _10789_, _10782_);
  or (_10791_, _10790_, _10678_);
  or (_10792_, _10696_, word_in[31]);
  and (_09635_, _10792_, _10791_);
  nor (_10793_, _07325_, _06794_);
  and (_10794_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_10795_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_10796_, _10795_, _10794_);
  and (_10797_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_10798_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_10799_, _10798_, _10797_);
  and (_10800_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_10801_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_10802_, _10801_, _10800_);
  and (_10803_, _10802_, _10799_);
  and (_10804_, _10803_, _10796_);
  nor (_10805_, _10804_, _08477_);
  nor (_10806_, _10805_, _10793_);
  nor (_09651_, _10806_, rst);
  not (_10807_, _07360_);
  not (_10808_, _08496_);
  not (_10809_, _08529_);
  and (_10810_, _10809_, _08512_);
  and (_10811_, _10810_, _10808_);
  and (_10812_, _10811_, _10807_);
  nor (_10813_, _08576_, _08463_);
  nor (_10814_, _08561_, _08545_);
  and (_10815_, _10814_, _10813_);
  and (_10816_, _10815_, _10812_);
  and (_10817_, _08561_, _08545_);
  and (_10818_, _10817_, _10813_);
  not (_10819_, _08512_);
  and (_10820_, _10819_, _08496_);
  and (_10821_, _10820_, _10809_);
  and (_10822_, _10821_, _10818_);
  nor (_10823_, _10822_, _10816_);
  and (_10824_, _08576_, _08463_);
  and (_10825_, _10824_, _10817_);
  and (_10826_, _10825_, _10812_);
  and (_10827_, _10813_, _08561_);
  and (_10828_, _10827_, _10812_);
  nor (_10829_, _10828_, _10826_);
  and (_10830_, _10829_, _10823_);
  and (_10831_, _10811_, _07360_);
  nor (_10832_, _08512_, _08496_);
  and (_10833_, _10832_, _10809_);
  and (_10834_, _10833_, _10807_);
  not (_10835_, _08576_);
  nor (_10836_, _10835_, _08463_);
  and (_10837_, _10836_, _08561_);
  and (_10838_, _10837_, _10834_);
  nor (_10839_, _10838_, _10831_);
  not (_10840_, _08545_);
  and (_10841_, _10824_, _10840_);
  and (_10842_, _10841_, _10821_);
  and (_10843_, _10821_, _08545_);
  and (_10844_, _10824_, _08561_);
  and (_10845_, _10844_, _10843_);
  nor (_10846_, _10845_, _10842_);
  and (_10847_, _10846_, _10839_);
  and (_10848_, _10847_, _10830_);
  and (_10849_, _10833_, _07360_);
  and (_10850_, _10835_, _08463_);
  and (_10851_, _10850_, _08561_);
  and (_10852_, _10851_, _10849_);
  not (_10853_, _10852_);
  not (_10854_, _08561_);
  and (_10855_, _10854_, _08463_);
  and (_10856_, _10855_, _10835_);
  and (_10857_, _10856_, _10812_);
  not (_10858_, _10857_);
  and (_10859_, _10824_, _10814_);
  and (_10860_, _10859_, _10812_);
  and (_10861_, _10825_, _08529_);
  nor (_10862_, _10861_, _10860_);
  and (_10863_, _10862_, _10858_);
  and (_10864_, _10863_, _10853_);
  and (_10865_, _10864_, _10848_);
  nor (_10866_, _10854_, _08545_);
  and (_10867_, _10866_, _10824_);
  not (_10868_, _10867_);
  and (_10869_, _08512_, _08496_);
  and (_10870_, _10869_, _10809_);
  and (_10871_, _10870_, _10807_);
  nor (_10872_, _10871_, _10812_);
  nor (_10873_, _10872_, _10868_);
  not (_10874_, _10873_);
  and (_10875_, _10854_, _08545_);
  and (_10876_, _10875_, _10850_);
  and (_10878_, _10876_, _08529_);
  and (_10879_, _10875_, _10813_);
  not (_10880_, _10879_);
  nor (_10881_, _10871_, _10833_);
  nor (_10882_, _10881_, _10880_);
  nor (_10883_, _10882_, _10878_);
  and (_10884_, _10883_, _10874_);
  not (_10885_, _10815_);
  nor (_10886_, _10881_, _10885_);
  and (_10887_, _10849_, _10836_);
  nor (_10888_, _10887_, _10886_);
  and (_10889_, _10866_, _10813_);
  nor (_10890_, _10869_, _10832_);
  nor (_10891_, _10890_, _08529_);
  and (_10892_, _10891_, _10889_);
  not (_10893_, _10859_);
  nor (_10894_, _10871_, _08529_);
  nor (_10895_, _10894_, _10893_);
  nor (_10896_, _10895_, _10892_);
  and (_10897_, _10896_, _10888_);
  and (_10898_, _10897_, _10884_);
  and (_10899_, _10898_, _10865_);
  nor (_10900_, _10859_, _10818_);
  not (_10901_, _10900_);
  and (_10902_, _10901_, _10849_);
  and (_10903_, _10836_, _10854_);
  and (_10904_, _10903_, _10871_);
  nor (_10905_, _10904_, _10902_);
  and (_10906_, _10876_, _10849_);
  not (_10907_, _10817_);
  not (_10908_, _10814_);
  and (_10909_, _10836_, _10908_);
  and (_10910_, _10909_, _10907_);
  and (_10911_, _10910_, _10812_);
  and (_10912_, _10833_, _10825_);
  and (_10913_, _10912_, _10807_);
  or (_10914_, _10913_, _10911_);
  nor (_10915_, _10914_, _10906_);
  and (_10916_, _10915_, _10905_);
  and (_10917_, _10870_, _07360_);
  and (_10918_, _10917_, _10815_);
  and (_10919_, _10875_, _10824_);
  and (_10920_, _10919_, _10812_);
  nor (_10921_, _10920_, _10918_);
  nor (_10922_, _10867_, _10818_);
  nor (_10923_, _10922_, _10809_);
  not (_10924_, _10871_);
  not (_10925_, _10876_);
  nor (_10926_, _10825_, _10818_);
  and (_10927_, _10926_, _10925_);
  nor (_10928_, _10927_, _10924_);
  nor (_10929_, _10928_, _10923_);
  and (_10930_, _10929_, _10921_);
  and (_10931_, _10849_, _10825_);
  and (_10932_, _10917_, _10879_);
  or (_10933_, _10932_, _10931_);
  and (_10934_, _10850_, _10814_);
  nor (_10935_, _10934_, _10919_);
  nor (_10936_, _10871_, _10849_);
  nor (_10937_, _10936_, _10935_);
  nor (_10938_, _10937_, _10933_);
  and (_10939_, _10836_, _10817_);
  or (_10940_, _10939_, _10879_);
  nand (_10941_, _10940_, _10812_);
  not (_10942_, _10834_);
  nor (_10943_, _10919_, _10818_);
  nor (_10944_, _10943_, _10942_);
  not (_10945_, _10944_);
  and (_10946_, _10945_, _10941_);
  and (_10947_, _10946_, _10938_);
  and (_10948_, _10947_, _10930_);
  and (_10949_, _10948_, _10916_);
  and (_10950_, _10949_, _10899_);
  nor (_10951_, _10861_, _10845_);
  and (_10952_, _10917_, _10889_);
  and (_10953_, _10939_, _10812_);
  nor (_10954_, _10953_, _10952_);
  and (_10955_, _10954_, _10951_);
  not (_10956_, _10933_);
  and (_10957_, _10956_, _10921_);
  and (_10958_, _10957_, _10955_);
  and (_10959_, _10958_, _10916_);
  not (_10960_, _10959_);
  nor (_10961_, _10960_, _10950_);
  nor (_10962_, _10961_, _07490_);
  nand (_10963_, _10962_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_10964_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  or (_10965_, _10962_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_10966_, _10965_, _10964_);
  and (_09655_, _10966_, _10963_);
  nor (_10967_, _07035_, _06810_);
  not (_10968_, _10967_);
  and (_10969_, _10968_, _09133_);
  and (_10970_, _10969_, _09115_);
  nor (_10971_, _10970_, _07262_);
  nor (_10972_, _08994_, _06982_);
  nand (_10973_, _10972_, _07127_);
  or (_10974_, _10973_, _07131_);
  and (_10975_, _10974_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_10976_, _10975_, _10971_);
  and (_09662_, _10976_, _06989_);
  and (_10977_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _06989_);
  and (_10978_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_10979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_10980_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_10981_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_10982_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_10983_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_10984_, _10983_, _10981_);
  and (_10985_, _10984_, _10982_);
  nor (_10986_, _10985_, _10981_);
  nor (_10987_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_10988_, _10987_, _10980_);
  not (_10990_, _10988_);
  nor (_10991_, _10990_, _10986_);
  nor (_10992_, _10991_, _10980_);
  not (_10993_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_10994_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not (_10995_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_10996_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_10997_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_10998_, _10997_, _10996_);
  and (_10999_, _10998_, _10995_);
  and (_11000_, _10999_, _10994_);
  and (_11001_, _11000_, _10993_);
  and (_11002_, _11001_, _10992_);
  nor (_11003_, _11002_, _10979_);
  and (_11004_, _11002_, _10979_);
  nor (_11006_, _11004_, _11003_);
  not (_11007_, _11006_);
  and (_11008_, _10999_, _10992_);
  and (_11009_, _11008_, _10994_);
  nor (_11010_, _11009_, _10993_);
  nor (_11011_, _11010_, _11002_);
  nor (_11012_, _11008_, _10994_);
  nor (_11013_, _11012_, _11009_);
  not (_11014_, _11013_);
  and (_11015_, _10998_, _10992_);
  nor (_11016_, _11015_, _10995_);
  nor (_11017_, _11016_, _11008_);
  not (_11018_, _11017_);
  and (_11019_, _10992_, _10997_);
  nor (_11020_, _11019_, _10996_);
  nor (_11021_, _11020_, _11015_);
  not (_11022_, _11021_);
  nor (_11023_, _10992_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_11024_, _10992_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_11025_, _11024_, _11023_);
  not (_11026_, _11025_);
  nor (_11027_, _10984_, _10982_);
  nor (_11028_, _11027_, _10985_);
  not (_11029_, _11028_);
  nor (_11030_, _11029_, _10950_);
  not (_11032_, _10961_);
  nor (_11033_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_11034_, _11033_, _10982_);
  and (_11035_, _11034_, _11032_);
  and (_11036_, _11029_, _10950_);
  nor (_11037_, _11036_, _11030_);
  and (_11038_, _11037_, _11035_);
  nor (_11039_, _11038_, _11030_);
  not (_11040_, _11039_);
  and (_11041_, _10990_, _10986_);
  nor (_11042_, _11041_, _10991_);
  and (_11043_, _11042_, _11040_);
  and (_11044_, _11043_, _11026_);
  and (_11045_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_11046_, _11045_, _10997_);
  nand (_11047_, _11046_, _11023_);
  or (_11048_, _11046_, _11023_);
  and (_11049_, _11048_, _11047_);
  and (_11050_, _11049_, _11044_);
  and (_11051_, _11050_, _11022_);
  and (_11052_, _11051_, _11018_);
  nand (_11053_, _11052_, _11014_);
  nor (_11054_, _11053_, _11011_);
  and (_11055_, _11054_, _11007_);
  nor (_11056_, _11054_, _11007_);
  nor (_11057_, _11056_, _11055_);
  or (_11058_, _11057_, _08477_);
  or (_11059_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_11060_, _11059_, _10964_);
  and (_11061_, _11060_, _11058_);
  or (_09669_, _11061_, _10978_);
  and (_11062_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_11063_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor (_11064_, _11063_, _11062_);
  and (_11065_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_11066_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_11067_, _11066_, _11065_);
  and (_11068_, _11067_, _11064_);
  and (_11069_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_11070_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor (_11071_, _11070_, _11069_);
  and (_11072_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_11073_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_11074_, _11073_, _11072_);
  and (_11075_, _11074_, _11071_);
  and (_11076_, _11075_, _11068_);
  nor (_11077_, _11076_, _07378_);
  and (_11078_, _09009_, _07378_);
  nor (_11079_, _11078_, _11077_);
  nor (_09677_, _11079_, rst);
  or (_11080_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  not (_11081_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand (_11082_, _07493_, _11081_);
  and (_11083_, _11082_, _06989_);
  and (_09687_, _11083_, _11080_);
  or (_11084_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  not (_11085_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand (_11086_, _07493_, _11085_);
  and (_11087_, _11086_, _06989_);
  and (_09691_, _11087_, _11084_);
  and (_11088_, _09891_, _08880_);
  and (_11089_, _09893_, _08822_);
  not (_11090_, _11089_);
  or (_11091_, _11090_, _09648_);
  and (_11092_, _09897_, _08726_);
  not (_11093_, _11092_);
  not (_11094_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_11095_, _10574_, _09902_);
  nor (_11096_, _11095_, _11094_);
  and (_11097_, _11095_, _09636_);
  or (_11098_, _11097_, _11096_);
  and (_11099_, _11098_, _11093_);
  and (_11100_, _11092_, word_in[8]);
  or (_11101_, _11100_, _11089_);
  or (_11102_, _11101_, _11099_);
  and (_11103_, _11102_, _11091_);
  or (_11104_, _11103_, _11088_);
  not (_11105_, _11088_);
  or (_11106_, _11105_, word_in[24]);
  and (_14649_, _11106_, _11104_);
  or (_11107_, _11090_, _09801_);
  not (_11108_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_11109_, _11095_, _11108_);
  and (_11110_, _11095_, _09660_);
  or (_11111_, _11110_, _11109_);
  and (_11112_, _11111_, _11093_);
  and (_11113_, _11092_, word_in[9]);
  or (_11114_, _11113_, _11089_);
  or (_11115_, _11114_, _11112_);
  and (_11116_, _11115_, _11107_);
  or (_11117_, _11116_, _11088_);
  or (_11118_, _11105_, word_in[25]);
  and (_14650_, _11118_, _11117_);
  or (_11119_, _11090_, _09816_);
  not (_11120_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_11121_, _11095_, _11120_);
  and (_11122_, _11095_, _09674_);
  or (_11123_, _11122_, _11121_);
  and (_11124_, _11123_, _11093_);
  and (_11125_, _11092_, word_in[10]);
  or (_11126_, _11125_, _11089_);
  or (_11127_, _11126_, _11124_);
  and (_11128_, _11127_, _11119_);
  and (_11129_, _11128_, _11105_);
  and (_11130_, _11088_, word_in[26]);
  or (_14651_, _11130_, _11129_);
  or (_11131_, _11090_, _09829_);
  not (_11132_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_11133_, _11095_, _11132_);
  and (_11134_, _11095_, _09690_);
  or (_11135_, _11134_, _11133_);
  and (_11136_, _11135_, _11093_);
  and (_11137_, _11092_, word_in[11]);
  or (_11138_, _11137_, _11089_);
  or (_11139_, _11138_, _11136_);
  and (_11140_, _11139_, _11131_);
  or (_11141_, _11140_, _11088_);
  or (_11142_, _11105_, word_in[27]);
  and (_14652_, _11142_, _11141_);
  or (_11143_, _11090_, _09842_);
  not (_11144_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_11145_, _11095_, _11144_);
  and (_11146_, _11095_, _09707_);
  or (_11147_, _11146_, _11145_);
  and (_11148_, _11147_, _11093_);
  and (_11149_, _11092_, word_in[12]);
  or (_11150_, _11149_, _11089_);
  or (_11151_, _11150_, _11148_);
  and (_11152_, _11151_, _11143_);
  or (_11153_, _11152_, _11088_);
  or (_11154_, _11105_, word_in[28]);
  and (_14653_, _11154_, _11153_);
  or (_11155_, _11090_, _09855_);
  not (_11156_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_11157_, _11095_, _11156_);
  and (_11158_, _11095_, _09722_);
  or (_11159_, _11158_, _11157_);
  and (_11160_, _11159_, _11093_);
  and (_11161_, _11092_, word_in[13]);
  or (_11162_, _11161_, _11089_);
  or (_11163_, _11162_, _11160_);
  and (_11164_, _11163_, _11155_);
  or (_11165_, _11164_, _11088_);
  or (_11166_, _11105_, word_in[29]);
  and (_14654_, _11166_, _11165_);
  or (_11167_, _11090_, _09871_);
  not (_11168_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_11169_, _11095_, _11168_);
  and (_11170_, _11095_, _09735_);
  or (_11171_, _11170_, _11169_);
  and (_11172_, _11171_, _11093_);
  and (_11173_, _11092_, word_in[14]);
  or (_11174_, _11173_, _11089_);
  or (_11175_, _11174_, _11172_);
  and (_11176_, _11175_, _11167_);
  or (_11177_, _11176_, _11088_);
  or (_11178_, _11105_, word_in[30]);
  and (_09711_, _11178_, _11177_);
  or (_11179_, _11090_, _08942_);
  nor (_11180_, _11095_, _08760_);
  and (_11181_, _11095_, _08953_);
  or (_11182_, _11181_, _11180_);
  and (_11183_, _11182_, _11093_);
  and (_11184_, _11092_, word_in[15]);
  or (_11185_, _11184_, _11089_);
  or (_11186_, _11185_, _11183_);
  and (_11187_, _11186_, _11179_);
  or (_11188_, _11187_, _11088_);
  or (_11189_, _11105_, word_in[31]);
  and (_14655_, _11189_, _11188_);
  and (_11190_, _07490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_11191_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_11192_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_11193_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_11194_, _11193_, _11192_);
  and (_11195_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_11196_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_11197_, _11196_, _11195_);
  and (_11198_, _11197_, _11194_);
  and (_11199_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_11201_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_11202_, _11201_, _11199_);
  and (_11203_, _11202_, _11198_);
  nor (_11204_, _11203_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11205_, _11204_, _11191_);
  nor (_11206_, _11205_, _07490_);
  nor (_11207_, _11206_, _11190_);
  nor (_09733_, _11207_, rst);
  nor (_11208_, _07325_, _06716_);
  and (_11209_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_11210_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_11211_, _11210_, _11209_);
  and (_11212_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_11213_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_11214_, _11213_, _11212_);
  and (_11215_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_11216_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_11217_, _11216_, _11215_);
  and (_11218_, _11217_, _11214_);
  and (_11219_, _11218_, _11211_);
  nor (_11220_, _11219_, _08477_);
  nor (_11221_, _11220_, _11208_);
  nor (_09747_, _11221_, rst);
  and (_11223_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  not (_11224_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_11225_, _07493_, _11224_);
  or (_11226_, _11225_, _11223_);
  and (_09779_, _11226_, _06989_);
  and (_11227_, _08945_, _08726_);
  not (_11229_, _11227_);
  not (_11230_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_11231_, _10574_, _08948_);
  nor (_11232_, _11231_, _11230_);
  and (_11233_, _11231_, _09636_);
  or (_11234_, _11233_, _11232_);
  and (_11235_, _11234_, _11229_);
  and (_11236_, _10023_, _08822_);
  and (_11237_, _11227_, word_in[8]);
  or (_11238_, _11237_, _11236_);
  or (_11239_, _11238_, _11235_);
  and (_11240_, _08935_, _09299_);
  not (_11241_, _11240_);
  not (_11242_, _11236_);
  or (_11243_, _11242_, _09648_);
  and (_11244_, _11243_, _11241_);
  and (_11245_, _11244_, _11239_);
  and (_11246_, _11240_, word_in[24]);
  or (_14656_, _11246_, _11245_);
  not (_11247_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_11248_, _11231_, _11247_);
  and (_11249_, _11231_, _09660_);
  or (_11250_, _11249_, _11248_);
  and (_11251_, _11250_, _11229_);
  and (_11252_, _11227_, word_in[9]);
  or (_11253_, _11252_, _11236_);
  or (_11254_, _11253_, _11251_);
  or (_11255_, _11242_, _09801_);
  and (_11256_, _11255_, _11241_);
  and (_11257_, _11256_, _11254_);
  and (_11258_, _11240_, word_in[25]);
  or (_14657_, _11258_, _11257_);
  not (_11260_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_11261_, _11231_, _11260_);
  and (_11262_, _11231_, _09674_);
  or (_11263_, _11262_, _11261_);
  and (_11264_, _11263_, _11229_);
  and (_11265_, _11227_, word_in[10]);
  or (_11266_, _11265_, _11236_);
  or (_11267_, _11266_, _11264_);
  or (_11269_, _11242_, _09816_);
  and (_11270_, _11269_, _11241_);
  and (_11271_, _11270_, _11267_);
  and (_11272_, _11240_, word_in[26]);
  or (_14658_, _11272_, _11271_);
  not (_11273_, _07493_);
  and (_11274_, _11045_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_11275_, _11274_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_11276_, _11275_, _11273_);
  and (_11277_, _11276_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_11278_, _11276_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_11279_, _11278_, _11277_);
  not (_11280_, _07412_);
  and (_11281_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_11282_, _07324_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_11283_, _11282_);
  or (_11284_, _08529_, _07327_);
  nor (_11285_, _07325_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_11286_, _11285_, _07362_);
  and (_11287_, _11286_, _11284_);
  nor (_11288_, _11287_, _09388_);
  and (_11289_, _11288_, _09547_);
  and (_11290_, _11289_, _07365_);
  or (_11291_, _08561_, _07327_);
  nor (_11292_, _07325_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_11293_, _11292_, _07362_);
  and (_11294_, _11293_, _11291_);
  not (_11295_, _11294_);
  or (_11296_, _08463_, _07327_);
  nor (_11297_, _07325_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_11298_, _11297_, _07362_);
  and (_11299_, _11298_, _11296_);
  nand (_11300_, _08576_, _07326_);
  nor (_11301_, _07325_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_11302_, _11301_, _07362_);
  and (_11303_, _11302_, _11300_);
  not (_11304_, _11303_);
  and (_11305_, _11304_, _11299_);
  and (_11306_, _11305_, _11295_);
  nor (_11308_, _08545_, _07327_);
  not (_11309_, _11308_);
  nor (_11310_, _07325_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_11311_, _11310_, _07362_);
  and (_11312_, _11311_, _11309_);
  and (_11313_, _11312_, _11306_);
  and (_11314_, _11313_, _11290_);
  not (_11315_, _11314_);
  not (_11316_, _11312_);
  and (_11317_, _11305_, _11294_);
  and (_11319_, _11317_, _11316_);
  and (_11320_, _11319_, _11290_);
  nor (_11321_, _11304_, _11299_);
  and (_11322_, _11321_, _11294_);
  and (_11324_, _11322_, _11312_);
  and (_11325_, _11324_, _11290_);
  nor (_11326_, _11325_, _11320_);
  and (_11327_, _11326_, _11315_);
  and (_11328_, _11316_, _11306_);
  nor (_11329_, _09547_, _07365_);
  not (_11330_, _11287_);
  and (_11331_, _11330_, _09388_);
  and (_11332_, _11331_, _11329_);
  and (_11333_, _11332_, _11328_);
  and (_11334_, _11332_, _11319_);
  nor (_11335_, _11334_, _11333_);
  and (_11336_, _11335_, _11327_);
  nor (_11337_, _11336_, _11283_);
  not (_11338_, _11337_);
  and (_11339_, _11329_, _11288_);
  not (_11340_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_11341_, \oc8051_top_1.oc8051_decoder1.state [1], _06406_);
  and (_11342_, _11341_, _11340_);
  and (_11343_, _11342_, _11321_);
  and (_11344_, _11343_, _11339_);
  not (_11345_, _07324_);
  nor (_11346_, _11335_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11347_, _11346_, _11345_);
  nor (_11348_, _11347_, _11344_);
  and (_11349_, _11348_, _11338_);
  nor (_11350_, _11349_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11351_, _11350_, _11281_);
  and (_11352_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11353_, _06406_, \oc8051_top_1.oc8051_decoder1.state [0]);
  nor (_11354_, _11303_, _11299_);
  and (_11355_, _11354_, _11295_);
  and (_11356_, _11355_, _11312_);
  and (_11358_, _11356_, _11339_);
  and (_11359_, _11354_, _11294_);
  and (_11360_, _11359_, _11339_);
  nor (_11361_, _11360_, _11358_);
  not (_11363_, _11361_);
  and (_11364_, _11321_, _11295_);
  and (_11365_, _11364_, _11339_);
  and (_11366_, _11365_, _11342_);
  nor (_11367_, _11366_, _11363_);
  nor (_11368_, _11367_, _11353_);
  and (_11369_, _11339_, _11321_);
  and (_11370_, _11369_, _11342_);
  not (_11371_, _11370_);
  nor (_11372_, _11371_, _11368_);
  nor (_11373_, _11304_, _11294_);
  and (_11374_, _11373_, _11299_);
  and (_11375_, _11374_, _11312_);
  and (_11376_, _11375_, _11339_);
  and (_11377_, _09547_, _09388_);
  nor (_11378_, _11287_, _11312_);
  and (_11379_, _11378_, _11377_);
  and (_11380_, _11379_, _11306_);
  nor (_11381_, _11380_, _11376_);
  and (_11382_, _11289_, _07383_);
  and (_11383_, _11359_, _11382_);
  and (_11385_, _11379_, _11322_);
  nor (_11386_, _11385_, _11383_);
  and (_11387_, _11379_, _11364_);
  and (_11388_, _11303_, _11294_);
  and (_11389_, _11388_, _11299_);
  and (_11390_, _11379_, _11389_);
  nor (_11391_, _11390_, _11387_);
  and (_11392_, _11391_, _11386_);
  and (_11393_, _11392_, _11381_);
  and (_11394_, _11377_, _11330_);
  and (_11395_, _11394_, _11374_);
  and (_11396_, _11394_, _11312_);
  and (_11397_, _11396_, _11306_);
  nor (_11398_, _11397_, _11395_);
  and (_11399_, _11317_, _11312_);
  and (_11400_, _11399_, _11394_);
  and (_11401_, _11355_, _11394_);
  nor (_11402_, _11401_, _11400_);
  and (_11403_, _11364_, _11312_);
  and (_11404_, _11403_, _11394_);
  and (_11405_, _11359_, _11394_);
  nor (_11406_, _11405_, _11404_);
  and (_11407_, _11406_, _11402_);
  and (_11408_, _11407_, _11398_);
  and (_11409_, _11408_, _11393_);
  and (_11410_, _11409_, _11327_);
  nor (_11411_, _11410_, _11283_);
  and (_11412_, _11341_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_11413_, _11412_, _11383_);
  or (_11414_, _11413_, _11411_);
  nor (_11415_, _11414_, _11372_);
  nor (_11416_, _11415_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11417_, _11416_, _11352_);
  not (_11418_, _11417_);
  and (_11419_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_11420_, _09547_);
  and (_11421_, _11420_, _07365_);
  and (_11422_, _11421_, _11331_);
  and (_11423_, _11422_, _11356_);
  not (_11424_, _11423_);
  and (_11425_, _11422_, _11375_);
  and (_11426_, _11399_, _11339_);
  nor (_11427_, _11426_, _11425_);
  and (_11428_, _11427_, _11424_);
  and (_11429_, _11382_, _11324_);
  and (_11430_, _11364_, _11316_);
  and (_11431_, _11430_, _11289_);
  nor (_11432_, _11431_, _11429_);
  and (_11433_, _11339_, _11319_);
  and (_11435_, _11430_, _11422_);
  nor (_11436_, _11435_, _11433_);
  and (_11437_, _11399_, _11382_);
  and (_11438_, _11374_, _11316_);
  and (_11439_, _11438_, _11382_);
  nor (_11440_, _11439_, _11437_);
  and (_11441_, _11440_, _11436_);
  and (_11442_, _11441_, _11432_);
  and (_11443_, _11442_, _11428_);
  not (_11444_, _11443_);
  nor (_11445_, _11403_, _11359_);
  not (_11446_, _11422_);
  nor (_11447_, _11446_, _11445_);
  or (_11448_, _11375_, _11313_);
  and (_11449_, _11448_, _11382_);
  or (_11450_, _11449_, _11447_);
  and (_11451_, _11322_, _11316_);
  and (_11452_, _11422_, _11451_);
  and (_11453_, _11438_, _11422_);
  nor (_11454_, _11453_, _11452_);
  and (_11455_, _11382_, _11328_);
  and (_11456_, _11403_, _11289_);
  nor (_11457_, _11456_, _11455_);
  nand (_11458_, _11457_, _11454_);
  or (_11459_, _11458_, _11450_);
  and (_11460_, _11451_, _11289_);
  and (_11461_, _11422_, _11328_);
  and (_11462_, _11394_, _11316_);
  and (_11463_, _11462_, _11317_);
  or (_11464_, _11463_, _11461_);
  or (_11466_, _11464_, _11460_);
  and (_11467_, _11389_, _11316_);
  and (_11468_, _11467_, _11422_);
  and (_11469_, _11422_, _11312_);
  and (_11470_, _11469_, _11305_);
  or (_11471_, _11470_, _11468_);
  and (_11472_, _11355_, _11316_);
  and (_11473_, _11472_, _11422_);
  and (_11474_, _11382_, _11319_);
  or (_11475_, _11474_, _11473_);
  or (_11476_, _11475_, _11471_);
  and (_11477_, _11374_, _11339_);
  nor (_11478_, _11330_, _11312_);
  and (_11479_, _11478_, _11305_);
  and (_11480_, _11479_, _11294_);
  or (_11481_, _11480_, _11477_);
  or (_11482_, _11481_, _11383_);
  or (_11483_, _11482_, _11363_);
  or (_11484_, _11483_, _11476_);
  or (_11485_, _11484_, _11466_);
  or (_11488_, _11485_, _11459_);
  nor (_11489_, _11488_, _11444_);
  nor (_11490_, _11489_, _11283_);
  nor (_11491_, _11490_, _11413_);
  and (_11492_, _11491_, _11371_);
  nor (_11493_, _11492_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11494_, _11493_, _11419_);
  and (_11495_, _11494_, _11418_);
  and (_11496_, _11495_, _11351_);
  and (_11497_, _11496_, _11280_);
  nor (_11498_, _11494_, _11418_);
  and (_11499_, _11351_, _11498_);
  nor (_11500_, _07325_, _06657_);
  and (_11501_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_11502_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_11503_, _11502_, _11501_);
  and (_11504_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_11505_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_11506_, _11505_, _11504_);
  and (_11507_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_11508_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_11509_, _11508_, _11507_);
  and (_11510_, _11509_, _11506_);
  and (_11511_, _11510_, _11503_);
  nor (_11512_, _11511_, _08477_);
  nor (_11513_, _11512_, _11500_);
  not (_11514_, _11513_);
  and (_11515_, _11514_, _11499_);
  nor (_11516_, _11515_, _11497_);
  nor (_11517_, _11494_, _11417_);
  and (_11518_, _11351_, _11517_);
  and (_11519_, _09239_, _07089_);
  not (_11520_, _11519_);
  nor (_11521_, _11520_, _07317_);
  and (_11522_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_11523_, _11521_, _11522_);
  and (_11524_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_11525_, _07106_, _06700_);
  not (_11526_, _11525_);
  and (_11527_, _11526_, _09213_);
  and (_11528_, _11527_, _09210_);
  and (_11529_, _11528_, _09202_);
  nor (_11530_, _11529_, _11520_);
  nor (_11531_, _11530_, _11524_);
  and (_11532_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_11533_, _11519_, _09009_);
  nor (_11534_, _11533_, _11532_);
  nor (_11535_, _11519_, _06508_);
  and (_11536_, _11519_, _09599_);
  nor (_11537_, _11536_, _11535_);
  and (_11538_, _11537_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_11539_, _11538_, _11534_);
  and (_11540_, _11539_, _11531_);
  and (_11541_, _11540_, _11523_);
  nor (_11542_, _11540_, _11523_);
  nor (_11543_, _11542_, _11541_);
  nor (_11545_, _11543_, _06409_);
  nor (_11546_, _11545_, _06438_);
  nor (_11547_, _11546_, _11519_);
  nor (_11548_, _11547_, _11521_);
  not (_11549_, _11548_);
  and (_11550_, _11549_, _11518_);
  not (_11551_, _07319_);
  and (_11552_, _11351_, _11417_);
  and (_11553_, _11552_, _11494_);
  and (_11554_, _11553_, _11551_);
  nor (_11555_, _11554_, _11550_);
  and (_11556_, _11555_, _11516_);
  nor (_11557_, _11556_, _06448_);
  and (_11558_, _11556_, _06448_);
  nor (_11559_, _11558_, _11557_);
  not (_11560_, _06499_);
  and (_11561_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_11562_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_11563_, _11562_, _11561_);
  and (_11564_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_11565_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor (_11566_, _11565_, _11564_);
  and (_11567_, _11566_, _11563_);
  and (_11568_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_11569_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_11570_, _11569_, _11568_);
  and (_11571_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_11572_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_11573_, _11572_, _11571_);
  and (_11574_, _11573_, _11570_);
  and (_11575_, _11574_, _11567_);
  nor (_11576_, _11575_, _07378_);
  not (_11577_, _07040_);
  and (_11578_, _07378_, _11577_);
  nor (_11579_, _11578_, _11576_);
  not (_11580_, _11579_);
  and (_11581_, _11496_, _11580_);
  not (_11582_, _11581_);
  and (_11583_, _11519_, _07040_);
  nor (_11584_, _11520_, _07260_);
  and (_11585_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_11586_, _11585_, _11584_);
  and (_11587_, _11586_, _11541_);
  and (_11588_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_11589_, _11520_, _07118_);
  nor (_11590_, _11589_, _11588_);
  and (_11591_, _11590_, _11587_);
  and (_11593_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_11594_, _11520_, _10970_);
  nor (_11595_, _11594_, _11593_);
  and (_11596_, _11595_, _11591_);
  nor (_11597_, _11519_, _06487_);
  nor (_11598_, _11597_, _11596_);
  and (_11599_, _11597_, _11596_);
  or (_11600_, _11599_, _11598_);
  nor (_11601_, _11600_, _06409_);
  nor (_11602_, _11519_, _06491_);
  not (_11603_, _11602_);
  nor (_11604_, _11603_, _11601_);
  nor (_11605_, _11604_, _11583_);
  and (_11606_, _11605_, _11517_);
  not (_11607_, _11606_);
  not (_11608_, _08479_);
  and (_11609_, _11498_, _11608_);
  not (_11610_, _11351_);
  nor (_11611_, _11610_, _11609_);
  and (_11612_, _11611_, _11607_);
  and (_11613_, _11612_, _11582_);
  nor (_11614_, _11613_, _11560_);
  and (_11615_, _11613_, _11560_);
  nor (_11616_, _11615_, _11614_);
  nor (_11617_, _11495_, _11351_);
  not (_11618_, _10806_);
  and (_11619_, _11499_, _11618_);
  nor (_11620_, _11619_, _11617_);
  nor (_11621_, _11595_, _11591_);
  nor (_11622_, _11621_, _11596_);
  nor (_11623_, _11622_, _06409_);
  nor (_11624_, _11623_, _06455_);
  nor (_11625_, _11624_, _11519_);
  nor (_11626_, _11625_, _11594_);
  not (_11627_, _11626_);
  and (_11628_, _11627_, _11518_);
  and (_11629_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_11630_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_11631_, _11630_, _11629_);
  and (_11632_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_11634_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor (_11635_, _11634_, _11632_);
  and (_11636_, _11635_, _11631_);
  and (_11637_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_11638_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_11639_, _11638_, _11637_);
  and (_11640_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_11641_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_11642_, _11641_, _11640_);
  and (_11643_, _11642_, _11639_);
  and (_11644_, _11643_, _11636_);
  nor (_11645_, _11644_, _07378_);
  not (_11646_, _10970_);
  and (_11647_, _11646_, _07378_);
  nor (_11648_, _11647_, _11645_);
  not (_11649_, _11648_);
  and (_11650_, _11649_, _11496_);
  nor (_11651_, _11650_, _11628_);
  and (_11652_, _11651_, _11620_);
  nor (_11653_, _11652_, _07452_);
  and (_11654_, _11652_, _07452_);
  nor (_11655_, _11654_, _11653_);
  and (_11656_, _11655_, _11616_);
  nor (_11657_, _07325_, _06600_);
  and (_11658_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_11659_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_11660_, _11659_, _11658_);
  and (_11661_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_11662_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_11663_, _11662_, _11661_);
  and (_11664_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_11665_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_11666_, _11665_, _11664_);
  and (_11667_, _11666_, _11663_);
  and (_11668_, _11667_, _11660_);
  nor (_11669_, _11668_, _08477_);
  nor (_11670_, _11669_, _11657_);
  not (_11671_, _11670_);
  and (_11672_, _11671_, _11499_);
  not (_11673_, _11498_);
  and (_11674_, _11617_, _11673_);
  nor (_11675_, _11674_, _11672_);
  nor (_11676_, _11590_, _11587_);
  nor (_11678_, _11676_, _11591_);
  nor (_11679_, _11678_, _06409_);
  nor (_11680_, _11679_, _06467_);
  nor (_11681_, _11680_, _11519_);
  nor (_11682_, _11681_, _11589_);
  not (_11683_, _11682_);
  and (_11684_, _11683_, _11518_);
  not (_11685_, _07450_);
  and (_11686_, _11496_, _11685_);
  nor (_11687_, _11686_, _11684_);
  and (_11688_, _11687_, _11675_);
  nor (_11689_, _11688_, _06478_);
  and (_11690_, _11688_, _06478_);
  nor (_11691_, _11690_, _11689_);
  nor (_11692_, _11586_, _11541_);
  nor (_11693_, _11692_, _11587_);
  nor (_11694_, _11693_, _06409_);
  nor (_11695_, _11694_, _06413_);
  nor (_11696_, _11695_, _11519_);
  nor (_11697_, _11696_, _11584_);
  not (_11698_, _11697_);
  and (_11699_, _11698_, _11518_);
  and (_11700_, _11610_, _11417_);
  nor (_11701_, _11700_, _11699_);
  not (_11702_, _07431_);
  and (_11703_, _11496_, _11702_);
  nor (_11704_, _07325_, _06628_);
  and (_11705_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_11706_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_11707_, _11706_, _11705_);
  and (_11708_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_11709_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_11710_, _11709_, _11708_);
  and (_11711_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_11712_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_11713_, _11712_, _11711_);
  and (_11714_, _11713_, _11710_);
  and (_11715_, _11714_, _11707_);
  nor (_11716_, _11715_, _08477_);
  nor (_11717_, _11716_, _11704_);
  not (_11718_, _11717_);
  and (_11719_, _11718_, _11499_);
  nor (_11720_, _11719_, _11703_);
  and (_11721_, _11553_, _07382_);
  not (_11722_, _11721_);
  and (_11723_, _11722_, _11720_);
  and (_11724_, _11723_, _11701_);
  nor (_11725_, _11724_, _07084_);
  and (_11726_, _11724_, _07084_);
  nor (_11727_, _11726_, _11725_);
  and (_11728_, _11727_, _11691_);
  and (_11729_, _11728_, _11656_);
  and (_11730_, _11729_, _11559_);
  not (_11731_, _11079_);
  and (_11732_, _11496_, _11731_);
  and (_11733_, _11495_, _11610_);
  nor (_11734_, _11538_, _11534_);
  nor (_11735_, _11734_, _11539_);
  nor (_11736_, _11735_, _06409_);
  nor (_11737_, _11736_, _06528_);
  nor (_11738_, _11737_, _11519_);
  nor (_11739_, _11738_, _11533_);
  not (_11740_, _11739_);
  and (_11741_, _11740_, _11518_);
  or (_11742_, _11741_, _11733_);
  and (_11743_, _11553_, _09547_);
  not (_11744_, _11221_);
  and (_11745_, _11499_, _11744_);
  or (_11746_, _11745_, _11743_);
  or (_11747_, _11746_, _11742_);
  nor (_11748_, _11747_, _11732_);
  nor (_11749_, _11748_, _06537_);
  and (_11750_, _11748_, _06537_);
  nor (_11751_, _11750_, _11749_);
  and (_11752_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_11753_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_11754_, _11753_, _11752_);
  and (_11755_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_11756_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_11757_, _11756_, _11755_);
  and (_11758_, _11757_, _11754_);
  and (_11759_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_11760_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_11761_, _11760_, _11759_);
  and (_11762_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_11763_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor (_11764_, _11763_, _11762_);
  and (_11765_, _11764_, _11761_);
  and (_11766_, _11765_, _11758_);
  nor (_11767_, _11766_, _07378_);
  and (_11768_, _09599_, _07378_);
  nor (_11769_, _11768_, _11767_);
  not (_11770_, _11769_);
  and (_11771_, _11770_, _11496_);
  nor (_11772_, _07325_, _06737_);
  and (_11773_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_11774_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_11775_, _11774_, _11773_);
  and (_11776_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_11777_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_11778_, _11777_, _11776_);
  and (_11779_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_11780_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_11781_, _11780_, _11779_);
  and (_11782_, _11781_, _11778_);
  and (_11783_, _11782_, _11775_);
  nor (_11784_, _11783_, _08477_);
  nor (_11785_, _11784_, _11772_);
  not (_11786_, _11785_);
  and (_11787_, _11786_, _11499_);
  nor (_11788_, _11787_, _11771_);
  nor (_11789_, _11537_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_11790_, _11789_, _11538_);
  nor (_11791_, _11790_, _06409_);
  nor (_11792_, _11791_, _06509_);
  nor (_11793_, _11792_, _11519_);
  nor (_11794_, _11793_, _11536_);
  not (_11795_, _11794_);
  and (_11796_, _11795_, _11518_);
  and (_11797_, _11553_, _07365_);
  nor (_11798_, _11797_, _11796_);
  and (_11799_, _11798_, _11788_);
  nor (_11800_, _11799_, _06514_);
  and (_11801_, _11799_, _06514_);
  or (_11802_, _11801_, _11800_);
  nor (_11803_, _11802_, _11751_);
  not (_11804_, _06484_);
  and (_11805_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_11806_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_11807_, _11806_, _11805_);
  and (_11808_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_11809_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor (_11810_, _11809_, _11808_);
  and (_11811_, _11810_, _11807_);
  and (_11812_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and (_11813_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_11814_, _11813_, _11812_);
  and (_11815_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_11816_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_11817_, _11816_, _11815_);
  and (_11818_, _11817_, _11814_);
  and (_11819_, _11818_, _11811_);
  nor (_11820_, _11819_, _07378_);
  not (_11821_, _11529_);
  and (_11822_, _11821_, _07378_);
  nor (_11823_, _11822_, _11820_);
  not (_11824_, _11823_);
  and (_11825_, _11824_, _11496_);
  nor (_11827_, _07325_, _06685_);
  and (_11828_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_11829_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_11830_, _11829_, _11828_);
  and (_11832_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_11833_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_11834_, _11833_, _11832_);
  and (_11835_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_11836_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_11837_, _11836_, _11835_);
  and (_11838_, _11837_, _11834_);
  and (_11839_, _11838_, _11830_);
  nor (_11840_, _11839_, _08477_);
  nor (_11841_, _11840_, _11827_);
  not (_11842_, _11841_);
  and (_11843_, _11842_, _11499_);
  nor (_11844_, _11843_, _11825_);
  nor (_11845_, _11539_, _11531_);
  nor (_11846_, _11845_, _11540_);
  nor (_11848_, _11846_, _06409_);
  nor (_11849_, _11848_, _06517_);
  nor (_11850_, _11849_, _11519_);
  nor (_11851_, _11850_, _11530_);
  not (_11852_, _11851_);
  and (_11853_, _11852_, _11518_);
  and (_11855_, _11553_, _09388_);
  nor (_11856_, _11855_, _11853_);
  and (_11857_, _11856_, _11844_);
  nor (_11858_, _11857_, _06525_);
  and (_11859_, _11857_, _06525_);
  nor (_11860_, _11859_, _11858_);
  nor (_11861_, _11860_, _11804_);
  and (_11862_, _11861_, _11803_);
  and (_11863_, _11862_, _11730_);
  nor (_11864_, _06499_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_11865_, _11864_, _11863_);
  not (_11866_, _11865_);
  not (_11867_, _11344_);
  and (_11868_, _11344_, _11295_);
  nor (_11869_, _11868_, _11363_);
  nor (_11870_, _11869_, _11353_);
  and (_11871_, _11870_, _11867_);
  nor (_11872_, _06984_, _06539_);
  and (_11873_, _11872_, _11730_);
  and (_11874_, _11873_, _11871_);
  not (_11875_, _11342_);
  not (_11876_, _06849_);
  and (_11877_, _06898_, _11876_);
  nor (_11878_, _06898_, _11876_);
  nor (_11879_, _11878_, _11877_);
  not (_11880_, _11879_);
  or (_11881_, _08089_, _06881_);
  nor (_11882_, _11881_, _06878_);
  and (_11883_, _11882_, _11867_);
  and (_11884_, _11883_, _08405_);
  nand (_11885_, _11884_, _08234_);
  nor (_11886_, _11885_, _11368_);
  not (_11887_, _08322_);
  and (_11888_, _09100_, _11887_);
  and (_11889_, _11888_, _11886_);
  and (_11890_, _11889_, _11880_);
  not (_11891_, _11890_);
  and (_11892_, _11868_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  not (_11894_, _11892_);
  nor (_11895_, _11870_, _11867_);
  nor (_11896_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_11897_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_11898_, _11897_, _11896_);
  nor (_11899_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_11900_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_11901_, _11900_, _11899_);
  and (_11902_, _11901_, _11898_);
  and (_11903_, _11902_, _11895_);
  and (_11904_, _11871_, _06776_);
  nor (_11905_, _11904_, _11903_);
  and (_11906_, _11905_, _11894_);
  and (_11907_, _11906_, _11891_);
  and (_11908_, _11331_, _11420_);
  and (_11909_, _11908_, _11399_);
  nor (_11910_, _11909_, _11425_);
  and (_11911_, _11287_, _11312_);
  and (_11912_, _11911_, _11374_);
  and (_11913_, _11360_, _11312_);
  nor (_11914_, _11913_, _11912_);
  and (_11915_, _11914_, _11910_);
  not (_11916_, _11339_);
  nor (_11917_, _11403_, _11324_);
  nor (_11918_, _11917_, _11916_);
  and (_11919_, _11911_, _11317_);
  nor (_11920_, _11919_, _11400_);
  not (_11921_, _11920_);
  nor (_11922_, _11921_, _11918_);
  and (_11923_, _11922_, _11915_);
  and (_11924_, _11923_, _11907_);
  or (_11925_, _11430_, _11451_);
  nand (_11926_, _11925_, _11339_);
  and (_11927_, _11359_, _11316_);
  and (_11928_, _11927_, _11339_);
  or (_11929_, _11928_, _11358_);
  nor (_11930_, _11907_, _11929_);
  and (_11931_, _11930_, _11926_);
  nor (_11932_, _11931_, _11924_);
  not (_11933_, _11932_);
  and (_11934_, _11290_, _11312_);
  and (_11935_, _11322_, _11934_);
  and (_11936_, _11328_, _11339_);
  nor (_11937_, _11936_, _11935_);
  and (_11938_, _11937_, _11933_);
  nor (_11939_, _11938_, _11875_);
  and (_11940_, _11421_, _11288_);
  and (_11941_, _11355_, _11382_);
  nor (_11942_, _11941_, _11940_);
  nor (_11943_, _11942_, _11283_);
  and (_11944_, _11383_, _11341_);
  nor (_11945_, _11944_, _11943_);
  not (_11946_, _11945_);
  nor (_11947_, _11946_, _11939_);
  nand (_11948_, _08041_, _08125_);
  and (_11949_, _11948_, _11895_);
  nor (_11950_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_11951_, _11950_);
  nor (_11952_, _06448_, _06463_);
  and (_11953_, _11952_, _07085_);
  and (_11954_, _11953_, _06500_);
  or (_11955_, _11954_, _11951_);
  nor (_11956_, _11955_, _07291_);
  not (_11957_, _11956_);
  and (_11958_, _11957_, _11868_);
  nor (_11959_, _11958_, _11949_);
  not (_11960_, _11959_);
  nor (_11961_, _11960_, _11947_);
  not (_11962_, _11961_);
  nor (_11963_, _11962_, _11874_);
  and (_11964_, _11963_, _11866_);
  nor (_11965_, _11964_, _11279_);
  not (_11966_, _09145_);
  and (_11968_, _11342_, _11325_);
  nor (_11969_, _11968_, _11943_);
  nand (_11970_, _11910_, _11361_);
  or (_11971_, _11970_, _11921_);
  and (_11972_, _11971_, _11342_);
  not (_11973_, _11972_);
  and (_11974_, _11941_, _11282_);
  nor (_11975_, _11974_, _11413_);
  and (_11976_, _11975_, _11973_);
  nor (_11977_, _11912_, _11369_);
  and (_11978_, _11977_, _11937_);
  nor (_11979_, _11978_, _11875_);
  not (_11980_, _11979_);
  nand (_11981_, _11360_, _11282_);
  and (_11982_, _11981_, _11973_);
  and (_11983_, _11982_, _11980_);
  and (_11984_, _11983_, _11976_);
  and (_11985_, _11984_, _11969_);
  or (_11986_, _11985_, _11968_);
  and (_11987_, _11986_, _11966_);
  not (_11988_, _11974_);
  not (_11989_, _11413_);
  and (_11990_, _11981_, _11989_);
  and (_11991_, _11990_, _11988_);
  and (_11992_, _11991_, _11973_);
  and (_11993_, _11992_, _11670_);
  nand (_11994_, _11991_, _11973_);
  and (_11995_, _07490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  and (_11996_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_11998_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_11999_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_12001_, _11999_, _11998_);
  and (_12002_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_12003_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_12004_, _12003_, _12002_);
  and (_12005_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_12006_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_12007_, _12006_, _12005_);
  and (_12008_, _12007_, _12004_);
  and (_12009_, _12008_, _12001_);
  nor (_12010_, _12009_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12011_, _12010_, _11996_);
  nor (_12012_, _12011_, _07490_);
  nor (_12013_, _12012_, _11995_);
  and (_12014_, _12013_, _11994_);
  nor (_12015_, _12014_, _11993_);
  and (_12016_, _12015_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_12017_, _12015_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_12018_, _12017_, _12016_);
  and (_12019_, _11992_, _11717_);
  and (_12020_, _07490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  and (_12021_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12022_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_12023_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_12024_, _12023_, _12022_);
  and (_12025_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_12026_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_12027_, _12026_, _12025_);
  and (_12028_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_12029_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_12030_, _12029_, _12028_);
  and (_12031_, _12030_, _12027_);
  and (_12032_, _12031_, _12024_);
  nor (_12033_, _12032_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12034_, _12033_, _12021_);
  nor (_12035_, _12034_, _07490_);
  nor (_12036_, _12035_, _12020_);
  and (_12037_, _12036_, _11994_);
  nor (_12038_, _12037_, _12019_);
  nand (_12040_, _12038_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_12041_, _11992_, _11513_);
  and (_12042_, _07490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_12043_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12044_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_12045_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_12046_, _12045_, _12044_);
  and (_12047_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_12048_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_12049_, _12048_, _12047_);
  and (_12050_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_12051_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_12053_, _12051_, _12050_);
  and (_12054_, _12053_, _12049_);
  and (_12055_, _12054_, _12046_);
  nor (_12056_, _12055_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12058_, _12056_, _12043_);
  nor (_12059_, _12058_, _07490_);
  nor (_12061_, _12059_, _12042_);
  and (_12062_, _12061_, _11994_);
  nor (_12063_, _12062_, _12041_);
  nor (_12064_, _12063_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_12065_, _12063_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_12066_, _11992_, _11841_);
  and (_12067_, _11994_, _11207_);
  nor (_12068_, _12067_, _12066_);
  and (_12069_, _12068_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_12070_, _11994_, _11744_);
  and (_12071_, _07490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_12072_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12073_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_12074_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_12076_, _12074_, _12073_);
  and (_12077_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_12078_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_12079_, _12078_, _12077_);
  and (_12080_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_12081_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_12083_, _12081_, _12080_);
  and (_12084_, _12083_, _12079_);
  and (_12086_, _12084_, _12076_);
  nor (_12087_, _12086_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12088_, _12087_, _12072_);
  nor (_12089_, _12088_, _07490_);
  nor (_12090_, _12089_, _12071_);
  not (_12091_, _12090_);
  or (_12092_, _12091_, _11992_);
  nand (_12093_, _12092_, _12070_);
  or (_12094_, _12093_, _06714_);
  or (_12095_, _11994_, _11786_);
  and (_12096_, _07490_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_12097_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12098_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_12099_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_12100_, _12099_, _12098_);
  and (_12101_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_12102_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_12103_, _12102_, _12101_);
  and (_12105_, _12103_, _12100_);
  and (_12106_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_12107_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_12108_, _12107_, _12106_);
  and (_12109_, _12108_, _12105_);
  nor (_12110_, _12109_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12111_, _12110_, _12097_);
  nor (_12112_, _12111_, _07490_);
  nor (_12113_, _12112_, _12096_);
  not (_12114_, _12113_);
  or (_12116_, _12114_, _11992_);
  and (_12117_, _12116_, _12095_);
  and (_12118_, _12117_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand (_12119_, _12093_, _06714_);
  and (_12120_, _12119_, _12094_);
  and (_12122_, _12120_, _12118_);
  not (_12123_, _12122_);
  nand (_12124_, _12123_, _12094_);
  nor (_12125_, _12068_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_12126_, _12125_, _12069_);
  and (_12127_, _12126_, _12124_);
  or (_12129_, _12127_, _12069_);
  nor (_12130_, _12129_, _12065_);
  nor (_12131_, _12130_, _12064_);
  or (_12132_, _12038_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_12134_, _12132_, _12040_);
  nand (_12135_, _12134_, _12131_);
  nand (_12136_, _12135_, _12040_);
  and (_12137_, _12136_, _12018_);
  or (_12138_, _12137_, _12016_);
  and (_12139_, _11992_, _10806_);
  and (_12140_, _07490_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and (_12141_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12142_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_12143_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_12144_, _12143_, _12142_);
  and (_12145_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_12146_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_12147_, _12146_, _12145_);
  and (_12148_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_12149_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_12150_, _12149_, _12148_);
  and (_12151_, _12150_, _12147_);
  and (_12152_, _12151_, _12144_);
  nor (_12153_, _12152_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12154_, _12153_, _12141_);
  nor (_12155_, _12154_, _07490_);
  nor (_12156_, _12155_, _12140_);
  and (_12157_, _12156_, _11994_);
  nor (_12158_, _12157_, _12139_);
  nand (_12159_, _12158_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_12161_, _12158_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_12162_, _12161_, _12159_);
  nand (_12163_, _12162_, _12138_);
  or (_12164_, _12162_, _12138_);
  nor (_12165_, _11979_, _11972_);
  and (_12166_, _11981_, _12165_);
  and (_12167_, _11342_, _11935_);
  nor (_12168_, _12167_, _11943_);
  nor (_12169_, _12168_, _11994_);
  nor (_12171_, _12169_, _12166_);
  and (_12172_, _12171_, _12164_);
  and (_12173_, _12172_, _12163_);
  nor (_12174_, _12156_, _11988_);
  and (_12175_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_12176_, _12169_, _12165_);
  and (_12177_, _12176_, _11618_);
  or (_12178_, _12177_, _12175_);
  or (_12179_, _12178_, _12174_);
  or (_12180_, _12179_, _12173_);
  or (_12181_, _12180_, _11987_);
  and (_12182_, _12181_, _11964_);
  or (_12183_, _12182_, _11965_);
  and (_09791_, _12183_, _06989_);
  and (_12184_, _11240_, word_in[27]);
  not (_12185_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_12186_, _11231_, _12185_);
  and (_12187_, _11231_, _09690_);
  or (_12188_, _12187_, _12186_);
  and (_12189_, _12188_, _11229_);
  and (_12190_, _11227_, word_in[11]);
  or (_12191_, _12190_, _11236_);
  or (_12192_, _12191_, _12189_);
  or (_12193_, _11242_, _09829_);
  and (_12194_, _12193_, _11241_);
  and (_12195_, _12194_, _12192_);
  or (_14659_, _12195_, _12184_);
  nor (_09795_, _11823_, rst);
  not (_12196_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_12197_, _11231_, _12196_);
  and (_12198_, _11231_, _09707_);
  or (_12199_, _12198_, _12197_);
  and (_12200_, _12199_, _11229_);
  and (_12201_, _11227_, word_in[12]);
  or (_12202_, _12201_, _11236_);
  or (_12203_, _12202_, _12200_);
  or (_12204_, _11242_, _09842_);
  and (_12205_, _12204_, _11241_);
  and (_12206_, _12205_, _12203_);
  and (_12207_, _11240_, word_in[28]);
  or (_14660_, _12207_, _12206_);
  not (_12209_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_12210_, _11231_, _12209_);
  and (_12212_, _11231_, _09722_);
  or (_12213_, _12212_, _12210_);
  and (_12215_, _12213_, _11229_);
  and (_12216_, _11227_, word_in[13]);
  or (_12217_, _12216_, _11236_);
  or (_12218_, _12217_, _12215_);
  or (_12219_, _11242_, _09855_);
  and (_12221_, _12219_, _11241_);
  and (_12222_, _12221_, _12218_);
  and (_12223_, _11240_, word_in[29]);
  or (_14661_, _12223_, _12222_);
  and (_12224_, _11240_, word_in[30]);
  not (_12225_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_12226_, _11231_, _12225_);
  and (_12227_, _11231_, _09735_);
  or (_12228_, _12227_, _12226_);
  and (_12230_, _12228_, _11229_);
  and (_12231_, _11227_, word_in[14]);
  or (_12232_, _12231_, _11236_);
  or (_12233_, _12232_, _12230_);
  or (_12234_, _11242_, _09871_);
  and (_12235_, _12234_, _11241_);
  and (_12236_, _12235_, _12233_);
  or (_14662_, _12236_, _12224_);
  or (_12237_, _07808_, _07803_);
  or (_12238_, _07794_, _07723_);
  nand (_12239_, _12238_, _12237_);
  or (_12240_, _12238_, _12237_);
  nand (_12241_, _12240_, _12239_);
  nand (_12242_, _12241_, _07814_);
  nand (_12243_, _07810_, _07802_);
  nand (_12244_, _12243_, _12242_);
  nand (_12245_, _12244_, _07024_);
  and (_12246_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_12247_, _12246_, _09090_);
  or (_12248_, _09090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_12249_, _12248_, _12247_);
  nand (_12250_, _12249_, _07027_);
  and (_12251_, _11879_, _06845_);
  not (_12252_, _12251_);
  nor (_12253_, _11876_, _06834_);
  and (_12254_, _11876_, _06834_);
  or (_12255_, _12254_, _12253_);
  nor (_12256_, _12255_, _06549_);
  nor (_12257_, _08245_, _06914_);
  nor (_12258_, _12257_, _06586_);
  and (_12259_, _12257_, _06586_);
  nor (_12260_, _12259_, _12258_);
  nor (_12261_, _12260_, _06918_);
  nor (_12262_, _08001_, _06810_);
  and (_12263_, _06926_, _06778_);
  nor (_12264_, _12263_, _12262_);
  and (_12265_, _06951_, _06957_);
  and (_12266_, _06949_, _06924_);
  nor (_12267_, _12266_, _12265_);
  and (_12268_, _12267_, _12264_);
  and (_12269_, _12268_, _07023_);
  and (_12270_, _12269_, _07020_);
  not (_12271_, _12270_);
  nor (_12272_, _12271_, _12261_);
  and (_12273_, _12272_, _07016_);
  not (_12274_, _12273_);
  nor (_12275_, _12274_, _12256_);
  and (_12276_, _12275_, _12252_);
  and (_12277_, _12276_, _12250_);
  nand (_12278_, _12277_, _12245_);
  nand (_12279_, _12278_, _08045_);
  nor (_12280_, _06539_, _06592_);
  nor (_12281_, _12280_, _06969_);
  nor (_12282_, _12281_, _08043_);
  nor (_12283_, _11948_, _06592_);
  or (_12284_, _12283_, _07699_);
  nor (_12285_, _12284_, _12282_);
  nand (_12286_, _12285_, _12279_);
  and (_12287_, _06951_, _06847_);
  and (_12288_, _06958_, _07003_);
  nor (_12289_, _09262_, _09104_);
  not (_12290_, _12289_);
  and (_12291_, _12290_, _09256_);
  nor (_12292_, _12291_, _06847_);
  and (_12293_, _12291_, _06847_);
  nor (_12294_, _12293_, _12292_);
  and (_12295_, _12294_, _06997_);
  nor (_12296_, _06778_, _06597_);
  nor (_12297_, _12296_, _06919_);
  nor (_12298_, _12297_, _06992_);
  or (_12299_, _12298_, _12295_);
  or (_12300_, _12299_, _12288_);
  and (_12301_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_12302_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_12303_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_12304_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _12303_);
  nor (_12305_, _12304_, _12302_);
  nand (_12306_, _12305_, _09275_);
  or (_12307_, _12305_, _09275_);
  and (_12308_, _12307_, _06548_);
  and (_12309_, _12308_, _12306_);
  and (_12310_, _09550_, _07027_);
  or (_12311_, _12310_, _12309_);
  or (_12312_, _12311_, _12301_);
  or (_12313_, _12312_, _12300_);
  or (_12314_, _12313_, _12287_);
  or (_12315_, _12314_, _07700_);
  and (_12316_, _12315_, _12286_);
  and (_09804_, _12316_, _06989_);
  and (_12317_, _11240_, word_in[31]);
  nor (_12318_, _11231_, _08663_);
  and (_12319_, _11231_, _08953_);
  or (_12320_, _12319_, _12318_);
  and (_12321_, _12320_, _11229_);
  and (_12322_, _11227_, word_in[15]);
  or (_12323_, _12322_, _11236_);
  or (_12324_, _12323_, _12321_);
  or (_12325_, _11242_, _08942_);
  and (_12326_, _12325_, _11241_);
  and (_12327_, _12326_, _12324_);
  or (_14663_, _12327_, _12317_);
  or (_12328_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand (_12329_, _07493_, _10755_);
  and (_12330_, _12329_, _06989_);
  and (_09812_, _12330_, _12328_);
  and (_12331_, _08939_, _08711_);
  and (_12332_, _08944_, _09447_);
  not (_12333_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_12334_, _09627_, _08950_);
  nor (_12335_, _12334_, _12333_);
  and (_12336_, _12334_, _09636_);
  or (_12337_, _12336_, _12335_);
  or (_12338_, _12337_, _12332_);
  not (_12339_, _12332_);
  or (_12340_, _12339_, word_in[8]);
  and (_12341_, _12340_, _12338_);
  or (_12342_, _12341_, _12331_);
  not (_12343_, _08879_);
  and (_12344_, _10150_, _12343_);
  and (_12345_, _12344_, _08740_);
  not (_12346_, _12345_);
  not (_12347_, _12331_);
  or (_12348_, _12347_, _09648_);
  and (_12349_, _12348_, _12346_);
  and (_12350_, _12349_, _12342_);
  and (_12351_, _12345_, _10171_);
  or (_09864_, _12351_, _12350_);
  not (_12352_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_12353_, _12334_, _12352_);
  and (_12354_, _12334_, word_in[1]);
  or (_12355_, _12354_, _12353_);
  and (_12356_, _12355_, _12339_);
  and (_12357_, _12332_, word_in[9]);
  or (_12358_, _12357_, _12356_);
  and (_12359_, _12358_, _12347_);
  and (_12360_, _12331_, _09801_);
  or (_12361_, _12360_, _12359_);
  and (_12362_, _12361_, _12346_);
  and (_12363_, _12345_, _09656_);
  or (_09867_, _12363_, _12362_);
  or (_12364_, _12347_, _09816_);
  not (_12365_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_12366_, _12334_, _12365_);
  and (_12367_, _12334_, _09674_);
  or (_12368_, _12367_, _12366_);
  or (_12369_, _12368_, _12332_);
  or (_12370_, _12339_, word_in[10]);
  and (_12371_, _12370_, _12369_);
  or (_12372_, _12371_, _12331_);
  and (_12374_, _12372_, _12364_);
  or (_12375_, _12374_, _12345_);
  or (_12376_, _12346_, _09685_);
  and (_09869_, _12376_, _12375_);
  or (_12377_, _12347_, _09829_);
  not (_12378_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_12379_, _12334_, _12378_);
  and (_12380_, _12334_, _09690_);
  or (_12381_, _12380_, _12379_);
  or (_12382_, _12381_, _12332_);
  or (_12383_, _12339_, word_in[11]);
  and (_12384_, _12383_, _12382_);
  or (_12385_, _12384_, _12331_);
  and (_12386_, _12385_, _12377_);
  or (_12388_, _12386_, _12345_);
  or (_12389_, _12346_, _09701_);
  and (_09874_, _12389_, _12388_);
  not (_12390_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_12391_, _12334_, _12390_);
  and (_12392_, _12334_, word_in[4]);
  or (_12393_, _12392_, _12391_);
  and (_12394_, _12393_, _12339_);
  and (_12395_, _12332_, word_in[12]);
  or (_12396_, _12395_, _12394_);
  or (_12397_, _12396_, _12331_);
  nor (_12398_, _12347_, _09842_);
  nor (_12399_, _12398_, _12345_);
  and (_12400_, _12399_, _12397_);
  and (_12401_, _12345_, _09703_);
  or (_09877_, _12401_, _12400_);
  or (_12402_, _12347_, _09855_);
  not (_12403_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_12404_, _12334_, _12403_);
  and (_12406_, _12334_, _09722_);
  or (_12407_, _12406_, _12404_);
  or (_12408_, _12407_, _12332_);
  or (_12409_, _12339_, word_in[13]);
  and (_12410_, _12409_, _12408_);
  or (_12411_, _12410_, _12331_);
  and (_12412_, _12411_, _12402_);
  or (_12413_, _12412_, _12345_);
  or (_12415_, _12346_, _09718_);
  and (_09880_, _12415_, _12413_);
  or (_12416_, _12347_, _09871_);
  not (_12417_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_12418_, _12334_, _12417_);
  and (_12419_, _12334_, _09735_);
  or (_12420_, _12419_, _12418_);
  or (_12421_, _12420_, _12332_);
  or (_12422_, _12339_, word_in[14]);
  and (_12424_, _12422_, _12421_);
  or (_12425_, _12424_, _12331_);
  and (_12426_, _12425_, _12416_);
  or (_12427_, _12426_, _12345_);
  or (_12428_, _12346_, _09745_);
  and (_14664_, _12428_, _12427_);
  nor (_12429_, _12334_, _08803_);
  and (_12430_, _12334_, word_in[7]);
  or (_12431_, _12430_, _12429_);
  and (_12432_, _12431_, _12339_);
  and (_12433_, _12332_, word_in[15]);
  or (_12434_, _12433_, _12432_);
  and (_12435_, _12434_, _12347_);
  and (_12436_, _12331_, _08942_);
  or (_12437_, _12436_, _12435_);
  and (_12438_, _12437_, _12346_);
  and (_12439_, _12345_, _10256_);
  or (_09885_, _12439_, _12438_);
  nor (_09919_, _11648_, rst);
  nor (_09922_, _11785_, rst);
  nor (_09929_, _11717_, rst);
  nor (_09936_, _12090_, rst);
  and (_12442_, _09768_, _08797_);
  not (_12443_, _12442_);
  or (_12444_, _12443_, word_in[8]);
  and (_12446_, _08939_, _08713_);
  not (_12447_, _12446_);
  not (_12448_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_12449_, _09772_, _08950_);
  nor (_12450_, _12449_, _12448_);
  and (_12451_, _12449_, _09636_);
  or (_12452_, _12451_, _12450_);
  or (_12453_, _12452_, _12442_);
  and (_12454_, _12453_, _12447_);
  and (_12455_, _12454_, _12444_);
  and (_12456_, _12344_, _08711_);
  and (_12457_, _12446_, _09648_);
  or (_12458_, _12457_, _12456_);
  or (_12459_, _12458_, _12455_);
  not (_12460_, _12456_);
  or (_12461_, _12460_, word_in[24]);
  and (_14665_, _12461_, _12459_);
  or (_12462_, _12443_, word_in[9]);
  not (_12463_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_12464_, _12449_, _12463_);
  and (_12465_, _12449_, _09660_);
  or (_12466_, _12465_, _12464_);
  or (_12467_, _12466_, _12442_);
  and (_12468_, _12467_, _12447_);
  and (_12469_, _12468_, _12462_);
  and (_12470_, _12446_, _09801_);
  or (_12471_, _12470_, _12456_);
  or (_12472_, _12471_, _12469_);
  or (_12473_, _12460_, word_in[25]);
  and (_09956_, _12473_, _12472_);
  not (_12474_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_12476_, _12449_, _12474_);
  and (_12477_, _12449_, _09674_);
  nor (_12479_, _12477_, _12476_);
  nor (_12480_, _12479_, _12442_);
  and (_12481_, _12442_, word_in[10]);
  or (_12482_, _12481_, _12480_);
  and (_12483_, _12482_, _12447_);
  and (_12484_, _12446_, _09816_);
  or (_12485_, _12484_, _12456_);
  or (_12486_, _12485_, _12483_);
  or (_12487_, _12460_, word_in[26]);
  and (_09961_, _12487_, _12486_);
  not (_12488_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_12489_, _12449_, _12488_);
  and (_12490_, _12449_, _09690_);
  nor (_12491_, _12490_, _12489_);
  nor (_12492_, _12491_, _12442_);
  and (_12493_, _12442_, word_in[11]);
  or (_12494_, _12493_, _12492_);
  and (_12495_, _12494_, _12447_);
  and (_12496_, _12446_, _09829_);
  or (_12497_, _12496_, _12456_);
  or (_12498_, _12497_, _12495_);
  or (_12499_, _12460_, word_in[27]);
  and (_09963_, _12499_, _12498_);
  or (_12500_, _12443_, word_in[12]);
  not (_12501_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_12502_, _12449_, _12501_);
  and (_12503_, _12449_, _09707_);
  or (_12504_, _12503_, _12502_);
  or (_12505_, _12504_, _12442_);
  and (_12506_, _12505_, _12447_);
  and (_12507_, _12506_, _12500_);
  and (_12508_, _12446_, _09842_);
  or (_12509_, _12508_, _12456_);
  or (_12510_, _12509_, _12507_);
  or (_12511_, _12460_, word_in[28]);
  and (_09967_, _12511_, _12510_);
  or (_12512_, _12443_, word_in[13]);
  not (_12513_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_12514_, _12449_, _12513_);
  and (_12515_, _12449_, _09722_);
  or (_12516_, _12515_, _12514_);
  or (_12517_, _12516_, _12442_);
  and (_12518_, _12517_, _12447_);
  and (_12519_, _12518_, _12512_);
  and (_12520_, _12446_, _09855_);
  or (_12521_, _12520_, _12456_);
  or (_12522_, _12521_, _12519_);
  or (_12523_, _12460_, word_in[29]);
  and (_09971_, _12523_, _12522_);
  not (_12524_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_12525_, _12449_, _12524_);
  and (_12526_, _12449_, _09735_);
  nor (_12527_, _12526_, _12525_);
  nor (_12528_, _12527_, _12442_);
  and (_12529_, _12442_, word_in[14]);
  or (_12530_, _12529_, _12528_);
  and (_12531_, _12530_, _12447_);
  and (_12532_, _12446_, _09871_);
  or (_12533_, _12532_, _12456_);
  or (_12534_, _12533_, _12531_);
  or (_12535_, _12460_, word_in[30]);
  and (_09973_, _12535_, _12534_);
  and (_09976_, t2_i, _06989_);
  or (_12536_, _12443_, word_in[15]);
  nor (_12537_, _12449_, _08669_);
  and (_12538_, _12449_, _08953_);
  or (_12539_, _12538_, _12537_);
  or (_12540_, _12539_, _12442_);
  and (_12541_, _12540_, _12447_);
  and (_12542_, _12541_, _12536_);
  and (_12543_, _12446_, _08942_);
  or (_12544_, _12543_, _12456_);
  or (_12545_, _12544_, _12542_);
  or (_12546_, _12460_, word_in[31]);
  and (_09978_, _12546_, _12545_);
  nor (_09999_, _12113_, rst);
  or (_12547_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  not (_12549_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nand (_12550_, _07493_, _12549_);
  and (_12551_, _12550_, _06989_);
  and (_10020_, _12551_, _12547_);
  and (_12552_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_12553_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  or (_12554_, _12553_, _12552_);
  and (_10025_, _12554_, _06989_);
  or (_12555_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not (_12556_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_12557_, _07493_, _12556_);
  and (_12558_, _12557_, _06989_);
  and (_10029_, _12558_, _12555_);
  and (_12559_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_12560_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or (_12561_, _12560_, _12559_);
  and (_10033_, _12561_, _06989_);
  or (_12562_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  nand (_12563_, _07493_, _10739_);
  and (_12564_, _12563_, _06989_);
  and (_10036_, _12564_, _12562_);
  and (_12566_, _12344_, _08713_);
  and (_12567_, _08939_, _08731_);
  not (_12568_, _12567_);
  or (_12569_, _12568_, _09648_);
  and (_12570_, _09897_, _08797_);
  not (_12571_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_12572_, _09902_, _08932_);
  nor (_12573_, _12572_, _12571_);
  and (_12574_, _12572_, _09636_);
  or (_12575_, _12574_, _12573_);
  or (_12576_, _12575_, _12570_);
  not (_12577_, _12570_);
  or (_12578_, _12577_, word_in[8]);
  and (_12579_, _12578_, _12576_);
  or (_12580_, _12579_, _12567_);
  and (_12581_, _12580_, _12569_);
  or (_12582_, _12581_, _12566_);
  not (_12583_, _12566_);
  or (_12584_, _12583_, word_in[24]);
  and (_10042_, _12584_, _12582_);
  or (_12585_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  nand (_12586_, _07493_, _10723_);
  and (_12587_, _12586_, _06989_);
  and (_10045_, _12587_, _12585_);
  or (_12588_, _12568_, _09801_);
  not (_12589_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_12590_, _12572_, _12589_);
  and (_12591_, _12572_, _09660_);
  or (_12592_, _12591_, _12590_);
  or (_12593_, _12592_, _12570_);
  or (_12594_, _12577_, word_in[9]);
  and (_12595_, _12594_, _12593_);
  or (_12596_, _12595_, _12567_);
  and (_12597_, _12596_, _12588_);
  or (_12598_, _12597_, _12566_);
  or (_12599_, _12583_, word_in[25]);
  and (_10047_, _12599_, _12598_);
  or (_12600_, _12568_, _09816_);
  not (_12601_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_12602_, _12572_, _12601_);
  and (_12603_, _12572_, _09674_);
  or (_12604_, _12603_, _12602_);
  or (_12605_, _12604_, _12570_);
  or (_12606_, _12577_, word_in[10]);
  and (_12607_, _12606_, _12605_);
  or (_12608_, _12607_, _12567_);
  and (_12609_, _12608_, _12600_);
  or (_12610_, _12609_, _12566_);
  or (_12611_, _12583_, word_in[26]);
  and (_10049_, _12611_, _12610_);
  or (_12612_, _12568_, _09829_);
  not (_12613_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_12614_, _12572_, _12613_);
  and (_12615_, _12572_, _09690_);
  or (_12616_, _12615_, _12614_);
  or (_12617_, _12616_, _12570_);
  or (_12618_, _12577_, word_in[11]);
  and (_12619_, _12618_, _12617_);
  or (_12620_, _12619_, _12567_);
  and (_12621_, _12620_, _12612_);
  and (_12622_, _12621_, _12583_);
  and (_12623_, _12566_, word_in[27]);
  or (_10051_, _12623_, _12622_);
  or (_12624_, _12568_, _09842_);
  not (_12625_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_12626_, _12572_, _12625_);
  and (_12627_, _12572_, _09707_);
  or (_12628_, _12627_, _12626_);
  or (_12629_, _12628_, _12570_);
  or (_12630_, _12577_, word_in[12]);
  and (_12631_, _12630_, _12629_);
  or (_12632_, _12631_, _12567_);
  and (_12633_, _12632_, _12624_);
  or (_12634_, _12633_, _12566_);
  or (_12635_, _12583_, word_in[28]);
  and (_10053_, _12635_, _12634_);
  or (_12636_, _12568_, _09855_);
  not (_12637_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_12638_, _12572_, _12637_);
  and (_12639_, _12572_, _09722_);
  or (_12640_, _12639_, _12638_);
  or (_12641_, _12640_, _12570_);
  or (_12642_, _12577_, word_in[13]);
  and (_12643_, _12642_, _12641_);
  or (_12644_, _12643_, _12567_);
  and (_12645_, _12644_, _12636_);
  and (_12646_, _12645_, _12583_);
  and (_12647_, _12566_, word_in[29]);
  or (_10055_, _12647_, _12646_);
  nor (_10056_, _11769_, rst);
  or (_12648_, _12568_, _09871_);
  not (_12649_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_12650_, _12572_, _12649_);
  and (_12651_, _12572_, _09735_);
  or (_12652_, _12651_, _12650_);
  or (_12653_, _12652_, _12570_);
  or (_12654_, _12577_, word_in[14]);
  and (_12656_, _12654_, _12653_);
  or (_12657_, _12656_, _12567_);
  and (_12658_, _12657_, _12648_);
  or (_12659_, _12658_, _12566_);
  or (_12660_, _12583_, word_in[30]);
  and (_10058_, _12660_, _12659_);
  nor (_12661_, _12572_, _08798_);
  and (_12662_, _12572_, _08953_);
  or (_12663_, _12662_, _12661_);
  and (_12664_, _12663_, _12577_);
  and (_12665_, _12570_, word_in[15]);
  or (_12666_, _12665_, _12664_);
  or (_12667_, _12666_, _12567_);
  or (_12668_, _12568_, _08942_);
  and (_12669_, _12668_, _12667_);
  and (_12670_, _12669_, _12583_);
  and (_12671_, _12566_, word_in[31]);
  or (_10062_, _12671_, _12670_);
  and (_12673_, _11045_, _08586_);
  nor (_12674_, _12673_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_12675_, _12674_, _11276_);
  nor (_12676_, _12675_, _11964_);
  and (_12677_, _11986_, _08268_);
  or (_12678_, _12136_, _12018_);
  not (_12679_, _12137_);
  and (_12680_, _12171_, _12679_);
  and (_12681_, _12680_, _12678_);
  and (_12682_, _12176_, _11671_);
  and (_12683_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_12684_, _12013_, _11988_);
  or (_12685_, _12684_, _12683_);
  or (_12686_, _12685_, _12682_);
  or (_12687_, _12686_, _12681_);
  or (_12688_, _12687_, _12677_);
  and (_12689_, _12688_, _11964_);
  or (_12690_, _12689_, _12676_);
  and (_10074_, _12690_, _06989_);
  not (_12691_, _11964_);
  and (_12692_, _12691_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_12694_, _11986_, _08123_);
  or (_12695_, _12117_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_12696_, _12118_);
  and (_12697_, _12171_, _12696_);
  and (_12698_, _12697_, _12695_);
  and (_12699_, _12114_, _11974_);
  and (_12700_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_12701_, _12176_, _11786_);
  or (_12702_, _12701_, _12700_);
  or (_12703_, _12702_, _12699_);
  or (_12704_, _12703_, _12698_);
  or (_12705_, _12704_, _12694_);
  and (_12706_, _12705_, _11964_);
  or (_12707_, _12706_, _12692_);
  and (_10079_, _12707_, _06989_);
  and (_12708_, _11275_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_12709_, _12708_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_12710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_12711_, _12710_, _12709_);
  and (_12712_, _12711_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_12713_, _12712_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_12714_, _12713_, _11273_);
  nor (_12715_, _12714_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_12716_, _12714_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_12717_, _12716_, _12715_);
  or (_12718_, _12717_, _11964_);
  and (_12719_, _12718_, _06989_);
  nand (_12720_, _11976_, _11981_);
  nor (_12721_, _12720_, _11969_);
  nor (_12722_, _12721_, _11983_);
  and (_12723_, _11992_, _08479_);
  and (_12724_, _07490_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_12725_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12726_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_12727_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_12728_, _12727_, _12726_);
  and (_12729_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_12730_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_12731_, _12730_, _12729_);
  and (_12732_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_12733_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_12734_, _12733_, _12732_);
  and (_12735_, _12734_, _12731_);
  and (_12736_, _12735_, _12728_);
  nor (_12737_, _12736_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12738_, _12737_, _12725_);
  nor (_12739_, _12738_, _07490_);
  nor (_12740_, _12739_, _12724_);
  and (_12741_, _12740_, _11994_);
  nor (_12742_, _12741_, _12723_);
  nor (_12743_, _12742_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_12744_, _12742_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand (_12745_, _12163_, _12159_);
  nor (_12746_, _12745_, _12744_);
  nor (_12747_, _12746_, _12743_);
  or (_12748_, _12747_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_12749_, _12748_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_12750_, _12749_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_12751_, _12750_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand (_12752_, _12751_, _12742_);
  not (_12753_, _12742_);
  and (_12754_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_12755_, _12754_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_12756_, _12755_, _12747_);
  nand (_12757_, _12756_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand (_12758_, _12757_, _12753_);
  and (_12759_, _12758_, _12752_);
  or (_12760_, _12759_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_12761_, _12759_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_12762_, _12761_, _12760_);
  and (_12763_, _12762_, _12722_);
  and (_12764_, _11863_, _11560_);
  and (_12765_, _12764_, _06980_);
  nor (_12766_, _11936_, _11325_);
  not (_12767_, _12766_);
  or (_12768_, _12767_, _11383_);
  nor (_12769_, _12768_, _11932_);
  nor (_12770_, _11342_, _11413_);
  nor (_12771_, _12770_, _12769_);
  nor (_12772_, _12771_, _11943_);
  and (_12773_, _11370_, _11368_);
  and (_12774_, _11957_, _12773_);
  or (_12775_, _12774_, _12772_);
  or (_12776_, _12775_, _12765_);
  and (_12777_, _11948_, _11372_);
  and (_12778_, _11371_, _11368_);
  and (_12779_, _12778_, _11873_);
  or (_12780_, _12779_, _12777_);
  or (_12781_, _12780_, _12776_);
  not (_12782_, _11969_);
  and (_12783_, _11984_, _12782_);
  and (_12784_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_12785_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_12786_, _12785_, _12784_);
  and (_12787_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_12788_, _12787_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_12789_, _12788_, _12755_);
  and (_12790_, _12789_, _12786_);
  and (_12791_, _12790_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_12792_, _12791_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_12793_, _12791_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_12794_, _12793_, _12792_);
  and (_12795_, _12794_, _12783_);
  and (_12796_, _11413_, _08346_);
  not (_12797_, _11968_);
  nor (_12798_, _12797_, _08307_);
  and (_12799_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_12800_, _11974_, _11718_);
  or (_12801_, _12800_, _12799_);
  or (_12802_, _12801_, _12798_);
  or (_12803_, _12802_, _12796_);
  or (_12804_, _12803_, _12795_);
  or (_12805_, _12804_, _12781_);
  or (_12806_, _12805_, _12763_);
  and (_10092_, _12806_, _12719_);
  and (_12807_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_12808_, _11053_, _11011_);
  nor (_12809_, _12808_, _11054_);
  or (_12811_, _12809_, _08477_);
  or (_12812_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_12813_, _12812_, _10964_);
  and (_12814_, _12813_, _12811_);
  or (_10098_, _12814_, _12807_);
  and (_12815_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_12816_, _11043_, _11026_);
  nor (_12817_, _12816_, _11044_);
  or (_12818_, _12817_, _08477_);
  or (_12819_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_12820_, _12819_, _10964_);
  and (_12821_, _12820_, _12818_);
  or (_10101_, _12821_, _12815_);
  and (_12822_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _06989_);
  nor (_12823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_12824_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and (_12825_, _12824_, _12823_);
  nor (_12826_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor (_12827_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_12828_, _12827_, _12826_);
  and (_12829_, _12828_, _12825_);
  and (_12830_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _06989_);
  and (_12831_, _12830_, _12829_);
  or (_10112_, _12831_, _12822_);
  nor (_10114_, _11670_, rst);
  not (_12833_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_12834_, _08951_, _12833_);
  and (_12835_, _08951_, word_in[0]);
  nor (_12836_, _12835_, _12834_);
  nor (_12837_, _12836_, _08946_);
  and (_12838_, _08946_, word_in[8]);
  or (_12839_, _12838_, _12837_);
  and (_12840_, _12839_, _08941_);
  and (_12841_, _09648_, _08940_);
  or (_12842_, _12841_, _12840_);
  and (_12843_, _12842_, _08964_);
  and (_12844_, _08936_, word_in[24]);
  or (_10126_, _12844_, _12843_);
  and (_12845_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _08578_);
  and (_12846_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_12847_, _12846_, _12845_);
  and (_10129_, _12847_, _06989_);
  not (_12848_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_12849_, _08951_, _12848_);
  and (_12850_, _08951_, word_in[1]);
  nor (_12852_, _12850_, _12849_);
  nor (_12853_, _12852_, _08946_);
  and (_12854_, _08946_, word_in[9]);
  or (_12855_, _12854_, _12853_);
  and (_12856_, _12855_, _08941_);
  and (_12857_, _09801_, _08940_);
  or (_12858_, _12857_, _12856_);
  and (_12859_, _12858_, _08964_);
  and (_12860_, _08936_, word_in[25]);
  or (_10131_, _12860_, _12859_);
  not (_12861_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_12862_, _08951_, _12861_);
  and (_12864_, _08951_, word_in[2]);
  or (_12865_, _12864_, _12862_);
  or (_12866_, _12865_, _08946_);
  or (_12867_, _08957_, word_in[10]);
  and (_12868_, _12867_, _12866_);
  or (_12869_, _12868_, _08940_);
  or (_12870_, _09816_, _08941_);
  and (_12871_, _12870_, _08964_);
  and (_12872_, _12871_, _12869_);
  and (_12873_, _09685_, _08936_);
  or (_10133_, _12873_, _12872_);
  not (_12874_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_12875_, _08951_, _12874_);
  and (_12876_, _08951_, word_in[3]);
  or (_12877_, _12876_, _12875_);
  or (_12878_, _12877_, _08946_);
  or (_12879_, _08957_, word_in[11]);
  and (_12880_, _12879_, _12878_);
  or (_12881_, _12880_, _08940_);
  or (_12882_, _09829_, _08941_);
  and (_12883_, _12882_, _08964_);
  and (_12884_, _12883_, _12881_);
  and (_12885_, _09701_, _08936_);
  or (_10135_, _12885_, _12884_);
  and (_12886_, _09842_, _08940_);
  not (_12887_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_12888_, _08951_, _12887_);
  and (_12889_, _08951_, word_in[4]);
  nor (_12890_, _12889_, _12888_);
  nor (_12891_, _12890_, _08946_);
  and (_12892_, _08946_, word_in[12]);
  or (_12893_, _12892_, _12891_);
  and (_12894_, _12893_, _08941_);
  or (_12895_, _12894_, _12886_);
  and (_12896_, _12895_, _08964_);
  and (_12897_, _08936_, word_in[28]);
  or (_10137_, _12897_, _12896_);
  and (_12898_, _09855_, _08940_);
  not (_12899_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_12900_, _08951_, _12899_);
  and (_12901_, _08951_, word_in[5]);
  nor (_12902_, _12901_, _12900_);
  nor (_12903_, _12902_, _08946_);
  and (_12904_, _08946_, word_in[13]);
  or (_12905_, _12904_, _12903_);
  and (_12906_, _12905_, _08941_);
  or (_12907_, _12906_, _12898_);
  and (_12908_, _12907_, _08964_);
  and (_12909_, _08936_, word_in[29]);
  or (_10139_, _12909_, _12908_);
  and (_12910_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_12911_, _07493_, _11085_);
  or (_12912_, _12911_, _12910_);
  and (_10142_, _12912_, _06989_);
  and (_12913_, _08951_, word_in[6]);
  not (_12914_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_12915_, _08951_, _12914_);
  nor (_12916_, _12915_, _12913_);
  nor (_12917_, _12916_, _08946_);
  and (_12918_, _08946_, word_in[14]);
  or (_12919_, _12918_, _12917_);
  or (_12920_, _12919_, _08940_);
  or (_12921_, _09871_, _08941_);
  and (_12922_, _12921_, _08964_);
  and (_12923_, _12922_, _12920_);
  and (_12924_, _08936_, word_in[30]);
  or (_10144_, _12924_, _12923_);
  or (_12925_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or (_12926_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_12927_, _12926_, _06989_);
  and (_10400_, _12927_, _12925_);
  and (_12928_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_12929_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_12930_, _12929_, _12928_);
  and (_10446_, _12930_, _06989_);
  or (_12931_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or (_12932_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and (_12933_, _12932_, _06989_);
  and (_10449_, _12933_, _12931_);
  or (_12934_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_12935_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_12936_, _12935_, _06989_);
  and (_10452_, _12936_, _12934_);
  and (_12937_, _08996_, _06981_);
  not (_12938_, _12937_);
  nor (_12939_, _12938_, _11529_);
  not (_12940_, _08996_);
  and (_12942_, _09606_, _12940_);
  nor (_12943_, _12942_, _06982_);
  or (_12944_, _09606_, _06982_);
  nand (_12945_, _12944_, _12943_);
  and (_12946_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or (_12947_, _12946_, _12939_);
  and (_10877_, _12947_, _06989_);
  and (_12948_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_12949_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_12950_, _08139_, _12949_);
  or (_12951_, _12950_, _12948_);
  and (_10989_, _12951_, _06989_);
  and (_12952_, _07134_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_12953_, _11529_, _09489_);
  or (_12954_, _12953_, _12952_);
  nand (_12955_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor (_12956_, _12955_, _07131_);
  or (_12957_, _12956_, _12954_);
  and (_11005_, _12957_, _06989_);
  not (_12958_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_12959_, _07123_, _12958_);
  and (_12960_, _09599_, _07123_);
  or (_12961_, _12960_, _06982_);
  or (_12962_, _12961_, _12959_);
  or (_12963_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_12964_, _12963_, _06989_);
  and (_11031_, _12964_, _12962_);
  and (_12966_, _08708_, word_in[0]);
  nand (_12967_, _08580_, _10685_);
  or (_12968_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_12969_, _12968_, _12967_);
  and (_12970_, _12969_, _08623_);
  nand (_12971_, _08580_, _11230_);
  or (_12972_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_12973_, _12972_, _12971_);
  and (_12974_, _12973_, _08606_);
  nand (_12975_, _08580_, _12448_);
  or (_12977_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_12978_, _12977_, _12975_);
  and (_12979_, _12978_, _08592_);
  or (_12980_, _12979_, _12974_);
  or (_12981_, _12980_, _12970_);
  nand (_12982_, _08580_, _12833_);
  or (_12983_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_12984_, _12983_, _12982_);
  and (_12985_, _12984_, _08613_);
  or (_12986_, _12985_, _08632_);
  or (_12987_, _12986_, _12981_);
  nand (_12988_, _08580_, _09771_);
  or (_12989_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_12990_, _12989_, _12988_);
  and (_12991_, _12990_, _08623_);
  nand (_12992_, _08580_, _10016_);
  or (_12993_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_12994_, _12993_, _12992_);
  and (_12995_, _12994_, _08606_);
  nand (_12996_, _08580_, _10263_);
  or (_12997_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_12998_, _12997_, _12996_);
  and (_12999_, _12998_, _08592_);
  or (_13000_, _12999_, _12995_);
  or (_13001_, _13000_, _12991_);
  nand (_13002_, _08580_, _10474_);
  or (_13003_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_13004_, _13003_, _13002_);
  and (_13005_, _13004_, _08613_);
  or (_13006_, _13005_, _08599_);
  or (_13007_, _13006_, _13001_);
  and (_13008_, _13007_, _12987_);
  and (_13009_, _13008_, _08656_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _13009_, _12966_);
  and (_13010_, _08708_, word_in[1]);
  nand (_13011_, _08580_, _11247_);
  or (_13012_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_13013_, _13012_, _13011_);
  and (_13014_, _13013_, _08606_);
  nand (_13015_, _08580_, _12463_);
  or (_13016_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_13017_, _13016_, _13015_);
  and (_13018_, _13017_, _08592_);
  nand (_13019_, _08580_, _10699_);
  or (_13020_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_13021_, _13020_, _13019_);
  and (_13022_, _13021_, _08623_);
  or (_13023_, _13022_, _13018_);
  or (_13024_, _13023_, _13014_);
  nand (_13025_, _08580_, _12848_);
  or (_13026_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_13027_, _13026_, _13025_);
  and (_13028_, _13027_, _08613_);
  or (_13029_, _13028_, _08632_);
  or (_13030_, _13029_, _13024_);
  nand (_13031_, _08580_, _10037_);
  or (_13032_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_13033_, _13032_, _13031_);
  and (_13034_, _13033_, _08606_);
  nand (_13035_, _08580_, _09792_);
  or (_13036_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_13037_, _13036_, _13035_);
  and (_13038_, _13037_, _08623_);
  nand (_13039_, _08580_, _10276_);
  or (_13040_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_13041_, _13040_, _13039_);
  and (_13042_, _13041_, _08592_);
  or (_13043_, _13042_, _13038_);
  or (_13044_, _13043_, _13034_);
  nand (_13045_, _08580_, _10489_);
  or (_13046_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_13047_, _13046_, _13045_);
  and (_13048_, _13047_, _08613_);
  or (_13049_, _13048_, _08599_);
  or (_13050_, _13049_, _13044_);
  and (_13051_, _13050_, _13030_);
  and (_13052_, _13051_, _08656_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _13052_, _13010_);
  and (_13053_, _08708_, word_in[2]);
  nand (_13054_, _08580_, _10710_);
  or (_13055_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_13056_, _13055_, _13054_);
  and (_13057_, _13056_, _08623_);
  nand (_13058_, _08580_, _11260_);
  or (_13059_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_13060_, _13059_, _13058_);
  and (_13061_, _13060_, _08606_);
  nand (_13062_, _08580_, _12474_);
  or (_13063_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_13064_, _13063_, _13062_);
  and (_13065_, _13064_, _08592_);
  or (_13066_, _13065_, _13061_);
  or (_13067_, _13066_, _13057_);
  nand (_13068_, _08580_, _12861_);
  or (_13069_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_13070_, _13069_, _13068_);
  and (_13071_, _13070_, _08613_);
  or (_13072_, _13071_, _08632_);
  or (_13073_, _13072_, _13067_);
  nand (_13074_, _08580_, _09807_);
  or (_13075_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_13076_, _13075_, _13074_);
  and (_13077_, _13076_, _08623_);
  nand (_13078_, _08580_, _10057_);
  or (_13079_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_13080_, _13079_, _13078_);
  and (_13081_, _13080_, _08606_);
  nand (_13082_, _08580_, _10290_);
  or (_13083_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_13084_, _13083_, _13082_);
  and (_13085_, _13084_, _08592_);
  or (_13086_, _13085_, _13081_);
  or (_13087_, _13086_, _13077_);
  nand (_13088_, _08580_, _10501_);
  or (_13089_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_13090_, _13089_, _13088_);
  and (_13091_, _13090_, _08613_);
  or (_13092_, _13091_, _08599_);
  or (_13094_, _13092_, _13087_);
  and (_13095_, _13094_, _13073_);
  and (_13096_, _13095_, _08656_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _13096_, _13053_);
  and (_13097_, _08708_, word_in[3]);
  nand (_13098_, _08580_, _10727_);
  or (_13099_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_13100_, _13099_, _13098_);
  and (_13101_, _13100_, _08623_);
  nand (_13102_, _08580_, _12185_);
  or (_13104_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_13105_, _13104_, _13102_);
  and (_13106_, _13105_, _08606_);
  nand (_13107_, _08580_, _12488_);
  or (_13108_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_13109_, _13108_, _13107_);
  and (_13110_, _13109_, _08592_);
  or (_13111_, _13110_, _13106_);
  or (_13112_, _13111_, _13101_);
  nand (_13113_, _08580_, _12874_);
  or (_13115_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_13116_, _13115_, _13113_);
  and (_13117_, _13116_, _08613_);
  or (_13119_, _13117_, _08632_);
  or (_13120_, _13119_, _13112_);
  nand (_13121_, _08580_, _09821_);
  or (_13122_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_13123_, _13122_, _13121_);
  and (_13124_, _13123_, _08623_);
  nand (_13125_, _08580_, _10072_);
  or (_13126_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_13127_, _13126_, _13125_);
  and (_13128_, _13127_, _08606_);
  nand (_13129_, _08580_, _10301_);
  or (_13130_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_13131_, _13130_, _13129_);
  and (_13132_, _13131_, _08592_);
  or (_13133_, _13132_, _13128_);
  or (_13134_, _13133_, _13124_);
  nand (_13135_, _08580_, _10512_);
  or (_13136_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_13138_, _13136_, _13135_);
  and (_13139_, _13138_, _08613_);
  or (_13140_, _13139_, _08599_);
  or (_13141_, _13140_, _13134_);
  and (_13142_, _13141_, _13120_);
  and (_13143_, _13142_, _08656_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _13143_, _13097_);
  and (_13144_, _08708_, word_in[4]);
  nand (_13145_, _08580_, _10743_);
  or (_13147_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_13148_, _13147_, _13145_);
  and (_13149_, _13148_, _08623_);
  nand (_13150_, _08580_, _12196_);
  or (_13151_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_13152_, _13151_, _13150_);
  and (_13153_, _13152_, _08606_);
  nand (_13155_, _08580_, _12501_);
  or (_13156_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_13158_, _13156_, _13155_);
  and (_13159_, _13158_, _08592_);
  or (_13160_, _13159_, _13153_);
  or (_13161_, _13160_, _13149_);
  nand (_13162_, _08580_, _12887_);
  or (_13163_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_13164_, _13163_, _13162_);
  and (_13165_, _13164_, _08613_);
  or (_13166_, _13165_, _08632_);
  or (_13167_, _13166_, _13161_);
  nand (_13168_, _08580_, _09834_);
  or (_13169_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_13170_, _13169_, _13168_);
  and (_13171_, _13170_, _08623_);
  nand (_13172_, _08580_, _10086_);
  or (_13173_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_13174_, _13173_, _13172_);
  and (_13175_, _13174_, _08606_);
  nand (_13176_, _08580_, _10315_);
  or (_13177_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_13178_, _13177_, _13176_);
  and (_13179_, _13178_, _08592_);
  or (_13180_, _13179_, _13175_);
  or (_13181_, _13180_, _13171_);
  nand (_13182_, _08580_, _10525_);
  or (_13183_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_13184_, _13183_, _13182_);
  and (_13185_, _13184_, _08613_);
  or (_13186_, _13185_, _08599_);
  or (_13187_, _13186_, _13181_);
  and (_13188_, _13187_, _13167_);
  and (_13189_, _13188_, _08656_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _13189_, _13144_);
  and (_13190_, _08708_, word_in[5]);
  nand (_13191_, _08580_, _10759_);
  or (_13192_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_13193_, _13192_, _13191_);
  and (_13194_, _13193_, _08623_);
  nand (_13195_, _08580_, _12209_);
  or (_13196_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_13197_, _13196_, _13195_);
  and (_13198_, _13197_, _08606_);
  nand (_13199_, _08580_, _12513_);
  or (_13200_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_13201_, _13200_, _13199_);
  and (_13202_, _13201_, _08592_);
  or (_13203_, _13202_, _13198_);
  or (_13204_, _13203_, _13194_);
  nand (_13205_, _08580_, _12899_);
  or (_13206_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_13208_, _13206_, _13205_);
  and (_13209_, _13208_, _08613_);
  or (_13210_, _13209_, _08632_);
  or (_13211_, _13210_, _13204_);
  nand (_13212_, _08580_, _09847_);
  or (_13213_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_13214_, _13213_, _13212_);
  and (_13215_, _13214_, _08623_);
  nand (_13216_, _08580_, _10100_);
  or (_13217_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_13218_, _13217_, _13216_);
  and (_13219_, _13218_, _08606_);
  nand (_13220_, _08580_, _10325_);
  or (_13221_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_13222_, _13221_, _13220_);
  and (_13223_, _13222_, _08592_);
  or (_13224_, _13223_, _13219_);
  or (_13226_, _13224_, _13215_);
  nand (_13227_, _08580_, _10537_);
  or (_13228_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_13229_, _13228_, _13227_);
  and (_13230_, _13229_, _08613_);
  or (_13231_, _13230_, _08599_);
  or (_13232_, _13231_, _13226_);
  and (_13233_, _13232_, _13211_);
  and (_13234_, _13233_, _08656_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _13234_, _13190_);
  and (_13235_, _08708_, word_in[6]);
  nand (_13236_, _08580_, _10771_);
  or (_13237_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_13238_, _13237_, _13236_);
  and (_13239_, _13238_, _08623_);
  nand (_13240_, _08580_, _12225_);
  or (_13241_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_13242_, _13241_, _13240_);
  and (_13243_, _13242_, _08606_);
  nand (_13244_, _08580_, _12524_);
  or (_13245_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_13246_, _13245_, _13244_);
  and (_13247_, _13246_, _08592_);
  or (_13248_, _13247_, _13243_);
  or (_13249_, _13248_, _13239_);
  nand (_13250_, _08580_, _12914_);
  or (_13251_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_13252_, _13251_, _13250_);
  and (_13253_, _13252_, _08613_);
  or (_13254_, _13253_, _08632_);
  or (_13255_, _13254_, _13249_);
  nand (_13256_, _08580_, _09860_);
  or (_13257_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_13258_, _13257_, _13256_);
  and (_13259_, _13258_, _08623_);
  nand (_13260_, _08580_, _10113_);
  or (_13261_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_13262_, _13261_, _13260_);
  and (_13263_, _13262_, _08606_);
  nand (_13264_, _08580_, _10338_);
  or (_13265_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_13266_, _13265_, _13264_);
  and (_13267_, _13266_, _08592_);
  or (_13268_, _13267_, _13263_);
  or (_13269_, _13268_, _13259_);
  nand (_13270_, _08580_, _10548_);
  or (_13271_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_13273_, _13271_, _13270_);
  and (_13274_, _13273_, _08613_);
  or (_13275_, _13274_, _08599_);
  or (_13276_, _13275_, _13269_);
  and (_13277_, _13276_, _13255_);
  and (_13278_, _13277_, _08656_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _13278_, _13235_);
  and (_13279_, _08757_, word_in[8]);
  nand (_13280_, _08580_, _09900_);
  or (_13281_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_13282_, _13281_, _13280_);
  and (_13283_, _13282_, _08759_);
  nand (_13284_, _08580_, _09625_);
  or (_13285_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_13286_, _13285_, _13284_);
  and (_13287_, _13286_, _08758_);
  or (_13288_, _13287_, _13283_);
  and (_13289_, _13288_, _08724_);
  nand (_13290_, _08580_, _11094_);
  or (_13291_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_13292_, _13291_, _13290_);
  and (_13293_, _13292_, _08759_);
  nand (_13294_, _08580_, _10573_);
  or (_13295_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_13296_, _13295_, _13294_);
  and (_13297_, _13296_, _08758_);
  or (_13298_, _13297_, _13293_);
  and (_13299_, _13298_, _08726_);
  nand (_13300_, _08580_, _10368_);
  or (_13301_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_13302_, _13301_, _13300_);
  and (_13303_, _13302_, _08759_);
  nand (_13304_, _08580_, _10158_);
  or (_13305_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_13306_, _13305_, _13304_);
  and (_13307_, _13306_, _08758_);
  or (_13308_, _13307_, _13303_);
  and (_13309_, _13308_, _08784_);
  nand (_13310_, _08580_, _12571_);
  or (_13311_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_13312_, _13311_, _13310_);
  and (_13313_, _13312_, _08759_);
  nand (_13314_, _08580_, _12333_);
  or (_13315_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_13316_, _13315_, _13314_);
  and (_13317_, _13316_, _08758_);
  or (_13318_, _13317_, _13313_);
  and (_13319_, _13318_, _08797_);
  or (_13320_, _13319_, _13309_);
  or (_13321_, _13320_, _13299_);
  nor (_13322_, _13321_, _13289_);
  nor (_13323_, _13322_, _08757_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _13323_, _13279_);
  and (_13324_, _08757_, word_in[9]);
  nand (_13325_, _08580_, _09916_);
  or (_13326_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_13327_, _13326_, _13325_);
  and (_13328_, _13327_, _08759_);
  nand (_13329_, _08580_, _09658_);
  or (_13330_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_13331_, _13330_, _13329_);
  and (_13332_, _13331_, _08758_);
  or (_13333_, _13332_, _13328_);
  and (_13334_, _13333_, _08724_);
  nand (_13335_, _08580_, _11108_);
  or (_13336_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_13337_, _13336_, _13335_);
  and (_13338_, _13337_, _08759_);
  nand (_13339_, _08580_, _10591_);
  or (_13340_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_13341_, _13340_, _13339_);
  and (_13342_, _13341_, _08758_);
  or (_13344_, _13342_, _13338_);
  and (_13345_, _13344_, _08726_);
  nand (_13346_, _08580_, _10382_);
  or (_13347_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_13348_, _13347_, _13346_);
  and (_13349_, _13348_, _08759_);
  nand (_13350_, _08580_, _10175_);
  or (_13351_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_13352_, _13351_, _13350_);
  and (_13353_, _13352_, _08758_);
  or (_13354_, _13353_, _13349_);
  and (_13355_, _13354_, _08784_);
  nand (_13356_, _08580_, _12589_);
  or (_13357_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_13358_, _13357_, _13356_);
  and (_13359_, _13358_, _08759_);
  nand (_13360_, _08580_, _12352_);
  or (_13361_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_13362_, _13361_, _13360_);
  and (_13363_, _13362_, _08758_);
  or (_13364_, _13363_, _13359_);
  and (_13366_, _13364_, _08797_);
  or (_13367_, _13366_, _13355_);
  or (_13368_, _13367_, _13345_);
  nor (_13369_, _13368_, _13334_);
  nor (_13370_, _13369_, _08757_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _13370_, _13324_);
  and (_13371_, _08757_, word_in[10]);
  nand (_13372_, _08580_, _09931_);
  or (_13373_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_13374_, _13373_, _13372_);
  and (_13375_, _13374_, _08759_);
  nand (_13376_, _08580_, _09672_);
  or (_13377_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and (_13378_, _13377_, _13376_);
  and (_13379_, _13378_, _08758_);
  or (_13380_, _13379_, _13375_);
  and (_13381_, _13380_, _08724_);
  nand (_13382_, _08580_, _11120_);
  or (_13383_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_13384_, _13383_, _13382_);
  and (_13385_, _13384_, _08759_);
  nand (_13386_, _08580_, _10603_);
  or (_13387_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_13388_, _13387_, _13386_);
  and (_13389_, _13388_, _08758_);
  or (_13390_, _13389_, _13385_);
  and (_13391_, _13390_, _08726_);
  nand (_13392_, _08580_, _10395_);
  or (_13393_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_13394_, _13393_, _13392_);
  and (_13395_, _13394_, _08759_);
  nand (_13396_, _08580_, _10187_);
  or (_13397_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_13398_, _13397_, _13396_);
  and (_13399_, _13398_, _08758_);
  or (_13400_, _13399_, _13395_);
  and (_13401_, _13400_, _08784_);
  nand (_13402_, _08580_, _12601_);
  or (_13403_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_13404_, _13403_, _13402_);
  and (_13405_, _13404_, _08759_);
  nand (_13406_, _08580_, _12365_);
  or (_13407_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_13408_, _13407_, _13406_);
  and (_13409_, _13408_, _08758_);
  or (_13410_, _13409_, _13405_);
  and (_13411_, _13410_, _08797_);
  or (_13412_, _13411_, _13401_);
  or (_13413_, _13412_, _13391_);
  nor (_13414_, _13413_, _13381_);
  nor (_13416_, _13414_, _08757_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _13416_, _13371_);
  and (_13417_, _08757_, word_in[11]);
  nand (_13418_, _08580_, _09944_);
  or (_13419_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_13420_, _13419_, _13418_);
  and (_13421_, _13420_, _08759_);
  nand (_13422_, _08580_, _09688_);
  or (_13424_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and (_13425_, _13424_, _13422_);
  and (_13426_, _13425_, _08758_);
  or (_13427_, _13426_, _13421_);
  and (_13428_, _13427_, _08724_);
  nand (_13429_, _08580_, _11132_);
  or (_13430_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_13431_, _13430_, _13429_);
  and (_13432_, _13431_, _08759_);
  nand (_13433_, _08580_, _10615_);
  or (_13434_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_13435_, _13434_, _13433_);
  and (_13436_, _13435_, _08758_);
  or (_13437_, _13436_, _13432_);
  and (_13438_, _13437_, _08726_);
  nand (_13439_, _08580_, _10407_);
  or (_13440_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_13441_, _13440_, _13439_);
  and (_13442_, _13441_, _08759_);
  nand (_13443_, _08580_, _10199_);
  or (_13444_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_13445_, _13444_, _13443_);
  and (_13447_, _13445_, _08758_);
  or (_13448_, _13447_, _13442_);
  and (_13449_, _13448_, _08784_);
  nand (_13450_, _08580_, _12613_);
  or (_13451_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_13452_, _13451_, _13450_);
  and (_13453_, _13452_, _08759_);
  nand (_13454_, _08580_, _12378_);
  or (_13455_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_13456_, _13455_, _13454_);
  and (_13457_, _13456_, _08758_);
  or (_13458_, _13457_, _13453_);
  and (_13459_, _13458_, _08797_);
  or (_13460_, _13459_, _13449_);
  or (_13461_, _13460_, _13438_);
  nor (_13462_, _13461_, _13428_);
  nor (_13464_, _13462_, _08757_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _13464_, _13417_);
  and (_13465_, _08757_, word_in[12]);
  nand (_13466_, _08580_, _09957_);
  or (_13467_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_13468_, _13467_, _13466_);
  and (_13469_, _13468_, _08759_);
  nand (_13470_, _08580_, _09705_);
  or (_13471_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_13472_, _13471_, _13470_);
  and (_13473_, _13472_, _08758_);
  or (_13474_, _13473_, _13469_);
  and (_13475_, _13474_, _08724_);
  nand (_13476_, _08580_, _11144_);
  or (_13477_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_13478_, _13477_, _13476_);
  and (_13479_, _13478_, _08759_);
  nand (_13480_, _08580_, _10627_);
  or (_13481_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_13482_, _13481_, _13480_);
  and (_13483_, _13482_, _08758_);
  or (_13484_, _13483_, _13479_);
  and (_13485_, _13484_, _08726_);
  nand (_13486_, _08580_, _10420_);
  or (_13487_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_13488_, _13487_, _13486_);
  and (_13489_, _13488_, _08759_);
  nand (_13490_, _08580_, _10212_);
  or (_13491_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_13492_, _13491_, _13490_);
  and (_13493_, _13492_, _08758_);
  or (_13494_, _13493_, _13489_);
  and (_13495_, _13494_, _08784_);
  nand (_13496_, _08580_, _12625_);
  or (_13497_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_13498_, _13497_, _13496_);
  and (_13499_, _13498_, _08759_);
  nand (_13500_, _08580_, _12390_);
  or (_13501_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_13502_, _13501_, _13500_);
  and (_13503_, _13502_, _08758_);
  or (_13504_, _13503_, _13499_);
  and (_13505_, _13504_, _08797_);
  or (_13506_, _13505_, _13495_);
  or (_13507_, _13506_, _13485_);
  nor (_13508_, _13507_, _13475_);
  nor (_13509_, _13508_, _08757_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _13509_, _13465_);
  and (_13510_, _08757_, word_in[13]);
  nand (_13511_, _08580_, _09974_);
  or (_13512_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_13513_, _13512_, _13511_);
  and (_13514_, _13513_, _08759_);
  nand (_13515_, _08580_, _09720_);
  or (_13516_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_13517_, _13516_, _13515_);
  and (_13518_, _13517_, _08758_);
  or (_13519_, _13518_, _13514_);
  and (_13520_, _13519_, _08724_);
  nand (_13521_, _08580_, _11156_);
  or (_13522_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_13523_, _13522_, _13521_);
  and (_13524_, _13523_, _08759_);
  nand (_13525_, _08580_, _10639_);
  or (_13526_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_13527_, _13526_, _13525_);
  and (_13528_, _13527_, _08758_);
  or (_13529_, _13528_, _13524_);
  and (_13530_, _13529_, _08726_);
  nand (_13531_, _08580_, _10431_);
  or (_13532_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_13533_, _13532_, _13531_);
  and (_13534_, _13533_, _08759_);
  nand (_13535_, _08580_, _10223_);
  or (_13536_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_13537_, _13536_, _13535_);
  and (_13538_, _13537_, _08758_);
  or (_13539_, _13538_, _13534_);
  and (_13540_, _13539_, _08784_);
  nand (_13541_, _08580_, _12637_);
  or (_13542_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_13543_, _13542_, _13541_);
  and (_13544_, _13543_, _08759_);
  nand (_13545_, _08580_, _12403_);
  or (_13546_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_13547_, _13546_, _13545_);
  and (_13548_, _13547_, _08758_);
  or (_13549_, _13548_, _13544_);
  and (_13550_, _13549_, _08797_);
  or (_13551_, _13550_, _13540_);
  or (_13552_, _13551_, _13530_);
  nor (_13553_, _13552_, _13520_);
  nor (_13554_, _13553_, _08757_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _13554_, _13510_);
  and (_13555_, _08757_, word_in[14]);
  nand (_13556_, _08580_, _09988_);
  or (_13557_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_13558_, _13557_, _13556_);
  and (_13559_, _13558_, _08759_);
  nand (_13560_, _08580_, _09732_);
  or (_13561_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_13562_, _13561_, _13560_);
  and (_13563_, _13562_, _08758_);
  or (_13564_, _13563_, _13559_);
  and (_13565_, _13564_, _08724_);
  nand (_13566_, _08580_, _11168_);
  or (_13567_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_13568_, _13567_, _13566_);
  and (_13569_, _13568_, _08759_);
  nand (_13570_, _08580_, _10652_);
  or (_13571_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_13572_, _13571_, _13570_);
  and (_13574_, _13572_, _08758_);
  or (_13575_, _13574_, _13569_);
  and (_13576_, _13575_, _08726_);
  nand (_13577_, _08580_, _10444_);
  or (_13578_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_13579_, _13578_, _13577_);
  and (_13581_, _13579_, _08759_);
  nand (_13582_, _08580_, _10235_);
  or (_13583_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_13584_, _13583_, _13582_);
  and (_13585_, _13584_, _08758_);
  or (_13586_, _13585_, _13581_);
  and (_13587_, _13586_, _08784_);
  nand (_13588_, _08580_, _12649_);
  or (_13589_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_13590_, _13589_, _13588_);
  and (_13591_, _13590_, _08759_);
  nand (_13593_, _08580_, _12417_);
  or (_13594_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_13595_, _13594_, _13593_);
  and (_13596_, _13595_, _08758_);
  or (_13598_, _13596_, _13591_);
  and (_13599_, _13598_, _08797_);
  or (_13600_, _13599_, _13587_);
  or (_13601_, _13600_, _13576_);
  nor (_13602_, _13601_, _13565_);
  nor (_13603_, _13602_, _08757_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _13603_, _13555_);
  and (_13604_, _08850_, word_in[16]);
  and (_13605_, _12998_, _08606_);
  and (_13606_, _12990_, _08613_);
  or (_13607_, _13606_, _13605_);
  and (_13608_, _13004_, _08592_);
  and (_13609_, _12994_, _08623_);
  or (_13610_, _13609_, _13608_);
  or (_13611_, _13610_, _13607_);
  or (_13612_, _13611_, _08821_);
  and (_13613_, _12978_, _08606_);
  and (_13614_, _12969_, _08613_);
  or (_13615_, _13614_, _13613_);
  and (_13616_, _12984_, _08592_);
  and (_13617_, _12973_, _08623_);
  or (_13618_, _13617_, _13616_);
  or (_13619_, _13618_, _13615_);
  or (_13620_, _13619_, _08860_);
  nand (_13621_, _13620_, _13612_);
  nor (_13622_, _13621_, _08850_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _13622_, _13604_);
  and (_13623_, _08850_, word_in[17]);
  and (_13624_, _13037_, _08613_);
  and (_13625_, _13047_, _08592_);
  or (_13626_, _13625_, _13624_);
  and (_13627_, _13041_, _08606_);
  and (_13628_, _13033_, _08623_);
  or (_13629_, _13628_, _13627_);
  or (_13630_, _13629_, _13626_);
  or (_13631_, _13630_, _08821_);
  and (_13632_, _13017_, _08606_);
  and (_13633_, _13021_, _08613_);
  or (_13634_, _13633_, _13632_);
  and (_13635_, _13027_, _08592_);
  and (_13636_, _13013_, _08623_);
  or (_13637_, _13636_, _13635_);
  or (_13638_, _13637_, _13634_);
  or (_13639_, _13638_, _08860_);
  nand (_13640_, _13639_, _13631_);
  nor (_13641_, _13640_, _08850_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _13641_, _13623_);
  and (_13642_, _08850_, word_in[18]);
  and (_13643_, _13084_, _08606_);
  and (_13644_, _13076_, _08613_);
  or (_13645_, _13644_, _13643_);
  and (_13646_, _13090_, _08592_);
  and (_13647_, _13080_, _08623_);
  or (_13648_, _13647_, _13646_);
  or (_13650_, _13648_, _13645_);
  or (_13652_, _13650_, _08821_);
  and (_13653_, _13064_, _08606_);
  and (_13654_, _13056_, _08613_);
  or (_13655_, _13654_, _13653_);
  and (_13656_, _13070_, _08592_);
  and (_13657_, _13060_, _08623_);
  or (_13658_, _13657_, _13656_);
  or (_13659_, _13658_, _13655_);
  or (_13660_, _13659_, _08860_);
  nand (_13661_, _13660_, _13652_);
  nor (_13662_, _13661_, _08850_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _13662_, _13642_);
  and (_13663_, _08850_, word_in[19]);
  and (_13664_, _13131_, _08606_);
  and (_13665_, _13123_, _08613_);
  or (_13666_, _13665_, _13664_);
  and (_13667_, _13138_, _08592_);
  and (_13668_, _13127_, _08623_);
  or (_13669_, _13668_, _13667_);
  or (_13670_, _13669_, _13666_);
  or (_13671_, _13670_, _08821_);
  and (_13672_, _13100_, _08613_);
  and (_13673_, _13116_, _08592_);
  or (_13674_, _13673_, _13672_);
  and (_13675_, _13109_, _08606_);
  and (_13676_, _13105_, _08623_);
  or (_13677_, _13676_, _13675_);
  or (_13678_, _13677_, _13674_);
  or (_13679_, _13678_, _08860_);
  nand (_13680_, _13679_, _13671_);
  nor (_13681_, _13680_, _08850_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _13681_, _13663_);
  and (_13682_, _08850_, word_in[20]);
  and (_13683_, _13178_, _08606_);
  and (_13684_, _13170_, _08613_);
  or (_13685_, _13684_, _13683_);
  and (_13686_, _13184_, _08592_);
  and (_13687_, _13174_, _08623_);
  or (_13688_, _13687_, _13686_);
  or (_13689_, _13688_, _13685_);
  or (_13690_, _13689_, _08821_);
  and (_13691_, _13158_, _08606_);
  and (_13692_, _13148_, _08613_);
  or (_13693_, _13692_, _13691_);
  and (_13694_, _13164_, _08592_);
  and (_13695_, _13152_, _08623_);
  or (_13696_, _13695_, _13694_);
  or (_13697_, _13696_, _13693_);
  or (_13698_, _13697_, _08860_);
  nand (_13699_, _13698_, _13690_);
  nor (_13700_, _13699_, _08850_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _13700_, _13682_);
  and (_13701_, _08850_, word_in[21]);
  and (_13702_, _13222_, _08606_);
  and (_13703_, _13214_, _08613_);
  or (_13704_, _13703_, _13702_);
  and (_13705_, _13229_, _08592_);
  and (_13706_, _13218_, _08623_);
  or (_13708_, _13706_, _13705_);
  or (_13709_, _13708_, _13704_);
  or (_13711_, _13709_, _08821_);
  and (_13712_, _13193_, _08613_);
  and (_13713_, _13208_, _08592_);
  or (_13714_, _13713_, _13712_);
  and (_13715_, _13201_, _08606_);
  and (_13716_, _13197_, _08623_);
  or (_13717_, _13716_, _13715_);
  or (_13718_, _13717_, _13714_);
  or (_13719_, _13718_, _08860_);
  nand (_13720_, _13719_, _13711_);
  nor (_13721_, _13720_, _08850_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _13721_, _13701_);
  and (_13722_, _08850_, word_in[22]);
  and (_13723_, _13258_, _08613_);
  and (_13724_, _13273_, _08592_);
  or (_13725_, _13724_, _13723_);
  and (_13726_, _13266_, _08606_);
  and (_13727_, _13262_, _08623_);
  or (_13728_, _13727_, _13726_);
  or (_13730_, _13728_, _13725_);
  or (_13731_, _13730_, _08821_);
  and (_13732_, _13246_, _08606_);
  and (_13733_, _13238_, _08613_);
  or (_13734_, _13733_, _13732_);
  and (_13736_, _13252_, _08592_);
  and (_13737_, _13242_, _08623_);
  or (_13738_, _13737_, _13736_);
  or (_13739_, _13738_, _13734_);
  or (_13740_, _13739_, _08860_);
  nand (_13741_, _13740_, _13731_);
  nor (_13742_, _13741_, _08850_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _13742_, _13722_);
  and (_13743_, _08908_, word_in[24]);
  and (_13744_, _13286_, _08759_);
  and (_13746_, _13282_, _08758_);
  or (_13747_, _13746_, _13744_);
  and (_13748_, _13747_, _08885_);
  and (_13749_, _13296_, _08759_);
  and (_13750_, _13292_, _08758_);
  or (_13751_, _13750_, _13749_);
  and (_13752_, _13751_, _08880_);
  and (_13753_, _13306_, _08759_);
  and (_13754_, _13302_, _08758_);
  or (_13755_, _13754_, _13753_);
  and (_13756_, _13755_, _08917_);
  and (_13757_, _13316_, _08759_);
  and (_13759_, _13312_, _08758_);
  or (_13760_, _13759_, _13757_);
  and (_13761_, _13760_, _08925_);
  or (_13762_, _13761_, _13756_);
  or (_13763_, _13762_, _13752_);
  nor (_13764_, _13763_, _13748_);
  nor (_13765_, _13764_, _08908_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _13765_, _13743_);
  and (_13767_, _08908_, word_in[25]);
  and (_13769_, _13331_, _08759_);
  and (_13770_, _13327_, _08758_);
  or (_13771_, _13770_, _13769_);
  and (_13772_, _13771_, _08885_);
  and (_13773_, _13341_, _08759_);
  and (_13774_, _13337_, _08758_);
  or (_13775_, _13774_, _13773_);
  and (_13776_, _13775_, _08880_);
  and (_13777_, _13352_, _08759_);
  and (_13778_, _13348_, _08758_);
  or (_13779_, _13778_, _13777_);
  and (_13780_, _13779_, _08917_);
  and (_13781_, _13362_, _08759_);
  and (_13782_, _13358_, _08758_);
  or (_13783_, _13782_, _13781_);
  and (_13784_, _13783_, _08925_);
  or (_13785_, _13784_, _13780_);
  or (_13786_, _13785_, _13776_);
  nor (_13787_, _13786_, _13772_);
  nor (_13789_, _13787_, _08908_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _13789_, _13767_);
  and (_13790_, _08908_, word_in[26]);
  and (_13791_, _13378_, _08759_);
  and (_13792_, _13374_, _08758_);
  or (_13793_, _13792_, _13791_);
  and (_13794_, _13793_, _08885_);
  and (_13795_, _13388_, _08759_);
  and (_13796_, _13384_, _08758_);
  or (_13797_, _13796_, _13795_);
  and (_13799_, _13797_, _08880_);
  and (_13800_, _13398_, _08759_);
  and (_13801_, _13394_, _08758_);
  or (_13803_, _13801_, _13800_);
  and (_13804_, _13803_, _08917_);
  and (_13805_, _13408_, _08759_);
  and (_13806_, _13404_, _08758_);
  or (_13807_, _13806_, _13805_);
  and (_13808_, _13807_, _08925_);
  or (_13810_, _13808_, _13804_);
  or (_13811_, _13810_, _13799_);
  nor (_13813_, _13811_, _13794_);
  nor (_13814_, _13813_, _08908_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _13814_, _13790_);
  and (_13816_, _08908_, word_in[27]);
  and (_13818_, _13435_, _08759_);
  and (_13819_, _13431_, _08758_);
  or (_13820_, _13819_, _13818_);
  and (_13821_, _13820_, _08880_);
  and (_13823_, _13425_, _08759_);
  and (_13824_, _13420_, _08758_);
  or (_13825_, _13824_, _13823_);
  and (_13826_, _13825_, _08885_);
  and (_13827_, _13445_, _08759_);
  and (_13828_, _13441_, _08758_);
  or (_13829_, _13828_, _13827_);
  and (_13830_, _13829_, _08917_);
  and (_13831_, _13456_, _08759_);
  and (_13832_, _13452_, _08758_);
  or (_13833_, _13832_, _13831_);
  and (_13834_, _13833_, _08925_);
  or (_13835_, _13834_, _13830_);
  or (_13836_, _13835_, _13826_);
  nor (_13837_, _13836_, _13821_);
  nor (_13838_, _13837_, _08908_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _13838_, _13816_);
  and (_13839_, _08908_, word_in[28]);
  and (_13840_, _13472_, _08759_);
  and (_13841_, _13468_, _08758_);
  or (_13842_, _13841_, _13840_);
  and (_13843_, _13842_, _08885_);
  and (_13844_, _13482_, _08759_);
  and (_13845_, _13478_, _08758_);
  or (_13846_, _13845_, _13844_);
  and (_13847_, _13846_, _08880_);
  and (_13848_, _13492_, _08759_);
  and (_13849_, _13488_, _08758_);
  or (_13850_, _13849_, _13848_);
  and (_13851_, _13850_, _08917_);
  and (_13852_, _13502_, _08759_);
  and (_13853_, _13498_, _08758_);
  or (_13854_, _13853_, _13852_);
  and (_13855_, _13854_, _08925_);
  or (_13856_, _13855_, _13851_);
  or (_13857_, _13856_, _13847_);
  nor (_13858_, _13857_, _13843_);
  nor (_13859_, _13858_, _08908_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _13859_, _13839_);
  and (_13860_, _08908_, word_in[29]);
  and (_13861_, _13517_, _08759_);
  and (_13862_, _13513_, _08758_);
  or (_13863_, _13862_, _13861_);
  and (_13864_, _13863_, _08885_);
  and (_13865_, _13527_, _08759_);
  and (_13866_, _13523_, _08758_);
  or (_13867_, _13866_, _13865_);
  and (_13868_, _13867_, _08880_);
  and (_13869_, _13537_, _08759_);
  and (_13870_, _13533_, _08758_);
  or (_13871_, _13870_, _13869_);
  and (_13873_, _13871_, _08917_);
  and (_13874_, _13547_, _08759_);
  and (_13875_, _13543_, _08758_);
  or (_13876_, _13875_, _13874_);
  and (_13877_, _13876_, _08925_);
  or (_13878_, _13877_, _13873_);
  or (_13879_, _13878_, _13868_);
  nor (_13880_, _13879_, _13864_);
  nor (_13881_, _13880_, _08908_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _13881_, _13860_);
  and (_13882_, _08908_, word_in[30]);
  and (_13883_, _13572_, _08759_);
  and (_13885_, _13568_, _08758_);
  or (_13886_, _13885_, _13883_);
  and (_13887_, _13886_, _08880_);
  and (_13888_, _13562_, _08759_);
  and (_13889_, _13558_, _08758_);
  or (_13890_, _13889_, _13888_);
  and (_13891_, _13890_, _08885_);
  and (_13892_, _13584_, _08759_);
  and (_13893_, _13579_, _08758_);
  or (_13894_, _13893_, _13892_);
  and (_13895_, _13894_, _08917_);
  and (_13896_, _13595_, _08759_);
  and (_13897_, _13590_, _08758_);
  or (_13898_, _13897_, _13896_);
  and (_13899_, _13898_, _08925_);
  or (_13900_, _13899_, _13895_);
  or (_13901_, _13900_, _13891_);
  nor (_13902_, _13901_, _13887_);
  nor (_13903_, _13902_, _08908_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _13903_, _13882_);
  and (_11200_, _08085_, _06989_);
  and (_11222_, _09182_, _06989_);
  and (_11228_, _07978_, _06989_);
  and (_11259_, _08231_, _06989_);
  and (_11268_, _08317_, _06989_);
  nor (_13904_, _07027_, _07662_);
  and (_13905_, _07027_, _07662_);
  or (_13906_, _13905_, _13904_);
  and (_11307_, _13906_, _06989_);
  and (_11318_, _07691_, _06989_);
  and (_11323_, _07684_, _06989_);
  and (_11357_, _08197_, _06989_);
  and (_11362_, _08302_, _06989_);
  and (_11384_, _08380_, _06989_);
  and (_11434_, _09280_, _06989_);
  or (_13909_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or (_13911_, _09516_, _09418_);
  and (_11465_, _13911_, _13909_);
  and (_11487_, _09349_, _06989_);
  or (_13912_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or (_13913_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_13915_, _13913_, _06989_);
  and (_11544_, _13915_, _13912_);
  and (_13916_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_13917_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_13918_, _13917_, _13916_);
  and (_11592_, _13918_, _06989_);
  and (_11633_, _08402_, _06989_);
  and (_13920_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_13921_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_13922_, _08139_, _13921_);
  or (_13923_, _13922_, _13920_);
  and (_11677_, _13923_, _06989_);
  and (_13924_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_13925_, _07493_, _11081_);
  or (_13926_, _13925_, _13924_);
  and (_11826_, _13926_, _06989_);
  or (_13927_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or (_13928_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and (_13929_, _13928_, _06989_);
  and (_11831_, _13929_, _13927_);
  and (_13930_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_13931_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or (_13932_, _13931_, _13930_);
  and (_11847_, _13932_, _06989_);
  or (_13933_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or (_13934_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_13935_, _13934_, _06989_);
  and (_11854_, _13935_, _13933_);
  nand (_13936_, _11529_, _10146_);
  or (_13937_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_13938_, _13937_, _06989_);
  and (_11893_, _13938_, _13936_);
  and (_11967_, _07816_, _06989_);
  and (_11997_, _08396_, _06989_);
  and (_12000_, _09179_, _06989_);
  nor (_13939_, _07262_, _07118_);
  and (_13940_, _07262_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or (_13941_, _13940_, _13939_);
  and (_12039_, _13941_, _06989_);
  and (_13942_, _09393_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_13943_, _13942_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_13944_, _13943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_13945_, _13944_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_13946_, _13945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or (_13947_, _13946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_13948_, _13946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_13949_, _13948_, _13947_);
  and (_13950_, _07453_, _07085_);
  and (_13951_, _06985_, _07089_);
  and (_13952_, _13951_, _13950_);
  nor (_13953_, _13952_, rst);
  and (_12052_, _13953_, _13949_);
  and (_13955_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_13956_, _07493_, _12556_);
  or (_13957_, _13956_, _13955_);
  and (_12057_, _13957_, _06989_);
  and (_13958_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_13959_, _13958_, _09392_);
  nor (_13960_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_13961_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_13962_, _13961_, _13960_);
  nor (_13963_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_13964_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor (_13965_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_13966_, _13965_, _13964_);
  and (_13967_, _13966_, _13963_);
  and (_13968_, _13967_, _13962_);
  not (_13969_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_13970_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_13971_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_13972_, _13971_, _13970_);
  and (_13973_, _13972_, _13969_);
  and (_13974_, _13973_, _13968_);
  not (_13975_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_13976_, _13972_, _13975_);
  or (_13977_, _13976_, _13974_);
  and (_13978_, _13977_, _13943_);
  nand (_13979_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_13980_, _13979_, _13942_);
  nor (_13981_, _13980_, _13978_);
  nor (_13982_, _13981_, _13959_);
  and (_13983_, _13968_, _13959_);
  or (_13984_, _13983_, _13982_);
  and (_12060_, _13984_, _13953_);
  and (_13985_, _07090_, _06983_);
  and (_13986_, _13985_, _13950_);
  nand (_13987_, _13974_, _13942_);
  nand (_13988_, _13987_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_13989_, _13988_, _13983_);
  or (_13990_, _13989_, _13986_);
  and (_12075_, _13990_, _06989_);
  not (_13991_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_13992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not (_13993_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_13994_, _07462_, _13993_);
  not (_13995_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_13996_, _13995_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_13997_, _13996_, _13994_);
  nor (_13998_, _13997_, _13992_);
  nand (_13999_, _13998_, _13991_);
  nor (_14000_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor (_14001_, _14000_, _13998_);
  nand (_14002_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_14003_, _14002_, _14001_);
  and (_14004_, _14003_, _06989_);
  and (_12082_, _14004_, _13999_);
  and (_12085_, _14001_, _06989_);
  and (_14005_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  not (_14007_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_14008_, _07493_, _14007_);
  or (_14010_, _14008_, _14005_);
  and (_12104_, _14010_, _06989_);
  and (_14011_, _09072_, _06539_);
  and (_14012_, _14011_, _07454_);
  or (_14013_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_14015_, _14013_, _06989_);
  and (_14016_, _09239_, _06539_);
  nand (_14017_, _14016_, _07040_);
  and (_12115_, _14017_, _14015_);
  and (_14018_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  not (_14020_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_14021_, _07493_, _14020_);
  or (_14023_, _14021_, _14018_);
  and (_12121_, _14023_, _06989_);
  nor (_14025_, _06447_, _06434_);
  and (_14026_, _06477_, _06463_);
  and (_14027_, _14026_, _06500_);
  and (_14028_, _14027_, _14025_);
  and (_14029_, _14028_, _06539_);
  nand (_14030_, _14029_, _06968_);
  and (_14031_, _13950_, _06986_);
  not (_14032_, _14031_);
  or (_14033_, _14029_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_14034_, _14033_, _14032_);
  and (_14035_, _14034_, _14030_);
  nor (_14036_, _14032_, _07040_);
  or (_14037_, _14036_, _14035_);
  and (_12128_, _14037_, _06989_);
  and (_12133_, _08212_, _06989_);
  and (_14038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_14039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_14040_, _07462_, _14039_);
  or (_14041_, _14040_, _13996_);
  nor (_14042_, _14041_, _14038_);
  or (_14043_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_14044_, _14043_, _06989_);
  nor (_12160_, _14044_, _14042_);
  nor (_12170_, _07461_, rst);
  or (_14045_, _09403_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  not (_14046_, rxd_i);
  nand (_14047_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _14046_);
  nand (_14048_, _14047_, _09403_);
  and (_14049_, _14048_, _09393_);
  and (_14050_, _14049_, _14045_);
  or (_14051_, _09414_, _09411_);
  or (_14052_, _14051_, _14050_);
  and (_12208_, _14052_, _09418_);
  and (_14053_, _09763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_14054_, _14053_, _09396_);
  and (_14055_, _09762_, _14054_);
  not (_14056_, _09395_);
  nor (_14057_, _14053_, _14056_);
  or (_14058_, _14057_, _09760_);
  and (_14060_, _14058_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_14061_, _14060_, _14055_);
  and (_12211_, _14061_, _06989_);
  and (_14062_, _09764_, _09397_);
  and (_14063_, _09762_, _14062_);
  nand (_14065_, _14063_, _14046_);
  or (_14066_, _14063_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_14067_, _14066_, _06989_);
  and (_12214_, _14067_, _14065_);
  not (_14068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor (_14069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _09405_);
  not (_14070_, _14069_);
  nor (_14071_, _09392_, _09389_);
  and (_14073_, _14071_, _14070_);
  and (_14074_, _14073_, _14056_);
  nor (_14076_, _14074_, _14068_);
  and (_14077_, _14074_, rxd_i);
  or (_14078_, _14077_, rst);
  or (_12220_, _14078_, _14076_);
  or (_14079_, _09420_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_14080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_14081_, _14080_, _09392_);
  or (_14083_, _14081_, _09395_);
  nand (_14084_, _14083_, _14079_);
  nand (_12229_, _14084_, _09418_);
  nand (_14086_, _07669_, _07027_);
  or (_14088_, _07027_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_14089_, _14088_, _06989_);
  and (_12373_, _14089_, _14086_);
  and (_12387_, _09086_, _06989_);
  and (_14091_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  not (_14092_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_14093_, _07493_, _14092_);
  or (_14094_, _14093_, _14091_);
  and (_12405_, _14094_, _06989_);
  or (_14095_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or (_14096_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_14097_, _14096_, _06989_);
  and (_12414_, _14097_, _14095_);
  and (_14098_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not (_14099_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_14100_, _07493_, _14099_);
  or (_14101_, _14100_, _14098_);
  and (_12423_, _14101_, _06989_);
  and (_14102_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_12440_, _14102_, _09477_);
  and (_14103_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  not (_14104_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_14106_, _07493_, _14104_);
  or (_14107_, _14106_, _14103_);
  and (_12441_, _14107_, _06989_);
  and (_14109_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  not (_14110_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_14112_, _07493_, _14110_);
  or (_14113_, _14112_, _14109_);
  and (_12445_, _14113_, _06989_);
  and (_14114_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_14116_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_14117_, _14116_, _14114_);
  and (_12475_, _14117_, _06989_);
  or (_14119_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_14120_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_14122_, _14120_, _06989_);
  and (_12478_, _14122_, _14119_);
  nor (_14124_, _07486_, _07260_);
  and (_14125_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or (_14126_, _14125_, _14124_);
  and (_12548_, _14126_, _06989_);
  nor (_14128_, _07486_, _07118_);
  and (_14129_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_14130_, _14129_, _14128_);
  and (_12655_, _14130_, _06989_);
  nor (_14131_, _12938_, _10970_);
  and (_14132_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_14133_, _14132_, _14131_);
  and (_12672_, _14133_, _06989_);
  nor (_14134_, _12938_, _07118_);
  and (_14135_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_14136_, _14135_, _14134_);
  and (_12693_, _14136_, _06989_);
  and (_14137_, _07262_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor (_14138_, _07262_, _07040_);
  or (_14140_, _14138_, _14137_);
  and (_12810_, _14140_, _06989_);
  and (_14141_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_12863_, _14141_, _09391_);
  and (_14143_, _07135_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_14144_, _09488_, _09009_);
  or (_14145_, _14144_, _14143_);
  and (_12941_, _14145_, _06989_);
  and (_12965_, _06989_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  not (_14146_, _09010_);
  and (_14147_, _14146_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor (_14148_, _14146_, _07317_);
  or (_14149_, _14148_, _14147_);
  and (_12976_, _14149_, _06989_);
  or (_14150_, _14056_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or (_14151_, _14150_, _09401_);
  and (_14152_, _14151_, _09481_);
  or (_14153_, _14152_, rxd_i);
  and (_14154_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], rxd_i);
  nor (_14155_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  and (_14156_, _14155_, _09395_);
  and (_14157_, _14156_, _09400_);
  nor (_14158_, _14157_, _09426_);
  and (_14159_, _14158_, _14153_);
  or (_14160_, _14159_, _09389_);
  nor (_14161_, _09420_, _09389_);
  or (_14162_, _14161_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_14163_, _14162_, _06989_);
  and (_13093_, _14163_, _14160_);
  and (_14164_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_14165_, _07493_, _12549_);
  or (_14166_, _14165_, _14164_);
  and (_13103_, _14166_, _06989_);
  and (_13114_, _06989_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  and (_13118_, _07643_, _06989_);
  and (_14167_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  not (_14168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_14169_, _07493_, _14168_);
  or (_14170_, _14169_, _14167_);
  and (_13137_, _14170_, _06989_);
  nand (_14171_, _10146_, _07260_);
  or (_14172_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_14173_, _14172_, _06989_);
  and (_13146_, _14173_, _14171_);
  and (_14174_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_14175_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_14176_, _14175_, _14174_);
  and (_13154_, _14176_, _06989_);
  nor (_14177_, _11529_, _09614_);
  and (_14178_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_14179_, _14178_, _06982_);
  or (_14180_, _14179_, _14177_);
  or (_14181_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_14182_, _14181_, _06989_);
  and (_13157_, _14182_, _14180_);
  and (_14183_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not (_14184_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_14185_, _07493_, _14184_);
  or (_14186_, _14185_, _14183_);
  and (_13207_, _14186_, _06989_);
  or (_14187_, _09607_, _06982_);
  or (_14188_, _14187_, _12943_);
  and (_14189_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_14190_, _08994_, _06981_);
  and (_14191_, _14190_, _11821_);
  or (_14192_, _14191_, _14189_);
  and (_13272_, _14192_, _06989_);
  and (_14193_, _07135_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor (_14194_, _09489_, _07040_);
  or (_14195_, _14194_, _14193_);
  and (_13343_, _14195_, _06989_);
  and (_14196_, _06538_, _06513_);
  and (_14197_, _14028_, _14196_);
  nand (_14198_, _14197_, _06968_);
  or (_14199_, _14197_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_14200_, _14199_, _14032_);
  and (_14201_, _14200_, _14198_);
  nor (_14202_, _14032_, _10970_);
  or (_14203_, _14202_, _14201_);
  and (_13365_, _14203_, _06989_);
  not (_14204_, _11799_);
  nor (_14205_, _14204_, _11748_);
  and (_14206_, _11724_, _11688_);
  not (_14207_, _11613_);
  and (_14208_, _11652_, _14207_);
  and (_14209_, _14208_, _14206_);
  and (_14210_, _11857_, _11556_);
  and (_14211_, _14210_, _14209_);
  and (_14212_, _14211_, _14205_);
  and (_14213_, _14212_, _09071_);
  nor (_14214_, _11652_, _11613_);
  and (_14215_, _14206_, _14214_);
  and (_14217_, _11799_, _11748_);
  nor (_14218_, _11857_, _11556_);
  and (_14219_, _14218_, _14217_);
  and (_14220_, _14219_, _14215_);
  and (_14221_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  not (_14222_, _11556_);
  and (_14223_, _11857_, _14222_);
  and (_14224_, _14217_, _14223_);
  and (_14226_, _14224_, _14215_);
  and (_14228_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_14229_, _14228_, _14221_);
  and (_14230_, _14223_, _14205_);
  and (_14231_, _14230_, _14215_);
  and (_14232_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_14233_, _14204_, _11748_);
  and (_14234_, _14233_, _14218_);
  and (_14235_, _14234_, _14215_);
  and (_14236_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_14237_, _14236_, _14232_);
  or (_14238_, _14237_, _14229_);
  and (_14239_, _14224_, _14209_);
  and (_14240_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_14241_, _11799_, _11748_);
  and (_14242_, _14241_, _14223_);
  and (_14243_, _14242_, _14215_);
  and (_14244_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_14245_, _14244_, _14240_);
  not (_14246_, _11688_);
  and (_14247_, _14208_, _14246_);
  and (_14248_, _14247_, _11724_);
  and (_14249_, _14248_, _14224_);
  and (_14250_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  not (_14251_, _11724_);
  and (_14252_, _14247_, _14251_);
  not (_14253_, _11857_);
  and (_14254_, _14241_, _14253_);
  and (_14256_, _14254_, _11556_);
  and (_14257_, _14256_, _14252_);
  and (_14258_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_14259_, _14258_, _14250_);
  or (_14260_, _14259_, _14245_);
  or (_14261_, _14260_, _14238_);
  and (_14262_, _14233_, _14223_);
  and (_14263_, _14262_, _14209_);
  and (_14265_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_14266_, _14242_, _14209_);
  and (_14267_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_14268_, _14267_, _14265_);
  and (_14269_, _14234_, _14209_);
  and (_14270_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_14271_, _14209_, _14230_);
  and (_14272_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_14273_, _14272_, _14270_);
  or (_14274_, _14273_, _14268_);
  and (_14275_, _14208_, _11688_);
  and (_14276_, _14275_, _14251_);
  and (_14277_, _14276_, _14224_);
  and (_14278_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_14279_, _14276_, _14262_);
  and (_14280_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or (_14281_, _14280_, _14278_);
  and (_14282_, _14219_, _14209_);
  and (_14283_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_14284_, _14256_, _14209_);
  and (_14285_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_14286_, _14285_, _14283_);
  or (_14287_, _14286_, _14281_);
  or (_14288_, _14287_, _14274_);
  or (_14289_, _14288_, _14261_);
  and (_14290_, _14217_, _14210_);
  and (_14291_, _14290_, _14251_);
  and (_14292_, _14214_, _14246_);
  and (_14293_, _14292_, _14291_);
  and (_14294_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_14295_, _14233_, _14210_);
  and (_14296_, _14295_, _14209_);
  and (_14297_, _14296_, _11627_);
  or (_14298_, _14297_, _14294_);
  and (_14299_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_14300_, _14241_, _14210_);
  and (_14301_, _14300_, _14209_);
  and (_14302_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_14303_, _14302_, _14299_);
  or (_14304_, _14303_, _14298_);
  and (_14305_, _14252_, _14290_);
  nor (_14306_, _11460_, _11401_);
  nor (_14307_, _11330_, _11299_);
  and (_14308_, _14307_, _11295_);
  nor (_14309_, _14308_, _11473_);
  nor (_14310_, _11912_, _11452_);
  and (_14311_, _14310_, _14309_);
  and (_14312_, _14311_, _14306_);
  and (_14313_, _11908_, _11403_);
  not (_14314_, _14313_);
  and (_14315_, _14314_, _11457_);
  and (_14316_, _11396_, _11364_);
  and (_14317_, _11478_, _11322_);
  nor (_14318_, _14317_, _14316_);
  and (_14319_, _11382_, _11375_);
  and (_14320_, _11462_, _11321_);
  nor (_14321_, _14320_, _14319_);
  and (_14322_, _14321_, _14318_);
  and (_14323_, _14322_, _14315_);
  and (_14324_, _14323_, _14312_);
  and (_14325_, _14324_, _11443_);
  nor (_14326_, _14325_, _11283_);
  or (_14327_, _14326_, p3_in[6]);
  not (_14328_, _14326_);
  or (_14329_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_14330_, _14329_, _14327_);
  and (_14331_, _14330_, _14305_);
  and (_14332_, _14290_, _11724_);
  and (_14333_, _14332_, _14247_);
  or (_14334_, _14326_, p2_in[6]);
  or (_14335_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_14336_, _14335_, _14334_);
  and (_14337_, _14336_, _14333_);
  or (_14338_, _14337_, _14331_);
  and (_14339_, _14290_, _14209_);
  or (_14340_, _14326_, p0_in[6]);
  or (_14341_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_14342_, _14341_, _14340_);
  and (_14343_, _14342_, _14339_);
  and (_14344_, _14291_, _14275_);
  or (_14345_, _14326_, p1_in[6]);
  or (_14346_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_14347_, _14346_, _14345_);
  and (_14348_, _14347_, _14344_);
  or (_14349_, _14348_, _14343_);
  or (_14350_, _14349_, _14338_);
  or (_14351_, _14350_, _14304_);
  and (_14352_, _14332_, _14292_);
  and (_14353_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_14354_, _14214_, _11688_);
  and (_14355_, _14291_, _14354_);
  and (_14356_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_14357_, _14356_, _14353_);
  or (_14358_, _14357_, _14351_);
  or (_14359_, _14358_, _14289_);
  and (_14360_, _14355_, _11951_);
  and (_14361_, _14352_, _07699_);
  and (_14362_, _14241_, _14211_);
  and (_14363_, _14362_, _09071_);
  or (_14364_, _14363_, _14361_);
  nor (_14365_, _14364_, _14360_);
  nor (_14366_, _14365_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_14367_, _14366_);
  and (_14368_, _14352_, _07705_);
  not (_14369_, _06500_);
  nor (_14370_, _14254_, _14369_);
  and (_14371_, _14370_, _11730_);
  nor (_14372_, _14371_, _14368_);
  and (_14373_, _14372_, _11866_);
  and (_14374_, _14373_, _14367_);
  and (_14375_, _14374_, _14359_);
  not (_14376_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  not (_14377_, _14374_);
  nor (_14378_, _14226_, _14220_);
  nor (_14379_, _14235_, _14231_);
  and (_14380_, _14379_, _14378_);
  nor (_14381_, _14243_, _14239_);
  nor (_14382_, _14257_, _14249_);
  and (_14383_, _14382_, _14381_);
  and (_14384_, _14383_, _14380_);
  nor (_14385_, _14266_, _14263_);
  nor (_14386_, _14271_, _14269_);
  and (_14387_, _14386_, _14385_);
  nor (_14388_, _14279_, _14277_);
  nor (_14389_, _14284_, _14282_);
  and (_14390_, _14389_, _14388_);
  and (_14391_, _14390_, _14387_);
  and (_14392_, _14391_, _14384_);
  nor (_14394_, _14355_, _14352_);
  and (_14395_, _14290_, _14208_);
  not (_14396_, _14395_);
  nor (_14397_, _14301_, _14212_);
  nor (_14398_, _14296_, _14293_);
  and (_14399_, _14398_, _14397_);
  and (_14400_, _14399_, _14396_);
  and (_14401_, _14400_, _14394_);
  and (_14402_, _14401_, _14392_);
  nor (_14404_, _14402_, _14377_);
  nor (_14405_, _14404_, _14376_);
  or (_14406_, _14405_, _14375_);
  or (_14407_, _14406_, _14213_);
  nand (_14408_, _14213_, _09145_);
  and (_14409_, _14408_, _06989_);
  and (_13423_, _14409_, _14407_);
  and (_14410_, _07262_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_14411_, _09009_, _07261_);
  or (_14412_, _14411_, _14410_);
  and (_13446_, _14412_, _06989_);
  and (_13463_, _07814_, _06989_);
  and (_14413_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_14414_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_14415_, _14414_, _14413_);
  and (_14416_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_14417_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_14418_, _14417_, _14416_);
  or (_14419_, _14418_, _14415_);
  and (_14420_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_14421_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or (_14422_, _14421_, _14420_);
  and (_14423_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_14424_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_14425_, _14424_, _14423_);
  or (_14426_, _14425_, _14422_);
  or (_14427_, _14426_, _14419_);
  and (_14428_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_14429_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_14430_, _14429_, _14428_);
  and (_14431_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_14432_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_14433_, _14432_, _14431_);
  or (_14434_, _14433_, _14430_);
  and (_14435_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_14436_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_14437_, _14436_, _14435_);
  and (_14438_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_14439_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_14440_, _14439_, _14438_);
  or (_14441_, _14440_, _14437_);
  or (_14442_, _14441_, _14434_);
  or (_14443_, _14442_, _14427_);
  and (_14444_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_14445_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_14446_, _14445_, _14444_);
  and (_14447_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_14448_, _14296_, _11549_);
  or (_14449_, _14448_, _14447_);
  or (_14450_, _14449_, _14446_);
  or (_14451_, _14326_, p2_in[3]);
  or (_14452_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_14453_, _14452_, _14451_);
  and (_14454_, _14453_, _14333_);
  or (_14455_, _14326_, p3_in[3]);
  or (_14457_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_14458_, _14457_, _14455_);
  and (_14459_, _14458_, _14305_);
  or (_14460_, _14459_, _14454_);
  or (_14461_, _14326_, p0_in[3]);
  or (_14462_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_14463_, _14462_, _14461_);
  and (_14464_, _14463_, _14339_);
  or (_14465_, _14326_, p1_in[3]);
  or (_14466_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_14467_, _14466_, _14465_);
  and (_14468_, _14467_, _14344_);
  or (_14469_, _14468_, _14464_);
  or (_14470_, _14469_, _14460_);
  or (_14471_, _14470_, _14450_);
  and (_14472_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_14473_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_14474_, _14473_, _14472_);
  or (_14475_, _14474_, _14471_);
  or (_14476_, _14475_, _14443_);
  not (_14477_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nor (_14478_, _14404_, _14477_);
  or (_14479_, _14478_, _14476_);
  or (_14480_, _14374_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_14481_, _14480_, _14479_);
  or (_14482_, _14481_, _14213_);
  not (_14483_, _14213_);
  or (_14484_, _14483_, _08433_);
  and (_14485_, _14484_, _06989_);
  and (_13573_, _14485_, _14482_);
  not (_14486_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nor (_14487_, _14404_, _14486_);
  nand (_14488_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  nand (_14489_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_14490_, _14489_, _14488_);
  nand (_14491_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand (_14492_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_14493_, _14492_, _14491_);
  and (_14494_, _14493_, _14490_);
  nand (_14495_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand (_14496_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_14497_, _14496_, _14495_);
  nand (_14498_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nand (_14499_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_14500_, _14499_, _14498_);
  and (_14501_, _14500_, _14497_);
  and (_14502_, _14501_, _14494_);
  nand (_14503_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand (_14504_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_14505_, _14504_, _14503_);
  nand (_14506_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand (_14507_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_14508_, _14507_, _14506_);
  and (_14509_, _14508_, _14505_);
  nand (_14510_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nand (_14511_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and (_14512_, _14511_, _14510_);
  nand (_14513_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_14514_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_14515_, _14514_, _14513_);
  and (_14516_, _14515_, _14512_);
  and (_14517_, _14516_, _14509_);
  and (_14518_, _14517_, _14502_);
  nand (_14519_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_14520_, _14296_, _11852_);
  and (_14521_, _14520_, _14519_);
  nand (_14522_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand (_14523_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_14524_, _14523_, _14522_);
  and (_14525_, _14524_, _14521_);
  nor (_14526_, _14326_, p0_in[2]);
  not (_14527_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_14528_, _14326_, _14527_);
  nor (_14529_, _14528_, _14526_);
  nand (_14530_, _14529_, _14339_);
  nor (_14531_, _14326_, p1_in[2]);
  not (_14532_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_14533_, _14326_, _14532_);
  nor (_14534_, _14533_, _14531_);
  nand (_14535_, _14534_, _14344_);
  and (_14536_, _14535_, _14530_);
  nor (_14537_, _14326_, p3_in[2]);
  not (_14538_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_14539_, _14326_, _14538_);
  nor (_14540_, _14539_, _14537_);
  nand (_14541_, _14540_, _14305_);
  or (_14542_, _14326_, p2_in[2]);
  or (_14543_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_14544_, _14543_, _14542_);
  nand (_14545_, _14544_, _14333_);
  and (_14546_, _14545_, _14541_);
  and (_14547_, _14546_, _14536_);
  and (_14548_, _14547_, _14525_);
  nand (_14549_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand (_14550_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_14551_, _14550_, _14549_);
  and (_14552_, _14551_, _14548_);
  nand (_14553_, _14552_, _14518_);
  nand (_14554_, _14553_, _14374_);
  nand (_14555_, _14554_, _14483_);
  or (_14556_, _14555_, _14487_);
  nand (_14557_, _14213_, _09227_);
  and (_14558_, _14557_, _06989_);
  and (_13580_, _14558_, _14556_);
  and (_14559_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_14560_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_14561_, _14560_, _14559_);
  and (_14562_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_14563_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_14564_, _14563_, _14562_);
  or (_14565_, _14564_, _14561_);
  and (_14566_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_14567_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_14568_, _14567_, _14566_);
  and (_14569_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_14570_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_14571_, _14570_, _14569_);
  or (_14573_, _14571_, _14568_);
  or (_14574_, _14573_, _14565_);
  and (_14575_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_14576_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_14577_, _14576_, _14575_);
  and (_14578_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_14579_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_14580_, _14579_, _14578_);
  or (_14581_, _14580_, _14577_);
  and (_14582_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_14584_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_14586_, _14584_, _14582_);
  and (_14587_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_14588_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_14589_, _14588_, _14587_);
  or (_14590_, _14589_, _14586_);
  or (_14591_, _14590_, _14581_);
  or (_14592_, _14591_, _14574_);
  and (_14593_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_14594_, _14296_, _11740_);
  or (_14595_, _14594_, _14593_);
  and (_14596_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_14597_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_14598_, _14597_, _14596_);
  or (_14599_, _14598_, _14595_);
  or (_14600_, _14326_, p0_in[1]);
  or (_14601_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_14602_, _14601_, _14600_);
  and (_14603_, _14602_, _14339_);
  or (_14604_, _14326_, p1_in[1]);
  or (_14605_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_14606_, _14605_, _14604_);
  and (_14608_, _14606_, _14344_);
  or (_14609_, _14608_, _14603_);
  or (_14610_, _14326_, p3_in[1]);
  or (_14611_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_14612_, _14611_, _14610_);
  and (_14613_, _14612_, _14305_);
  or (_14614_, _14326_, p2_in[1]);
  or (_14615_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_14616_, _14615_, _14614_);
  and (_14617_, _14616_, _14333_);
  or (_14618_, _14617_, _14613_);
  or (_14619_, _14618_, _14609_);
  or (_14620_, _14619_, _14599_);
  and (_14621_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_14622_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_14623_, _14622_, _14621_);
  or (_14624_, _14623_, _14620_);
  or (_14625_, _14624_, _14592_);
  not (_14626_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nor (_14627_, _14404_, _14626_);
  or (_14628_, _14627_, _14625_);
  or (_14629_, _14374_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_14630_, _14629_, _14628_);
  or (_14631_, _14630_, _14213_);
  or (_14632_, _14483_, _08030_);
  and (_14633_, _14632_, _06989_);
  and (_13592_, _14633_, _14631_);
  and (_14634_, _07135_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_14635_, _09489_, _07317_);
  or (_14636_, _14635_, _14634_);
  and (_13597_, _14636_, _06989_);
  or (_14637_, _12278_, _09077_);
  or (_14638_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_14639_, _14638_, _06989_);
  and (_13649_, _14639_, _14637_);
  and (_14640_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_14641_, _12278_, _09292_);
  or (_00001_, _14641_, _14640_);
  or (_00002_, _00001_, _09071_);
  or (_00003_, _12314_, _09369_);
  and (_00004_, _00003_, _06989_);
  and (_13651_, _00004_, _00002_);
  and (_00005_, _13951_, _07454_);
  or (_00006_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_00007_, _00006_, _06989_);
  nand (_00008_, _00005_, _11529_);
  and (_13707_, _00008_, _00007_);
  and (_00010_, _13985_, _07454_);
  nand (_00011_, _00010_, _09008_);
  or (_00012_, _00010_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00013_, _00012_, _06989_);
  and (_13710_, _00013_, _00011_);
  or (_00014_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_00015_, _00014_, _06989_);
  nand (_00016_, _00005_, _07317_);
  and (_13729_, _00016_, _00015_);
  or (_00017_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_00019_, _00017_, _06989_);
  nand (_00020_, _00005_, _07260_);
  and (_13735_, _00020_, _00019_);
  nand (_00021_, _00010_, _09598_);
  or (_00022_, _00010_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00023_, _00022_, _06989_);
  and (_13745_, _00023_, _00021_);
  and (_00025_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_13758_, _00025_, _09434_);
  and (_00027_, _07454_, _07045_);
  nand (_00029_, _00027_, _07118_);
  and (_00030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00032_, _00030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00033_, _00032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_00034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_00035_, _00034_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_00036_, t0_i);
  and (_00037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_00038_, _00037_, _00036_);
  or (_00039_, _00038_, _00035_);
  and (_00040_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_00041_, _00040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_00042_, _00041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_00043_, _00042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_00044_, _00043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_00045_, _00044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_00046_, _00045_, _00033_);
  and (_00047_, _00046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_00049_, _00047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_00051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_00052_, _00051_);
  and (_00053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00054_, _00053_, _00033_);
  and (_00056_, _00054_, _00045_);
  nor (_00057_, _00056_, _00052_);
  and (_00058_, _00057_, _00049_);
  not (_00059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor (_00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _00059_);
  and (_00061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _00059_);
  or (_00062_, _00061_, _00060_);
  not (_00063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_00065_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_00066_, _00065_, _00064_);
  and (_00067_, _00066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_00068_, _00067_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_00069_, _00068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00070_, _00069_, _00040_);
  and (_00071_, _00070_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_00072_, _00071_, _00033_);
  and (_00073_, _00072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00074_, _00073_, _00059_);
  nor (_00075_, _00074_, _00063_);
  and (_00076_, _00074_, _00063_);
  or (_00077_, _00076_, _00075_);
  and (_00078_, _00077_, _00062_);
  and (_00079_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_00080_, _00079_, _00033_);
  and (_00081_, _00080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_00082_, _00081_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00083_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00084_, _00080_, _00053_);
  not (_00085_, _00084_);
  and (_00086_, _00085_, _00083_);
  and (_00087_, _00086_, _00082_);
  or (_00088_, _00087_, _00078_);
  or (_00089_, _00088_, _00058_);
  or (_00090_, _00089_, _00027_);
  and (_00091_, _09075_, _06985_);
  not (_00092_, _00091_);
  and (_00093_, _00092_, _00090_);
  and (_00094_, _00093_, _00029_);
  and (_00095_, _00091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_00096_, _00095_, _00094_);
  and (_13766_, _00096_, _06989_);
  not (_00097_, _00027_);
  nor (_00098_, _00097_, _10970_);
  and (_00099_, _00056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_00100_, _00056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_00101_, _00100_, _00051_);
  nor (_00102_, _00101_, _00099_);
  and (_00103_, _00054_, _00071_);
  or (_00104_, _00103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00105_, _00103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_00106_, _00105_);
  and (_00107_, _00106_, _00061_);
  and (_00108_, _00107_, _00104_);
  and (_00109_, _00080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00110_, _00109_, _00053_);
  or (_00112_, _00110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_00114_, _00110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00115_, _00114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00116_, _00115_, _00112_);
  or (_00118_, _00116_, _00108_);
  nor (_00120_, _00118_, _00102_);
  nor (_00122_, _00120_, _00027_);
  or (_00124_, _00122_, _00091_);
  or (_00125_, _00124_, _00098_);
  or (_00126_, _00092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00127_, _00126_, _06989_);
  and (_13768_, _00127_, _00125_);
  and (_00129_, _00071_, _00059_);
  nor (_00131_, _00129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_00132_, _00129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_00133_, _00132_, _00131_);
  and (_00134_, _00133_, _00062_);
  and (_00135_, _00079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_00137_, _00079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_00139_, _00137_, _00083_);
  nor (_00141_, _00139_, _00135_);
  and (_00142_, _00045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_00143_, _00045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_00144_, _00143_, _00142_);
  and (_00145_, _00144_, _00051_);
  or (_00146_, _00145_, _00141_);
  or (_00147_, _00146_, _00134_);
  or (_00149_, _00147_, _00027_);
  and (_00150_, _00027_, _09598_);
  nor (_00151_, _00150_, _00091_);
  and (_00152_, _00151_, _00149_);
  and (_00153_, _00091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_00154_, _00153_, _00152_);
  and (_13788_, _00154_, _06989_);
  nand (_00155_, _00091_, _10970_);
  or (_00156_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00157_, _00045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_00158_, _00157_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_00159_, _00051_, _00070_);
  or (_00161_, _00159_, _00027_);
  and (_00163_, _00161_, _00158_);
  and (_00164_, _00051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00166_, _00165_, _00040_);
  and (_00167_, _00166_, _00067_);
  and (_00168_, _00167_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_00169_, _00168_, _00060_);
  and (_00170_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_00171_, _00170_, _00164_);
  or (_00172_, _00171_, _00163_);
  and (_00173_, _00172_, _00156_);
  or (_00174_, _00173_, _00091_);
  and (_00175_, _00174_, _06989_);
  and (_13798_, _00175_, _00155_);
  and (_00176_, _00052_, _00045_);
  nand (_00177_, _00176_, _00097_);
  and (_00178_, _00177_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not (_00180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_00182_, _00176_, _00180_);
  and (_00183_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_00184_, _00183_, _00182_);
  nor (_00185_, _00184_, _00027_);
  or (_00186_, _00185_, _00178_);
  and (_00187_, _00186_, _00092_);
  nor (_00189_, _00092_, _07118_);
  or (_00190_, _00189_, _00187_);
  and (_13802_, _00190_, _06989_);
  nand (_00191_, _00027_, _11529_);
  and (_00192_, _00071_, _00030_);
  or (_00193_, _00192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_00194_, _00168_, _00032_);
  and (_00195_, _00194_, _00061_);
  and (_00196_, _00195_, _00193_);
  not (_00197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00198_, _00067_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_00199_, _00040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00200_, _00199_, _00198_);
  and (_00201_, _00200_, _00197_);
  nor (_00202_, _00200_, _00197_);
  or (_00203_, _00202_, _00201_);
  and (_00204_, _00203_, _00051_);
  and (_00205_, _00079_, _00030_);
  and (_00206_, _00205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nor (_00207_, _00206_, _00197_);
  and (_00208_, _00206_, _00197_);
  or (_00209_, _00208_, _00207_);
  and (_00210_, _00209_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_00211_, _00210_, _00204_);
  or (_00212_, _00211_, _00196_);
  nor (_00214_, _00212_, _00027_);
  nor (_00215_, _00214_, _00091_);
  and (_00216_, _00215_, _00191_);
  and (_00217_, _00091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_00218_, _00217_, _00216_);
  and (_13809_, _00218_, _06989_);
  nand (_00220_, _00027_, _07260_);
  or (_00221_, _00046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_00223_, _00221_, _00051_);
  nor (_00224_, _00223_, _00047_);
  or (_00225_, _00072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_00226_, _00073_);
  and (_00227_, _00226_, _00061_);
  and (_00229_, _00227_, _00225_);
  or (_00231_, _00109_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00232_, _00231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand (_00233_, _00081_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_00234_, _00233_, _00232_);
  or (_00235_, _00234_, _00229_);
  or (_00236_, _00235_, _00224_);
  nor (_00237_, _00236_, _00027_);
  nor (_00238_, _00237_, _00091_);
  and (_00239_, _00238_, _00220_);
  and (_00240_, _00091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_00241_, _00240_, _00239_);
  and (_13812_, _00241_, _06989_);
  nand (_00242_, _00027_, _07317_);
  nand (_00243_, _00045_, _00030_);
  nor (_00244_, _00243_, _00197_);
  or (_00245_, _00244_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_00246_, _00244_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00247_, _00051_, _00246_);
  and (_00248_, _00247_, _00245_);
  and (_00249_, _00079_, _00032_);
  or (_00251_, _00249_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_00253_, _00080_);
  and (_00255_, _00083_, _00253_);
  and (_00257_, _00255_, _00251_);
  and (_00259_, _00129_, _00032_);
  or (_00260_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_00262_, _00072_);
  or (_00263_, _00262_, _00060_);
  and (_00264_, _00263_, _00062_);
  and (_00265_, _00264_, _00260_);
  or (_00266_, _00265_, _00257_);
  or (_00267_, _00266_, _00248_);
  or (_00268_, _00267_, _00027_);
  and (_00269_, _00268_, _00242_);
  or (_00270_, _00269_, _00091_);
  or (_00271_, _00092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00273_, _00271_, _06989_);
  and (_13815_, _00273_, _00270_);
  or (_00274_, _00132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_00276_, _00192_);
  or (_00277_, _00276_, _00060_);
  and (_00278_, _00277_, _00062_);
  and (_00279_, _00278_, _00274_);
  or (_00280_, _00135_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_00281_, _00205_);
  and (_00282_, _00083_, _00281_);
  and (_00283_, _00282_, _00280_);
  or (_00284_, _00142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00285_, _00051_, _00243_);
  and (_00286_, _00285_, _00284_);
  or (_00287_, _00286_, _00283_);
  or (_00288_, _00287_, _00279_);
  or (_00290_, _00288_, _00027_);
  nand (_00291_, _00027_, _09008_);
  and (_00292_, _00291_, _00290_);
  or (_00293_, _00292_, _00091_);
  or (_00294_, _00092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00295_, _00294_, _06989_);
  and (_13817_, _00295_, _00293_);
  and (_00296_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00297_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or (_00298_, _00297_, _00296_);
  and (_13822_, _00298_, _06989_);
  and (_00299_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00300_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or (_00301_, _00300_, _00299_);
  and (_13872_, _00301_, _06989_);
  nand (_00302_, _00044_, _00097_);
  and (_00303_, _00302_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nand (_00304_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_00305_, _00043_);
  or (_00306_, _00305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_00307_, _00306_, _00304_);
  nor (_00308_, _00307_, _00027_);
  or (_00309_, _00308_, _00303_);
  and (_00311_, _00309_, _00092_);
  nor (_00312_, _00092_, _07317_);
  or (_00313_, _00312_, _00311_);
  and (_13907_, _00313_, _06989_);
  or (_00314_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_00315_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_00316_, _00044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nand (_00317_, _00045_, _00097_);
  and (_00319_, _00317_, _00316_);
  or (_00320_, _00319_, _00315_);
  and (_00322_, _00320_, _00314_);
  or (_00323_, _00322_, _00091_);
  nand (_00324_, _00091_, _07260_);
  and (_00326_, _00324_, _06989_);
  and (_13908_, _00326_, _00323_);
  or (_00328_, _00305_, _00027_);
  and (_00329_, _00328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nand (_00330_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_00331_, _00305_, _00042_);
  and (_00332_, _00331_, _00330_);
  nor (_00333_, _00332_, _00027_);
  or (_00335_, _00333_, _00329_);
  and (_00336_, _00335_, _00092_);
  nor (_00337_, _00092_, _11529_);
  or (_00338_, _00337_, _00336_);
  and (_13910_, _00338_, _06989_);
  or (_00339_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00340_, _00339_, _06989_);
  nand (_00341_, _00005_, _10970_);
  and (_13914_, _00341_, _00340_);
  or (_00342_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00343_, _00342_, _06989_);
  nand (_00344_, _00005_, _07118_);
  and (_13919_, _00344_, _00343_);
  and (_00346_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00347_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  or (_00349_, _00347_, _00346_);
  and (_13954_, _00349_, _06989_);
  or (_00350_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_00351_, _00040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_00352_, _00351_, _00041_);
  and (_00353_, _00071_, _00060_);
  and (_00354_, _00353_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_00355_, _00354_, _00352_);
  or (_00356_, _00355_, _00027_);
  and (_00357_, _00356_, _00350_);
  or (_00358_, _00357_, _00091_);
  nand (_00359_, _00091_, _09598_);
  and (_00360_, _00359_, _06989_);
  and (_14006_, _00360_, _00358_);
  nor (_00361_, _00041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_00362_, _00361_, _00042_);
  and (_00363_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_00364_, _00363_, _00362_);
  nor (_00365_, _00364_, _00027_);
  and (_00366_, _00027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_00367_, _00366_, _00365_);
  and (_00368_, _00367_, _00092_);
  and (_00369_, _00091_, _09009_);
  or (_00370_, _00369_, _00368_);
  and (_14009_, _00370_, _06989_);
  nand (_00371_, _10146_, _07040_);
  or (_00372_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_00373_, _00372_, _06989_);
  and (_14014_, _00373_, _00371_);
  and (_00374_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_00375_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or (_00376_, _00375_, _00374_);
  and (_14019_, _00376_, _06989_);
  nor (_00377_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_14022_, _00377_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_00378_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00379_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or (_00380_, _00379_, _00378_);
  and (_14024_, _00380_, _06989_);
  and (_00381_, _07454_, _07049_);
  not (_00382_, _00381_);
  nor (_00383_, _00382_, _10970_);
  nor (_00384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_00385_, _00384_);
  and (_00386_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00388_, _00386_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not (_00389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_00390_, _00389_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  not (_00391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00392_, _00391_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_00393_, t1_i);
  and (_00394_, _00393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00395_, _00394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or (_00396_, _00395_, _00392_);
  and (_00397_, _00396_, _00390_);
  and (_00398_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_00400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_00401_, _00400_, _00399_);
  and (_00402_, _00401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00403_, _00402_, _00398_);
  and (_00404_, _00403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00405_, _00404_, _00397_);
  and (_00406_, _00405_, _00388_);
  and (_00407_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00408_, _00407_, _00385_);
  not (_00409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _00409_);
  not (_00411_, _00410_);
  and (_00412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_00413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_00414_, _00413_, _00412_);
  and (_00415_, _00414_, _00401_);
  and (_00416_, _00415_, _00398_);
  and (_00417_, _00416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00418_, _00417_, _00397_);
  and (_00419_, _00418_, _00388_);
  and (_00420_, _00419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00421_, _00420_, _00411_);
  or (_00422_, _00421_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00423_, _00412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_00424_, _00421_, _00423_);
  or (_00425_, _00424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_00426_, _00425_, _00422_);
  or (_00427_, _00426_, _00408_);
  or (_00428_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_00429_, _09560_, _07454_);
  nor (_00430_, _00429_, _00381_);
  and (_00431_, _00430_, _00428_);
  and (_00432_, _00431_, _00427_);
  and (_00433_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_00434_, _00433_, _00432_);
  or (_00435_, _00434_, _00383_);
  and (_14059_, _00435_, _06989_);
  nor (_00436_, _00382_, _07118_);
  not (_00437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00438_, _00402_, _00397_);
  and (_00439_, _00423_, _00438_);
  and (_00440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00441_, _00440_, _00398_);
  and (_00443_, _00441_, _00410_);
  and (_00444_, _00443_, _00439_);
  and (_00446_, _00403_, _00397_);
  and (_00447_, _00440_, _00446_);
  and (_00448_, _00447_, _00384_);
  nor (_00449_, _00448_, _00444_);
  or (_00450_, _00449_, _00437_);
  nor (_00451_, _00450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_00452_, _00450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_00454_, _00452_, _00451_);
  and (_00455_, _00454_, _00430_);
  and (_00456_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_00458_, _00456_, _00455_);
  or (_00459_, _00458_, _00436_);
  and (_14064_, _00459_, _06989_);
  nor (_00460_, _00382_, _07317_);
  and (_00461_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_00462_, _00418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_00463_, _00418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00464_, _00463_, _00462_);
  and (_00466_, _00464_, _00410_);
  not (_00467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00468_, _00384_, _00467_);
  nor (_00469_, _00446_, _00385_);
  or (_00470_, _00469_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_00471_, _00470_, _00468_);
  and (_00472_, _00471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand (_00473_, _00405_, _00384_);
  nor (_00474_, _00473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_00475_, _00474_, _00472_);
  or (_00476_, _00475_, _00466_);
  and (_00477_, _00476_, _00430_);
  or (_00478_, _00477_, _00461_);
  or (_00479_, _00478_, _00460_);
  and (_14072_, _00479_, _06989_);
  nor (_00480_, _00382_, _07260_);
  nand (_00481_, _00449_, _00437_);
  and (_00482_, _00481_, _00450_);
  and (_00483_, _00482_, _00430_);
  and (_00484_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_00485_, _00484_, _00483_);
  or (_00486_, _00485_, _00480_);
  and (_14075_, _00486_, _06989_);
  not (_00487_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_00488_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and (_00489_, _00488_, _00487_);
  and (_00490_, _00489_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor (_00491_, _00488_, _00487_);
  or (_00492_, _00491_, _00489_);
  nand (_00493_, _00492_, _06989_);
  nor (_14082_, _00493_, _00490_);
  and (_00495_, _09529_, _07454_);
  and (_00496_, _00495_, _06983_);
  and (_00497_, _00438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00498_, _00497_, _00423_);
  nand (_00499_, _00498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_00500_, _00498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00501_, _00500_, _00410_);
  and (_00503_, _00501_, _00499_);
  and (_00504_, _00497_, _00469_);
  or (_00505_, _00504_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00506_, _00505_, _00470_);
  nor (_00507_, _00506_, _00503_);
  or (_00508_, _00507_, _00381_);
  or (_00509_, _00382_, _09008_);
  and (_00510_, _00509_, _00508_);
  nor (_00511_, _00510_, _00496_);
  and (_00512_, _00496_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_00513_, _00512_, _00511_);
  and (_14085_, _00513_, _06989_);
  or (_00514_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor (_00515_, _00488_, rst);
  and (_14087_, _00515_, _00514_);
  nor (_00516_, _00382_, _11529_);
  nor (_00517_, _00418_, _00411_);
  or (_00518_, _00517_, _00471_);
  and (_00519_, _00518_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00520_, _00410_, _00467_);
  and (_00521_, _00520_, _00423_);
  or (_00522_, _00521_, _00468_);
  and (_00523_, _00522_, _00446_);
  or (_00524_, _00523_, _00519_);
  and (_00525_, _00524_, _00430_);
  and (_00526_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_00527_, _00526_, _00525_);
  or (_00528_, _00527_, _00516_);
  and (_14090_, _00528_, _06989_);
  and (_00530_, _09530_, _07454_);
  nand (_00531_, _00530_, _07118_);
  and (_00532_, _00438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  not (_00533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_00534_, _00533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_00535_, _00534_, _00410_);
  nor (_00536_, _00438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_00537_, _00536_, _00535_);
  nor (_00538_, _00537_, _00532_);
  and (_00539_, _00534_, _00439_);
  and (_00540_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_00541_, _00540_, _00538_);
  nor (_00542_, _00541_, _00381_);
  nor (_00543_, _00535_, _00381_);
  not (_00544_, _00543_);
  and (_00545_, _00544_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or (_00546_, _00545_, _00542_);
  or (_00547_, _00546_, _00530_);
  and (_00548_, _00547_, _06989_);
  and (_14105_, _00548_, _00531_);
  and (_00549_, _00532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_00550_, _00532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_00551_, _00550_, _00549_);
  nand (_00552_, _00551_, _00543_);
  or (_00553_, _00543_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_00554_, _00553_, _00552_);
  and (_00555_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_00556_, _00555_, _00429_);
  and (_00557_, _00556_, _00382_);
  or (_00558_, _00557_, _00554_);
  and (_00559_, _00558_, _06989_);
  nand (_00560_, _00530_, _10970_);
  and (_14108_, _00560_, _00559_);
  nand (_00561_, _00530_, _07260_);
  and (_00562_, _00397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_00563_, _00562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_00564_, _00563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_00565_, _00564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_00566_, _00565_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00567_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_00568_, _00567_, _00438_);
  and (_00569_, _00568_, _00566_);
  and (_00571_, _00534_, _00397_);
  and (_00572_, _00571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00573_, _00572_, _00415_);
  nor (_00574_, _00573_, _00569_);
  nor (_00576_, _00574_, _00381_);
  or (_00577_, _00567_, _00381_);
  and (_00578_, _00577_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or (_00579_, _00578_, _00576_);
  or (_00580_, _00579_, _00530_);
  and (_00581_, _00580_, _06989_);
  and (_14111_, _00581_, _00561_);
  and (_00582_, _00577_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_00583_, _00563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor (_00584_, _00564_, _00567_);
  and (_00585_, _00584_, _00583_);
  and (_00586_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_00587_, _00586_, _00585_);
  nor (_00589_, _00587_, _00381_);
  or (_00590_, _00589_, _00582_);
  or (_00591_, _00590_, _00530_);
  nand (_00592_, _00530_, _11529_);
  and (_00593_, _00592_, _06989_);
  and (_14115_, _00593_, _00591_);
  not (_00594_, _00496_);
  and (_00595_, _00577_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_00597_, _00564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_00598_, _00565_, _00567_);
  and (_00599_, _00598_, _00597_);
  and (_00600_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_00601_, _00600_, _00599_);
  nor (_00602_, _00601_, _00381_);
  or (_00603_, _00602_, _00595_);
  and (_00604_, _00603_, _00594_);
  nor (_00605_, _00594_, _07317_);
  or (_00606_, _00605_, _00604_);
  and (_14118_, _00606_, _06989_);
  and (_00607_, _00577_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_00608_, _00562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor (_00609_, _00563_, _00567_);
  and (_00610_, _00609_, _00608_);
  and (_00611_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_00612_, _00611_, _00610_);
  nor (_00613_, _00612_, _00381_);
  or (_00614_, _00613_, _00530_);
  or (_00615_, _00614_, _00607_);
  nand (_00616_, _00530_, _09008_);
  and (_00617_, _00616_, _06989_);
  and (_14121_, _00617_, _00615_);
  and (_00618_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_00619_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_00620_, _08139_, _00619_);
  or (_00621_, _00620_, _00618_);
  and (_14123_, _00621_, _06989_);
  or (_00622_, _00439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_00623_, _00498_, _00411_);
  and (_00624_, _00623_, _00622_);
  or (_00625_, _00438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_00627_, _00497_, _00385_);
  or (_00628_, _00627_, _00626_);
  and (_00629_, _00628_, _00625_);
  nor (_00630_, _00629_, _00624_);
  and (_00631_, _00630_, _00430_);
  nand (_00632_, _00381_, _09598_);
  not (_00633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand (_00634_, _00530_, _00633_);
  and (_00635_, _00634_, _06989_);
  nand (_00636_, _00635_, _00632_);
  nor (_14127_, _00636_, _00631_);
  and (_00637_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_14139_, _00637_, _09441_);
  nor (_14216_, _11613_, rst);
  and (_00640_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_00641_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_00642_, _00641_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_00643_, _00641_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_00644_, _00643_, _00642_);
  or (_00645_, _00644_, _00640_);
  and (_14225_, _00645_, _06989_);
  not (_00646_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  nor (_00648_, _00640_, _00646_);
  nor (_00649_, _00648_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_00650_, _00648_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_00651_, _00650_, _00649_);
  nor (_14227_, _00651_, rst);
  and (_00652_, _00640_, _00646_);
  nor (_00653_, _00652_, _00648_);
  and (_14255_, _00653_, _06989_);
  and (_00654_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_00655_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_00656_, _08139_, _00655_);
  or (_00657_, _00656_, _00654_);
  and (_14264_, _00657_, _06989_);
  or (_00658_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not (_00659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_00660_, _08139_, _00659_);
  and (_00661_, _00660_, _06989_);
  and (_14403_, _00661_, _00658_);
  not (_00662_, _00567_);
  and (_00664_, _00662_, _00397_);
  nand (_00665_, _00664_, _00382_);
  and (_00666_, _00665_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  not (_00668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_00669_, _00664_, _00668_);
  and (_00670_, _00534_, _00498_);
  nor (_00671_, _00670_, _00669_);
  nor (_00672_, _00671_, _00381_);
  or (_00673_, _00672_, _00666_);
  or (_00674_, _00673_, _00530_);
  nand (_00675_, _00530_, _09598_);
  and (_00676_, _00675_, _06989_);
  and (_14456_, _00676_, _00674_);
  nand (_00677_, _10146_, _09008_);
  or (_00678_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_00680_, _00678_, _06989_);
  and (_14572_, _00680_, _00677_);
  and (_00682_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not (_00683_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_00684_, _08139_, _00683_);
  or (_00685_, _00684_, _00682_);
  and (_14583_, _00685_, _06989_);
  or (_00686_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not (_00687_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_00688_, _08139_, _00687_);
  and (_00689_, _00688_, _06989_);
  and (_14585_, _00689_, _00686_);
  and (_00690_, _08036_, _07084_);
  and (_00691_, _00690_, _14026_);
  and (_00692_, _00691_, _06539_);
  nand (_00693_, _00692_, _06968_);
  or (_00694_, _00692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_00695_, _00694_, _06485_);
  and (_00696_, _00695_, _00693_);
  and (_00697_, _13950_, _07125_);
  nand (_00698_, _00697_, _07040_);
  or (_00699_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_00700_, _00699_, _06983_);
  and (_00701_, _00700_, _00698_);
  not (_00702_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor (_00703_, _06484_, _00702_);
  or (_00704_, _00703_, rst);
  or (_00706_, _00704_, _00701_);
  or (_14607_, _00706_, _00696_);
  and (_00707_, _09022_, _06500_);
  and (_00708_, _00707_, _14025_);
  and (_00709_, _00708_, _14196_);
  nand (_00710_, _00709_, _06968_);
  or (_00711_, _00709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nor (_00712_, _06477_, _06434_);
  and (_00713_, _00712_, _07453_);
  and (_00714_, _00713_, _14011_);
  not (_00715_, _00714_);
  and (_00716_, _00715_, _00711_);
  and (_00717_, _00716_, _00710_);
  nor (_00718_, _00715_, _10970_);
  or (_00719_, _00718_, _00717_);
  and (_00009_, _00719_, _06989_);
  and (_00720_, _08037_, _14026_);
  and (_00721_, _00720_, _06539_);
  nand (_00722_, _00721_, _06968_);
  or (_00723_, _00721_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_00724_, _00723_, _06485_);
  and (_00725_, _00724_, _00722_);
  and (_00726_, _07454_, _07125_);
  nand (_00727_, _00726_, _07040_);
  or (_00728_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_00729_, _00728_, _06983_);
  and (_00730_, _00729_, _00727_);
  not (_00731_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor (_00732_, _06484_, _00731_);
  or (_00733_, _00732_, rst);
  or (_00734_, _00733_, _00730_);
  or (_00018_, _00734_, _00725_);
  and (_00735_, _00708_, _07048_);
  nand (_00736_, _00735_, _06968_);
  or (_00737_, _00735_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_00738_, _00737_, _00715_);
  and (_00739_, _00738_, _00736_);
  nor (_00740_, _00715_, _07118_);
  or (_00741_, _00740_, _00739_);
  and (_00024_, _00741_, _06989_);
  and (_00742_, _00708_, _07044_);
  nand (_00743_, _00742_, _06968_);
  or (_00744_, _00742_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_00745_, _00744_, _00715_);
  and (_00746_, _00745_, _00743_);
  nor (_00747_, _00715_, _07260_);
  or (_00748_, _00747_, _00746_);
  and (_00026_, _00748_, _06989_);
  or (_00749_, _08435_, _07043_);
  nor (_00750_, _00749_, _07217_);
  or (_00751_, _00750_, _08437_);
  and (_00752_, _00751_, _00708_);
  nand (_00753_, _00708_, _06525_);
  and (_00754_, _00753_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_00755_, _00754_, _00714_);
  or (_00756_, _00755_, _00752_);
  nand (_00757_, _00714_, _07317_);
  and (_00758_, _00757_, _06989_);
  and (_00028_, _00758_, _00756_);
  not (_00759_, _09074_);
  nor (_00760_, _06968_, _00759_);
  and (_00761_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_00762_, _00761_, _00760_);
  and (_00763_, _00762_, _00708_);
  not (_00764_, _00749_);
  nand (_00765_, _00708_, _00764_);
  and (_00766_, _00765_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_00767_, _00766_, _00714_);
  or (_00768_, _00767_, _00763_);
  nand (_00769_, _00714_, _11529_);
  and (_00770_, _00769_, _06989_);
  and (_00031_, _00770_, _00768_);
  and (_00771_, _00708_, _07089_);
  or (_00772_, _00771_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_00773_, _00772_, _00715_);
  nand (_00774_, _00771_, _06968_);
  and (_00775_, _00774_, _00773_);
  nor (_00776_, _00715_, _09008_);
  or (_00777_, _00776_, _00775_);
  and (_00048_, _00777_, _06989_);
  and (_00778_, _00708_, _06979_);
  or (_00779_, _00778_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_00780_, _00779_, _00715_);
  nand (_00781_, _00778_, _06968_);
  and (_00782_, _00781_, _00780_);
  and (_00783_, _00714_, _09599_);
  or (_00784_, _00783_, _00782_);
  and (_00050_, _00784_, _06989_);
  or (_00785_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  nand (_00786_, _07493_, _07495_);
  and (_00787_, _00786_, _06989_);
  and (_00055_, _00787_, _00785_);
  not (_00788_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nor (_00789_, _00749_, _00788_);
  or (_00790_, _00789_, _08437_);
  and (_00791_, _00707_, _06449_);
  and (_00792_, _00791_, _00790_);
  and (_00793_, _09029_, _06986_);
  and (_00795_, _00791_, _06525_);
  nor (_00796_, _00795_, _00788_);
  or (_00797_, _00796_, _00793_);
  or (_00798_, _00797_, _00792_);
  nand (_00799_, _00793_, _07317_);
  and (_00800_, _00799_, _06989_);
  and (_00111_, _00800_, _00798_);
  and (_00801_, _00791_, _14196_);
  nand (_00802_, _00801_, _06968_);
  not (_00803_, _00793_);
  or (_00804_, _00801_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_00805_, _00804_, _00803_);
  and (_00806_, _00805_, _00802_);
  nor (_00807_, _00803_, _10970_);
  or (_00808_, _00807_, _00806_);
  and (_00113_, _00808_, _06989_);
  and (_00809_, _00791_, _07048_);
  nand (_00810_, _00809_, _06968_);
  or (_00811_, _00809_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_00812_, _00811_, _00803_);
  and (_00813_, _00812_, _00810_);
  nor (_00814_, _00803_, _07118_);
  or (_00815_, _00814_, _00813_);
  and (_00117_, _00815_, _06989_);
  and (_00816_, _00791_, _08349_);
  nor (_00817_, _06978_, _06525_);
  not (_00818_, _00791_);
  or (_00819_, _00818_, _00817_);
  or (_00820_, _00819_, _00795_);
  and (_00821_, _00820_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_00822_, _00821_, _00793_);
  or (_00823_, _00822_, _00816_);
  nand (_00824_, _00793_, _07260_);
  and (_00825_, _00824_, _06989_);
  and (_00119_, _00825_, _00823_);
  and (_00826_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _08578_);
  and (_00827_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_00828_, _00827_, _00826_);
  and (_00121_, _00828_, _06989_);
  and (_00829_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_00830_, _00829_, _00760_);
  and (_00831_, _00830_, _00791_);
  nand (_00832_, _00791_, _00764_);
  and (_00833_, _00832_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_00834_, _00833_, _00793_);
  or (_00835_, _00834_, _00831_);
  nand (_00836_, _00793_, _11529_);
  and (_00837_, _00836_, _06989_);
  and (_00123_, _00837_, _00835_);
  and (_00838_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _08578_);
  and (_00839_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00840_, _00839_, _00838_);
  and (_00128_, _00840_, _06989_);
  and (_00841_, _08578_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_00842_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_00843_, _00842_, _00841_);
  and (_00130_, _00843_, _06989_);
  and (_00844_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _08578_);
  and (_00845_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00846_, _00845_, _00844_);
  and (_00136_, _00846_, _06989_);
  and (_00847_, _00791_, _07089_);
  or (_00848_, _00847_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_00849_, _00848_, _00803_);
  nand (_00850_, _00847_, _06968_);
  and (_00851_, _00850_, _00849_);
  nor (_00852_, _00803_, _09008_);
  or (_00853_, _00852_, _00851_);
  and (_00138_, _00853_, _06989_);
  and (_00854_, _00791_, _06979_);
  or (_00855_, _00854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_00856_, _00855_, _00803_);
  nand (_00857_, _00854_, _06968_);
  and (_00858_, _00857_, _00856_);
  and (_00859_, _00793_, _09599_);
  or (_00860_, _00859_, _00858_);
  and (_00140_, _00860_, _06989_);
  and (_00861_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _08578_);
  and (_00862_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00863_, _00862_, _00861_);
  and (_00148_, _00863_, _06989_);
  and (_00864_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _08578_);
  and (_00865_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00866_, _00865_, _00864_);
  and (_00160_, _00866_, _06989_);
  and (_00867_, _14027_, _06449_);
  and (_00868_, _00867_, _07044_);
  nand (_00869_, _00868_, _06968_);
  or (_00870_, _00868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_00871_, _00870_, _07460_);
  and (_00872_, _00871_, _00869_);
  nor (_00873_, _07460_, _07260_);
  or (_00874_, _00873_, _00872_);
  and (_00162_, _00874_, _06989_);
  and (_00875_, _00867_, _09074_);
  nand (_00876_, _00875_, _06968_);
  or (_00877_, _00875_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_00878_, _00877_, _07460_);
  and (_00879_, _00878_, _00876_);
  nor (_00880_, _11529_, _07460_);
  or (_00881_, _00880_, _00879_);
  and (_00179_, _00881_, _06989_);
  and (_00882_, _00867_, _06979_);
  or (_00883_, _00882_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_00884_, _00883_, _07460_);
  nand (_00885_, _00882_, _06968_);
  and (_00886_, _00885_, _00884_);
  and (_00887_, _09599_, _07459_);
  or (_00888_, _00887_, _00886_);
  and (_00181_, _00888_, _06989_);
  and (_00889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_00890_, _00889_, _09510_);
  and (_00188_, _00890_, _06989_);
  nor (_00891_, _14042_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_00892_, _00891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_00893_, _00891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_00894_, _00893_, _06989_);
  and (_00213_, _00894_, _00892_);
  nor (_00895_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_00896_, _00895_, _09393_);
  and (_00897_, _00896_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not (_00898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor (_00899_, _00896_, _00898_);
  or (_00900_, _00899_, _00897_);
  or (_00901_, _00900_, _14028_);
  or (_00902_, _09074_, _00898_);
  nand (_00903_, _00902_, _14028_);
  or (_00904_, _00903_, _00760_);
  and (_00905_, _00904_, _00901_);
  or (_00906_, _00905_, _14031_);
  nand (_00907_, _14031_, _11529_);
  and (_00908_, _00907_, _06989_);
  and (_00219_, _00908_, _00906_);
  nor (_00909_, _07161_, _07166_);
  nand (_00910_, _00909_, _07274_);
  and (_00911_, _00909_, _07196_);
  or (_00912_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and (_00913_, _00912_, _06989_);
  and (_00222_, _00913_, _00910_);
  nand (_00914_, _07277_, _07274_);
  and (_00915_, _07277_, _07196_);
  or (_00916_, _00915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and (_00917_, _00916_, _06989_);
  and (_00228_, _00917_, _00914_);
  and (_00918_, _13972_, _13943_);
  nor (_00919_, _00918_, _13959_);
  and (_00920_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_00921_, _00920_, _13953_);
  and (_00922_, _13952_, _06989_);
  and (_00923_, _00922_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_00230_, _00923_, _00921_);
  nor (_00924_, _11413_, rst);
  and (_00250_, _00924_, _11964_);
  or (_00925_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00926_, _00925_, _07202_);
  or (_00927_, _00926_, _07208_);
  and (_00928_, _07212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_00929_, _00928_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00930_, _07215_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_00931_, _00930_, _07218_);
  and (_00932_, _00931_, _00929_);
  nand (_00933_, _07474_, _07218_);
  nand (_00934_, _00933_, _07207_);
  or (_00935_, _00934_, _00932_);
  and (_00936_, _00935_, _00927_);
  and (_00937_, _07474_, _07201_);
  or (_00938_, _00937_, _07222_);
  or (_00939_, _00938_, _00936_);
  not (_00940_, _07222_);
  or (_00941_, _00940_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00942_, _00941_, _00939_);
  and (_00943_, _00942_, _07197_);
  and (_00944_, _00925_, _07187_);
  or (_00945_, _00944_, _07194_);
  and (_00946_, _07175_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_00947_, _00946_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00948_, _07179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_00949_, _00948_, _07182_);
  and (_00950_, _00949_, _00947_);
  nand (_00951_, _07474_, _07182_);
  nand (_00952_, _00951_, _07193_);
  or (_00953_, _00952_, _00950_);
  and (_00954_, _00953_, _00945_);
  and (_00955_, _07474_, _07186_);
  or (_00956_, _00955_, _00954_);
  and (_00957_, _00956_, _07196_);
  or (_00958_, _00957_, _07161_);
  or (_00959_, _00958_, _00943_);
  or (_00960_, _07164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00961_, _00960_, _06989_);
  and (_00252_, _00961_, _00959_);
  not (_00962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_00963_, _00928_, _00962_);
  nand (_00964_, _00963_, _00931_);
  or (_00965_, _07465_, _07219_);
  and (_00966_, _00965_, _00964_);
  or (_00967_, _00966_, _07206_);
  not (_00968_, _07204_);
  not (_00969_, _07206_);
  or (_00970_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_00971_, _00970_, _00969_);
  and (_00972_, _00971_, _00968_);
  and (_00973_, _00972_, _00967_);
  and (_00974_, _07465_, _07204_);
  or (_00975_, _00974_, _07201_);
  or (_00976_, _00975_, _00973_);
  or (_00977_, _00970_, _07202_);
  nand (_00978_, _00977_, _00976_);
  nand (_00979_, _00978_, _07274_);
  not (_00980_, _07189_);
  or (_00981_, _07465_, _00980_);
  or (_00982_, _00946_, _00962_);
  nand (_00983_, _00982_, _00949_);
  not (_00984_, _07191_);
  or (_00985_, _07465_, _07183_);
  and (_00986_, _00985_, _00984_);
  and (_00987_, _00986_, _00983_);
  and (_00988_, _00970_, _07191_);
  or (_00989_, _00988_, _07189_);
  or (_00990_, _00989_, _00987_);
  and (_00991_, _00990_, _00981_);
  or (_00992_, _00991_, _07186_);
  or (_00993_, _00970_, _07187_);
  and (_00994_, _00993_, _00992_);
  or (_00995_, _00994_, _07197_);
  and (_00996_, _00995_, _00979_);
  or (_00997_, _00996_, _07161_);
  nor (_00998_, _07223_, _07161_);
  or (_00999_, _00998_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_01001_, _00999_, _06989_);
  and (_00254_, _01001_, _00997_);
  or (_01002_, _00642_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_00256_, _01002_, _06989_);
  nor (_00258_, _12740_, rst);
  nand (_01003_, _11351_, _06989_);
  nor (_00261_, _01003_, _11417_);
  or (_01004_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01005_, _01004_, _07202_);
  or (_01006_, _01005_, _07208_);
  and (_01007_, _07212_, _07166_);
  or (_01008_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01009_, _07215_, _07166_);
  nor (_01010_, _01009_, _07218_);
  and (_01011_, _01010_, _01008_);
  nand (_01012_, _07473_, _07218_);
  nand (_01013_, _01012_, _07207_);
  or (_01014_, _01013_, _01011_);
  and (_01015_, _01014_, _01006_);
  and (_01016_, _07473_, _07201_);
  or (_01017_, _01016_, _07222_);
  or (_01018_, _01017_, _01015_);
  or (_01019_, _00940_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01020_, _01019_, _01018_);
  and (_01021_, _01020_, _07197_);
  and (_01022_, _01004_, _07187_);
  or (_01024_, _01022_, _07194_);
  and (_01025_, _07175_, _07166_);
  or (_01026_, _01025_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01027_, _07179_, _07166_);
  nor (_01028_, _01027_, _07182_);
  and (_01029_, _01028_, _01026_);
  nand (_01030_, _07473_, _07182_);
  nand (_01031_, _01030_, _07193_);
  or (_01032_, _01031_, _01029_);
  and (_01033_, _01032_, _01024_);
  and (_01034_, _07473_, _07186_);
  or (_01035_, _01034_, _01033_);
  and (_01036_, _01035_, _07196_);
  or (_01037_, _01036_, _07161_);
  or (_01038_, _01037_, _01021_);
  or (_01039_, _07164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_01040_, _01039_, _06989_);
  and (_00272_, _01040_, _01038_);
  nor (_01041_, _07196_, _07161_);
  and (_01042_, _07222_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not (_01043_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_01044_, _01007_, _01043_);
  nand (_01045_, _01044_, _01010_);
  or (_01046_, _07464_, _07219_);
  and (_01047_, _01046_, _01045_);
  or (_01048_, _01047_, _07206_);
  or (_01049_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_01050_, _01049_, _00969_);
  and (_01051_, _01050_, _00968_);
  and (_01052_, _01051_, _01048_);
  and (_01053_, _07464_, _07204_);
  or (_01054_, _01053_, _07201_);
  or (_01055_, _01054_, _01052_);
  nor (_01056_, _01049_, _07202_);
  nor (_01057_, _01056_, _07222_);
  and (_01058_, _01057_, _01055_);
  or (_01059_, _01058_, _01042_);
  and (_01060_, _01059_, _01041_);
  or (_01061_, _07189_, _07182_);
  or (_01062_, _01061_, _07175_);
  and (_01063_, _01062_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_01064_, _01063_, _07179_);
  nand (_01065_, _07182_, _07166_);
  and (_01066_, _01065_, _01064_);
  or (_01067_, _01066_, _07191_);
  nand (_01068_, _07189_, _07166_);
  and (_01069_, _01068_, _01067_);
  or (_01070_, _07186_, _07161_);
  or (_01071_, _01070_, _01069_);
  or (_01072_, _07277_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_01073_, \oc8051_top_1.oc8051_memory_interface1.reti , _07165_);
  or (_01074_, _01073_, _07170_);
  and (_01075_, _01074_, _01072_);
  and (_01076_, _01075_, _01071_);
  or (_01077_, _01076_, _01060_);
  and (_00275_, _01077_, _06989_);
  nand (_01078_, _07277_, _07223_);
  or (_01079_, _01041_, _07166_);
  and (_01080_, _01079_, _06989_);
  and (_00289_, _01080_, _01078_);
  and (_01081_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _06989_);
  and (_00310_, _01081_, _07161_);
  nor (_01082_, _07216_, _07199_);
  and (_01083_, _07219_, _07208_);
  nand (_01084_, _01083_, _01082_);
  nor (_01085_, _01084_, _07196_);
  and (_01086_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  or (_01087_, _07182_, _07161_);
  nor (_01088_, _01087_, _07171_);
  not (_01089_, _07194_);
  nor (_01090_, _01089_, _07180_);
  and (_01091_, _01090_, _01088_);
  or (_01092_, _01091_, _01086_);
  or (_01093_, _01092_, _01085_);
  and (_00318_, _01093_, _06989_);
  or (_01094_, _07218_, _07206_);
  and (_01095_, _07216_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_01096_, _01095_, _01094_);
  and (_01097_, _01096_, _00968_);
  and (_01098_, _07274_, _07202_);
  and (_01099_, _01098_, _01097_);
  or (_01100_, _07191_, _07182_);
  and (_01101_, _07180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_01102_, _01101_, _01100_);
  and (_01103_, _01102_, _00980_);
  and (_01104_, _07196_, _07187_);
  and (_01105_, _01104_, _01103_);
  or (_01106_, _01105_, _07161_);
  or (_01107_, _01106_, _01099_);
  or (_01108_, _07164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_01109_, _01108_, _06989_);
  and (_00321_, _01109_, _01107_);
  nor (_01110_, _07212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_01111_, _01110_, _07215_);
  or (_01112_, _01111_, _07218_);
  and (_01113_, _01112_, _00969_);
  or (_01114_, _01113_, _07204_);
  and (_01115_, _01114_, _01098_);
  nor (_01116_, _07175_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_01117_, _01116_, _07179_);
  or (_01118_, _01117_, _07182_);
  and (_01119_, _01118_, _00984_);
  or (_01120_, _01119_, _07189_);
  and (_01121_, _01120_, _01104_);
  or (_01122_, _01121_, _07161_);
  or (_01123_, _01122_, _01115_);
  or (_01124_, _07164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01125_, _01124_, _06989_);
  and (_00325_, _01125_, _01123_);
  and (_00327_, _12822_, _07161_);
  and (_01126_, _14028_, _07048_);
  nand (_01127_, _01126_, _06968_);
  or (_01128_, _01126_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_01129_, _01128_, _14032_);
  and (_01130_, _01129_, _01127_);
  nor (_01131_, _14032_, _07118_);
  or (_01132_, _01131_, _01130_);
  and (_00334_, _01132_, _06989_);
  and (_01133_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_01134_, _01133_, _00998_);
  and (_00345_, _01134_, _06989_);
  and (_01135_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_01136_, _01135_, _00998_);
  and (_00348_, _01136_, _06989_);
  or (_01137_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  nand (_01138_, _07493_, _09525_);
  and (_01139_, _01138_, _06989_);
  and (_00387_, _01139_, _01137_);
  and (_01140_, _12937_, _09009_);
  and (_01141_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or (_01142_, _01141_, _01140_);
  and (_00442_, _01142_, _06989_);
  or (_01143_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  not (_01144_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_01145_, _08139_, _01144_);
  and (_01146_, _01145_, _06989_);
  and (_00445_, _01146_, _01143_);
  and (_01147_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_00453_, _01147_, _09459_);
  or (_01148_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  not (_01149_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_01150_, _08139_, _01149_);
  and (_01151_, _01150_, _06989_);
  and (_00457_, _01151_, _01148_);
  and (_01152_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_00465_, _01152_, _09466_);
  nor (_01153_, _12938_, _07317_);
  and (_01154_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_01155_, _01154_, _01153_);
  and (_00494_, _01155_, _06989_);
  and (_01156_, _00690_, _09022_);
  and (_01157_, _01156_, _06539_);
  nand (_01158_, _01157_, _06968_);
  or (_01159_, _01157_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_01160_, _01159_, _06485_);
  and (_01161_, _01160_, _01158_);
  and (_01162_, _00713_, _07125_);
  not (_01163_, _01162_);
  nor (_01164_, _01163_, _07040_);
  not (_01165_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor (_01166_, _01162_, _01165_);
  or (_01167_, _01166_, _01164_);
  and (_01168_, _01167_, _06983_);
  nor (_01169_, _06484_, _01165_);
  or (_01170_, _01169_, rst);
  or (_01171_, _01170_, _01168_);
  or (_00502_, _01171_, _01161_);
  and (_01172_, _14190_, _07429_);
  and (_01173_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or (_01174_, _01173_, _01172_);
  and (_00529_, _01174_, _06989_);
  and (_01175_, _14028_, _08349_);
  not (_01176_, _14028_);
  or (_01177_, _00817_, _01176_);
  and (_01179_, _14028_, _06525_);
  or (_01180_, _01179_, _01177_);
  and (_01181_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_01182_, _01181_, _14031_);
  or (_01183_, _01182_, _01175_);
  nand (_01184_, _14031_, _07260_);
  and (_01185_, _01184_, _06989_);
  and (_00570_, _01185_, _01183_);
  or (_01186_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not (_01188_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_01189_, _08139_, _01188_);
  and (_01190_, _01189_, _06989_);
  and (_00575_, _01190_, _01186_);
  or (_01191_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  not (_01192_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_01193_, _08139_, _01192_);
  and (_01194_, _01193_, _06989_);
  and (_00588_, _01194_, _01191_);
  nor (_00596_, _11513_, rst);
  and (_01195_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_01196_, _08139_, _01192_);
  or (_01197_, _01196_, _01195_);
  and (_00638_, _01197_, _06989_);
  not (_01198_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor (_01199_, _00749_, _01198_);
  or (_01200_, _01199_, _08437_);
  and (_01202_, _01200_, _14028_);
  nor (_01203_, _01179_, _01198_);
  or (_01204_, _01203_, _14031_);
  or (_01205_, _01204_, _01202_);
  nand (_01206_, _14031_, _07317_);
  and (_01207_, _01206_, _06989_);
  and (_00639_, _01207_, _01205_);
  nor (_01209_, _10961_, _07335_);
  nor (_01210_, _10950_, _07349_);
  and (_01211_, _10950_, _07349_);
  nor (_01212_, _01211_, _01210_);
  and (_01213_, _01212_, _01209_);
  nor (_01214_, _01212_, _01209_);
  nor (_01215_, _01214_, _01213_);
  or (_01216_, _01215_, _07490_);
  or (_01217_, _07325_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01218_, _01217_, _10964_);
  and (_00647_, _01218_, _01216_);
  or (_01219_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  not (_01220_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_01221_, _08139_, _01220_);
  and (_01222_, _01221_, _06989_);
  and (_00663_, _01222_, _01219_);
  and (_01223_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_01224_, _08139_, _01220_);
  or (_01225_, _01224_, _01223_);
  and (_00667_, _01225_, _06989_);
  or (_01226_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  not (_01227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_01228_, _08139_, _01227_);
  and (_01229_, _01228_, _06989_);
  and (_00679_, _01229_, _01226_);
  and (_01230_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_01231_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_01232_, _08139_, _01231_);
  or (_01233_, _01232_, _01230_);
  and (_00681_, _01233_, _06989_);
  or (_01234_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand (_01235_, _07493_, _14104_);
  and (_01236_, _01235_, _06989_);
  and (_00705_, _01236_, _01234_);
  nor (_01237_, _13945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_01238_, _01237_, _13946_);
  and (_00794_, _01238_, _13953_);
  and (_01239_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_01241_, _01239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_01000_, _01241_, _06989_);
  and (_01242_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_01243_, _01242_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_01023_, _01243_, _06989_);
  not (_01244_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nor (_01245_, _14404_, _01244_);
  nand (_01246_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand (_01247_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_01248_, _01247_, _01246_);
  nand (_01249_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nand (_01251_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_01252_, _01251_, _01249_);
  and (_01253_, _01252_, _01248_);
  nand (_01254_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  nand (_01255_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_01256_, _01255_, _01254_);
  nand (_01257_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nand (_01258_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_01259_, _01258_, _01257_);
  and (_01260_, _01259_, _01256_);
  and (_01261_, _01260_, _01253_);
  nand (_01262_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nand (_01263_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_01264_, _01263_, _01262_);
  nand (_01265_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand (_01266_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_01267_, _01266_, _01265_);
  and (_01268_, _01267_, _01264_);
  nand (_01269_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  nand (_01270_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_01271_, _01270_, _01269_);
  nand (_01272_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  nand (_01273_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_01274_, _01273_, _01272_);
  and (_01275_, _01274_, _01271_);
  and (_01276_, _01275_, _01268_);
  and (_01277_, _01276_, _01261_);
  nand (_01278_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand (_01279_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and (_01280_, _01279_, _01278_);
  nand (_01281_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_01282_, _14296_, _11683_);
  and (_01283_, _01282_, _01281_);
  and (_01284_, _01283_, _01280_);
  nor (_01285_, _14326_, p0_in[5]);
  not (_01286_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01287_, _14326_, _01286_);
  nor (_01288_, _01287_, _01285_);
  nand (_01289_, _01288_, _14339_);
  nor (_01290_, _14326_, p1_in[5]);
  not (_01291_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_01292_, _14326_, _01291_);
  nor (_01293_, _01292_, _01290_);
  nand (_01294_, _01293_, _14344_);
  and (_01295_, _01294_, _01289_);
  or (_01296_, _14326_, p2_in[5]);
  or (_01297_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_01298_, _01297_, _01296_);
  nand (_01299_, _01298_, _14333_);
  nor (_01300_, _14326_, p3_in[5]);
  not (_01301_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_01302_, _14326_, _01301_);
  nor (_01303_, _01302_, _01300_);
  nand (_01304_, _01303_, _14305_);
  and (_01305_, _01304_, _01299_);
  and (_01306_, _01305_, _01295_);
  and (_01307_, _01306_, _01284_);
  nand (_01308_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand (_01309_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01310_, _01309_, _01308_);
  and (_01311_, _01310_, _01307_);
  nand (_01312_, _01311_, _01277_);
  and (_01313_, _01312_, _14374_);
  or (_01314_, _01313_, _14213_);
  or (_01315_, _01314_, _01245_);
  or (_01316_, _14483_, _08268_);
  and (_01317_, _01316_, _06989_);
  and (_01187_, _01317_, _01315_);
  and (_01318_, _00690_, _08038_);
  nand (_01319_, _01318_, _06979_);
  or (_01320_, _01319_, _08268_);
  not (_01321_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_01322_, _01319_, _01321_);
  and (_01323_, _01322_, _06983_);
  and (_01324_, _01323_, _01320_);
  nor (_01325_, _06484_, _01321_);
  and (_01326_, _01318_, _07048_);
  nand (_01327_, _01326_, _06968_);
  or (_01328_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01329_, _01328_, _06485_);
  and (_01330_, _01329_, _01327_);
  or (_01331_, _01330_, _01325_);
  or (_01332_, _01331_, _01324_);
  and (_01201_, _01332_, _06989_);
  nor (_01333_, _11529_, _07262_);
  and (_01334_, _10974_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or (_01335_, _01334_, _01333_);
  and (_01208_, _01335_, _06989_);
  and (_01336_, _09599_, _09488_);
  and (_01337_, _09489_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or (_01338_, _01337_, _01336_);
  and (_01240_, _01338_, _06989_);
  and (_01339_, _09599_, _09605_);
  and (_01340_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or (_01341_, _01340_, _06982_);
  or (_01342_, _01341_, _01339_);
  or (_01343_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_01344_, _01343_, _06989_);
  and (_01250_, _01344_, _01342_);
  and (_01345_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not (_01346_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_01347_, _08139_, _01346_);
  or (_01348_, _01347_, _01345_);
  and (_01627_, _01348_, _06989_);
  and (_01349_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_01350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_01351_, _08139_, _01350_);
  or (_01352_, _01351_, _01349_);
  and (_01629_, _01352_, _06989_);
  or (_01353_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_01354_, _01353_, _14028_);
  nand (_01355_, _08032_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_01356_, _01355_, _14028_);
  or (_01357_, _01356_, _08033_);
  and (_01358_, _01357_, _01354_);
  or (_01359_, _01358_, _14031_);
  nand (_01360_, _14031_, _09008_);
  and (_01361_, _01360_, _06989_);
  and (_01649_, _01361_, _01359_);
  and (_01363_, _14190_, _07410_);
  and (_01364_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_01365_, _01364_, _01363_);
  and (_01662_, _01365_, _06989_);
  nor (_01366_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_01367_, _01366_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  not (_01368_, _01367_);
  or (_01369_, _01368_, _08433_);
  or (_01370_, _01367_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_01371_, _01370_, _06989_);
  and (_01669_, _01371_, _01369_);
  not (_01372_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_01373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01372_);
  or (_01374_, _01373_, _09392_);
  and (_01375_, _01374_, _00895_);
  or (_01376_, _01375_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_01377_, _01376_, _14028_);
  or (_01378_, _06979_, _09407_);
  nand (_01379_, _01378_, _14028_);
  or (_01380_, _01379_, _08127_);
  and (_01381_, _01380_, _01377_);
  or (_01382_, _01381_, _14031_);
  nand (_01383_, _14031_, _09598_);
  and (_01384_, _01383_, _06989_);
  and (_01673_, _01384_, _01382_);
  and (_01385_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_01386_, _01385_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_01695_, _01386_, _06989_);
  and (_01387_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_01388_, _01387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_01697_, _01388_, _06989_);
  nand (_01389_, _01367_, _09227_);
  or (_01390_, _01367_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_01391_, _01390_, _06989_);
  and (_01711_, _01391_, _01389_);
  and (_01392_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_01393_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or (_01394_, _01393_, _01392_);
  and (_01721_, _01394_, _06989_);
  and (_01395_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_01396_, _01395_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_01732_, _01396_, _06989_);
  and (_01397_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_01398_, _01397_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01734_, _01398_, _06989_);
  or (_01399_, _01368_, _08030_);
  or (_01400_, _01367_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_01401_, _01400_, _06989_);
  and (_01762_, _01401_, _01399_);
  and (_01402_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_01403_, _14190_, _11646_);
  or (_01404_, _01403_, _01402_);
  and (_01770_, _01404_, _06989_);
  and (_01405_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_01406_, _07486_, _07040_);
  or (_01407_, _01406_, _01405_);
  and (_01800_, _01407_, _06989_);
  or (_01408_, _01368_, _08123_);
  or (_01409_, _01367_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_01410_, _01409_, _06989_);
  and (_01803_, _01410_, _01408_);
  and (_01411_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_01412_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or (_01413_, _01412_, _01411_);
  and (_01817_, _01413_, _06989_);
  nor (_01821_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  not (_01414_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nor (_01415_, _14404_, _01414_);
  nand (_01416_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand (_01417_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_01418_, _01417_, _01416_);
  nand (_01419_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nand (_01420_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_01421_, _01420_, _01419_);
  and (_01422_, _01421_, _01418_);
  nand (_01423_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand (_01424_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_01425_, _01424_, _01423_);
  nand (_01426_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand (_01427_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_01428_, _01427_, _01426_);
  and (_01429_, _01428_, _01425_);
  and (_01430_, _01429_, _01422_);
  nand (_01431_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nand (_01432_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_01433_, _01432_, _01431_);
  nand (_01434_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_01435_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_01436_, _01435_, _01434_);
  and (_01437_, _01436_, _01433_);
  nand (_01438_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand (_01439_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and (_01440_, _01439_, _01438_);
  nand (_01441_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand (_01442_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_01443_, _01442_, _01441_);
  and (_01444_, _01443_, _01440_);
  and (_01445_, _01444_, _01437_);
  and (_01446_, _01445_, _01430_);
  nand (_01447_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_01448_, _14296_, _11698_);
  and (_01449_, _01448_, _01447_);
  nand (_01450_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand (_01451_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_01452_, _01451_, _01450_);
  and (_01453_, _01452_, _01449_);
  nor (_01454_, _14326_, p1_in[4]);
  not (_01455_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_01456_, _14326_, _01455_);
  nor (_01457_, _01456_, _01454_);
  nand (_01458_, _01457_, _14344_);
  nor (_01459_, _14326_, p0_in[4]);
  not (_01460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_01461_, _14326_, _01460_);
  nor (_01462_, _01461_, _01459_);
  nand (_01463_, _01462_, _14339_);
  and (_01464_, _01463_, _01458_);
  nor (_01465_, _14326_, p3_in[4]);
  not (_01466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_01467_, _14326_, _01466_);
  nor (_01468_, _01467_, _01465_);
  nand (_01469_, _01468_, _14305_);
  nor (_01470_, _14326_, p2_in[4]);
  not (_01471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_01472_, _14326_, _01471_);
  nor (_01473_, _01472_, _01470_);
  nand (_01474_, _01473_, _14333_);
  and (_01475_, _01474_, _01469_);
  and (_01476_, _01475_, _01464_);
  and (_01477_, _01476_, _01453_);
  nand (_01478_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand (_01479_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_01480_, _01479_, _01478_);
  and (_01481_, _01480_, _01477_);
  nand (_01482_, _01481_, _01446_);
  nand (_01483_, _01482_, _14374_);
  nand (_01484_, _01483_, _14483_);
  or (_01485_, _01484_, _01415_);
  or (_01486_, _14483_, _08346_);
  and (_01487_, _01486_, _06989_);
  and (_01823_, _01487_, _01485_);
  nand (_01488_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_01489_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_01490_, _01489_, _01488_);
  nand (_01491_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_01492_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_01493_, _01492_, _01491_);
  and (_01494_, _01493_, _01490_);
  nand (_01495_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand (_01496_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_01497_, _01496_, _01495_);
  nand (_01498_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand (_01499_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_01500_, _01499_, _01498_);
  and (_01501_, _01500_, _01497_);
  and (_01502_, _01501_, _01494_);
  nand (_01503_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand (_01504_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_01505_, _01504_, _01503_);
  nand (_01506_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand (_01507_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_01508_, _01507_, _01506_);
  and (_01509_, _01508_, _01505_);
  nand (_01510_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_01511_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and (_01512_, _01511_, _01510_);
  nand (_01513_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_01514_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_01515_, _01514_, _01513_);
  and (_01516_, _01515_, _01512_);
  and (_01517_, _01516_, _01509_);
  and (_01518_, _01517_, _01502_);
  nand (_01519_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand (_01520_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and (_01521_, _01520_, _01519_);
  nand (_01522_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_01523_, _14296_, _11795_);
  and (_01524_, _01523_, _01522_);
  and (_01525_, _01524_, _01521_);
  nor (_01527_, _14326_, p2_in[0]);
  not (_01528_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_01529_, _14326_, _01528_);
  nor (_01530_, _01529_, _01527_);
  nand (_01531_, _01530_, _14333_);
  nor (_01532_, _14326_, p3_in[0]);
  not (_01533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_01534_, _14326_, _01533_);
  nor (_01535_, _01534_, _01532_);
  nand (_01536_, _01535_, _14305_);
  and (_01537_, _01536_, _01531_);
  nor (_01538_, _14326_, p0_in[0]);
  not (_01539_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_01540_, _14326_, _01539_);
  nor (_01541_, _01540_, _01538_);
  nand (_01542_, _01541_, _14339_);
  nor (_01543_, _14326_, p1_in[0]);
  not (_01544_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_01545_, _14326_, _01544_);
  nor (_01546_, _01545_, _01543_);
  nand (_01547_, _01546_, _14344_);
  and (_01548_, _01547_, _01542_);
  and (_01549_, _01548_, _01537_);
  and (_01550_, _01549_, _01525_);
  nand (_01551_, _08359_, _08279_);
  or (_01552_, _08359_, _08279_);
  nand (_01553_, _01552_, _01551_);
  or (_01554_, _09145_, _07710_);
  not (_01555_, _14196_);
  nor (_01556_, _06968_, _01555_);
  nor (_01557_, _14196_, _06813_);
  nor (_01558_, _01557_, _01556_);
  nor (_01559_, _01558_, _08043_);
  nor (_01560_, _11948_, _06813_);
  or (_01561_, _01560_, _07699_);
  nor (_01562_, _01561_, _01559_);
  nand (_01563_, _01562_, _01554_);
  and (_01564_, _09285_, _07699_);
  not (_01565_, _01564_);
  and (_01566_, _01565_, _01563_);
  or (_01567_, _01566_, _12316_);
  nand (_01568_, _01566_, _12316_);
  and (_01569_, _01568_, _01567_);
  nand (_01570_, _01569_, _01553_);
  or (_01571_, _01569_, _01553_);
  nand (_01572_, _01571_, _01570_);
  nand (_01573_, _08138_, _08052_);
  or (_01574_, _08138_, _08052_);
  nand (_01575_, _01574_, _01573_);
  or (_01576_, _09227_, _07710_);
  nor (_01577_, _09074_, _06703_);
  nor (_01578_, _01577_, _00760_);
  nor (_01579_, _01578_, _08043_);
  nor (_01580_, _11948_, _06703_);
  or (_01581_, _01580_, _07699_);
  nor (_01582_, _01581_, _01579_);
  nand (_01583_, _01582_, _01576_);
  and (_01584_, _09356_, _07699_);
  not (_01585_, _01584_);
  and (_01586_, _01585_, _01583_);
  or (_01587_, _01586_, _08447_);
  nand (_01588_, _01586_, _08447_);
  and (_01589_, _01588_, _01587_);
  nand (_01590_, _01589_, _01575_);
  or (_01591_, _01589_, _01575_);
  nand (_01592_, _01591_, _01590_);
  nand (_01593_, _01592_, _01572_);
  or (_01594_, _01592_, _01572_);
  and (_01595_, _01594_, _01593_);
  nand (_01596_, _01595_, _14355_);
  nand (_01597_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_01598_, _01597_, _01596_);
  and (_01599_, _01598_, _01550_);
  and (_01600_, _01599_, _01518_);
  nor (_01601_, _01600_, _14377_);
  not (_01602_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nor (_01603_, _14404_, _01602_);
  or (_01604_, _01603_, _14213_);
  or (_01605_, _01604_, _01601_);
  or (_01606_, _14483_, _08123_);
  and (_01607_, _01606_, _06989_);
  and (_01825_, _01607_, _01605_);
  and (_01608_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_01609_, _08139_, _00687_);
  or (_01610_, _01609_, _01608_);
  and (_01835_, _01610_, _06989_);
  not (_01611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_01612_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01613_, _11004_, _01612_);
  and (_01614_, _01613_, _01611_);
  nor (_01615_, _01613_, _01611_);
  nor (_01616_, _01615_, _01614_);
  not (_01617_, _01616_);
  nor (_01618_, _11004_, _01612_);
  or (_01619_, _01618_, _01613_);
  and (_01620_, _01619_, _11055_);
  and (_01621_, _01620_, _01617_);
  nor (_01622_, _01620_, _01617_);
  nor (_01623_, _01622_, _01621_);
  or (_01624_, _01623_, _08477_);
  or (_01625_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01626_, _01625_, _10964_);
  and (_01628_, _01626_, _01624_);
  and (_01630_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_01860_, _01630_, _01628_);
  not (_01631_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_01632_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_01633_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_01634_, _01614_, _01633_);
  and (_01635_, _01634_, _01632_);
  nor (_01636_, _01635_, _01631_);
  and (_01637_, _01635_, _01631_);
  nor (_01638_, _01637_, _01636_);
  not (_01639_, _01638_);
  nor (_01640_, _01634_, _01632_);
  or (_01641_, _01640_, _01635_);
  nor (_01642_, _01614_, _01633_);
  nor (_01643_, _01642_, _01634_);
  not (_01644_, _01643_);
  and (_01645_, _01644_, _01621_);
  and (_01646_, _01645_, _01641_);
  and (_01647_, _01646_, _01639_);
  nor (_01648_, _01646_, _01639_);
  nor (_01650_, _01648_, _01647_);
  or (_01651_, _01650_, _08477_);
  or (_01652_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01653_, _01652_, _10964_);
  and (_01654_, _01653_, _01651_);
  and (_01655_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01865_, _01655_, _01654_);
  nor (_01656_, _01645_, _01641_);
  nor (_01657_, _01656_, _01646_);
  or (_01658_, _01657_, _08477_);
  or (_01659_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01660_, _01659_, _10964_);
  and (_01661_, _01660_, _01658_);
  and (_01663_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_01870_, _01663_, _01661_);
  nor (_01664_, _13943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_01665_, _01664_, _13944_);
  and (_01896_, _01665_, _13953_);
  and (_01666_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_01667_, _08139_, _00659_);
  or (_01668_, _01667_, _01666_);
  and (_02001_, _01668_, _06989_);
  nor (_01670_, _01644_, _01621_);
  nor (_01671_, _01670_, _01645_);
  or (_01672_, _01671_, _08477_);
  or (_01674_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01675_, _01674_, _10964_);
  and (_01676_, _01675_, _01672_);
  and (_01677_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_02024_, _01677_, _01676_);
  nor (_01678_, _01619_, _11055_);
  nor (_01679_, _01678_, _01620_);
  or (_01680_, _01679_, _08477_);
  or (_01681_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01682_, _01681_, _10964_);
  and (_01683_, _01682_, _01680_);
  and (_01684_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_02056_, _01684_, _01683_);
  and (_01685_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_01686_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_01687_, _08139_, _01686_);
  or (_01688_, _01687_, _01685_);
  and (_02058_, _01688_, _06989_);
  or (_01689_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_01690_, _08139_, _08171_);
  and (_01691_, _01690_, _06989_);
  and (_02100_, _01691_, _01689_);
  or (_01692_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_01693_, _01692_, _06989_);
  nand (_01694_, _14016_, _07118_);
  and (_02185_, _01694_, _01693_);
  or (_01696_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_01698_, _01696_, _06989_);
  nand (_01699_, _14016_, _10970_);
  and (_02212_, _01699_, _01698_);
  or (_01700_, _09760_, _09398_);
  or (_01701_, _09762_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_01702_, _01701_, _06989_);
  and (_02225_, _01702_, _01700_);
  or (_01703_, _14055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand (_01704_, _14055_, _14046_);
  and (_01705_, _01704_, _06989_);
  and (_02284_, _01705_, _01703_);
  or (_01706_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_01707_, _01706_, _06989_);
  nand (_01708_, _14016_, _07260_);
  and (_02286_, _01708_, _01707_);
  nor (_01709_, _10970_, _09489_);
  nor (_01710_, _07131_, _06982_);
  or (_01712_, _01710_, _07134_);
  and (_01713_, _01712_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or (_01714_, _01713_, _01709_);
  and (_02294_, _01714_, _06989_);
  nor (_01715_, _07260_, _09614_);
  and (_01716_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_01717_, _01716_, _06982_);
  or (_01718_, _01717_, _01715_);
  or (_01719_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_01720_, _01719_, _06989_);
  and (_02297_, _01720_, _01718_);
  or (_01722_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_01723_, _01722_, _06989_);
  nand (_01724_, _14016_, _07317_);
  and (_02300_, _01724_, _01723_);
  and (_02542_, _01566_, _06989_);
  or (_01725_, _01319_, _08433_);
  not (_01726_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_01727_, _01319_, _01726_);
  and (_01728_, _01727_, _06983_);
  and (_01729_, _01728_, _01725_);
  nor (_01730_, _06484_, _01726_);
  nand (_01731_, _01318_, _06525_);
  and (_01733_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_01735_, _00749_, _01726_);
  or (_01736_, _01735_, _08437_);
  and (_01737_, _01736_, _01318_);
  or (_01738_, _01737_, _01733_);
  and (_01739_, _01738_, _06485_);
  or (_01740_, _01739_, _01730_);
  or (_01741_, _01740_, _01729_);
  and (_02563_, _01741_, _06989_);
  and (_02576_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _06989_);
  or (_01742_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand (_01743_, _07493_, _14099_);
  and (_01744_, _01743_, _06989_);
  and (_02578_, _01744_, _01742_);
  or (_01745_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or (_01746_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and (_01747_, _01746_, _06989_);
  and (_02597_, _01747_, _01745_);
  or (_01748_, _01319_, _08346_);
  not (_01749_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_01750_, _01319_, _01749_);
  and (_01751_, _01750_, _06983_);
  and (_01752_, _01751_, _01748_);
  nor (_01753_, _06484_, _01749_);
  and (_01754_, _01318_, _07044_);
  nand (_01755_, _01754_, _06968_);
  or (_01756_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01757_, _01756_, _06485_);
  and (_01758_, _01757_, _01755_);
  or (_01759_, _01758_, _01753_);
  or (_01760_, _01759_, _01752_);
  and (_02622_, _01760_, _06989_);
  and (_01761_, _09599_, _07261_);
  and (_01763_, _10974_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  or (_01764_, _01763_, _01761_);
  and (_02650_, _01764_, _06989_);
  or (_01765_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_01766_, _01765_, _06989_);
  nand (_01767_, _00005_, _07040_);
  and (_02668_, _01767_, _01766_);
  nand (_01768_, _00027_, _07040_);
  and (_01769_, _00105_, _00059_);
  or (_01771_, _01769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_01772_, _01769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_01773_, _01772_, _01771_);
  and (_01774_, _01773_, _00062_);
  and (_01775_, _00084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_01776_, _01775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01777_, _01775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_01778_, _01777_, _00083_);
  nor (_01779_, _01778_, _01776_);
  or (_01780_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_01781_, _01780_, _00051_);
  and (_01782_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_01783_, _01782_, _01781_);
  or (_01784_, _01783_, _01779_);
  or (_01785_, _01784_, _01774_);
  or (_01786_, _01785_, _00027_);
  and (_01787_, _01786_, _00092_);
  and (_01788_, _01787_, _01768_);
  and (_01789_, _00091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01790_, _01789_, _01788_);
  and (_02671_, _01790_, _06989_);
  not (_01791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_01792_, _00079_, _01791_);
  or (_01793_, _01792_, _01776_);
  and (_01794_, _01793_, _00083_);
  or (_01795_, _00027_, rst);
  nor (_01796_, _01795_, _00091_);
  and (_02677_, _01796_, _01794_);
  nand (_01797_, _00091_, _07040_);
  and (_01798_, _00353_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_01799_, _00052_, _00070_);
  nand (_01801_, _01799_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_01802_, _01799_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_01804_, _01802_, _01801_);
  or (_01805_, _01804_, _01798_);
  or (_01806_, _01805_, _00027_);
  or (_01807_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_01808_, _01807_, _01806_);
  or (_01809_, _01808_, _00091_);
  and (_01810_, _01809_, _06989_);
  and (_02680_, _01810_, _01797_);
  not (_01811_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_01812_, _00040_, _01811_);
  or (_01813_, _01812_, _01782_);
  and (_01814_, _01813_, _00051_);
  and (_01815_, _00105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01816_, _01815_, _01812_);
  and (_01818_, _01816_, _00061_);
  or (_01819_, _01812_, _00071_);
  and (_01820_, _01819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_01822_, _01820_, _01818_);
  or (_01824_, _01822_, _01814_);
  and (_02683_, _01824_, _01796_);
  not (_01826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_01827_, _00397_, _01826_);
  and (_01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_01829_, _01828_, _00419_);
  or (_01830_, _01829_, _01827_);
  and (_01831_, _01830_, _00410_);
  nand (_01832_, _00397_, _00533_);
  and (_01833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_01834_, _01833_, _01832_);
  or (_01836_, _01834_, _00539_);
  and (_01837_, _01828_, _00406_);
  or (_01838_, _01837_, _01827_);
  and (_01839_, _01838_, _00384_);
  or (_01840_, _01839_, _01836_);
  or (_01841_, _01840_, _01831_);
  and (_01842_, _00430_, _06989_);
  and (_02684_, _01842_, _01841_);
  and (_02689_, t0_i, _06989_);
  nor (_01843_, _00382_, _07040_);
  and (_01844_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_01845_, _00407_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_01846_, _00407_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_01847_, _01846_, _01845_);
  and (_01848_, _01847_, _00384_);
  and (_01849_, _00422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_01850_, _00420_, _00410_);
  nor (_01851_, _01850_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_01852_, _01851_, _01849_);
  or (_01853_, _01852_, _01848_);
  and (_01854_, _01853_, _00430_);
  or (_01855_, _01854_, _01844_);
  or (_01856_, _01855_, _01843_);
  and (_02692_, _01856_, _06989_);
  or (_01857_, _00549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_01858_, _00535_, _00439_);
  and (_01859_, _01858_, _01857_);
  and (_01861_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_01862_, _01861_, _01859_);
  and (_01863_, _01862_, _00430_);
  not (_01864_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or (_01866_, _00429_, _01864_);
  nor (_01867_, _01866_, _00543_);
  or (_01868_, _01867_, _01863_);
  nor (_01869_, _00594_, _07040_);
  or (_01871_, _01869_, _01868_);
  and (_02695_, _01871_, _06989_);
  and (_02698_, t1_i, _06989_);
  nand (_01872_, _14012_, _11529_);
  or (_01873_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_01874_, _01873_, _06989_);
  and (_02703_, _01874_, _01872_);
  nand (_01875_, _14012_, _09008_);
  or (_01876_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_01877_, _01876_, _06989_);
  and (_02705_, _01877_, _01875_);
  nand (_01878_, _14012_, _09598_);
  or (_01879_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_01880_, _01879_, _06989_);
  and (_02723_, _01880_, _01878_);
  nand (_01881_, _12937_, _07040_);
  or (_01882_, _12937_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_01883_, _01882_, _06989_);
  and (_02737_, _01883_, _01881_);
  or (_01884_, _01319_, _11966_);
  not (_01885_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_01886_, _01319_, _01885_);
  and (_01887_, _01886_, _06983_);
  and (_01888_, _01887_, _01884_);
  nor (_01889_, _06484_, _01885_);
  and (_01890_, _01318_, _14196_);
  nand (_01891_, _01890_, _06968_);
  or (_01892_, _01890_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01893_, _01892_, _06485_);
  and (_01894_, _01893_, _01891_);
  or (_01895_, _01894_, _01889_);
  or (_01897_, _01895_, _01888_);
  and (_02756_, _01897_, _06989_);
  not (_01898_, _09227_);
  or (_01899_, _01319_, _01898_);
  not (_01900_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_01901_, _01319_, _01900_);
  and (_01902_, _01901_, _06983_);
  and (_01903_, _01902_, _01899_);
  nor (_01904_, _06484_, _01900_);
  nand (_01905_, _01318_, _00764_);
  and (_01906_, _01905_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_01907_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_01908_, _01907_, _00760_);
  and (_01909_, _01908_, _01318_);
  or (_01910_, _01909_, _01906_);
  and (_01911_, _01910_, _06485_);
  or (_01912_, _01911_, _01904_);
  or (_01913_, _01912_, _01903_);
  and (_02759_, _01913_, _06989_);
  or (_01914_, _01319_, _08030_);
  not (_01915_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_01916_, _01319_, _01915_);
  and (_01917_, _01916_, _06983_);
  and (_01918_, _01917_, _01914_);
  nor (_01919_, _06484_, _01915_);
  and (_01920_, _01318_, _07089_);
  nand (_01921_, _01920_, _06968_);
  or (_01922_, _01920_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_01923_, _01922_, _06485_);
  and (_01924_, _01923_, _01921_);
  or (_01925_, _01924_, _01919_);
  or (_01926_, _01925_, _01918_);
  and (_02805_, _01926_, _06989_);
  and (_01927_, _01156_, _07089_);
  nand (_01928_, _01927_, _06968_);
  or (_01929_, _01927_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_01930_, _01929_, _06485_);
  and (_01931_, _01930_, _01928_);
  nor (_01932_, _01163_, _09008_);
  and (_01933_, _01163_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_01934_, _01933_, _01932_);
  and (_01935_, _01934_, _06983_);
  and (_01936_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_01937_, _01936_, rst);
  or (_01938_, _01937_, _01935_);
  or (_02899_, _01938_, _01931_);
  and (_01939_, _01156_, _07048_);
  nand (_01940_, _01939_, _06968_);
  or (_01941_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_01942_, _01941_, _06485_);
  and (_01943_, _01942_, _01940_);
  nor (_01944_, _01163_, _07118_);
  nor (_01945_, _01162_, _01301_);
  or (_01946_, _01945_, _01944_);
  and (_01947_, _01946_, _06983_);
  nor (_01948_, _06484_, _01301_);
  or (_01949_, _01948_, rst);
  or (_01950_, _01949_, _01947_);
  or (_02900_, _01950_, _01943_);
  and (_01951_, _09023_, _07089_);
  nand (_01952_, _01951_, _06968_);
  or (_01953_, _01951_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_01954_, _01953_, _06485_);
  and (_01955_, _01954_, _01952_);
  nor (_01956_, _09031_, _09008_);
  and (_01957_, _09031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_01958_, _01957_, _01956_);
  and (_01959_, _01958_, _06983_);
  and (_01960_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_01961_, _01960_, rst);
  or (_01962_, _01961_, _01959_);
  or (_02903_, _01962_, _01955_);
  and (_01963_, _09023_, _07048_);
  nand (_01964_, _01963_, _06968_);
  or (_01965_, _01963_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_01966_, _01965_, _06485_);
  and (_01967_, _01966_, _01964_);
  nor (_01968_, _09031_, _07118_);
  and (_01969_, _09031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_01970_, _01969_, _01968_);
  and (_01971_, _01970_, _06983_);
  and (_01972_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_01973_, _01972_, rst);
  or (_01974_, _01973_, _01971_);
  or (_02905_, _01974_, _01967_);
  and (_01975_, _00691_, _09074_);
  nand (_01976_, _01975_, _06968_);
  or (_01977_, _01975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_01978_, _01977_, _06485_);
  and (_01979_, _01978_, _01976_);
  nand (_01980_, _11529_, _00697_);
  or (_01981_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_01982_, _01981_, _06983_);
  and (_01983_, _01982_, _01980_);
  nor (_01984_, _06484_, _14532_);
  or (_01985_, _01984_, rst);
  or (_01986_, _01985_, _01983_);
  or (_02907_, _01986_, _01979_);
  and (_01987_, _00720_, _07048_);
  nand (_01988_, _01987_, _06968_);
  or (_01989_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01990_, _01989_, _06485_);
  and (_01991_, _01990_, _01988_);
  nand (_01992_, _00726_, _07118_);
  or (_01993_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01994_, _01993_, _06983_);
  and (_01995_, _01994_, _01992_);
  nor (_01996_, _06484_, _01286_);
  or (_01997_, _01996_, rst);
  or (_01998_, _01997_, _01995_);
  or (_02909_, _01998_, _01991_);
  and (_01999_, _00720_, _07089_);
  nand (_02000_, _01999_, _06968_);
  or (_02002_, _01999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_02003_, _02002_, _06485_);
  and (_02004_, _02003_, _02000_);
  nand (_02005_, _00726_, _09008_);
  or (_02006_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_02007_, _02006_, _06983_);
  and (_02008_, _02007_, _02005_);
  and (_02009_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_02010_, _02009_, rst);
  or (_02011_, _02010_, _02008_);
  or (_02911_, _02011_, _02004_);
  and (_02012_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_02013_, _08139_, _01227_);
  or (_02014_, _02013_, _02012_);
  and (_02922_, _02014_, _06989_);
  nand (_02015_, _01162_, _06968_);
  or (_02016_, _01162_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_02017_, _02016_, _06485_);
  and (_02018_, _02017_, _02015_);
  and (_02019_, _01162_, _09599_);
  nor (_02020_, _01162_, _01533_);
  or (_02021_, _02020_, _02019_);
  and (_02022_, _02021_, _06983_);
  nor (_02023_, _06484_, _01533_);
  or (_02025_, _02023_, rst);
  or (_02026_, _02025_, _02022_);
  or (_02928_, _02026_, _02018_);
  and (_02027_, _01156_, _08436_);
  nand (_02028_, _02027_, _06968_);
  or (_02029_, _02027_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_02030_, _02029_, _06485_);
  and (_02031_, _02030_, _02028_);
  nor (_02032_, _01163_, _07317_);
  and (_02033_, _01163_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_02034_, _02033_, _02032_);
  and (_02035_, _02034_, _06983_);
  and (_02036_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_02037_, _02036_, rst);
  or (_02038_, _02037_, _02035_);
  or (_02930_, _02038_, _02031_);
  and (_02039_, _00691_, _14196_);
  nand (_02040_, _02039_, _06968_);
  or (_02041_, _02039_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_02042_, _02041_, _06485_);
  and (_02043_, _02042_, _02040_);
  nand (_02044_, _10970_, _00697_);
  or (_02045_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_02046_, _02045_, _06983_);
  and (_02047_, _02046_, _02044_);
  and (_02048_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_02049_, _02048_, rst);
  or (_02050_, _02049_, _02047_);
  or (_02933_, _02050_, _02043_);
  and (_02051_, _00691_, _06979_);
  nand (_02052_, _02051_, _06968_);
  or (_02053_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_02054_, _02053_, _06485_);
  and (_02055_, _02054_, _02052_);
  nand (_02057_, _09598_, _00697_);
  and (_02059_, _02053_, _06983_);
  and (_02060_, _02059_, _02057_);
  nor (_02061_, _06484_, _01544_);
  or (_02062_, _02061_, rst);
  or (_02063_, _02062_, _02060_);
  or (_02935_, _02063_, _02055_);
  or (_02064_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_02065_, _02064_, _06485_);
  and (_02066_, _00720_, _06979_);
  nand (_02067_, _02066_, _06968_);
  and (_02068_, _02067_, _02065_);
  nand (_02069_, _09598_, _00726_);
  and (_02070_, _02064_, _06983_);
  and (_02071_, _02070_, _02069_);
  nor (_02072_, _06484_, _01539_);
  or (_02073_, _02072_, rst);
  or (_02074_, _02073_, _02071_);
  or (_02937_, _02074_, _02068_);
  nand (_02075_, _00720_, _06525_);
  and (_02076_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_02077_, _00764_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_02078_, _02077_, _08437_);
  and (_02079_, _02078_, _00720_);
  or (_02080_, _02079_, _02076_);
  and (_02081_, _02080_, _06485_);
  nand (_02082_, _00726_, _07317_);
  or (_02083_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_02084_, _02083_, _06983_);
  and (_02085_, _02084_, _02082_);
  and (_02086_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_02087_, _02086_, rst);
  or (_02088_, _02087_, _02085_);
  or (_02939_, _02088_, _02081_);
  and (_02089_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_02090_, _08139_, _01144_);
  or (_02091_, _02090_, _02089_);
  and (_02962_, _02091_, _06989_);
  and (_02092_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_02093_, _08139_, _01149_);
  or (_02094_, _02093_, _02092_);
  and (_02965_, _02094_, _06989_);
  and (_03047_, _01586_, _06989_);
  and (_02095_, _00691_, _07048_);
  nand (_02096_, _02095_, _06968_);
  or (_02097_, _02095_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_02098_, _02097_, _06485_);
  and (_02099_, _02098_, _02096_);
  nand (_02101_, _00697_, _07118_);
  or (_02102_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_02103_, _02102_, _06983_);
  and (_02104_, _02103_, _02101_);
  nor (_02105_, _06484_, _01291_);
  or (_02106_, _02105_, rst);
  or (_02107_, _02106_, _02104_);
  or (_03053_, _02107_, _02099_);
  and (_02108_, _00691_, _07044_);
  nand (_02109_, _02108_, _06968_);
  or (_02110_, _02108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_02111_, _02110_, _06485_);
  and (_02112_, _02111_, _02109_);
  nand (_02113_, _00697_, _07260_);
  or (_02114_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_02115_, _02114_, _06983_);
  and (_02116_, _02115_, _02113_);
  nor (_02117_, _06484_, _01455_);
  or (_02118_, _02117_, rst);
  or (_02119_, _02118_, _02116_);
  or (_03055_, _02119_, _02112_);
  and (_02120_, _09023_, _07044_);
  nand (_02121_, _02120_, _06968_);
  or (_02122_, _02120_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_02123_, _02122_, _06485_);
  and (_02124_, _02123_, _02121_);
  nor (_02125_, _09031_, _07260_);
  nor (_02126_, _09030_, _01471_);
  or (_02127_, _02126_, _02125_);
  and (_02128_, _02127_, _06983_);
  nor (_02129_, _06484_, _01471_);
  or (_02130_, _02129_, rst);
  or (_02131_, _02130_, _02128_);
  or (_03057_, _02131_, _02124_);
  and (_02132_, _09023_, _08436_);
  nand (_02133_, _02132_, _06968_);
  or (_02134_, _02132_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_02135_, _02134_, _06485_);
  and (_02136_, _02135_, _02133_);
  nor (_02137_, _09031_, _07317_);
  and (_02138_, _09031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_02139_, _02138_, _02137_);
  and (_02140_, _02139_, _06983_);
  and (_02141_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_02142_, _02141_, rst);
  or (_02143_, _02142_, _02140_);
  or (_03058_, _02143_, _02136_);
  nand (_02144_, _12937_, _09598_);
  or (_02145_, _12937_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_02146_, _02145_, _02144_);
  and (_03072_, _02146_, _06989_);
  and (_02147_, _00720_, _14196_);
  nand (_02148_, _02147_, _06968_);
  or (_02149_, _02147_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02150_, _02149_, _06485_);
  and (_02151_, _02150_, _02148_);
  nand (_02152_, _10970_, _00726_);
  or (_02153_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02154_, _02153_, _06983_);
  and (_02155_, _02154_, _02152_);
  and (_02156_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_02157_, _02156_, rst);
  or (_02158_, _02157_, _02155_);
  or (_03077_, _02158_, _02151_);
  and (_02159_, _00720_, _07044_);
  nand (_02160_, _02159_, _06968_);
  or (_02161_, _02159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02162_, _02161_, _06485_);
  and (_02163_, _02162_, _02160_);
  nand (_02164_, _00726_, _07260_);
  or (_02165_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02166_, _02165_, _06983_);
  and (_02167_, _02166_, _02164_);
  nor (_02168_, _06484_, _01460_);
  or (_02169_, _02168_, rst);
  or (_02170_, _02169_, _02167_);
  or (_03079_, _02170_, _02163_);
  nand (_02171_, _00720_, _00764_);
  and (_02172_, _02171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02173_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_02174_, _02173_, _00760_);
  and (_02175_, _02174_, _00720_);
  or (_02176_, _02175_, _02172_);
  and (_02177_, _02176_, _06485_);
  nand (_02178_, _11529_, _00726_);
  or (_02179_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02180_, _02179_, _06983_);
  and (_02181_, _02180_, _02178_);
  nor (_02182_, _06484_, _14527_);
  or (_02183_, _02182_, rst);
  or (_02184_, _02183_, _02181_);
  or (_03081_, _02184_, _02177_);
  and (_02186_, _00691_, _08436_);
  nand (_02187_, _02186_, _06968_);
  or (_02188_, _02186_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02189_, _02188_, _06485_);
  and (_02190_, _02189_, _02187_);
  nand (_02191_, _00697_, _07317_);
  or (_02192_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02193_, _02192_, _06983_);
  and (_02194_, _02193_, _02191_);
  and (_02195_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_02196_, _02195_, rst);
  or (_02197_, _02196_, _02194_);
  or (_03083_, _02197_, _02190_);
  and (_02198_, _09023_, _14196_);
  nand (_02199_, _02198_, _06968_);
  or (_02200_, _02198_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_02201_, _02200_, _06485_);
  and (_02202_, _02201_, _02199_);
  nor (_02203_, _10970_, _09031_);
  and (_02204_, _09031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02205_, _02204_, _02203_);
  and (_02206_, _02205_, _06983_);
  and (_02207_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02208_, _02207_, rst);
  or (_02209_, _02208_, _02206_);
  or (_03085_, _02209_, _02202_);
  and (_02210_, _00691_, _07089_);
  nand (_02211_, _02210_, _06968_);
  or (_02213_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_02214_, _02213_, _06485_);
  and (_02215_, _02214_, _02211_);
  nand (_02216_, _00697_, _09008_);
  or (_02217_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_02218_, _02217_, _06983_);
  and (_02219_, _02218_, _02216_);
  and (_02220_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_02221_, _02220_, rst);
  or (_02222_, _02221_, _02219_);
  or (_03087_, _02222_, _02215_);
  and (_02223_, _09023_, _09074_);
  nand (_02224_, _02223_, _06968_);
  or (_02226_, _02223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_02227_, _02226_, _06485_);
  and (_02228_, _02227_, _02224_);
  nor (_02229_, _11529_, _09031_);
  and (_02230_, _09031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02231_, _02230_, _02229_);
  and (_02232_, _02231_, _06983_);
  and (_02233_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02234_, _02233_, rst);
  or (_02235_, _02234_, _02232_);
  or (_03089_, _02235_, _02228_);
  nand (_02236_, _09030_, _06968_);
  or (_02237_, _09030_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_02238_, _02237_, _06485_);
  and (_02239_, _02238_, _02236_);
  and (_02240_, _09599_, _09030_);
  nor (_02241_, _09030_, _01528_);
  or (_02242_, _02241_, _02240_);
  and (_02243_, _02242_, _06983_);
  nor (_02244_, _06484_, _01528_);
  or (_02245_, _02244_, rst);
  or (_02246_, _02245_, _02243_);
  or (_03091_, _02246_, _02239_);
  and (_02247_, _01156_, _14196_);
  nand (_02248_, _02247_, _06968_);
  or (_02249_, _02247_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_02250_, _02249_, _06485_);
  and (_02251_, _02250_, _02248_);
  nor (_02252_, _01163_, _10970_);
  and (_02253_, _01163_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_02254_, _02253_, _02252_);
  and (_02255_, _02254_, _06983_);
  and (_02256_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_02257_, _02256_, rst);
  or (_02258_, _02257_, _02255_);
  or (_03093_, _02258_, _02251_);
  and (_02259_, _01156_, _07044_);
  nand (_02260_, _02259_, _06968_);
  or (_02261_, _02259_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_02262_, _02261_, _06485_);
  and (_02263_, _02262_, _02260_);
  nor (_02264_, _01163_, _07260_);
  nor (_02265_, _01162_, _01466_);
  or (_02266_, _02265_, _02264_);
  and (_02267_, _02266_, _06983_);
  nor (_02268_, _06484_, _01466_);
  or (_02269_, _02268_, rst);
  or (_02270_, _02269_, _02267_);
  or (_03095_, _02270_, _02263_);
  and (_02271_, _01156_, _09074_);
  nand (_02272_, _02271_, _06968_);
  or (_02273_, _02271_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_02274_, _02273_, _06485_);
  and (_02275_, _02274_, _02272_);
  nor (_02276_, _01163_, _11529_);
  nor (_02277_, _01162_, _14538_);
  or (_02278_, _02277_, _02276_);
  and (_02279_, _02278_, _06983_);
  nor (_02280_, _06484_, _14538_);
  or (_02281_, _02280_, rst);
  or (_02282_, _02281_, _02279_);
  or (_03098_, _02282_, _02275_);
  and (_02283_, _11954_, _07048_);
  or (_02285_, _02283_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_02287_, _02285_, _07292_);
  nand (_02288_, _02283_, _06968_);
  and (_02289_, _02288_, _02287_);
  nor (_02290_, _07292_, _07118_);
  or (_02291_, _02290_, _02289_);
  and (_03127_, _02291_, _06989_);
  and (_03135_, _01367_, _06989_);
  and (_03420_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _06989_);
  and (_02292_, _03420_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_03146_, _02292_, _03135_);
  or (_02293_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand (_02295_, _07493_, _14110_);
  and (_02296_, _02295_, _06989_);
  and (_03150_, _02296_, _02293_);
  nand (_02298_, _07321_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_03156_, _02298_, _06989_);
  nand (_02299_, _11951_, _06968_);
  nor (_02301_, _11951_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_02302_, _02301_, _11954_);
  and (_02303_, _02302_, _02299_);
  or (_02304_, _02303_, _07291_);
  and (_02305_, _06540_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_02306_, _02305_, _06969_);
  and (_02307_, _02306_, _11954_);
  or (_02308_, _02307_, _02304_);
  nand (_02309_, _07291_, _07040_);
  and (_02310_, _02309_, _06989_);
  and (_03209_, _02310_, _02308_);
  and (_03313_, _08080_, _06989_);
  nor (_02311_, _07493_, _07490_);
  nor (_02312_, _01213_, _01210_);
  nor (_02313_, _02312_, _07490_);
  and (_02314_, _02313_, _07331_);
  nor (_02315_, _02313_, _07331_);
  nor (_02316_, _02315_, _02314_);
  nor (_02317_, _02316_, _02311_);
  and (_02318_, _07350_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_02319_, _02318_, _02311_);
  nor (_02320_, _02319_, _10959_);
  or (_02321_, _02320_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02322_, _02321_, _02317_);
  and (_03315_, _02322_, _06989_);
  nor (_02323_, _12938_, _07260_);
  and (_02324_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or (_02325_, _02324_, _02323_);
  and (_03327_, _02325_, _06989_);
  and (_02326_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_02327_, _02326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_03329_, _02327_, _06989_);
  nor (_02328_, _12829_, rst);
  not (_02329_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nand (_02330_, _07325_, _02329_);
  and (_03350_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _06989_);
  and (_02331_, _03350_, _02330_);
  or (_03331_, _02331_, _02328_);
  and (_02332_, _14190_, _09599_);
  and (_02333_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or (_02334_, _02333_, _02332_);
  and (_03345_, _02334_, _06989_);
  and (_02335_, _14146_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_02336_, _14146_, _07260_);
  or (_02337_, _02336_, _02335_);
  and (_03354_, _02337_, _06989_);
  and (_02338_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_02339_, _14190_, _09009_);
  or (_02340_, _02339_, _02338_);
  and (_03364_, _02340_, _06989_);
  nor (_02341_, _11042_, _11040_);
  nor (_02342_, _02341_, _11043_);
  or (_02343_, _02342_, _08477_);
  or (_02344_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_02345_, _02344_, _10964_);
  and (_02346_, _02345_, _02343_);
  and (_02347_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_03372_, _02347_, _02346_);
  nor (_02348_, _11037_, _11035_);
  nor (_02349_, _02348_, _11038_);
  or (_02350_, _02349_, _08477_);
  or (_02351_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_02352_, _02351_, _10964_);
  and (_02353_, _02352_, _02350_);
  and (_02354_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_03374_, _02354_, _02353_);
  nor (_02355_, _11034_, _11032_);
  nor (_02356_, _02355_, _11035_);
  or (_02357_, _02356_, _08477_);
  or (_02358_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_02359_, _02358_, _10964_);
  and (_02360_, _02359_, _02357_);
  and (_02361_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_03399_, _02361_, _02360_);
  not (_02362_, _00653_);
  and (_02363_, _02362_, _00651_);
  and (_02364_, _00256_, _00645_);
  and (_03413_, _02364_, _02363_);
  nor (_02365_, _13944_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_02366_, _02365_, _13945_);
  and (_03422_, _02366_, _13953_);
  and (_02367_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _08578_);
  and (_02368_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_02369_, _02368_, _02367_);
  and (_03428_, _02369_, _06989_);
  and (_02370_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_02371_, _14190_, _07119_);
  or (_02372_, _02371_, _02370_);
  and (_03439_, _02372_, _06989_);
  and (_02373_, _08525_, _08459_);
  and (_02374_, _02373_, _08557_);
  not (_02375_, _08542_);
  and (_02376_, _02375_, _08509_);
  and (_02377_, _02376_, _08572_);
  and (_02378_, _07326_, _06989_);
  and (_02379_, _02378_, _08492_);
  and (_02380_, _02379_, _07356_);
  and (_02381_, _02380_, _02377_);
  and (_03444_, _02381_, _02374_);
  and (_02382_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor (_02383_, _10970_, _07486_);
  or (_02384_, _02383_, _02382_);
  and (_03447_, _02384_, _06989_);
  and (_03456_, _11518_, _06989_);
  and (_03475_, _11605_, _06989_);
  and (_02385_, _14058_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02386_, _09763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_02387_, _02386_, _14057_);
  or (_02388_, _02387_, _02385_);
  and (_03479_, _02388_, _06989_);
  and (_02389_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or (_02390_, _00909_, _07278_);
  nand (_02391_, _07209_, _07166_);
  or (_02392_, _02391_, _07196_);
  and (_02393_, _02392_, _02390_);
  or (_02394_, _02393_, _02389_);
  and (_02395_, _07271_, _07269_);
  or (_02396_, _02395_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_02397_, _07470_, rst);
  and (_02398_, _02397_, _02396_);
  and (_03486_, _02398_, _02394_);
  or (_02399_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  nand (_02400_, _07493_, _11224_);
  and (_02401_, _02400_, _06989_);
  and (_03489_, _02401_, _02399_);
  and (_02402_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_02403_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or (_02404_, _02403_, _02402_);
  and (_03512_, _02404_, _06989_);
  and (_02405_, _11908_, _11359_);
  and (_02406_, _11911_, _11364_);
  and (_02407_, _11359_, _11287_);
  or (_02408_, _02407_, _02406_);
  and (_02409_, _11911_, _11306_);
  or (_02410_, _02409_, _11405_);
  or (_02411_, _02410_, _02408_);
  or (_02412_, _02411_, _02405_);
  and (_02413_, _11339_, _11313_);
  and (_02414_, _11332_, _11430_);
  or (_02415_, _02414_, _11435_);
  or (_02416_, _02415_, _02413_);
  or (_02417_, _11332_, _11478_);
  and (_02418_, _02417_, _11389_);
  and (_02419_, _11354_, _11290_);
  or (_02420_, _02419_, _02418_);
  or (_02421_, _02420_, _02416_);
  and (_02422_, _11908_, _11451_);
  and (_02423_, _11908_, _11313_);
  or (_02424_, _02423_, _02422_);
  or (_02425_, _02424_, _11385_);
  and (_02426_, _11430_, _11287_);
  or (_02427_, _02426_, _11468_);
  or (_02428_, _02427_, _11404_);
  or (_02429_, _02428_, _02425_);
  or (_02430_, _02429_, _02421_);
  and (_02431_, _11332_, _11472_);
  and (_02432_, _11332_, _11356_);
  and (_02433_, _11332_, _11375_);
  or (_02434_, _02433_, _02432_);
  or (_02435_, _02434_, _02431_);
  or (_02436_, _14313_, _11320_);
  and (_02437_, _11332_, _11324_);
  or (_02438_, _02437_, _14317_);
  not (_02439_, _11397_);
  nand (_02440_, _02439_, _11391_);
  or (_02441_, _02440_, _02438_);
  or (_02442_, _02441_, _02436_);
  or (_02443_, _02442_, _02435_);
  or (_02444_, _02443_, _02430_);
  or (_02445_, _02444_, _02412_);
  and (_02446_, _02445_, _07325_);
  and (_02447_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_02448_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_02449_, _11353_, _02448_);
  and (_02450_, _11290_, _11306_);
  not (_02451_, _11467_);
  nor (_02452_, _11339_, _11289_);
  nor (_02453_, _02452_, _02451_);
  nor (_02454_, _02453_, _02450_);
  not (_02455_, _02454_);
  and (_02456_, _02455_, _02449_);
  or (_02457_, _02456_, _02447_);
  or (_02458_, _02457_, _02446_);
  and (_03518_, _02458_, _06989_);
  and (_02459_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_02460_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  or (_02461_, _02460_, _02459_);
  and (_03521_, _02461_, _06989_);
  nor (_03539_, _11579_, rst);
  and (_02462_, \oc8051_top_1.oc8051_sfr1.wait_data , _06989_);
  and (_02463_, _02462_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_02464_, _02422_, _07383_);
  and (_02465_, _11925_, _11382_);
  or (_02466_, _02465_, _02464_);
  and (_02467_, _11478_, _11373_);
  or (_02468_, _02467_, _14317_);
  or (_02469_, _11467_, _11359_);
  and (_02470_, _02469_, _11332_);
  or (_02471_, _02470_, _02468_);
  or (_02472_, _02471_, _02466_);
  or (_02473_, _14320_, _11395_);
  and (_02474_, _02450_, _11316_);
  or (_02475_, _02474_, _02473_);
  and (_02476_, _14313_, _07383_);
  and (_02477_, _02423_, _07383_);
  or (_02478_, _02477_, _02476_);
  or (_02479_, _02478_, _02475_);
  and (_02480_, _11332_, _11399_);
  or (_02481_, _11919_, _02480_);
  nor (_02482_, _02481_, _11400_);
  nand (_02483_, _02482_, _11454_);
  or (_02484_, _02483_, _02416_);
  or (_02485_, _02484_, _02479_);
  or (_02486_, _02485_, _02472_);
  and (_02487_, _07325_, _06989_);
  and (_02488_, _02487_, _02486_);
  or (_03541_, _02488_, _02463_);
  nor (_03549_, _07294_, rst);
  and (_02489_, _11358_, _11342_);
  not (_02490_, _11335_);
  and (_02491_, _02490_, _02449_);
  and (_02492_, _11941_, _11312_);
  and (_02493_, _11940_, _11312_);
  or (_02494_, _02493_, _02492_);
  and (_02495_, _02494_, _11342_);
  or (_02496_, _02495_, _02491_);
  or (_02497_, _02496_, _02489_);
  and (_02498_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_02499_, _11478_, _11306_);
  or (_02500_, _02499_, _11456_);
  and (_02501_, _11925_, _11289_);
  or (_02502_, _02501_, _11449_);
  or (_02503_, _11473_, _11425_);
  or (_02504_, _02503_, _02492_);
  or (_02505_, _02504_, _02502_);
  and (_02506_, _11469_, _11388_);
  or (_02507_, _11461_, _11453_);
  or (_02508_, _02507_, _02506_);
  nor (_02509_, _11477_, _11423_);
  nand (_02510_, _02509_, _11440_);
  or (_02511_, _02510_, _02508_);
  or (_02512_, _02511_, _02505_);
  or (_02513_, _02493_, _11380_);
  or (_02514_, _02513_, _02512_);
  or (_02515_, _02514_, _02500_);
  and (_02516_, _02515_, _07325_);
  or (_02517_, _02516_, _02498_);
  or (_02518_, _02517_, _02497_);
  and (_03557_, _02518_, _06989_);
  and (_02519_, _06894_, _06845_);
  and (_02520_, _06790_, _06548_);
  and (_02521_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand (_02522_, _06951_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_02523_, _02522_, _02521_);
  or (_02524_, _02523_, _02520_);
  or (_02525_, _02524_, _02519_);
  nor (_02526_, _02521_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_02527_, _02526_, _11954_);
  and (_02528_, _02527_, _02525_);
  or (_02529_, _02528_, _07291_);
  nor (_02530_, _14196_, _08412_);
  or (_02531_, _02530_, _01556_);
  and (_02532_, _02531_, _11954_);
  or (_02533_, _02532_, _02529_);
  nand (_02534_, _10970_, _07291_);
  and (_02535_, _02534_, _06989_);
  and (_03561_, _02535_, _02533_);
  and (_02536_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02537_, _02536_, _02496_);
  nor (_02538_, _11942_, _11316_);
  and (_02539_, _11477_, _11316_);
  and (_02540_, _11394_, _11319_);
  and (_02541_, _11396_, _11388_);
  or (_02543_, _02541_, _11401_);
  or (_02544_, _02543_, _02540_);
  or (_02545_, _02544_, _02539_);
  or (_02546_, _02545_, _11395_);
  or (_02547_, _02546_, _02538_);
  and (_02548_, _02547_, _07325_);
  or (_02549_, _02548_, _02537_);
  and (_03566_, _02549_, _06989_);
  and (_02550_, _11332_, _11451_);
  or (_02551_, _02550_, _02414_);
  or (_02552_, _02408_, _02419_);
  and (_02553_, _11389_, _11312_);
  and (_02554_, _02553_, _11422_);
  or (_02555_, _02541_, _02493_);
  or (_02556_, _02555_, _02554_);
  and (_02557_, _11403_, _11382_);
  or (_02558_, _02437_, _02557_);
  or (_02559_, _02558_, _02556_);
  or (_02560_, _02559_, _02552_);
  or (_02561_, _02560_, _02551_);
  or (_02562_, _02410_, _11404_);
  and (_02564_, _11911_, _11388_);
  or (_02565_, _11397_, _11325_);
  or (_02566_, _02565_, _02564_);
  and (_02567_, _11356_, _11382_);
  and (_02568_, _11908_, _11927_);
  or (_02569_, _02568_, _02567_);
  or (_02570_, _02569_, _02566_);
  or (_02571_, _02570_, _02562_);
  or (_02572_, _02571_, _02561_);
  and (_02573_, _11332_, _11438_);
  or (_02574_, _02573_, _02423_);
  and (_02575_, _11359_, _11312_);
  and (_02577_, _02575_, _11908_);
  or (_02579_, _02577_, _14313_);
  or (_02580_, _02579_, _02574_);
  and (_02581_, _11332_, _11467_);
  or (_02582_, _02581_, _11909_);
  and (_02583_, _02553_, _11332_);
  or (_02584_, _02583_, _11333_);
  or (_02585_, _02584_, _02582_);
  or (_02586_, _02585_, _02435_);
  or (_02587_, _02450_, _11334_);
  or (_02588_, _02587_, _02586_);
  or (_02589_, _02588_, _02580_);
  or (_02590_, _02589_, _02572_);
  and (_02591_, _02590_, _07325_);
  and (_02592_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_02593_, _02456_, _11347_);
  or (_02594_, _02593_, _02592_);
  or (_02595_, _02594_, _02591_);
  and (_03579_, _02595_, _06989_);
  or (_02596_, _02553_, _11324_);
  and (_02598_, _02596_, _11422_);
  or (_02599_, _02565_, _02598_);
  and (_02600_, _11451_, _11290_);
  and (_02601_, _11430_, _11290_);
  or (_02602_, _02601_, _02600_);
  or (_02603_, _02602_, _11456_);
  or (_02604_, _02603_, _02599_);
  and (_02605_, _02541_, _11299_);
  or (_02606_, _02605_, _02413_);
  and (_02607_, _02553_, _11287_);
  or (_02608_, _02607_, _02606_);
  or (_02609_, _11334_, _11314_);
  or (_02610_, _02609_, _02562_);
  or (_02611_, _02610_, _02608_);
  or (_02612_, _02611_, _02604_);
  or (_02613_, _02574_, _11447_);
  or (_02614_, _02613_, _02586_);
  or (_02615_, _02614_, _02612_);
  or (_02616_, _02615_, _02552_);
  and (_02617_, _02616_, _07325_);
  and (_02618_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or (_02619_, _02618_, _02593_);
  or (_02620_, _02619_, _02617_);
  and (_03598_, _02620_, _06989_);
  nand (_02621_, _01555_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_02623_, _02621_, _06501_);
  or (_02624_, _02623_, _01556_);
  not (_02625_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_02626_, _07075_, _02625_);
  or (_02627_, _02626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_02628_, _02627_, _06501_);
  and (_02629_, _02628_, _02624_);
  or (_02630_, _02629_, _06987_);
  nand (_02631_, _10970_, _06987_);
  and (_02632_, _02631_, _06989_);
  and (_03617_, _02632_, _02630_);
  and (_02633_, _07048_, _06501_);
  nand (_02634_, _02633_, _06968_);
  not (_02635_, _06987_);
  or (_02636_, _02633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_02637_, _02636_, _02635_);
  and (_02638_, _02637_, _02634_);
  nor (_02639_, _07118_, _02635_);
  or (_02640_, _02639_, _02638_);
  and (_03619_, _02640_, _06989_);
  and (_02641_, _07044_, _06501_);
  nand (_02642_, _02641_, _06968_);
  or (_02643_, _02641_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_02644_, _02643_, _02635_);
  and (_02645_, _02644_, _02642_);
  nor (_02646_, _07260_, _02635_);
  or (_02647_, _02646_, _02645_);
  and (_03622_, _02647_, _06989_);
  nor (_03634_, _11349_, rst);
  nand (_02648_, _02487_, _11389_);
  or (_03636_, _02648_, _02452_);
  and (_02649_, _10851_, _10812_);
  and (_02651_, _10841_, _10834_);
  and (_02652_, _10824_, _10854_);
  and (_02653_, _10917_, _02652_);
  or (_02654_, _02653_, _02651_);
  or (_02655_, _02654_, _02649_);
  or (_02656_, _10904_, _10860_);
  and (_02657_, _10917_, _10818_);
  and (_02658_, _10870_, _10851_);
  or (_02659_, _02658_, _02657_);
  or (_02660_, _02659_, _02656_);
  nor (_02661_, _02660_, _02655_);
  nand (_02662_, _02661_, _10941_);
  and (_02663_, _10871_, _10837_);
  not (_02664_, _10906_);
  nand (_02665_, _10951_, _02664_);
  or (_02666_, _02665_, _02663_);
  or (_02667_, _10912_, _10831_);
  or (_02669_, _10828_, _10816_);
  or (_02670_, _02669_, _02667_);
  or (_02672_, _10911_, _10878_);
  or (_02673_, _02672_, _02670_);
  or (_02674_, _02673_, _02666_);
  or (_02675_, _02674_, _02662_);
  and (_02676_, _02675_, _07326_);
  and (_02678_, _07323_, _06406_);
  and (_02679_, _02678_, _11340_);
  nor (_02681_, _02679_, _02448_);
  or (_02682_, _02681_, rst);
  or (_03638_, _02682_, _02676_);
  or (_02685_, _08463_, _11345_);
  or (_02686_, _07324_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_02687_, _02686_, _06989_);
  and (_03641_, _02687_, _02685_);
  and (_02688_, _02462_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_02690_, _11375_, _11289_);
  and (_02691_, _11438_, _11290_);
  or (_02693_, _02691_, _02581_);
  or (_02694_, _02693_, _02690_);
  or (_02696_, _11439_, _11369_);
  and (_02697_, _11360_, _11316_);
  or (_02699_, _11936_, _02697_);
  or (_02700_, _02699_, _02696_);
  or (_02701_, _11913_, _11358_);
  or (_02702_, _02701_, _02474_);
  or (_02704_, _02702_, _02700_);
  or (_02706_, _02704_, _02694_);
  and (_02707_, _02706_, _02487_);
  or (_03643_, _02707_, _02688_);
  or (_02708_, _02413_, _11320_);
  and (_02709_, _11908_, _11438_);
  and (_02710_, _11478_, _11374_);
  or (_02711_, _02710_, _11395_);
  or (_02712_, _02711_, _02709_);
  or (_02713_, _02712_, _02708_);
  and (_02714_, _02713_, _07325_);
  and (_02715_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02716_, _02715_, _02491_);
  or (_02717_, _02716_, _02714_);
  and (_03645_, _02717_, _06989_);
  and (_02718_, _02462_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_02719_, _11908_, _11356_);
  or (_02720_, _02503_, _02431_);
  or (_02721_, _02720_, _02719_);
  not (_02722_, _11402_);
  and (_02724_, _11355_, _11287_);
  or (_02725_, _02724_, _11912_);
  or (_02726_, _02725_, _02722_);
  or (_02727_, _02481_, _02477_);
  or (_02728_, _02727_, _02708_);
  or (_02729_, _02728_, _02726_);
  or (_02730_, _02729_, _02721_);
  and (_02731_, _02730_, _02487_);
  or (_03648_, _02731_, _02718_);
  or (_02732_, _11052_, _11014_);
  and (_02733_, _02732_, _11053_);
  or (_02734_, _02733_, _08477_);
  or (_02735_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_02736_, _02735_, _10964_);
  and (_02738_, _02736_, _02734_);
  and (_02739_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_03651_, _02739_, _02738_);
  and (_02740_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_02741_, _11461_, _07325_);
  or (_02742_, _02741_, _02740_);
  or (_02743_, _02742_, _02491_);
  and (_03655_, _02743_, _06989_);
  or (_02744_, _02494_, _02474_);
  and (_02745_, _02744_, _11282_);
  or (_02746_, _02456_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02747_, _02746_, _02495_);
  or (_02748_, _02747_, _02745_);
  or (_02749_, _06406_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_02750_, _02749_, _06989_);
  and (_03657_, _02750_, _02748_);
  and (_02751_, _02462_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_02752_, _11355_, _11374_);
  and (_02753_, _02752_, _11911_);
  or (_02754_, _11425_, _11320_);
  or (_02755_, _02754_, _02753_);
  or (_02757_, _02690_, _02719_);
  and (_02758_, _11438_, _11394_);
  and (_02760_, _11356_, _11394_);
  or (_02761_, _02760_, _02758_);
  or (_02762_, _02761_, _02757_);
  or (_02763_, _02710_, _11437_);
  or (_02764_, _11474_, _11453_);
  or (_02765_, _02764_, _02763_);
  or (_02766_, _02765_, _02762_);
  or (_02767_, _02766_, _02755_);
  and (_02768_, _02767_, _02487_);
  or (_03659_, _02768_, _02751_);
  and (_02769_, _02462_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  not (_02770_, _11432_);
  or (_02771_, _02414_, _02770_);
  or (_02772_, _02709_, _02422_);
  or (_02773_, _02419_, _11426_);
  or (_02774_, _02773_, _02772_);
  nand (_02775_, _14306_, _11436_);
  or (_02776_, _02775_, _02774_);
  or (_02777_, _02776_, _02771_);
  or (_02778_, _02473_, _02468_);
  or (_02779_, _02778_, _02725_);
  or (_02780_, _02779_, _02721_);
  or (_02781_, _02780_, _02777_);
  and (_02782_, _02781_, _02487_);
  or (_03662_, _02782_, _02769_);
  or (_02783_, _02405_, _02407_);
  or (_02784_, _02410_, _11397_);
  or (_02785_, _02784_, _02783_);
  or (_02786_, _02785_, _02423_);
  and (_02787_, _02786_, _07325_);
  and (_02788_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02789_, _02788_, _11346_);
  or (_02790_, _02789_, _02787_);
  and (_03664_, _02790_, _06989_);
  or (_02791_, _11456_, _11380_);
  or (_02792_, _02725_, _02711_);
  or (_02793_, _02493_, _11479_);
  or (_02794_, _02793_, _02564_);
  or (_02795_, _02794_, _02792_);
  or (_02796_, _02795_, _02791_);
  or (_02797_, _02796_, _02512_);
  or (_02798_, _02797_, _02544_);
  and (_02799_, _02798_, _07325_);
  and (_02800_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02801_, _02800_, _02497_);
  or (_02802_, _02801_, _02799_);
  and (_03666_, _02802_, _06989_);
  and (_02803_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_02804_, _02803_, _09580_);
  and (_02806_, _07071_, _07054_);
  or (_02807_, _02806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand (_02808_, _07071_, _07055_);
  and (_02809_, _02808_, _02807_);
  or (_02810_, _02809_, _02804_);
  and (_02811_, _02810_, _09574_);
  and (_02812_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_02813_, _02812_, _07046_);
  or (_02814_, _02813_, _02811_);
  nand (_02815_, _07260_, _07046_);
  and (_02816_, _02815_, _09590_);
  and (_02817_, _02816_, _02814_);
  and (_02818_, _07050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_02819_, _02818_, _02817_);
  and (_03669_, _02819_, _06989_);
  and (_02820_, _07071_, _07053_);
  nor (_02821_, _02820_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_02822_, _02821_, _02806_);
  and (_02823_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_02824_, _02823_, _09580_);
  or (_02825_, _02824_, _02822_);
  and (_02826_, _02825_, _09574_);
  and (_02827_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_02828_, _02827_, _07046_);
  or (_02829_, _02828_, _02826_);
  nand (_02830_, _07317_, _07046_);
  and (_02831_, _02830_, _09590_);
  and (_02832_, _02831_, _02829_);
  and (_02833_, _07050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_02834_, _02833_, _02832_);
  and (_03672_, _02834_, _06989_);
  and (_02835_, _07071_, _07052_);
  nor (_02836_, _02835_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_02837_, _02836_, _02820_);
  and (_02838_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_02839_, _02838_, _09580_);
  or (_02840_, _02839_, _02837_);
  and (_02841_, _02840_, _09574_);
  and (_02842_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_02843_, _02842_, _07046_);
  or (_02844_, _02843_, _02841_);
  nand (_02845_, _11529_, _07046_);
  and (_02846_, _02845_, _09590_);
  and (_02847_, _02846_, _02844_);
  and (_02848_, _07050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_02849_, _02848_, _02847_);
  and (_03675_, _02849_, _06989_);
  and (_02850_, _07071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor (_02851_, _02850_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor (_02852_, _02851_, _02835_);
  and (_02853_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_02854_, _02853_, _09580_);
  or (_02855_, _02854_, _02852_);
  and (_02856_, _02855_, _09574_);
  and (_02857_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_02858_, _02857_, _07046_);
  or (_02859_, _02858_, _02856_);
  nand (_02860_, _09008_, _07046_);
  and (_02861_, _02860_, _09590_);
  and (_02862_, _02861_, _02859_);
  and (_02863_, _07050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_02864_, _02863_, _02862_);
  and (_03679_, _02864_, _06989_);
  or (_02865_, _11051_, _11018_);
  nor (_02866_, _11052_, _08477_);
  and (_02867_, _02866_, _02865_);
  nor (_02868_, _08476_, _06798_);
  or (_02869_, _02868_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02870_, _02869_, _02867_);
  or (_02871_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _02329_);
  and (_02872_, _02871_, _06989_);
  and (_03682_, _02872_, _02870_);
  or (_02873_, _01319_, _08123_);
  not (_02874_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_02875_, _01319_, _02874_);
  and (_02876_, _02875_, _06983_);
  and (_02877_, _02876_, _02873_);
  nor (_02878_, _06484_, _02874_);
  or (_02879_, _01319_, _08126_);
  and (_02880_, _02875_, _06485_);
  and (_02881_, _02880_, _02879_);
  or (_02882_, _02881_, _02878_);
  or (_02883_, _02882_, _02877_);
  and (_03687_, _02883_, _06989_);
  not (_02884_, _02487_);
  or (_03693_, _02884_, _02454_);
  and (_02885_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_02886_, _02885_, _07066_);
  nand (_02887_, _02886_, _02850_);
  or (_02888_, _07071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_02889_, _02888_, _09574_);
  and (_02890_, _02889_, _02887_);
  and (_02891_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_02892_, _02891_, _07046_);
  or (_02893_, _02892_, _02890_);
  nand (_02894_, _09598_, _07046_);
  and (_02895_, _02894_, _02893_);
  or (_02896_, _02895_, _07050_);
  or (_02897_, _09590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_02898_, _02897_, _06989_);
  and (_03698_, _02898_, _02896_);
  or (_02901_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand (_02902_, _07493_, _14007_);
  and (_02904_, _02902_, _06989_);
  and (_03706_, _02904_, _02901_);
  or (_02906_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand (_02908_, _07493_, _14020_);
  and (_02910_, _02908_, _06989_);
  and (_03712_, _02910_, _02906_);
  and (_02912_, _11389_, _11339_);
  nor (_02913_, _02912_, _02450_);
  or (_03715_, _02913_, _02884_);
  and (_02914_, _02462_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_02915_, _11433_, _11429_);
  or (_02916_, _11455_, _11426_);
  or (_02917_, _02916_, _02915_);
  and (_02918_, _02407_, _11312_);
  and (_02919_, _11399_, _11290_);
  and (_02920_, _11405_, _11312_);
  or (_02921_, _02920_, _02919_);
  or (_02923_, _02921_, _02918_);
  or (_02924_, _02923_, _02755_);
  or (_02925_, _02924_, _02917_);
  or (_02926_, _02434_, _11423_);
  and (_02927_, _02752_, _11934_);
  or (_02929_, _02710_, _02409_);
  and (_02931_, _11359_, _11934_);
  or (_02932_, _02931_, _02929_);
  or (_02934_, _02932_, _02927_);
  and (_02936_, _02405_, _11312_);
  or (_02938_, _02936_, _02423_);
  or (_02940_, _02938_, _02761_);
  and (_02941_, _11394_, _11313_);
  or (_02942_, _11453_, _02941_);
  or (_02943_, _02942_, _11449_);
  or (_02944_, _02943_, _02940_);
  or (_02945_, _02944_, _02934_);
  or (_02946_, _02945_, _02926_);
  or (_02947_, _02946_, _02925_);
  and (_02948_, _02947_, _02487_);
  or (_03719_, _02948_, _02914_);
  or (_02949_, _02663_, _02651_);
  or (_02950_, _02653_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_02951_, _02950_, _02949_);
  and (_02952_, _02951_, _02679_);
  nor (_02953_, _02678_, _11340_);
  or (_02954_, _02953_, rst);
  or (_03721_, _02954_, _02952_);
  nor (_02955_, _11050_, _11022_);
  nor (_02956_, _02955_, _11051_);
  or (_02957_, _02956_, _08477_);
  or (_02958_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_02959_, _02958_, _10964_);
  and (_02960_, _02959_, _02957_);
  and (_02961_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_03723_, _02961_, _02960_);
  and (_02963_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not (_02964_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_02966_, _01637_, _02964_);
  and (_02967_, _01637_, _02964_);
  nor (_02968_, _02967_, _02966_);
  and (_02969_, _02968_, _01647_);
  nor (_02970_, _02968_, _01647_);
  or (_02971_, _02970_, _02969_);
  or (_02972_, _02971_, _08477_);
  or (_02973_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_02974_, _02973_, _10964_);
  and (_02975_, _02974_, _02972_);
  or (_03726_, _02975_, _02963_);
  and (_02976_, _12716_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_02977_, _02976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_02978_, _02977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_02979_, _02977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_02980_, _02979_, _02978_);
  or (_02981_, _02980_, _11964_);
  and (_02982_, _02981_, _06989_);
  and (_02983_, _12278_, _11413_);
  and (_02984_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_02985_, _11974_, _11608_);
  or (_02986_, _02985_, _02984_);
  and (_02987_, _12314_, _11968_);
  or (_02988_, _02987_, _02986_);
  or (_02989_, _02988_, _02983_);
  or (_02990_, _12751_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_02991_, _02990_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_02992_, _02991_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_02993_, _02992_, _12742_);
  or (_02994_, _12757_, _08182_);
  nor (_02995_, _02994_, _08187_);
  nand (_02996_, _02995_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_02997_, _02996_, _12753_);
  nand (_02998_, _02997_, _02993_);
  nand (_02999_, _02998_, _12303_);
  or (_03000_, _02998_, _12303_);
  and (_03001_, _03000_, _02999_);
  and (_03002_, _03001_, _12722_);
  or (_03003_, _03002_, _02989_);
  and (_03004_, _12793_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_03005_, _03004_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_03006_, _03005_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_03007_, _03005_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_03008_, _03007_, _03006_);
  and (_03009_, _03008_, _12783_);
  or (_03010_, _03009_, _12781_);
  or (_03011_, _03010_, _03003_);
  and (_03742_, _03011_, _02982_);
  and (_03755_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _06989_);
  nor (_03758_, _12156_, rst);
  nand (_03012_, _10970_, _09531_);
  not (_03013_, _09537_);
  and (_03014_, _03013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_03015_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_03016_, _03015_, _03014_);
  or (_03017_, _03016_, _09531_);
  and (_03018_, _03017_, _06989_);
  and (_03761_, _03018_, _03012_);
  nand (_03019_, _10146_, _09598_);
  or (_03020_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_03021_, _03020_, _06989_);
  and (_03764_, _03021_, _03019_);
  nor (_03766_, _11492_, rst);
  or (_03022_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_03023_, _03013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_03024_, _03023_, _03022_);
  or (_03025_, _03024_, _09561_);
  nand (_03026_, _09561_, _09008_);
  and (_03027_, _03026_, _06989_);
  and (_03791_, _03027_, _03025_);
  and (_03028_, _11954_, _07044_);
  or (_03029_, _03028_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03030_, _03029_, _07292_);
  nand (_03031_, _03028_, _06968_);
  and (_03032_, _03031_, _03030_);
  or (_03033_, _03032_, _07293_);
  and (_03793_, _03033_, _06989_);
  nor (_03795_, _11415_, rst);
  nand (_03034_, _09531_, _07118_);
  and (_03035_, _03013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_03036_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_03037_, _03036_, _03035_);
  or (_03038_, _03037_, _09531_);
  and (_03039_, _03038_, _06989_);
  and (_03799_, _03039_, _03034_);
  nand (_03040_, _09531_, _07260_);
  and (_03041_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_03042_, _03013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_03043_, _03042_, _03041_);
  or (_03044_, _03043_, _09531_);
  and (_03045_, _03044_, _06989_);
  and (_03802_, _03045_, _03040_);
  not (_03046_, _09561_);
  or (_03048_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  not (_03049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand (_03050_, _09537_, _03049_);
  and (_03051_, _03050_, _03048_);
  and (_03052_, _03051_, _03046_);
  nor (_03054_, _03046_, _07317_);
  or (_03056_, _03054_, _03052_);
  and (_03805_, _03056_, _06989_);
  nor (_03808_, _12013_, rst);
  nor (_03810_, _12036_, rst);
  and (_03059_, _02462_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_03060_, _02568_, _02709_);
  or (_03061_, _03060_, _11395_);
  nand (_03062_, _02575_, _11290_);
  nand (_03063_, _03062_, _11326_);
  or (_03064_, _03063_, _03061_);
  or (_03065_, _02587_, _02408_);
  or (_03066_, _03065_, _02579_);
  nand (_03067_, _11457_, _11406_);
  or (_03068_, _02467_, _11387_);
  or (_03069_, _03068_, _02433_);
  and (_03070_, _11356_, _11290_);
  or (_03071_, _03070_, _11435_);
  or (_03073_, _03071_, _03069_);
  or (_03074_, _03073_, _03067_);
  or (_03075_, _03074_, _03066_);
  or (_03076_, _03075_, _03064_);
  not (_03078_, _11429_);
  and (_03080_, _11430_, _11382_);
  nor (_03082_, _03080_, _02601_);
  and (_03084_, _03082_, _03078_);
  not (_03086_, _03084_);
  or (_03088_, _02414_, _03086_);
  or (_03090_, _03088_, _11283_);
  or (_03092_, _03090_, _03076_);
  or (_03094_, _11334_, _11282_);
  nor (_03096_, \oc8051_top_1.oc8051_sfr1.wait_data , rst);
  and (_03097_, _03096_, _03094_);
  and (_03099_, _03097_, _03092_);
  or (_03815_, _03099_, _03059_);
  or (_03100_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_03101_, _03013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_03102_, _03101_, _03100_);
  or (_03103_, _03102_, _09531_);
  nand (_03104_, _11529_, _09531_);
  and (_03105_, _03104_, _06989_);
  and (_03821_, _03105_, _03103_);
  and (_03106_, _11954_, _08436_);
  or (_03107_, _03106_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_03108_, _03107_, _07292_);
  nand (_03109_, _03106_, _06968_);
  and (_03110_, _03109_, _03108_);
  or (_03111_, _03110_, _07318_);
  and (_03825_, _03111_, _06989_);
  or (_03112_, _07360_, _11345_);
  or (_03113_, _07324_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_03114_, _03113_, _06989_);
  and (_03829_, _03114_, _03112_);
  nor (_03115_, _11049_, _11044_);
  nor (_03116_, _03115_, _11050_);
  or (_03117_, _03116_, _08477_);
  or (_03118_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_03119_, _03118_, _10964_);
  and (_03120_, _03119_, _03117_);
  and (_03121_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_03831_, _03121_, _03120_);
  or (_03122_, _08496_, _11345_);
  or (_03123_, _07324_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_03124_, _03123_, _06989_);
  and (_03833_, _03124_, _03122_);
  nand (_03125_, _08512_, _07324_);
  or (_03126_, _07324_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_03128_, _03126_, _06989_);
  and (_03835_, _03128_, _03125_);
  or (_03129_, _08529_, _11345_);
  or (_03130_, _07324_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_03131_, _03130_, _06989_);
  and (_03837_, _03131_, _03129_);
  or (_03132_, _08545_, _11345_);
  or (_03133_, _07324_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_03134_, _03133_, _06989_);
  and (_03839_, _03134_, _03132_);
  or (_03136_, _08561_, _11345_);
  or (_03137_, _07324_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_03138_, _03137_, _06989_);
  and (_03841_, _03138_, _03136_);
  nand (_03139_, _08576_, _07324_);
  or (_03140_, _07324_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_03141_, _03140_, _06989_);
  and (_03854_, _03141_, _03139_);
  or (_03142_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not (_03143_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_03144_, _09537_, _03143_);
  and (_03145_, _03144_, _03142_);
  or (_03147_, _03145_, _09561_);
  nand (_03148_, _09598_, _09561_);
  and (_03149_, _03148_, _06989_);
  and (_03862_, _03149_, _03147_);
  or (_03151_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03152_, _08085_, _07978_);
  or (_03153_, _03152_, _09182_);
  or (_03154_, _03153_, _08402_);
  or (_03155_, _03154_, _08231_);
  or (_03157_, _03155_, _09092_);
  and (_03158_, _03157_, _07027_);
  and (_03159_, _06898_, _06848_);
  not (_03160_, _06898_);
  and (_03161_, _06900_, _03160_);
  or (_03162_, _03161_, _03159_);
  and (_03163_, _03162_, _06845_);
  nand (_03164_, _06834_, _06599_);
  and (_03165_, _06837_, _06548_);
  and (_03166_, _03165_, _03164_);
  and (_03167_, _07024_, _06652_);
  and (_03168_, _03167_, _06622_);
  and (_03169_, _03168_, _07634_);
  nand (_03170_, _03169_, _08152_);
  nand (_03171_, _03170_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_03172_, _03171_, _03166_);
  nor (_03173_, _03172_, _03163_);
  and (_03174_, _03173_, _08318_);
  nand (_03175_, _03174_, _12250_);
  or (_03176_, _03175_, _03158_);
  and (_03177_, _03176_, _03151_);
  or (_03178_, _03177_, _11954_);
  not (_03179_, _11954_);
  and (_03180_, _00759_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03181_, _03180_, _03179_);
  or (_03182_, _03181_, _00760_);
  and (_03183_, _03182_, _03178_);
  or (_03184_, _03183_, _07291_);
  nand (_03185_, _11529_, _07291_);
  and (_03186_, _03185_, _06989_);
  and (_03864_, _03186_, _03184_);
  or (_03187_, _02583_, _11437_);
  or (_03188_, _03187_, _02919_);
  or (_03189_, _03188_, _02726_);
  not (_03190_, _14315_);
  or (_03191_, _02720_, _03190_);
  or (_03192_, _03191_, _03189_);
  or (_03193_, _02941_, _11395_);
  or (_03194_, _02709_, _02423_);
  or (_03195_, _03194_, _03193_);
  or (_03196_, _02929_, _02582_);
  or (_03197_, _03196_, _03195_);
  and (_03198_, _11359_, _11290_);
  or (_03199_, _02719_, _02406_);
  or (_03200_, _03199_, _03198_);
  or (_03201_, _11334_, _11433_);
  or (_03202_, _11919_, _14316_);
  or (_03203_, _03202_, _03201_);
  or (_03204_, _03203_, _03200_);
  or (_03205_, _03204_, _03197_);
  or (_03206_, _03205_, _03192_);
  and (_03207_, _03206_, _03097_);
  and (_03208_, _02462_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  or (_03869_, _03208_, _03207_);
  and (_03210_, _11954_, _07089_);
  or (_03211_, _03210_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03212_, _03211_, _07292_);
  nand (_03213_, _03210_, _06968_);
  and (_03214_, _03213_, _03212_);
  nor (_03215_, _09008_, _07292_);
  or (_03216_, _03215_, _03214_);
  and (_03873_, _03216_, _06989_);
  and (_03217_, _11355_, _11290_);
  or (_03218_, _02406_, _14313_);
  or (_03219_, _03218_, _03217_);
  or (_03220_, _03219_, _02720_);
  or (_03221_, _03188_, _02792_);
  or (_03222_, _03221_, _03220_);
  or (_03223_, _11456_, _11401_);
  or (_03224_, _11453_, _14316_);
  or (_03225_, _03224_, _03223_);
  or (_03226_, _03225_, _02916_);
  or (_03227_, _03226_, _02926_);
  or (_03228_, _03227_, _03222_);
  and (_03229_, _03228_, _07325_);
  and (_03230_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_03231_, _11333_, _06406_);
  or (_03232_, _03231_, _03230_);
  or (_03233_, _03232_, _03229_);
  and (_03879_, _03233_, _06989_);
  nand (_03234_, _09536_, _07317_);
  and (_03235_, _09534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_03236_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_03237_, _03236_, _03235_);
  or (_03238_, _03237_, _09536_);
  and (_03239_, _03238_, _09552_);
  and (_03240_, _03239_, _03234_);
  and (_03241_, _09531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_03242_, _03241_, _03240_);
  and (_03917_, _03242_, _06989_);
  not (_03243_, _09536_);
  or (_03244_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  not (_03245_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand (_03246_, _09533_, _03245_);
  nand (_03247_, _03246_, _03244_);
  nand (_03248_, _03247_, _03243_);
  nand (_03249_, _10970_, _09536_);
  and (_03250_, _03249_, _03248_);
  or (_03251_, _03250_, _09561_);
  not (_03252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nand (_03253_, _09561_, _03252_);
  and (_03254_, _03253_, _06989_);
  and (_03920_, _03254_, _03251_);
  nand (_03255_, _09536_, _07118_);
  not (_03256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor (_03257_, _09533_, _03256_);
  and (_03258_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_03259_, _03258_, _03257_);
  or (_03260_, _03259_, _09536_);
  and (_03261_, _03260_, _09552_);
  and (_03262_, _03261_, _03255_);
  and (_03263_, _09531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_03264_, _03263_, _03262_);
  and (_03926_, _03264_, _06989_);
  nand (_03265_, _09536_, _07260_);
  and (_03266_, _09534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_03267_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_03268_, _03267_, _03266_);
  or (_03269_, _03268_, _09536_);
  and (_03270_, _03269_, _09552_);
  and (_03271_, _03270_, _03265_);
  and (_03272_, _09531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_03273_, _03272_, _03271_);
  and (_03929_, _03273_, _06989_);
  nand (_03274_, _11529_, _09536_);
  and (_03275_, _09534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_03276_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_03277_, _03276_, _03275_);
  or (_03278_, _03277_, _09536_);
  and (_03279_, _03278_, _09552_);
  and (_03280_, _03279_, _03274_);
  and (_03281_, _09531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_03282_, _03281_, _03280_);
  and (_03942_, _03282_, _06989_);
  and (_03283_, _08999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_03284_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_03285_, _03284_, _09002_);
  and (_03286_, _11821_, _09010_);
  or (_03287_, _03286_, _03285_);
  or (_03288_, _03287_, _03283_);
  and (_03957_, _03288_, _06989_);
  nand (_03289_, _09536_, _09008_);
  or (_03290_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_03291_, _09534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_03292_, _03291_, _03290_);
  or (_03293_, _03292_, _09536_);
  and (_03294_, _03293_, _09552_);
  and (_03295_, _03294_, _03289_);
  and (_03296_, _09531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_03297_, _03296_, _03295_);
  and (_03966_, _03297_, _06989_);
  nand (_03298_, _09598_, _09536_);
  or (_03299_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_03300_, _09534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_03301_, _03300_, _03299_);
  or (_03302_, _03301_, _09536_);
  and (_03303_, _03302_, _03298_);
  or (_03304_, _03303_, _09561_);
  or (_03305_, _03046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_03306_, _03305_, _06989_);
  and (_03971_, _03306_, _03304_);
  or (_03307_, _08994_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand (_03308_, _08994_, _07040_);
  and (_03309_, _03308_, _03307_);
  or (_03310_, _03309_, _06982_);
  or (_03311_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and (_03312_, _03311_, _06989_);
  and (_03992_, _03312_, _03310_);
  and (_03314_, _02462_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor (_03316_, _11909_, _11474_);
  nand (_03317_, _03316_, _11920_);
  or (_03318_, _02931_, _02927_);
  or (_03319_, _03318_, _03317_);
  or (_03320_, _02433_, _02423_);
  or (_03321_, _02919_, _02691_);
  or (_03322_, _03321_, _03320_);
  or (_03323_, _03322_, _02785_);
  or (_03324_, _03323_, _02917_);
  or (_03325_, _03324_, _03319_);
  and (_03326_, _03325_, _02487_);
  or (_03995_, _03326_, _03314_);
  nor (_03328_, _14146_, _07118_);
  and (_03330_, _08999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_03332_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and (_03333_, _03332_, _09002_);
  or (_03334_, _03333_, _03330_);
  or (_03335_, _03334_, _03328_);
  and (_04003_, _03335_, _06989_);
  nor (_04007_, _12061_, rst);
  nor (_03336_, _09614_, _07040_);
  and (_03337_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_03338_, _03337_, _06982_);
  or (_03339_, _03338_, _03336_);
  or (_03340_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_03341_, _03340_, _06989_);
  and (_04034_, _03341_, _03339_);
  or (_03342_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand (_03343_, _07493_, _14092_);
  and (_03344_, _03343_, _06989_);
  and (_04059_, _03344_, _03342_);
  and (_03346_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_03347_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  or (_03348_, _03347_, _03346_);
  and (_04061_, _03348_, _06989_);
  and (_03349_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_03351_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  or (_03352_, _03351_, _03349_);
  and (_04068_, _03352_, _06989_);
  and (_04086_, _06989_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  and (_03353_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_03355_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_03356_, _03355_, _06989_);
  nor (_04099_, _03356_, _03353_);
  and (_04104_, _08314_, _06989_);
  and (_03357_, _09610_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_03358_, _11529_, _07486_);
  and (_03359_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_03360_, _03359_, _09615_);
  or (_03361_, _03360_, _03358_);
  or (_03362_, _03361_, _03357_);
  and (_04112_, _03362_, _06989_);
  and (_03363_, _11277_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_03365_, _03363_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_03366_, _03365_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_03367_, _03366_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_03368_, _03367_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand (_03369_, _03367_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_03370_, _03369_, _03368_);
  or (_03371_, _03370_, _11964_);
  and (_03373_, _03371_, _06989_);
  and (_03375_, _12750_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_03376_, _03375_, _12752_);
  or (_03377_, _12756_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_03378_, _03377_, _12757_);
  or (_03379_, _03378_, _12742_);
  and (_03380_, _03379_, _12722_);
  and (_03381_, _03380_, _03376_);
  nor (_03382_, _12790_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_03383_, _03382_, _12791_);
  and (_03384_, _03383_, _12783_);
  and (_03385_, _11413_, _08433_);
  nor (_03386_, _12797_, _08385_);
  and (_03387_, _11974_, _11514_);
  and (_03388_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_03389_, _03388_, _03387_);
  or (_03390_, _03389_, _03386_);
  or (_03391_, _03390_, _03385_);
  or (_03392_, _03391_, _03384_);
  or (_03393_, _03392_, _12781_);
  or (_03394_, _03393_, _03381_);
  and (_04114_, _03394_, _03373_);
  nand (_03395_, _10970_, _10146_);
  or (_03396_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_03397_, _03396_, _06989_);
  and (_04117_, _03397_, _03395_);
  nor (_03398_, _03366_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_03400_, _03398_, _03367_);
  or (_03401_, _03400_, _11964_);
  and (_03402_, _03401_, _06989_);
  nor (_03403_, _12797_, _09356_);
  nor (_03404_, _11989_, _09227_);
  and (_03405_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_03406_, _11974_, _11842_);
  and (_03407_, _12176_, _08463_);
  or (_03408_, _03407_, _03406_);
  or (_03409_, _03408_, _03405_);
  or (_03410_, _03409_, _03404_);
  or (_03411_, _03410_, _03403_);
  and (_03412_, _12749_, _12742_);
  and (_03414_, _12754_, _12747_);
  nor (_03415_, _03414_, _12742_);
  or (_03416_, _03415_, _03412_);
  nand (_03417_, _03416_, _08175_);
  or (_03418_, _03416_, _08175_);
  and (_03419_, _03418_, _03417_);
  and (_03421_, _03419_, _12722_);
  or (_03423_, _03421_, _03411_);
  or (_03424_, _03423_, _12781_);
  and (_04122_, _03424_, _03402_);
  nor (_03425_, _03365_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_03426_, _03425_, _03366_);
  or (_03427_, _03426_, _11964_);
  and (_03429_, _03427_, _06989_);
  and (_03430_, _12747_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_03431_, _03430_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_03432_, _03431_, _03415_);
  nand (_03433_, _12748_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_03434_, _03433_, _12749_);
  and (_03435_, _03434_, _12742_);
  or (_03436_, _03435_, _03432_);
  and (_03437_, _03436_, _12722_);
  and (_03438_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_03440_, _11974_, _11744_);
  or (_03441_, _03440_, _03438_);
  nor (_03442_, _12797_, _07696_);
  or (_03443_, _03442_, _03441_);
  and (_03445_, _11413_, _08030_);
  and (_03446_, _12783_, _10835_);
  or (_03448_, _03446_, _03445_);
  or (_03449_, _03448_, _03443_);
  or (_03450_, _03449_, _03437_);
  or (_03451_, _03450_, _12781_);
  and (_04130_, _03451_, _03429_);
  nor (_03452_, _03363_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_03453_, _03452_, _03365_);
  or (_03454_, _03453_, _11964_);
  and (_03455_, _03454_, _06989_);
  and (_03457_, _11413_, _08123_);
  nand (_03458_, _12747_, _07646_);
  or (_03459_, _12747_, _07646_);
  and (_03460_, _03459_, _03458_);
  and (_03461_, _03460_, _12742_);
  nor (_03462_, _03460_, _12742_);
  or (_03463_, _03462_, _03461_);
  and (_03464_, _03463_, _12171_);
  and (_03465_, _12167_, _08075_);
  and (_03466_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_03467_, _11974_, _11786_);
  or (_03468_, _03467_, _03466_);
  and (_03469_, _12176_, _08561_);
  nor (_03470_, _03469_, _03468_);
  nand (_03471_, _03470_, _11964_);
  or (_03472_, _03471_, _03465_);
  or (_03473_, _03472_, _03464_);
  or (_03474_, _03473_, _03457_);
  and (_04134_, _03474_, _03455_);
  nor (_03476_, _11277_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_03477_, _03476_, _03363_);
  or (_03478_, _03477_, _11964_);
  and (_03480_, _03478_, _06989_);
  and (_03481_, _12278_, _11986_);
  and (_03482_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_03483_, _12740_, _11988_);
  and (_03484_, _12783_, _11608_);
  or (_03485_, _03484_, _03483_);
  or (_03487_, _03485_, _03482_);
  or (_03488_, _12744_, _12743_);
  not (_03490_, _03488_);
  nand (_03491_, _03490_, _12745_);
  or (_03492_, _03490_, _12745_);
  and (_03493_, _03492_, _12722_);
  and (_03494_, _03493_, _03491_);
  or (_03495_, _03494_, _03487_);
  or (_03496_, _03495_, _03481_);
  or (_03497_, _03496_, _12781_);
  and (_04137_, _03497_, _03480_);
  not (_03498_, _00919_);
  and (_03499_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_03500_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_03501_, _03500_, _03499_);
  and (_03502_, _03501_, _13953_);
  and (_03503_, _13952_, _09393_);
  or (_03504_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _13995_);
  and (_03505_, _03504_, _06989_);
  and (_03506_, _03505_, _03503_);
  or (_04187_, _03506_, _03502_);
  nor (_03507_, _03353_, _07526_);
  and (_03508_, _03353_, _07526_);
  or (_03509_, _03508_, _03507_);
  and (_04196_, _03509_, _06989_);
  and (_04199_, _12244_, _06989_);
  and (_04206_, _06989_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor (_03510_, _14146_, _07040_);
  and (_03511_, _08999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_03513_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and (_03514_, _03513_, _09002_);
  or (_03515_, _03514_, _03511_);
  or (_03516_, _03515_, _03510_);
  and (_04207_, _03516_, _06989_);
  or (_03517_, _09605_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nand (_03519_, _09008_, _09605_);
  and (_03520_, _03519_, _03517_);
  or (_03522_, _03520_, _06982_);
  or (_03523_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_03524_, _03523_, _06989_);
  and (_04211_, _03524_, _03522_);
  nor (_03525_, _07317_, _09614_);
  and (_03526_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_03527_, _03526_, _06982_);
  or (_03528_, _03527_, _03525_);
  or (_03529_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_03530_, _03529_, _06989_);
  and (_04214_, _03530_, _03528_);
  nor (_03531_, _10970_, _09614_);
  and (_03532_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_03533_, _03532_, _06982_);
  or (_03534_, _03533_, _03531_);
  or (_03535_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_03536_, _03535_, _06989_);
  and (_04216_, _03536_, _03534_);
  nor (_03537_, _11724_, _14222_);
  and (_03538_, _03537_, _14354_);
  or (_03540_, _01595_, _14253_);
  or (_03542_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03543_, _03542_, _14217_);
  and (_03544_, _03543_, _03540_);
  and (_03545_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_03546_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_03547_, _03546_, _03545_);
  and (_03548_, _03547_, _14241_);
  nor (_03550_, _11857_, _08412_);
  and (_03551_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03552_, _03551_, _03550_);
  and (_03553_, _03552_, _14205_);
  and (_03554_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_03555_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_03556_, _03555_, _03554_);
  and (_03558_, _03556_, _14233_);
  or (_03559_, _03558_, _03553_);
  or (_03560_, _03559_, _03548_);
  or (_03562_, _03560_, _03544_);
  and (_03563_, _03562_, _03538_);
  and (_03564_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_03565_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03567_, _03565_, _03564_);
  and (_03568_, _03567_, _14233_);
  and (_03569_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_03570_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_03571_, _03570_, _03569_);
  and (_03572_, _03571_, _14205_);
  and (_03573_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_03574_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_03575_, _03574_, _03573_);
  and (_03576_, _03575_, _14217_);
  or (_03577_, _03576_, _03572_);
  and (_03578_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03580_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_03581_, _03580_, _03578_);
  and (_03582_, _03581_, _14241_);
  or (_03583_, _03582_, _03577_);
  or (_03584_, _03583_, _03568_);
  and (_03585_, _03584_, _14209_);
  and (_03586_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03587_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_03588_, _03587_, _03586_);
  and (_03589_, _03588_, _14241_);
  and (_03590_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_03591_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_03592_, _03591_, _03590_);
  and (_03593_, _03592_, _14205_);
  nor (_03594_, _11857_, _07176_);
  and (_03595_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_03596_, _03595_, _03594_);
  and (_03597_, _03596_, _14217_);
  or (_03599_, _03597_, _03593_);
  nor (_03600_, _11857_, _07172_);
  and (_03601_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_03602_, _03601_, _03600_);
  and (_03603_, _03602_, _14233_);
  or (_03604_, _03603_, _03599_);
  or (_03605_, _03604_, _03589_);
  and (_03606_, _03605_, _14248_);
  nor (_03607_, _11857_, _07213_);
  and (_03608_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_03609_, _03608_, _03607_);
  and (_03610_, _03609_, _14217_);
  and (_03611_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_03612_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_03613_, _03612_, _03611_);
  and (_03614_, _03613_, _14241_);
  or (_03615_, _03614_, _03610_);
  and (_03616_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_03618_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_03620_, _03618_, _03616_);
  and (_03621_, _03620_, _14205_);
  and (_03623_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor (_03624_, _11857_, _07211_);
  or (_03625_, _03624_, _03623_);
  and (_03626_, _03625_, _14233_);
  or (_03627_, _03626_, _03621_);
  or (_03628_, _03627_, _03615_);
  and (_03629_, _03628_, _14252_);
  or (_03630_, _03629_, _03606_);
  or (_03631_, _03630_, _03585_);
  and (_03632_, _03631_, _14222_);
  and (_03633_, _14209_, _11556_);
  nor (_03635_, _14326_, p0_in[7]);
  and (_03637_, _14326_, _00731_);
  nor (_03639_, _03637_, _03635_);
  and (_03640_, _03639_, _14253_);
  and (_03642_, _14463_, _11857_);
  or (_03644_, _03642_, _03640_);
  and (_03646_, _03644_, _14241_);
  and (_03647_, _14602_, _11857_);
  and (_03649_, _01288_, _14253_);
  or (_03650_, _03649_, _03647_);
  and (_03652_, _03650_, _14233_);
  and (_03653_, _14529_, _11857_);
  and (_03654_, _14342_, _14253_);
  or (_03656_, _03654_, _03653_);
  and (_03658_, _03656_, _14205_);
  and (_03660_, _01462_, _14253_);
  and (_03661_, _01541_, _11857_);
  or (_03663_, _03661_, _03660_);
  and (_03665_, _03663_, _14217_);
  or (_03667_, _03665_, _03658_);
  or (_03668_, _03667_, _03652_);
  or (_03670_, _03668_, _03646_);
  and (_03671_, _03670_, _03633_);
  and (_03673_, _11724_, _11556_);
  and (_03674_, _03673_, _14292_);
  nor (_03676_, _11857_, _06649_);
  and (_03677_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03678_, _03677_, _03676_);
  and (_03680_, _03678_, _14217_);
  nor (_03681_, _11857_, _06813_);
  and (_03683_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03684_, _03683_, _03681_);
  and (_03685_, _03684_, _14205_);
  or (_03686_, _03685_, _03680_);
  nor (_03688_, _11857_, _06619_);
  and (_03689_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_03690_, _03689_, _03688_);
  and (_03691_, _03690_, _14233_);
  nor (_03692_, _11857_, _06592_);
  and (_03694_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_03695_, _03694_, _03692_);
  and (_03696_, _03695_, _14241_);
  or (_03697_, _03696_, _03691_);
  or (_03699_, _03697_, _03686_);
  and (_03700_, _03699_, _03674_);
  or (_03701_, _03700_, _03671_);
  and (_03702_, _11863_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_03703_, _14214_, _14222_);
  and (_03704_, _03703_, _14206_);
  and (_03705_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_03707_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_03708_, _03707_, _03705_);
  and (_03709_, _03708_, _14205_);
  nor (_03710_, _11857_, _13993_);
  and (_03711_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_03713_, _03711_, _03710_);
  and (_03714_, _03713_, _14217_);
  or (_03716_, _03714_, _03709_);
  and (_03717_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor (_03718_, _11857_, _06970_);
  or (_03720_, _03718_, _03717_);
  and (_03722_, _03720_, _14241_);
  nor (_03724_, _11857_, _14039_);
  and (_03725_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_03727_, _03725_, _03724_);
  and (_03728_, _03727_, _14233_);
  or (_03729_, _03728_, _03722_);
  or (_03730_, _03729_, _03716_);
  and (_03731_, _03730_, _03704_);
  or (_03732_, _03731_, _03702_);
  or (_03733_, _03732_, _03701_);
  and (_03734_, _01535_, _11857_);
  and (_03735_, _01468_, _14253_);
  or (_03736_, _03735_, _03734_);
  and (_03737_, _03736_, _14217_);
  and (_03738_, _14612_, _11857_);
  and (_03739_, _01303_, _14253_);
  or (_03740_, _03739_, _03738_);
  and (_03741_, _03740_, _14233_);
  or (_03743_, _03741_, _11724_);
  or (_03744_, _03743_, _03737_);
  and (_03745_, _14540_, _14205_);
  and (_03746_, _14458_, _14241_);
  or (_03747_, _03746_, _03745_);
  and (_03748_, _03747_, _11857_);
  and (_03749_, _14330_, _14205_);
  nor (_03750_, _14326_, p3_in[7]);
  and (_03751_, _14326_, _01165_);
  nor (_03752_, _03751_, _03750_);
  and (_03753_, _03752_, _14241_);
  or (_03754_, _03753_, _03749_);
  and (_03756_, _03754_, _14253_);
  or (_03757_, _03756_, _03748_);
  or (_03759_, _03757_, _03744_);
  and (_03760_, _14247_, _11556_);
  and (_03762_, _14544_, _11857_);
  and (_03763_, _14336_, _14253_);
  or (_03765_, _03763_, _03762_);
  and (_03767_, _03765_, _14205_);
  and (_03768_, _14616_, _11857_);
  and (_03769_, _01298_, _14253_);
  or (_03770_, _03769_, _03768_);
  and (_03771_, _03770_, _14233_);
  or (_03772_, _03771_, _14251_);
  or (_03773_, _03772_, _03767_);
  and (_03774_, _14453_, _14241_);
  and (_03775_, _01530_, _14217_);
  or (_03776_, _03775_, _03774_);
  and (_03777_, _03776_, _11857_);
  nor (_03778_, _14326_, p2_in[7]);
  and (_03779_, _14326_, _09033_);
  nor (_03780_, _03779_, _03778_);
  and (_03781_, _03780_, _14241_);
  and (_03782_, _01473_, _14217_);
  or (_03783_, _03782_, _03781_);
  and (_03784_, _03783_, _14253_);
  or (_03785_, _03784_, _03777_);
  or (_03786_, _03785_, _03773_);
  and (_03787_, _03786_, _03760_);
  and (_03788_, _03787_, _03759_);
  nor (_03789_, _11857_, _01372_);
  and (_03790_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03792_, _03790_, _03789_);
  and (_03794_, _03792_, _14233_);
  or (_03796_, _03794_, _11556_);
  and (_03797_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_03798_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_03800_, _03798_, _03797_);
  and (_03801_, _03800_, _14205_);
  nor (_03803_, _11857_, _09405_);
  and (_03804_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_03806_, _03804_, _03803_);
  and (_03807_, _03806_, _14217_);
  and (_03809_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor (_03811_, _11857_, _13995_);
  or (_03812_, _03811_, _03809_);
  and (_03813_, _03812_, _14241_);
  or (_03814_, _03813_, _03807_);
  or (_03816_, _03814_, _03801_);
  or (_03817_, _03816_, _03796_);
  and (_03818_, _14534_, _11857_);
  and (_03819_, _14347_, _14253_);
  or (_03820_, _03819_, _03818_);
  and (_03822_, _03820_, _14205_);
  and (_03823_, _14606_, _11857_);
  and (_03824_, _01293_, _14253_);
  or (_03826_, _03824_, _03823_);
  and (_03827_, _03826_, _14233_);
  or (_03828_, _03827_, _14222_);
  or (_03830_, _03828_, _03822_);
  nor (_03832_, _14326_, p1_in[7]);
  and (_03834_, _14326_, _00702_);
  nor (_03836_, _03834_, _03832_);
  and (_03838_, _03836_, _14241_);
  and (_03840_, _01457_, _14217_);
  or (_03842_, _03840_, _03838_);
  and (_03843_, _03842_, _14253_);
  and (_03844_, _14467_, _14241_);
  and (_03845_, _01546_, _14217_);
  or (_03846_, _03845_, _03844_);
  and (_03847_, _03846_, _11857_);
  or (_03848_, _03847_, _03843_);
  or (_03849_, _03848_, _03830_);
  and (_03850_, _03849_, _14276_);
  and (_03851_, _03850_, _03817_);
  and (_03852_, _03537_, _14292_);
  nor (_03853_, _03852_, _03538_);
  nor (_03855_, _03704_, _03674_);
  and (_03856_, _03855_, _03853_);
  nor (_03857_, _14275_, _14222_);
  nor (_03858_, _14208_, _11556_);
  or (_03859_, _03858_, _03857_);
  not (_03860_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_03861_, _03760_, _03860_);
  and (_03863_, _03861_, _03859_);
  and (_03865_, _03863_, _03856_);
  nor (_03866_, _11857_, _01749_);
  and (_03867_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_03868_, _03867_, _03866_);
  and (_03870_, _03868_, _14217_);
  nor (_03871_, _11857_, _01885_);
  and (_03872_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_03874_, _03872_, _03871_);
  and (_03875_, _03874_, _14205_);
  or (_03876_, _03875_, _03870_);
  nor (_03877_, _11857_, _01321_);
  and (_03878_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_03880_, _03878_, _03877_);
  and (_03881_, _03880_, _14233_);
  not (_03882_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor (_03883_, _11857_, _03882_);
  and (_03884_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_03885_, _03884_, _03883_);
  and (_03886_, _03885_, _14241_);
  or (_03887_, _03886_, _03881_);
  or (_03888_, _03887_, _03876_);
  and (_03889_, _03888_, _03852_);
  or (_03890_, _03889_, _03865_);
  or (_03891_, _03890_, _03851_);
  or (_03892_, _03891_, _03788_);
  or (_03893_, _03892_, _03733_);
  or (_03894_, _03893_, _03632_);
  or (_03895_, _03894_, _03563_);
  and (_03896_, _03674_, _07705_);
  nor (_03897_, _03896_, _11873_);
  nand (_03898_, _03702_, _06968_);
  and (_03899_, _03898_, _03897_);
  and (_03900_, _03899_, _03895_);
  and (_03901_, _11857_, _09009_);
  nor (_03902_, _11857_, _07118_);
  or (_03903_, _03902_, _03901_);
  and (_03904_, _03903_, _14233_);
  and (_03905_, _11857_, _11821_);
  nor (_03906_, _11857_, _10970_);
  or (_03907_, _03906_, _03905_);
  and (_03908_, _03907_, _14205_);
  nor (_03909_, _11857_, _07260_);
  and (_03910_, _11857_, _09599_);
  or (_03911_, _03910_, _03909_);
  and (_03912_, _03911_, _14217_);
  or (_03913_, _03912_, _03908_);
  nor (_03914_, _11857_, _07040_);
  and (_03915_, _11857_, _07410_);
  or (_03916_, _03915_, _03914_);
  and (_03918_, _03916_, _14241_);
  or (_03919_, _03918_, _03913_);
  nor (_03921_, _03919_, _03904_);
  nor (_03922_, _03921_, _03897_);
  or (_03923_, _03922_, _03900_);
  and (_04219_, _03923_, _06989_);
  nor (_03924_, _00489_, rst);
  or (_03925_, _00488_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand (_03927_, _00488_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03928_, _03927_, _03925_);
  and (_04224_, _03928_, _03924_);
  and (_04227_, _00490_, _06989_);
  nor (_03930_, _02976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_03931_, _03930_, _02977_);
  or (_03932_, _03931_, _11964_);
  and (_03933_, _03932_, _06989_);
  and (_03934_, _02995_, _09270_);
  nor (_03935_, _02995_, _09270_);
  or (_03936_, _03935_, _03934_);
  and (_03937_, _03936_, _12753_);
  nand (_03938_, _02991_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_03939_, _03938_, _02992_);
  and (_03940_, _03939_, _12742_);
  or (_03941_, _03940_, _03937_);
  and (_03943_, _03941_, _12722_);
  nor (_03944_, _03004_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_03945_, _03944_, _03005_);
  and (_03946_, _03945_, _12783_);
  nor (_03947_, _11989_, _09145_);
  nor (_03948_, _12797_, _09285_);
  and (_03949_, _11974_, _11618_);
  and (_03950_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_03951_, _03950_, _03949_);
  or (_03952_, _03951_, _03948_);
  or (_03953_, _03952_, _03947_);
  or (_03954_, _03953_, _03946_);
  or (_03955_, _03954_, _12781_);
  or (_03956_, _03955_, _03943_);
  and (_04233_, _03956_, _03933_);
  nor (_03958_, _12716_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_03959_, _03958_, _02976_);
  or (_03960_, _03959_, _11964_);
  and (_03961_, _03960_, _06989_);
  or (_03962_, _12793_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_03963_, _03004_);
  and (_03964_, _03963_, _12783_);
  and (_03965_, _03964_, _03962_);
  and (_03967_, _11413_, _08268_);
  nor (_03968_, _12797_, _08202_);
  and (_03969_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_03970_, _11974_, _11671_);
  or (_03972_, _03970_, _03969_);
  or (_03973_, _03972_, _03968_);
  or (_03974_, _03973_, _03967_);
  or (_03975_, _02990_, _12753_);
  or (_03976_, _02994_, _12742_);
  and (_03977_, _03976_, _03975_);
  nand (_03978_, _03977_, _08187_);
  or (_03979_, _03977_, _08187_);
  and (_03980_, _03979_, _03978_);
  and (_03981_, _03980_, _12722_);
  or (_03982_, _03981_, _03974_);
  or (_03983_, _03982_, _03965_);
  or (_03984_, _03983_, _12781_);
  and (_04236_, _03984_, _03961_);
  and (_03986_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_03987_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_03988_, _03987_, _03986_);
  or (_03989_, _03988_, _13986_);
  and (_03990_, _03989_, _06989_);
  nand (_03991_, _03503_, _07040_);
  and (_04282_, _03991_, _03990_);
  or (_03993_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand (_03994_, _07493_, _14184_);
  and (_03996_, _03994_, _06989_);
  and (_04306_, _03996_, _03993_);
  and (_03997_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_03998_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_03999_, _03998_, _03997_);
  and (_04000_, _03999_, _13953_);
  nand (_04001_, _09392_, _07040_);
  nand (_04002_, _10970_, _09393_);
  and (_04004_, _04002_, _00922_);
  and (_04005_, _04004_, _04001_);
  or (_04334_, _04005_, _04000_);
  and (_04006_, _13952_, _09392_);
  and (_04008_, _04006_, _11646_);
  and (_04009_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_04010_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_04011_, _04010_, _04009_);
  nor (_04012_, _04011_, _13986_);
  and (_04013_, _03503_, _07119_);
  or (_04014_, _04013_, _04012_);
  or (_04015_, _04014_, _04008_);
  and (_04339_, _04015_, _06989_);
  not (_04016_, _11353_);
  and (_04017_, _02701_, _04016_);
  nor (_04018_, _02697_, _11474_);
  nand (_04019_, _04018_, _11440_);
  or (_04020_, _04019_, _11449_);
  or (_04021_, _04020_, _02917_);
  and (_04022_, _04021_, _11282_);
  or (_04023_, _04022_, _04017_);
  and (_04353_, _04023_, _06989_);
  nor (_04024_, _14213_, rst);
  and (_04025_, _12278_, _06989_);
  or (_04026_, _04025_, _04024_);
  not (_04027_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nor (_04028_, _14404_, _04027_);
  nand (_04029_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_04030_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_04031_, _04030_, _04029_);
  nand (_04032_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nand (_04033_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_04035_, _04033_, _04032_);
  and (_04036_, _04035_, _04031_);
  nand (_04037_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nand (_04038_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_04039_, _04038_, _04037_);
  nand (_04040_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nand (_04041_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_04042_, _04041_, _04040_);
  and (_04043_, _04042_, _04039_);
  and (_04044_, _04043_, _04036_);
  nand (_04045_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  nand (_04046_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_04047_, _04046_, _04045_);
  nand (_04048_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_04049_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_04050_, _04049_, _04048_);
  and (_04051_, _04050_, _04047_);
  nand (_04052_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nand (_04053_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_04054_, _04053_, _04052_);
  nand (_04055_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_04056_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_04057_, _04056_, _04055_);
  and (_04058_, _04057_, _04054_);
  and (_04060_, _04058_, _04051_);
  and (_04062_, _04060_, _04044_);
  nand (_04063_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand (_04064_, _14296_, _11605_);
  and (_04065_, _04064_, _04063_);
  nand (_04066_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand (_04067_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and (_04069_, _04067_, _04066_);
  and (_04070_, _04069_, _04065_);
  nand (_04071_, _03780_, _14333_);
  nand (_04072_, _03752_, _14305_);
  and (_04073_, _04072_, _04071_);
  nand (_04074_, _03639_, _14339_);
  nand (_04075_, _03836_, _14344_);
  and (_04076_, _04075_, _04074_);
  and (_04077_, _04076_, _04073_);
  and (_04078_, _04077_, _04070_);
  nand (_04079_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand (_04080_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_04081_, _04080_, _04079_);
  and (_04082_, _04081_, _04078_);
  nand (_04083_, _04082_, _04062_);
  nand (_04084_, _04083_, _14374_);
  nand (_04085_, _04084_, _14483_);
  or (_04087_, _04085_, _04028_);
  and (_04355_, _04087_, _04026_);
  or (_04088_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand (_04089_, _07493_, _14168_);
  and (_04090_, _04089_, _06989_);
  and (_04360_, _04090_, _04088_);
  or (_04091_, _01319_, _12278_);
  nand (_04092_, _01319_, _03882_);
  and (_04093_, _04092_, _06983_);
  and (_04094_, _04093_, _04091_);
  nor (_04095_, _06484_, _03882_);
  and (_04096_, _01318_, _06539_);
  nand (_04097_, _04096_, _06968_);
  or (_04098_, _04096_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_04100_, _04098_, _06485_);
  and (_04101_, _04100_, _04097_);
  or (_04102_, _04101_, _04095_);
  or (_04103_, _04102_, _04094_);
  and (_04485_, _04103_, _06989_);
  nor (_04487_, _11841_, rst);
  nor (_04105_, _09614_, _07118_);
  and (_04106_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_04107_, _04106_, _06982_);
  or (_04108_, _04107_, _04105_);
  or (_04109_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_04110_, _04109_, _06989_);
  and (_04524_, _04110_, _04108_);
  nand (_04111_, _06513_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_04113_, _04111_, _06538_);
  or (_04115_, _04113_, _01556_);
  and (_04116_, _04115_, _00867_);
  nand (_04118_, _00867_, _06513_);
  and (_04119_, _04118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_04120_, _04119_, _07459_);
  or (_04121_, _04120_, _04116_);
  nand (_04123_, _10970_, _07459_);
  and (_04124_, _04123_, _06989_);
  and (_04527_, _04124_, _04121_);
  and (_04125_, _00791_, _06539_);
  nand (_04126_, _04125_, _06968_);
  or (_04127_, _04125_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_04128_, _04127_, _00803_);
  and (_04129_, _04128_, _04126_);
  nor (_04131_, _00803_, _07040_);
  or (_04132_, _04131_, _04129_);
  and (_04529_, _04132_, _06989_);
  and (_04133_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_04135_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or (_04136_, _04135_, _04133_);
  and (_04532_, _04136_, _06989_);
  and (_04138_, _00708_, _06539_);
  nand (_04139_, _04138_, _06968_);
  or (_04140_, _04138_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_04141_, _04140_, _00715_);
  and (_04142_, _04141_, _04139_);
  nor (_04143_, _00715_, _07040_);
  or (_04144_, _04143_, _04142_);
  and (_04539_, _04144_, _06989_);
  and (_04145_, _08436_, _06501_);
  nand (_04146_, _04145_, _06968_);
  or (_04147_, _04145_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_04148_, _04147_, _02635_);
  and (_04149_, _04148_, _04146_);
  nor (_04150_, _07317_, _02635_);
  or (_04151_, _04150_, _04149_);
  and (_04544_, _04151_, _06989_);
  and (_04152_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_04153_, _04152_, _00760_);
  and (_04154_, _04153_, _06501_);
  nand (_04155_, _00764_, _06501_);
  and (_04156_, _04155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_04157_, _04156_, _06987_);
  or (_04158_, _04157_, _04154_);
  nand (_04159_, _11529_, _06987_);
  and (_04160_, _04159_, _06989_);
  and (_04547_, _04160_, _04158_);
  and (_04161_, _07089_, _06501_);
  nand (_04162_, _04161_, _06968_);
  or (_04163_, _04161_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_04164_, _04163_, _02635_);
  and (_04165_, _04164_, _04162_);
  nor (_04166_, _09008_, _02635_);
  or (_04167_, _04166_, _04165_);
  and (_04550_, _04167_, _06989_);
  and (_04168_, _06979_, _06501_);
  nand (_04169_, _04168_, _06968_);
  or (_04170_, _04168_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_04171_, _04170_, _02635_);
  and (_04172_, _04171_, _04169_);
  and (_04173_, _09599_, _06987_);
  or (_04174_, _04173_, _04172_);
  and (_04555_, _04174_, _06989_);
  and (_04175_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_04176_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor (_04177_, _04176_, _04175_);
  nor (_04178_, _04177_, _13986_);
  and (_04179_, _03503_, _07429_);
  or (_04180_, _04179_, _04178_);
  and (_04181_, _13986_, _09392_);
  and (_04182_, _04181_, _07119_);
  or (_04183_, _04182_, _04180_);
  and (_04557_, _04183_, _06989_);
  and (_04184_, _04006_, _07429_);
  and (_04185_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_04186_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_04188_, _04186_, _04185_);
  nor (_04189_, _04188_, _13986_);
  and (_04190_, _03503_, _07410_);
  or (_04191_, _04190_, _04189_);
  or (_04192_, _04191_, _04184_);
  and (_04560_, _04192_, _06989_);
  and (_04193_, _04006_, _07410_);
  and (_04194_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_04195_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_04197_, _04195_, _04194_);
  nor (_04198_, _04197_, _13986_);
  and (_04200_, _03503_, _11821_);
  or (_04201_, _04200_, _04198_);
  or (_04202_, _04201_, _04193_);
  and (_04563_, _04202_, _06989_);
  and (_04203_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_04204_, _08139_, _01188_);
  or (_04205_, _04204_, _04203_);
  and (_04566_, _04205_, _06989_);
  and (_04208_, _11986_, _08346_);
  or (_04209_, _12134_, _12131_);
  and (_04210_, _12171_, _12135_);
  and (_04212_, _04210_, _04209_);
  nor (_04213_, _12036_, _11988_);
  and (_04215_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_04217_, _12176_, _11718_);
  or (_04218_, _04217_, _04215_);
  or (_04220_, _04218_, _04213_);
  nor (_04221_, _04220_, _04212_);
  nand (_04222_, _04221_, _11964_);
  or (_04223_, _04222_, _04208_);
  nor (_04225_, _08595_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_04226_, _04225_, _12673_);
  or (_04228_, _04226_, _11964_);
  and (_04229_, _04228_, _06989_);
  and (_04568_, _04229_, _04223_);
  and (_04570_, _04024_, _14377_);
  or (_04230_, _11964_, _08596_);
  and (_04231_, _11986_, _08433_);
  and (_04232_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_04234_, _12061_, _11988_);
  and (_04235_, _12783_, _11514_);
  or (_04237_, _04235_, _04234_);
  or (_04238_, _04237_, _04232_);
  or (_04239_, _12064_, _12065_);
  nor (_04240_, _04239_, _12129_);
  and (_04241_, _04239_, _12129_);
  or (_04242_, _04241_, _04240_);
  and (_04243_, _04242_, _12722_);
  or (_04244_, _04243_, _04238_);
  or (_04245_, _04244_, _04231_);
  or (_04246_, _04245_, _12781_);
  and (_04247_, _04246_, _06989_);
  and (_04572_, _04247_, _04230_);
  and (_04248_, _12691_, _08588_);
  and (_04249_, _11986_, _01898_);
  and (_04250_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_04251_, _11988_, _11207_);
  and (_04252_, _12783_, _11842_);
  or (_04253_, _04252_, _04251_);
  or (_04254_, _04253_, _04250_);
  nor (_04255_, _12126_, _12124_);
  nor (_04256_, _04255_, _12127_);
  and (_04257_, _04256_, _12722_);
  or (_04258_, _04257_, _04254_);
  or (_04259_, _04258_, _04249_);
  and (_04260_, _04259_, _11964_);
  or (_04261_, _04260_, _04248_);
  and (_04582_, _04261_, _06989_);
  and (_04262_, _12691_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_04263_, _11986_, _08030_);
  or (_04264_, _12120_, _12118_);
  and (_04265_, _12171_, _12123_);
  and (_04266_, _04265_, _04264_);
  and (_04267_, _12091_, _11974_);
  and (_04268_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_04269_, _12176_, _11744_);
  or (_04270_, _04269_, _04268_);
  or (_04271_, _04270_, _04267_);
  or (_04272_, _04271_, _04266_);
  or (_04273_, _04272_, _04263_);
  and (_04274_, _04273_, _11964_);
  or (_04275_, _04274_, _04262_);
  and (_04585_, _04275_, _06989_);
  and (_04276_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_04277_, _04276_, _09580_);
  nor (_04278_, _07140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor (_04279_, _04278_, _07141_);
  or (_04280_, _04279_, _04277_);
  and (_04281_, _04280_, _09574_);
  and (_04283_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_04284_, _04283_, _07046_);
  or (_04285_, _04284_, _04281_);
  not (_04286_, _07046_);
  or (_04287_, _04286_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_04288_, _04287_, _09590_);
  and (_04289_, _04288_, _04285_);
  nor (_04290_, _10970_, _09590_);
  or (_04291_, _04290_, _04289_);
  and (_04592_, _04291_, _06989_);
  nor (_04292_, _07118_, _09590_);
  and (_04293_, _07071_, _07063_);
  nor (_04294_, _04293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor (_04295_, _04294_, _07140_);
  or (_04296_, _04295_, _07077_);
  and (_04297_, _07147_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_04298_, _04297_, _07066_);
  or (_04299_, _04298_, _04296_);
  or (_04300_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_04301_, _04300_, _07051_);
  and (_04302_, _04301_, _04299_);
  and (_04303_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_04304_, _04303_, _04302_);
  or (_04305_, _04304_, _04292_);
  and (_04594_, _04305_, _06989_);
  nand (_04799_, _11794_, _06989_);
  nand (_04801_, _11739_, _06989_);
  nand (_04805_, _11851_, _06989_);
  nor (_04813_, _11548_, rst);
  nor (_04815_, _11697_, rst);
  nor (_04817_, _11682_, rst);
  nor (_04819_, _11626_, rst);
  nor (_04307_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not (_04308_, _04307_);
  and (_04309_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_04310_, _04309_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04311_, _04309_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04312_, _04311_, _04310_);
  not (_04313_, _04312_);
  and (_04314_, _04310_, _01350_);
  nor (_04315_, _04310_, _01350_);
  nor (_04316_, _04315_, _04314_);
  nor (_04317_, _04316_, _08593_);
  and (_04318_, _04316_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_04319_, _04318_, _04317_);
  nor (_04320_, _04319_, _04313_);
  and (_04321_, _04316_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_04322_, _04316_, _08621_);
  nor (_04323_, _04322_, _04321_);
  nor (_04324_, _04323_, _04312_);
  nor (_04325_, _04324_, _04320_);
  nor (_04326_, _04325_, _04308_);
  and (_04327_, _13921_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not (_04328_, _04327_);
  not (_04329_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor (_04330_, _04316_, _04329_);
  and (_04331_, _04316_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_04332_, _04331_, _04330_);
  nor (_04333_, _04332_, _04313_);
  and (_04335_, _04316_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_04336_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_04337_, _04316_, _04336_);
  nor (_04338_, _04337_, _04335_);
  nor (_04340_, _04338_, _04312_);
  nor (_04341_, _04340_, _04333_);
  nor (_04342_, _04341_, _04328_);
  nor (_04343_, _04342_, _04326_);
  not (_04344_, _04309_);
  nor (_04345_, _04316_, _08647_);
  and (_04346_, _04316_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_04347_, _04346_, _04345_);
  nor (_04348_, _04347_, _04313_);
  and (_04349_, _04316_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_04350_, _04316_, _09234_);
  nor (_04351_, _04350_, _04349_);
  nor (_04352_, _04351_, _04312_);
  nor (_04354_, _04352_, _04348_);
  nor (_04356_, _04354_, _04344_);
  and (_04357_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _12949_);
  not (_04358_, _04357_);
  not (_04359_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor (_04361_, _04316_, _04359_);
  and (_04362_, _04316_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_04363_, _04362_, _04361_);
  nor (_04364_, _04363_, _04313_);
  and (_04365_, _04316_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not (_04366_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_04367_, _04316_, _04366_);
  nor (_04368_, _04367_, _04365_);
  nor (_04369_, _04368_, _04312_);
  nor (_04370_, _04369_, _04364_);
  nor (_04371_, _04370_, _04358_);
  nor (_04372_, _04371_, _04356_);
  and (_04373_, _04372_, _04343_);
  and (_04374_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_04375_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_04376_, _04375_, _04374_);
  and (_04377_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_04378_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_04379_, _04378_, _04377_);
  and (_04380_, _04379_, _04376_);
  and (_04381_, _04380_, _04313_);
  not (_04382_, _04316_);
  and (_04383_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_04384_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_04385_, _04384_, _04383_);
  and (_04386_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_04387_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_04388_, _04387_, _04386_);
  and (_04389_, _04388_, _04385_);
  and (_04390_, _04389_, _04312_);
  or (_04391_, _04390_, _04382_);
  nor (_04392_, _04391_, _04381_);
  and (_04393_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_04394_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_04395_, _04394_, _04393_);
  and (_04396_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_04397_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_04398_, _04397_, _04396_);
  and (_04399_, _04398_, _04395_);
  nor (_04400_, _04399_, _04312_);
  and (_04401_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_04402_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_04403_, _04402_, _04401_);
  and (_04404_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_04405_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_04406_, _04405_, _04404_);
  and (_04407_, _04406_, _04403_);
  nor (_04408_, _04407_, _04313_);
  or (_04409_, _04408_, _04400_);
  and (_04410_, _04409_, _04382_);
  nor (_04411_, _04410_, _04392_);
  nor (_04412_, _04411_, _04373_);
  or (_04413_, _04412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_04414_, _04412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04415_, _04414_, _04413_);
  not (_04416_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_04417_, _04373_);
  and (_04418_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_04419_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_04420_, _04419_, _04418_);
  and (_04421_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_04422_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_04423_, _04422_, _04421_);
  and (_04424_, _04423_, _04420_);
  and (_04425_, _04424_, _04313_);
  and (_04426_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_04427_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_04428_, _04427_, _04426_);
  and (_04429_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_04430_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_04431_, _04430_, _04429_);
  and (_04432_, _04431_, _04428_);
  and (_04433_, _04432_, _04312_);
  nor (_04434_, _04433_, _04425_);
  nor (_04435_, _04434_, _04382_);
  and (_04436_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_04437_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_04438_, _04437_, _04436_);
  and (_04439_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_04440_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_04441_, _04440_, _04439_);
  and (_04442_, _04441_, _04438_);
  and (_04443_, _04442_, _04313_);
  and (_04444_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_04445_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_04446_, _04445_, _04444_);
  and (_04447_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_04448_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_04449_, _04448_, _04447_);
  and (_04450_, _04449_, _04446_);
  and (_04451_, _04450_, _04312_);
  nor (_04452_, _04451_, _04443_);
  nor (_04453_, _04452_, _04316_);
  nor (_04454_, _04453_, _04435_);
  and (_04455_, _04454_, _04417_);
  and (_04456_, _04455_, _04416_);
  nor (_04457_, _04455_, _04416_);
  or (_04458_, _04457_, _04456_);
  or (_04459_, _04458_, _04415_);
  and (_04460_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_04461_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_04462_, _04461_, _04460_);
  and (_04463_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_04464_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_04465_, _04464_, _04463_);
  and (_04466_, _04465_, _04462_);
  and (_04467_, _04466_, _04313_);
  and (_04468_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_04469_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_04470_, _04469_, _04468_);
  and (_04471_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_04472_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_04473_, _04472_, _04471_);
  and (_04474_, _04473_, _04470_);
  and (_04475_, _04474_, _04312_);
  nor (_04476_, _04475_, _04467_);
  nor (_04477_, _04476_, _04382_);
  and (_04478_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_04479_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_04480_, _04479_, _04478_);
  and (_04481_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_04482_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_04483_, _04482_, _04481_);
  and (_04484_, _04483_, _04480_);
  and (_04486_, _04484_, _04313_);
  and (_04488_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_04489_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_04490_, _04489_, _04488_);
  and (_04491_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_04492_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_04493_, _04492_, _04491_);
  and (_04494_, _04493_, _04490_);
  and (_04495_, _04494_, _04312_);
  nor (_04496_, _04495_, _04486_);
  nor (_04497_, _04496_, _04316_);
  nor (_04498_, _04497_, _04477_);
  and (_04499_, _04498_, _04417_);
  or (_04500_, _04499_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_04501_, _04499_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04502_, _04501_, _04500_);
  not (_04503_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04504_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_04505_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_04506_, _04505_, _04504_);
  and (_04507_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_04508_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_04509_, _04508_, _04507_);
  and (_04510_, _04509_, _04506_);
  and (_04511_, _04510_, _04313_);
  and (_04512_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_04513_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_04514_, _04513_, _04512_);
  and (_04515_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_04516_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_04517_, _04516_, _04515_);
  and (_04518_, _04517_, _04514_);
  and (_04519_, _04518_, _04312_);
  or (_04520_, _04519_, _04382_);
  nor (_04521_, _04520_, _04511_);
  and (_04522_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_04523_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_04525_, _04523_, _04522_);
  and (_04526_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_04528_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_04530_, _04528_, _04526_);
  and (_04531_, _04530_, _04525_);
  nor (_04533_, _04531_, _04312_);
  and (_04534_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_04535_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_04536_, _04535_, _04534_);
  and (_04537_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_04538_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_04540_, _04538_, _04537_);
  and (_04541_, _04540_, _04536_);
  nor (_04542_, _04541_, _04313_);
  or (_04543_, _04542_, _04533_);
  and (_04545_, _04543_, _04382_);
  nor (_04546_, _04545_, _04521_);
  nor (_04548_, _04546_, _04373_);
  nor (_04549_, _04548_, _04503_);
  and (_04551_, _04548_, _04503_);
  or (_04552_, _04551_, _04549_);
  or (_04553_, _04552_, _04502_);
  or (_04554_, _04553_, _04459_);
  and (_04556_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_04558_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_04559_, _04558_, _04556_);
  and (_04561_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_04562_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_04564_, _04562_, _04561_);
  and (_04565_, _04564_, _04559_);
  and (_04567_, _04565_, _04313_);
  and (_04569_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_04571_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_04573_, _04571_, _04569_);
  and (_04574_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_04575_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_04576_, _04575_, _04574_);
  and (_04577_, _04576_, _04573_);
  and (_04578_, _04577_, _04312_);
  or (_04579_, _04578_, _04316_);
  nor (_04580_, _04579_, _04567_);
  and (_04581_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_04583_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_04584_, _04583_, _04581_);
  and (_04586_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_04587_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_04588_, _04587_, _04586_);
  and (_04589_, _04588_, _04584_);
  nor (_04590_, _04589_, _04312_);
  and (_04591_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_04593_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_04595_, _04593_, _04591_);
  and (_04596_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_04597_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_04598_, _04597_, _04596_);
  and (_04599_, _04598_, _04595_);
  nor (_04600_, _04599_, _04313_);
  or (_04601_, _04600_, _04590_);
  and (_04602_, _04601_, _04316_);
  nor (_04603_, _04602_, _04580_);
  nor (_04604_, _04603_, _04373_);
  or (_04605_, _04604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_04606_, _04604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_04607_, _04606_, _04605_);
  not (_04608_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_04609_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_04610_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_04611_, _04610_, _04609_);
  and (_04612_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_04613_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_04614_, _04613_, _04612_);
  and (_04615_, _04614_, _04611_);
  and (_04616_, _04615_, _04313_);
  and (_04617_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_04618_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_04619_, _04618_, _04617_);
  and (_04620_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_04621_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_04622_, _04621_, _04620_);
  and (_04623_, _04622_, _04619_);
  and (_04624_, _04623_, _04312_);
  or (_04625_, _04624_, _04382_);
  nor (_04626_, _04625_, _04616_);
  and (_04627_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_04628_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_04629_, _04628_, _04627_);
  and (_04630_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_04631_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_04632_, _04631_, _04630_);
  and (_04633_, _04632_, _04629_);
  and (_04634_, _04633_, _04313_);
  and (_04635_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_04636_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_04637_, _04636_, _04635_);
  and (_04638_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_04639_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_04640_, _04639_, _04638_);
  and (_04641_, _04640_, _04637_);
  and (_04642_, _04641_, _04312_);
  or (_04643_, _04642_, _04316_);
  nor (_04644_, _04643_, _04634_);
  nor (_04645_, _04644_, _04626_);
  nor (_04646_, _04645_, _04373_);
  and (_04647_, _04646_, _04608_);
  nor (_04648_, _04646_, _04608_);
  or (_04649_, _04648_, _04647_);
  or (_04650_, _04649_, _04607_);
  and (_04651_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_04652_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_04653_, _04652_, _04651_);
  and (_04654_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_04655_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_04656_, _04655_, _04654_);
  and (_04657_, _04656_, _04653_);
  and (_04658_, _04657_, _04313_);
  and (_04659_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_04660_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_04661_, _04660_, _04659_);
  and (_04662_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_04663_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_04664_, _04663_, _04662_);
  and (_04665_, _04664_, _04661_);
  and (_04666_, _04665_, _04312_);
  or (_04667_, _04666_, _04382_);
  nor (_04668_, _04667_, _04658_);
  and (_04669_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_04670_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor (_04671_, _04670_, _04669_);
  and (_04672_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_04673_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_04674_, _04673_, _04672_);
  and (_04675_, _04674_, _04671_);
  and (_04676_, _04675_, _04313_);
  and (_04677_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_04678_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_04679_, _04678_, _04677_);
  and (_04680_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_04681_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_04682_, _04681_, _04680_);
  and (_04683_, _04682_, _04679_);
  and (_04684_, _04683_, _04312_);
  or (_04685_, _04684_, _04316_);
  nor (_04686_, _04685_, _04676_);
  nor (_04687_, _04686_, _04668_);
  nor (_04688_, _04687_, _04373_);
  nor (_04689_, _04688_, _01149_);
  and (_04690_, _04688_, _01149_);
  or (_04691_, _04690_, _04689_);
  and (_04692_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_04693_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_04694_, _04693_, _04692_);
  and (_04695_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_04696_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_04697_, _04696_, _04695_);
  and (_04698_, _04697_, _04694_);
  and (_04699_, _04698_, _04313_);
  and (_04700_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_04701_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_04702_, _04701_, _04700_);
  and (_04703_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_04704_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_04705_, _04704_, _04703_);
  and (_04706_, _04705_, _04702_);
  and (_04707_, _04706_, _04312_);
  or (_04708_, _04707_, _04316_);
  nor (_04709_, _04708_, _04699_);
  and (_04710_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_04711_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_04712_, _04711_, _04710_);
  and (_04713_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_04714_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_04715_, _04714_, _04713_);
  and (_04716_, _04715_, _04712_);
  nor (_04717_, _04716_, _04312_);
  and (_04718_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_04719_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_04720_, _04719_, _04718_);
  and (_04721_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_04722_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_04723_, _04722_, _04721_);
  and (_04724_, _04723_, _04720_);
  nor (_04725_, _04724_, _04313_);
  or (_04726_, _04725_, _04717_);
  and (_04727_, _04726_, _04316_);
  nor (_04728_, _04727_, _04709_);
  nor (_04729_, _04728_, _04373_);
  nor (_04730_, _04729_, _01188_);
  and (_04731_, _04729_, _01188_);
  or (_04732_, _04731_, _04730_);
  or (_04733_, _04732_, _04691_);
  or (_04734_, _04733_, _04650_);
  or (_04735_, _04734_, _04554_);
  and (_04736_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04737_, _04736_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04738_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_04739_, _04738_, _04737_);
  and (_04740_, _04739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and (_04741_, _04740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_04742_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_04743_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_04744_, _04743_, _04742_);
  and (_04745_, _04744_, _04741_);
  and (_04746_, _04745_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_04747_, _04746_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_04748_, _04747_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and (_04749_, _04748_, _00655_);
  nor (_04750_, _04748_, _00655_);
  or (_04751_, _04750_, _04749_);
  nor (_04752_, _04751_, _00619_);
  and (_04753_, _04751_, _00619_);
  or (_04754_, _04753_, _04752_);
  and (_04755_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_04756_, _04755_, _04738_);
  and (_04757_, _04756_, _04737_);
  and (_04758_, _04757_, _04744_);
  and (_04759_, _04758_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_04760_, _04759_, _00683_);
  and (_04761_, _04759_, _00683_);
  or (_04762_, _04761_, _04760_);
  nor (_04763_, _04762_, _01686_);
  and (_04764_, _04762_, _01686_);
  or (_04765_, _04764_, _04763_);
  nor (_04766_, _04745_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_04767_, _04766_, _04746_);
  or (_04768_, _04767_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_04769_, _04767_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and (_04770_, _04769_, _04768_);
  or (_04771_, _04770_, _04765_);
  nor (_04772_, _04747_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04773_, _04772_, _04748_);
  or (_04774_, _04773_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_04775_, _04773_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_04776_, _04775_, _04774_);
  or (_04777_, _04776_, _04771_);
  or (_04778_, _04777_, _04754_);
  and (_04779_, _12949_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04780_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08593_);
  nor (_04781_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_04782_, _04781_, _04780_);
  and (_04783_, _04782_, _04779_);
  nor (_04784_, _04783_, _13921_);
  nor (_04785_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_04786_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04329_);
  or (_04787_, _04786_, _01231_);
  nor (_04788_, _04787_, _04785_);
  and (_04789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04336_);
  nor (_04790_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_04791_, _04790_, _04789_);
  and (_04792_, _04791_, _01231_);
  nor (_04793_, _04792_, _04788_);
  nor (_04794_, _04793_, _12949_);
  nor (_04795_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04796_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_04797_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08621_);
  nor (_04798_, _04797_, _04796_);
  and (_04800_, _04798_, _04795_);
  nor (_04802_, _04800_, _04794_);
  and (_04803_, _04802_, _04784_);
  nor (_04804_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_04806_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04359_);
  or (_04807_, _04806_, _01231_);
  nor (_04808_, _04807_, _04804_);
  and (_04809_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04366_);
  nor (_04810_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_04811_, _04810_, _04809_);
  and (_04812_, _04811_, _01231_);
  nor (_04814_, _04812_, _04808_);
  nor (_04816_, _04814_, _12949_);
  nor (_04818_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_04820_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _09234_);
  nor (_04821_, _04820_, _04818_);
  and (_04822_, _04821_, _04795_);
  and (_04823_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08647_);
  nor (_04824_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_04825_, _04824_, _04823_);
  and (_04826_, _04825_, _04779_);
  or (_04827_, _04826_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_04828_, _04827_, _04822_);
  nor (_04829_, _04828_, _04816_);
  nor (_04830_, _04829_, _04803_);
  nor (_04831_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04832_, _09847_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04833_, _04832_, _04831_);
  and (_04834_, _04833_, _04795_);
  nor (_04836_, _04834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_04837_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04838_, _10325_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04839_, _04838_, _04837_);
  and (_04840_, _04839_, _04779_);
  not (_04841_, _04840_);
  nor (_04842_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04844_, _10100_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04845_, _04844_, _04842_);
  and (_04846_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _01231_);
  and (_04847_, _04846_, _04845_);
  nor (_04849_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04850_, _10537_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04851_, _04850_, _04849_);
  and (_04852_, _04851_, _04736_);
  nor (_04853_, _04852_, _04847_);
  and (_04854_, _04853_, _04841_);
  and (_04855_, _04854_, _04836_);
  nor (_04856_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04857_, _10759_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04858_, _04857_, _04856_);
  and (_04859_, _04858_, _04795_);
  nor (_04860_, _04859_, _01350_);
  nor (_04861_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04862_, _12513_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04863_, _04862_, _04861_);
  and (_04864_, _04863_, _04779_);
  not (_04865_, _04864_);
  nor (_04866_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04867_, _12209_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04868_, _04867_, _04866_);
  and (_04869_, _04868_, _04846_);
  nor (_04870_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04871_, _12899_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04873_, _04871_, _04870_);
  and (_04874_, _04873_, _04736_);
  nor (_04875_, _04874_, _04869_);
  and (_04876_, _04875_, _04865_);
  and (_04877_, _04876_, _04860_);
  nor (_04878_, _04877_, _04855_);
  and (_04879_, _04878_, _04830_);
  nor (_04880_, _04879_, _01144_);
  and (_04881_, _04879_, _01144_);
  or (_04882_, _04881_, _04880_);
  nor (_04883_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04884_, _10113_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04885_, _04884_, _04883_);
  and (_04886_, _04885_, _04846_);
  nor (_04887_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04888_, _10338_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04890_, _04888_, _04887_);
  and (_04891_, _04890_, _04779_);
  nor (_04892_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04893_, _09860_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04894_, _04893_, _04892_);
  and (_04895_, _04894_, _04795_);
  nor (_04897_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04898_, _10548_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04899_, _04898_, _04897_);
  and (_04900_, _04899_, _04736_);
  or (_04901_, _04900_, _04895_);
  or (_04902_, _04901_, _04891_);
  or (_04903_, _04902_, _04886_);
  and (_04904_, _04903_, _01350_);
  nor (_04905_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04906_, _12225_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04907_, _04906_, _04905_);
  and (_04908_, _04907_, _04846_);
  nor (_04910_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04911_, _12524_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04912_, _04911_, _04910_);
  and (_04913_, _04912_, _04779_);
  nor (_04914_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04915_, _10771_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04917_, _04915_, _04914_);
  and (_04918_, _04917_, _04795_);
  nor (_04919_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_04921_, _12914_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04923_, _04921_, _04919_);
  and (_04925_, _04923_, _04736_);
  or (_04926_, _04925_, _04918_);
  or (_04927_, _04926_, _04913_);
  or (_04928_, _04927_, _04908_);
  and (_04929_, _04928_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_04930_, _04929_, _04904_);
  and (_04931_, _04930_, _04830_);
  nor (_04932_, _04931_, _01227_);
  and (_04933_, _04931_, _01227_);
  or (_04934_, _04933_, _04932_);
  or (_04935_, _04934_, _04882_);
  and (_04936_, _04741_, _04742_);
  and (_04937_, _04936_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_04938_, _04937_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_04939_, _04937_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_04940_, _04939_, _04938_);
  nor (_04942_, _04940_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_04944_, _04940_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_04946_, _04944_, _04942_);
  nor (_04947_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_04948_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08682_);
  nor (_04949_, _04948_, _04947_);
  and (_04950_, _04949_, _04846_);
  nor (_04951_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_04952_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08687_);
  nor (_04953_, _04952_, _04951_);
  and (_04954_, _04953_, _04736_);
  nor (_04955_, _04954_, _04950_);
  nor (_04956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_04957_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08693_);
  nor (_04958_, _04957_, _04956_);
  and (_04959_, _04958_, _04779_);
  nor (_04960_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_04961_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08698_);
  nor (_04962_, _04961_, _04960_);
  and (_04963_, _04962_, _04795_);
  nor (_04964_, _04963_, _04959_);
  and (_04965_, _04964_, _04955_);
  nor (_04966_, _04965_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_04967_, _04966_);
  nor (_04968_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_04969_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08663_);
  nor (_04970_, _04969_, _04968_);
  and (_04971_, _04970_, _04846_);
  nor (_04972_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_04973_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08669_);
  nor (_04974_, _04973_, _04972_);
  and (_04975_, _04974_, _04779_);
  nor (_04976_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_04977_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08674_);
  nor (_04979_, _04977_, _04976_);
  and (_04980_, _04979_, _04795_);
  nor (_04981_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_04982_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08657_);
  nor (_04983_, _04982_, _04981_);
  and (_04984_, _04983_, _04736_);
  or (_04985_, _04984_, _04980_);
  or (_04986_, _04985_, _04975_);
  nor (_04987_, _04986_, _04971_);
  or (_04988_, _04987_, _01350_);
  and (_04989_, _04988_, _04967_);
  not (_04991_, _04989_);
  and (_04992_, _04991_, _04830_);
  nor (_04993_, _04992_, _01220_);
  and (_04994_, _04992_, _01220_);
  or (_04995_, _04994_, _04993_);
  or (_04996_, _04995_, _04946_);
  or (_04997_, _04996_, _04935_);
  or (_04998_, _04997_, _04778_);
  or (_04999_, _04998_, _04735_);
  or (_05000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  not (_05001_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_05003_, _05001_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_05004_, _05003_, _05000_);
  and (_05005_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _04503_);
  and (_05006_, _05005_, _05004_);
  or (_05007_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05008_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05009_, _05001_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_05010_, _05009_, _05008_);
  and (_05011_, _05010_, _05007_);
  or (_05012_, _05011_, _05006_);
  not (_05013_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_05014_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_05015_, _05014_, _04503_);
  nor (_05016_, _05015_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_05017_, _05015_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_05019_, _05017_, _05016_);
  and (_05020_, _05019_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_05021_, _05014_, _04503_);
  nor (_05022_, _05021_, _05015_);
  or (_05023_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _08615_);
  nand (_05024_, _05023_, _05022_);
  or (_05025_, _05024_, _05020_);
  and (_05026_, _05025_, _05013_);
  nand (_05027_, _05019_, _04336_);
  or (_05028_, _05019_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_05029_, _05028_, _05027_);
  or (_05030_, _05022_, _05029_);
  and (_05031_, _05030_, _05026_);
  or (_05032_, _05031_, _05012_);
  and (_05034_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05035_, _05001_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05036_, _05035_, _05034_);
  and (_05037_, _05036_, _04503_);
  and (_05038_, _05001_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_05039_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_05040_, _05039_, _05038_);
  and (_05041_, _05040_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05042_, _05041_, _05037_);
  and (_05043_, _05042_, _05013_);
  and (_05044_, _05008_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_05045_, _05044_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_05046_, _05044_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_05047_, _05046_, _05045_);
  nand (_05048_, _05047_, _08593_);
  and (_05049_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_05050_, _05049_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_05051_, _05050_, _05044_);
  and (_05052_, _05051_, _05000_);
  and (_05053_, _05052_, _05048_);
  nand (_05054_, _05047_, _08621_);
  not (_05055_, _05051_);
  or (_05056_, _05047_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_05057_, _05056_, _05055_);
  and (_05058_, _05057_, _05054_);
  or (_05059_, _05058_, _05053_);
  and (_05060_, _05059_, _05043_);
  nand (_05061_, _05047_, _04329_);
  or (_05062_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_05063_, _05062_, _05051_);
  and (_05064_, _05063_, _05061_);
  nand (_05065_, _05047_, _04336_);
  or (_05066_, _05047_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_05067_, _05066_, _05055_);
  and (_05068_, _05067_, _05065_);
  or (_05069_, _05068_, _05064_);
  and (_05070_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_05071_, _05001_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_05072_, _05071_, _04503_);
  or (_05073_, _05072_, _05070_);
  or (_05074_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_05075_, _05001_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_05076_, _05075_, _05074_);
  or (_05077_, _05076_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05078_, _05077_, _05073_);
  and (_05079_, _05078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_05080_, _05040_, _05005_);
  or (_05081_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05082_, _05001_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05083_, _05082_, _05008_);
  and (_05084_, _05083_, _05081_);
  or (_05085_, _05084_, _05080_);
  and (_05086_, _05085_, _05079_);
  and (_05087_, _05086_, _05069_);
  or (_05088_, _05087_, _05060_);
  or (_05089_, _05085_, _05078_);
  and (_05090_, _05089_, _04416_);
  and (_05091_, _05090_, _05088_);
  and (_05092_, _05091_, _05032_);
  or (_05093_, _05013_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_05094_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05095_, _05094_, _05093_);
  or (_05096_, _05095_, _05019_);
  or (_05097_, _05013_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_05098_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_05099_, _05098_, _05097_);
  and (_05100_, _05099_, _05019_);
  nor (_05101_, _05100_, _05022_);
  and (_05102_, _05101_, _05096_);
  and (_05103_, _05019_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_05104_, _05038_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_05105_, _05104_, _05103_);
  and (_05106_, _05019_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_05107_, _05071_, _05013_);
  or (_05108_, _05107_, _05106_);
  and (_05109_, _05108_, _05022_);
  and (_05110_, _05109_, _05105_);
  or (_05111_, _05110_, _05102_);
  nand (_05112_, _05047_, _04359_);
  or (_05113_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_05114_, _05113_, _05112_);
  or (_05115_, _05114_, _05055_);
  or (_05116_, _05047_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_05117_, _05047_, _04366_);
  and (_05118_, _05117_, _05116_);
  or (_05119_, _05118_, _05051_);
  and (_05120_, _05119_, _05115_);
  or (_05121_, _05120_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_05122_, _05047_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_05123_, _05047_, _08639_);
  or (_05124_, _05123_, _05122_);
  and (_05125_, _05124_, _05055_);
  nand (_05126_, _05047_, _08647_);
  or (_05127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_05128_, _05127_, _05051_);
  and (_05129_, _05128_, _05126_);
  or (_05130_, _05129_, _05013_);
  or (_05131_, _05130_, _05125_);
  or (_05132_, _05001_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_05133_, _05062_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05134_, _05133_, _05132_);
  or (_05135_, _05001_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_05136_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_05137_, _05136_, _04503_);
  and (_05138_, _05137_, _05135_);
  or (_05139_, _05138_, _05134_);
  and (_05140_, _05139_, _05049_);
  and (_05141_, _05013_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_05142_, _05004_, _04503_);
  or (_05143_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05144_, _05001_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05145_, _05144_, _05143_);
  or (_05146_, _05145_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05147_, _05146_, _05142_);
  and (_05148_, _05147_, _05141_);
  or (_05149_, _05148_, _05140_);
  and (_05150_, _05139_, _05013_);
  or (_05151_, _05150_, _05012_);
  and (_05152_, _05151_, _05149_);
  and (_05153_, _05152_, _05131_);
  and (_05154_, _05153_, _05121_);
  and (_05155_, _05154_, _05111_);
  or (_05156_, _05155_, _05092_);
  nor (_05157_, _04307_, _01231_);
  and (_05158_, _04795_, _13921_);
  nor (_05159_, _05158_, _05157_);
  and (_05160_, _05157_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_05161_, _05157_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_05162_, _05161_, _05160_);
  and (_05163_, _05162_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_05164_, _05162_, _08967_);
  or (_05165_, _05164_, _05163_);
  and (_05166_, _05165_, _04327_);
  or (_05167_, _05166_, _05159_);
  and (_05168_, _05162_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_05169_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_05170_, _05162_, _05169_);
  or (_05171_, _05170_, _05168_);
  and (_05172_, _05171_, _04309_);
  and (_05173_, _05162_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05174_, _05162_, _08608_);
  or (_05175_, _05174_, _05173_);
  and (_05176_, _05175_, _04307_);
  and (_05177_, _05162_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_05178_, _05162_, _08639_);
  or (_05179_, _05178_, _05177_);
  and (_05180_, _05179_, _04357_);
  or (_05181_, _05180_, _05176_);
  or (_05182_, _05181_, _05172_);
  or (_05183_, _05182_, _05167_);
  or (_05184_, _05162_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_05185_, _04780_, _04328_);
  nand (_05186_, _05185_, _05184_);
  nand (_05187_, _05186_, _05159_);
  or (_05188_, _05162_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_05189_, _04806_, _04344_);
  and (_05190_, _05189_, _05188_);
  or (_05191_, _05162_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_05192_, _04786_, _04308_);
  and (_05193_, _05192_, _05191_);
  or (_05194_, _05162_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_05195_, _04823_, _04358_);
  and (_05196_, _05195_, _05194_);
  or (_05197_, _05196_, _05193_);
  or (_05198_, _05197_, _05190_);
  or (_05199_, _05198_, _05187_);
  nor (_05200_, _04793_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_05201_, _04846_, _04782_);
  nor (_05202_, _05201_, _13921_);
  not (_05203_, _05202_);
  nor (_05204_, _05203_, _05200_);
  nor (_05205_, _04814_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_05206_, _04846_, _04825_);
  nor (_05207_, _05206_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not (_05208_, _05207_);
  nor (_05209_, _05208_, _05205_);
  nor (_05210_, _05209_, _05204_);
  not (_05211_, _05210_);
  or (_05212_, _01350_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_05213_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_05214_, _05213_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05215_, _05214_, _05212_);
  and (_05216_, _05215_, _04327_);
  and (_05217_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08967_);
  nor (_05218_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_05219_, _05218_, _05217_);
  and (_05220_, _05219_, _04310_);
  nor (_05221_, _05220_, _05216_);
  and (_05222_, _05221_, _05211_);
  not (_05223_, _08139_);
  nor (_05224_, _05223_, first_instr);
  nand (_05225_, _05224_, _04830_);
  nor (_05226_, _05225_, _05222_);
  and (_05227_, _05226_, _05199_);
  and (_05228_, _05227_, _05183_);
  and (_05229_, _05228_, _04417_);
  and (_05230_, _05229_, _05156_);
  nor (_05231_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05232_, _10057_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05233_, _05232_, _05231_);
  and (_05234_, _05233_, _04846_);
  nor (_05235_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05236_, _10290_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05237_, _05236_, _05235_);
  and (_05238_, _05237_, _04779_);
  nor (_05239_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05240_, _09807_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05241_, _05240_, _05239_);
  and (_05242_, _05241_, _04795_);
  nor (_05243_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05244_, _10501_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05245_, _05244_, _05243_);
  and (_05246_, _05245_, _04736_);
  or (_05247_, _05246_, _05242_);
  or (_05248_, _05247_, _05238_);
  or (_05249_, _05248_, _05234_);
  and (_05250_, _05249_, _01350_);
  nor (_05251_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05252_, _11260_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05253_, _05252_, _05251_);
  and (_05254_, _05253_, _04846_);
  nor (_05255_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05256_, _12474_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05257_, _05256_, _05255_);
  and (_05258_, _05257_, _04779_);
  nor (_05259_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05260_, _10710_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05261_, _05260_, _05259_);
  and (_05262_, _05261_, _04795_);
  nor (_05263_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05264_, _12861_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05265_, _05264_, _05263_);
  and (_05266_, _05265_, _04736_);
  or (_05267_, _05266_, _05262_);
  or (_05268_, _05267_, _05258_);
  or (_05269_, _05268_, _05254_);
  and (_05270_, _05269_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_05271_, _05270_, _05250_);
  and (_05272_, _05271_, _04830_);
  nor (_05273_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05274_, _10072_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05275_, _05274_, _05273_);
  and (_05276_, _05275_, _04846_);
  nor (_05277_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05278_, _10301_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05279_, _05278_, _05277_);
  and (_05280_, _05279_, _04779_);
  nor (_05281_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05282_, _09821_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05283_, _05282_, _05281_);
  and (_05284_, _05283_, _04795_);
  nor (_05285_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05286_, _10512_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05287_, _05286_, _05285_);
  and (_05288_, _05287_, _04736_);
  or (_05289_, _05288_, _05284_);
  or (_05290_, _05289_, _05280_);
  or (_05291_, _05290_, _05276_);
  and (_05292_, _05291_, _01350_);
  nor (_05293_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05294_, _12185_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05295_, _05294_, _05293_);
  and (_05296_, _05295_, _04846_);
  nor (_05297_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05298_, _12488_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05299_, _05298_, _05297_);
  and (_05300_, _05299_, _04779_);
  nor (_05301_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05302_, _10727_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05303_, _05302_, _05301_);
  and (_05304_, _05303_, _04795_);
  nor (_05305_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05306_, _12874_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05307_, _05306_, _05305_);
  and (_05308_, _05307_, _04736_);
  or (_05309_, _05308_, _05304_);
  or (_05310_, _05309_, _05300_);
  or (_05311_, _05310_, _05296_);
  and (_05312_, _05311_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_05313_, _05312_, _05292_);
  and (_05314_, _05313_, _04830_);
  nor (_05315_, _05314_, _05272_);
  nor (_05316_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05317_, _10474_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05318_, _05317_, _05316_);
  and (_05319_, _05318_, _04736_);
  nor (_05320_, _05319_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_05321_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05322_, _09771_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05323_, _05322_, _05321_);
  and (_05324_, _05323_, _04795_);
  not (_05325_, _05324_);
  nor (_05326_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05327_, _10016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05328_, _05327_, _05326_);
  and (_05329_, _05328_, _04846_);
  nor (_05330_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05331_, _10263_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05332_, _05331_, _05330_);
  and (_05333_, _05332_, _04779_);
  nor (_05334_, _05333_, _05329_);
  and (_05335_, _05334_, _05325_);
  and (_05336_, _05335_, _05320_);
  nor (_05337_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05338_, _12833_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05339_, _05338_, _05337_);
  and (_05340_, _05339_, _04736_);
  nor (_05341_, _05340_, _01350_);
  nor (_05342_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05343_, _10685_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05344_, _05343_, _05342_);
  and (_05345_, _05344_, _04795_);
  not (_05346_, _05345_);
  nor (_05347_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05348_, _11230_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05349_, _05348_, _05347_);
  and (_05350_, _05349_, _04846_);
  nor (_05351_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05352_, _12448_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05353_, _05352_, _05351_);
  and (_05354_, _05353_, _04779_);
  nor (_05355_, _05354_, _05350_);
  and (_05356_, _05355_, _05346_);
  and (_05357_, _05356_, _05341_);
  nor (_05358_, _05357_, _05336_);
  and (_05359_, _05358_, _04830_);
  not (_05360_, _05359_);
  nor (_05361_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05362_, _10037_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05363_, _05362_, _05361_);
  and (_05364_, _05363_, _04846_);
  nor (_05365_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05366_, _10276_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05367_, _05366_, _05365_);
  and (_05368_, _05367_, _04779_);
  nor (_05369_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05370_, _09792_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05371_, _05370_, _05369_);
  and (_05372_, _05371_, _04795_);
  nor (_05373_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05374_, _10489_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05375_, _05374_, _05373_);
  and (_05376_, _05375_, _04736_);
  or (_05377_, _05376_, _05372_);
  or (_05378_, _05377_, _05368_);
  or (_05379_, _05378_, _05364_);
  and (_05380_, _05379_, _01350_);
  nor (_05381_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05382_, _11247_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05383_, _05382_, _05381_);
  and (_05384_, _05383_, _04846_);
  nor (_05385_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05386_, _12463_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05387_, _05386_, _05385_);
  and (_05388_, _05387_, _04779_);
  nor (_05389_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05390_, _10699_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05391_, _05390_, _05389_);
  and (_05392_, _05391_, _04795_);
  nor (_05393_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05394_, _12848_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05395_, _05394_, _05393_);
  and (_05396_, _05395_, _04736_);
  or (_05397_, _05396_, _05392_);
  or (_05398_, _05397_, _05388_);
  or (_05399_, _05398_, _05384_);
  and (_05400_, _05399_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_05401_, _05400_, _05380_);
  nor (_05402_, _05401_, _05360_);
  and (_05403_, _05402_, _05315_);
  and (_05404_, _05403_, _05230_);
  and (property_invalid_ajmp, _05404_, _04999_);
  and (_05405_, _04736_, _01350_);
  nor (_05406_, _04736_, _01350_);
  nor (_05407_, _05406_, _05405_);
  not (_05408_, _05407_);
  and (_05409_, _04846_, _04839_);
  or (_05410_, _05409_, _05408_);
  and (_05411_, _04833_, _04736_);
  and (_05412_, _04845_, _04795_);
  and (_05413_, _04851_, _04779_);
  or (_05414_, _05413_, _05412_);
  or (_05415_, _05414_, _05411_);
  or (_05416_, _05415_, _05410_);
  and (_05417_, _04863_, _04846_);
  or (_05418_, _05417_, _05407_);
  and (_05419_, _04858_, _04736_);
  and (_05420_, _04868_, _04795_);
  and (_05421_, _04873_, _04779_);
  or (_05422_, _05421_, _05420_);
  or (_05423_, _05422_, _05419_);
  or (_05424_, _05423_, _05418_);
  nand (_05425_, _05424_, _05416_);
  nor (_05426_, _05425_, _05222_);
  nand (_05427_, _05426_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or (_05428_, _05426_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_05429_, _05428_, _05427_);
  nor (_05430_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05431_, _10315_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05432_, _05431_, _05430_);
  and (_05433_, _05432_, _04846_);
  or (_05434_, _05433_, _05408_);
  nor (_05435_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05436_, _09834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05437_, _05436_, _05435_);
  and (_05438_, _05437_, _04736_);
  nor (_05439_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05440_, _10086_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05441_, _05440_, _05439_);
  and (_05442_, _05441_, _04795_);
  nor (_05443_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05444_, _10525_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05445_, _05444_, _05443_);
  and (_05446_, _05445_, _04779_);
  or (_05447_, _05446_, _05442_);
  or (_05448_, _05447_, _05438_);
  or (_05449_, _05448_, _05434_);
  nor (_05450_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05451_, _12501_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05452_, _05451_, _05450_);
  and (_05453_, _05452_, _04846_);
  or (_05454_, _05453_, _05407_);
  nor (_05455_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05456_, _10743_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05457_, _05456_, _05455_);
  and (_05458_, _05457_, _04736_);
  nor (_05459_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05460_, _12196_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05461_, _05460_, _05459_);
  and (_05462_, _05461_, _04795_);
  nor (_05463_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05464_, _12887_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05465_, _05464_, _05463_);
  and (_05466_, _05465_, _04779_);
  or (_05467_, _05466_, _05462_);
  or (_05468_, _05467_, _05458_);
  or (_05469_, _05468_, _05454_);
  nand (_05470_, _05469_, _05449_);
  nor (_05471_, _05470_, _05222_);
  nand (_05472_, _05471_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_05473_, _05471_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_05474_, _05473_, _05472_);
  or (_05475_, _05474_, _05429_);
  and (_05476_, _04958_, _04846_);
  or (_05477_, _05476_, _05408_);
  and (_05478_, _04962_, _04736_);
  and (_05479_, _04949_, _04795_);
  and (_05480_, _04953_, _04779_);
  or (_05481_, _05480_, _05479_);
  or (_05482_, _05481_, _05478_);
  or (_05483_, _05482_, _05477_);
  and (_05484_, _04974_, _04846_);
  or (_05485_, _05484_, _05407_);
  and (_05486_, _04979_, _04736_);
  and (_05487_, _04970_, _04795_);
  and (_05488_, _04983_, _04779_);
  or (_05489_, _05488_, _05487_);
  or (_05490_, _05489_, _05486_);
  or (_05491_, _05490_, _05485_);
  nand (_05492_, _05491_, _05483_);
  nor (_05493_, _05492_, _05222_);
  nor (_05494_, _05493_, _01149_);
  and (_05495_, _05493_, _01149_);
  or (_05496_, _05495_, _05494_);
  not (_05497_, _05222_);
  and (_05498_, _04907_, _04795_);
  and (_05499_, _04923_, _04779_);
  and (_05500_, _04912_, _04846_);
  and (_05501_, _04917_, _04736_);
  or (_05502_, _05501_, _05500_);
  or (_05503_, _05502_, _05499_);
  or (_05504_, _05503_, _05498_);
  and (_05505_, _05504_, _05408_);
  and (_05506_, _04885_, _04795_);
  and (_05507_, _04899_, _04779_);
  and (_05508_, _04894_, _04736_);
  and (_05509_, _04890_, _04846_);
  or (_05510_, _05509_, _05508_);
  or (_05511_, _05510_, _05507_);
  or (_05512_, _05511_, _05506_);
  and (_05513_, _05512_, _05407_);
  or (_05514_, _05513_, _05505_);
  and (_05515_, _05514_, _05497_);
  and (_05516_, _05515_, _01188_);
  nor (_05517_, _05515_, _01188_);
  or (_05518_, _05517_, _05516_);
  or (_05519_, _05518_, _05496_);
  or (_05520_, _05519_, _05475_);
  and (_05521_, _05349_, _04795_);
  and (_05522_, _05339_, _04779_);
  and (_05523_, _05344_, _04736_);
  and (_05524_, _05353_, _04846_);
  or (_05525_, _05524_, _05523_);
  or (_05526_, _05525_, _05522_);
  or (_05527_, _05526_, _05521_);
  and (_05528_, _05527_, _05408_);
  and (_05529_, _05328_, _04795_);
  and (_05530_, _05318_, _04779_);
  and (_05531_, _05323_, _04736_);
  and (_05532_, _05332_, _04846_);
  or (_05533_, _05532_, _05531_);
  or (_05534_, _05533_, _05530_);
  or (_05535_, _05534_, _05529_);
  and (_05536_, _05535_, _05407_);
  or (_05537_, _05536_, _05528_);
  and (_05538_, _05537_, _05497_);
  nand (_05539_, _05538_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_05540_, _05538_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and (_05541_, _05540_, _05539_);
  and (_05542_, _05367_, _04846_);
  and (_05543_, _05375_, _04779_);
  and (_05544_, _05371_, _04736_);
  or (_05545_, _05544_, _05543_);
  or (_05546_, _05545_, _05542_);
  and (_05547_, _05363_, _04795_);
  or (_05548_, _05547_, _05408_);
  or (_05549_, _05548_, _05546_);
  and (_05550_, _05387_, _04846_);
  or (_05551_, _05550_, _05407_);
  and (_05552_, _05391_, _04736_);
  and (_05553_, _05383_, _04795_);
  and (_05554_, _05395_, _04779_);
  or (_05555_, _05554_, _05553_);
  or (_05556_, _05555_, _05552_);
  or (_05557_, _05556_, _05551_);
  nand (_05558_, _05557_, _05549_);
  nor (_05559_, _05558_, _05222_);
  nor (_05560_, _05559_, _05013_);
  and (_05561_, _05559_, _05013_);
  or (_05562_, _05561_, _05560_);
  or (_05563_, _05562_, _05541_);
  and (_05564_, _05253_, _04795_);
  and (_05565_, _05265_, _04779_);
  and (_05566_, _05261_, _04736_);
  and (_05567_, _05257_, _04846_);
  or (_05568_, _05567_, _05566_);
  or (_05569_, _05568_, _05565_);
  or (_05570_, _05569_, _05564_);
  and (_05571_, _05570_, _05408_);
  and (_05572_, _05233_, _04795_);
  and (_05573_, _05245_, _04779_);
  and (_05574_, _05237_, _04846_);
  and (_05575_, _05241_, _04736_);
  or (_05576_, _05575_, _05574_);
  or (_05577_, _05576_, _05573_);
  or (_05578_, _05577_, _05572_);
  and (_05579_, _05578_, _05407_);
  or (_05580_, _05579_, _05571_);
  and (_05581_, _05580_, _05497_);
  nand (_05582_, _05581_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05583_, _05581_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05584_, _05583_, _05582_);
  and (_05585_, _05279_, _04846_);
  or (_05586_, _05585_, _05408_);
  and (_05587_, _05283_, _04736_);
  and (_05588_, _05275_, _04795_);
  and (_05589_, _05287_, _04779_);
  or (_05590_, _05589_, _05588_);
  or (_05591_, _05590_, _05587_);
  or (_05592_, _05591_, _05586_);
  and (_05593_, _05295_, _04795_);
  and (_05594_, _05299_, _04846_);
  or (_05595_, _05594_, _05593_);
  and (_05596_, _05303_, _04736_);
  and (_05597_, _05307_, _04779_);
  or (_05598_, _05597_, _05407_);
  or (_05599_, _05598_, _05596_);
  or (_05600_, _05599_, _05595_);
  nand (_05601_, _05600_, _05592_);
  nor (_05602_, _05601_, _05222_);
  nand (_05603_, _05602_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_05604_, _05602_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_05605_, _05604_, _05603_);
  or (_05606_, _05605_, _05584_);
  or (_05607_, _05606_, _05563_);
  or (_05608_, _05607_, _05520_);
  or (_05609_, _04412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_05610_, _04412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_05611_, _05610_, _05609_);
  and (_05612_, _04455_, _01144_);
  nor (_05613_, _04455_, _01144_);
  or (_05614_, _05613_, _05612_);
  or (_05615_, _05614_, _05611_);
  or (_05616_, _04499_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_05617_, _04499_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_05618_, _05617_, _05616_);
  nor (_05619_, _04548_, _01220_);
  and (_05620_, _04548_, _01220_);
  or (_05621_, _05620_, _05619_);
  or (_05622_, _05621_, _05618_);
  or (_05623_, _05622_, _05615_);
  or (_05624_, _04604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_05625_, _04604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_05626_, _05625_, _05624_);
  nor (_05627_, _04646_, _00687_);
  and (_05628_, _04646_, _00687_);
  or (_05629_, _05628_, _05627_);
  or (_05630_, _05629_, _05626_);
  and (_05631_, _04729_, _00659_);
  nor (_05632_, _04729_, _00659_);
  or (_05633_, _05632_, _05631_);
  and (_05634_, _04688_, _00619_);
  nor (_05635_, _04688_, _00619_);
  or (_05636_, _05635_, _05634_);
  or (_05637_, _05636_, _05633_);
  or (_05638_, _05637_, _05630_);
  or (_05639_, _05638_, _05623_);
  or (_05640_, _05639_, _05608_);
  nor (_05641_, _04992_, _04931_);
  not (_05642_, _04879_);
  and (_05643_, _05401_, _04830_);
  and (_05644_, _05360_, _05315_);
  and (_05645_, _05644_, _05643_);
  and (_05646_, _05645_, _05642_);
  and (_05647_, _05646_, _05641_);
  and (_05648_, _05647_, _05230_);
  and (property_invalid_ljmp, _05648_, _05640_);
  and (_05649_, _04688_, _04773_);
  nor (_05650_, _04688_, _04773_);
  nor (_05651_, _05650_, _05649_);
  and (_05652_, _04688_, _04762_);
  nor (_05653_, _04688_, _04762_);
  and (_05654_, _04688_, _04767_);
  and (_05655_, _04940_, _04688_);
  nor (_05656_, _04940_, _04688_);
  nor (_05657_, _04936_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_05658_, _05657_, _04937_);
  and (_05659_, _05658_, _04688_);
  nor (_05660_, _05658_, _04688_);
  nor (_05661_, _05660_, _05659_);
  and (_05662_, _04741_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_05663_, _05662_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_05664_, _05663_, _04936_);
  and (_05665_, _05664_, _04688_);
  nor (_05666_, _05664_, _04688_);
  nor (_05667_, _04741_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_05668_, _05667_, _05662_);
  and (_05669_, _05668_, _04688_);
  nor (_05670_, _04740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_05671_, _05670_, _04741_);
  and (_05672_, _05671_, _04688_);
  nor (_05673_, _05671_, _04688_);
  nor (_05674_, _04739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_05675_, _05674_, _04740_);
  and (_05676_, _05675_, _04729_);
  nor (_05677_, _05675_, _04729_);
  nor (_05678_, _05677_, _05676_);
  not (_05679_, _05678_);
  and (_05680_, _04737_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_05681_, _05680_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_05682_, _05681_, _04739_);
  and (_05683_, _05682_, _04604_);
  nor (_05684_, _05682_, _04604_);
  nor (_05685_, _05684_, _05683_);
  not (_05686_, _05685_);
  nor (_05687_, _04737_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_05688_, _05687_, _05680_);
  and (_05689_, _05688_, _04646_);
  and (_05690_, _04499_, _05408_);
  nor (_05691_, _04499_, _05408_);
  nor (_05692_, _04846_, _04779_);
  not (_05693_, _05692_);
  and (_05694_, _05693_, _04548_);
  and (_05695_, _04412_, _12949_);
  and (_05696_, _04455_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05697_, _04412_, _12949_);
  nor (_05698_, _05697_, _05695_);
  and (_05699_, _05698_, _05696_);
  nor (_05700_, _05699_, _05695_);
  nor (_05701_, _05693_, _04548_);
  nor (_05702_, _05701_, _05694_);
  not (_05703_, _05702_);
  nor (_05704_, _05703_, _05700_);
  nor (_05705_, _05704_, _05694_);
  nor (_05706_, _05705_, _05691_);
  nor (_05707_, _05706_, _05690_);
  nor (_05708_, _05688_, _04646_);
  nor (_05709_, _05708_, _05689_);
  not (_05710_, _05709_);
  nor (_05711_, _05710_, _05707_);
  nor (_05712_, _05711_, _05689_);
  nor (_05713_, _05712_, _05686_);
  nor (_05714_, _05713_, _05683_);
  nor (_05715_, _05714_, _05679_);
  nor (_05716_, _05715_, _05676_);
  nor (_05717_, _05716_, _05673_);
  or (_05718_, _05717_, _05672_);
  nor (_05719_, _05668_, _04688_);
  nor (_05720_, _05719_, _05669_);
  and (_05721_, _05720_, _05718_);
  nor (_05722_, _05721_, _05669_);
  nor (_05723_, _05722_, _05666_);
  or (_05724_, _05723_, _05665_);
  and (_05725_, _05724_, _05661_);
  nor (_05726_, _05725_, _05659_);
  nor (_05727_, _05726_, _05656_);
  or (_05728_, _05727_, _05655_);
  nor (_05729_, _04688_, _04767_);
  nor (_05730_, _05729_, _05654_);
  and (_05731_, _05730_, _05728_);
  nor (_05732_, _05731_, _05654_);
  nor (_05733_, _05732_, _05653_);
  or (_05734_, _05733_, _05652_);
  and (_05735_, _05734_, _05651_);
  nor (_05736_, _05735_, _05649_);
  and (_05737_, _04688_, _04751_);
  nor (_05738_, _04688_, _04751_);
  or (_05739_, _05738_, _05737_);
  and (_05740_, _05739_, _05736_);
  nor (_05741_, _05739_, _05736_);
  or (_05742_, _05741_, _05740_);
  nor (_05743_, _05742_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and (_05744_, _05742_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_05745_, _05734_, _05651_);
  nor (_05746_, _05745_, _05735_);
  nor (_05747_, _05746_, _00659_);
  and (_05748_, _05746_, _00659_);
  not (_05749_, _05732_);
  not (_05750_, _04688_);
  nand (_05751_, _05750_, _04765_);
  or (_05752_, _05750_, _04765_);
  and (_05753_, _05752_, _05751_);
  nor (_05754_, _05753_, _05749_);
  not (_05755_, _04946_);
  and (_05756_, _05755_, _04688_);
  nor (_05757_, _05755_, _04688_);
  nor (_05758_, _05757_, _05756_);
  or (_05759_, _05758_, _05726_);
  nand (_05760_, _05758_, _05726_);
  and (_05761_, _05760_, _05759_);
  nor (_05762_, _05724_, _05661_);
  nor (_05763_, _05762_, _05725_);
  nor (_05764_, _05763_, _01220_);
  and (_05765_, _05763_, _01220_);
  nor (_05766_, _05720_, _05718_);
  nor (_05767_, _05766_, _05721_);
  and (_05768_, _05767_, _01144_);
  nor (_05769_, _05672_, _05673_);
  nor (_05770_, _05769_, _05716_);
  and (_05771_, _05769_, _05716_);
  nor (_05772_, _05771_, _05770_);
  and (_05773_, _05772_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_05774_, _05772_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_05775_, _05714_, _05679_);
  nor (_05776_, _05775_, _05715_);
  and (_05777_, _05776_, _01188_);
  nor (_05778_, _05776_, _01188_);
  and (_05779_, _05712_, _05686_);
  nor (_05780_, _05779_, _05713_);
  nor (_05781_, _05780_, _01192_);
  and (_05782_, _05780_, _01192_);
  and (_05783_, _05710_, _05707_);
  nor (_05784_, _05783_, _05711_);
  nor (_05785_, _05784_, _04608_);
  nor (_05786_, _05691_, _05690_);
  and (_05787_, _05786_, _05705_);
  nor (_05788_, _05786_, _05705_);
  nor (_05789_, _05788_, _05787_);
  and (_05790_, _05789_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_05791_, _05789_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_05792_, _05703_, _05700_);
  nor (_05793_, _05792_, _05704_);
  and (_05794_, _05793_, _04503_);
  nor (_05795_, _05698_, _05696_);
  nor (_05796_, _05795_, _05699_);
  nor (_05797_, _05796_, _05013_);
  and (_05798_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05799_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_05800_, _05799_, _05798_);
  not (_05801_, _05800_);
  nand (_05802_, _05801_, _04455_);
  or (_05803_, _05801_, _04455_);
  and (_05804_, _05803_, _05802_);
  and (_05805_, _05796_, _05013_);
  or (_05806_, _05805_, _05804_);
  or (_05807_, _05806_, _05797_);
  nor (_05808_, _05793_, _04503_);
  or (_05809_, _05808_, _05807_);
  or (_05810_, _05809_, _05794_);
  or (_05811_, _05810_, _05791_);
  or (_05812_, _05811_, _05790_);
  and (_05813_, _05784_, _04608_);
  or (_05814_, _05813_, _05812_);
  or (_05815_, _05814_, _05785_);
  or (_05816_, _05815_, _05782_);
  or (_05817_, _05816_, _05781_);
  or (_05818_, _05817_, _05778_);
  or (_05819_, _05818_, _05777_);
  or (_05820_, _05819_, _05774_);
  or (_05821_, _05820_, _05773_);
  or (_05822_, _05821_, _05768_);
  or (_05823_, _05664_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_05824_, _05664_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_05825_, _05824_, _05823_);
  or (_05826_, _05825_, _04688_);
  nand (_05827_, _05825_, _04688_);
  and (_05828_, _05827_, _05826_);
  and (_05829_, _05828_, _05722_);
  nor (_05830_, _05767_, _01144_);
  nor (_05831_, _05828_, _05722_);
  or (_05832_, _05831_, _05830_);
  or (_05833_, _05832_, _05829_);
  or (_05834_, _05833_, _05822_);
  or (_05835_, _05834_, _05765_);
  or (_05836_, _05835_, _05764_);
  or (_05837_, _05836_, _05761_);
  or (_05838_, _05837_, _05754_);
  nor (_05839_, _05730_, _05728_);
  nor (_05840_, _05839_, _05731_);
  nor (_05841_, _05840_, _00687_);
  and (_05842_, _05753_, _05749_);
  and (_05843_, _05840_, _00687_);
  or (_05844_, _05843_, _05842_);
  or (_05845_, _05844_, _05841_);
  or (_05846_, _05845_, _05838_);
  or (_05847_, _05846_, _05748_);
  or (_05848_, _05847_, _05747_);
  or (_05849_, _05848_, _05744_);
  or (_05850_, _05849_, _05743_);
  not (_05851_, _04931_);
  and (_05852_, _04992_, _05851_);
  and (_05853_, _05445_, _04736_);
  nor (_05854_, _05853_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_05855_, _05437_, _04795_);
  not (_05856_, _05855_);
  and (_05857_, _05441_, _04846_);
  and (_05858_, _05432_, _04779_);
  nor (_05859_, _05858_, _05857_);
  and (_05860_, _05859_, _05856_);
  and (_05861_, _05860_, _05854_);
  and (_05862_, _05465_, _04736_);
  nor (_05863_, _05862_, _01350_);
  and (_05864_, _05461_, _04846_);
  not (_05865_, _05864_);
  and (_05866_, _05452_, _04779_);
  and (_05867_, _05457_, _04795_);
  nor (_05868_, _05867_, _05866_);
  and (_05869_, _05868_, _05865_);
  and (_05870_, _05869_, _05863_);
  or (_05871_, _05870_, _05861_);
  not (_05872_, _05871_);
  and (_05873_, _05872_, _04830_);
  nor (_05874_, _05873_, _04879_);
  nor (_05875_, _05643_, _05359_);
  and (_05876_, _05875_, _05315_);
  and (_05877_, _05876_, _05874_);
  and (_05878_, _05877_, _05852_);
  and (_05879_, _05878_, _05230_);
  and (property_invalid_sjmp, _05879_, _05850_);
  and (_05880_, _07455_, _07454_);
  nand (_05881_, _05880_, _08436_);
  nor (_05882_, _05881_, _06968_);
  and (_05883_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand (_05884_, _07467_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor (_05885_, _07475_, _07165_);
  not (_05886_, _05885_);
  or (_05887_, _05886_, _07472_);
  or (_05888_, _05887_, _05884_);
  and (_05889_, _05888_, _05883_);
  and (_05890_, _05889_, _05881_);
  or (_05891_, _05890_, _07459_);
  or (_05892_, _05891_, _05882_);
  nand (_05893_, _07459_, _07317_);
  and (_05894_, _05893_, _06989_);
  and (_04835_, _05894_, _05892_);
  not (_05895_, _04992_);
  nor (_05896_, _05401_, _05313_);
  and (_05897_, _05896_, _05272_);
  and (_05898_, _05897_, _05359_);
  and (_05899_, _04930_, _04878_);
  and (_05900_, _05899_, _05898_);
  and (_05901_, _05900_, _05873_);
  and (_05902_, _05643_, _05359_);
  and (_05903_, _05902_, _05315_);
  not (_05904_, _04878_);
  or (_05905_, _05871_, _05904_);
  and (_05906_, _05905_, _04931_);
  and (_05907_, _05906_, _05903_);
  or (_05908_, _05907_, _05901_);
  and (_05909_, _05908_, _05895_);
  and (_05910_, _05876_, _05873_);
  not (_05911_, _05873_);
  and (_05912_, _05898_, _05911_);
  or (_05913_, _05912_, _05910_);
  and (_05914_, _05852_, _05904_);
  and (_05915_, _05914_, _05913_);
  or (_05916_, _05915_, _05909_);
  and (_05917_, _05160_, _04756_);
  and (_05918_, _05917_, _04742_);
  and (_05919_, _05918_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_05920_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_05921_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_05922_, _05921_, _05920_);
  or (_05923_, _05922_, _05919_);
  nand (_05924_, _05922_, _05919_);
  and (_05925_, _05924_, _05923_);
  and (_05926_, _05160_, _04738_);
  and (_05927_, _05926_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_05928_, _05926_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_05929_, _05928_, _05927_);
  nor (_05930_, _05929_, _01188_);
  nor (_05931_, _05918_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_05932_, _05931_, _05919_);
  nor (_05933_, _05932_, _01220_);
  or (_05934_, _05933_, _05930_);
  or (_05935_, _05934_, _05925_);
  and (_05936_, _05917_, _04744_);
  and (_05937_, _05936_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_05938_, _05936_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_05939_, _05938_, _05937_);
  and (_05940_, _05939_, _00687_);
  and (_05941_, _05929_, _01188_);
  or (_05942_, _05941_, _05940_);
  and (_05943_, _05917_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_05944_, _05943_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_05945_, _05943_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_05946_, _05945_, _05944_);
  and (_05947_, _05946_, _01227_);
  and (_05948_, _05932_, _01220_);
  or (_05949_, _05948_, _05947_);
  or (_05950_, _05949_, _05942_);
  nor (_05951_, _05162_, _05001_);
  and (_05952_, _05162_, _05001_);
  or (_05953_, _05952_, _05951_);
  and (_05954_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_05955_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_05956_, _05955_, _05954_);
  nand (_05957_, _05956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_05958_, _05956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05959_, _05958_, _05957_);
  nand (_05960_, _05959_, _05801_);
  or (_05961_, _05159_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_05962_, _05159_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05963_, _05962_, _05961_);
  or (_05964_, _05963_, _05960_);
  or (_05965_, _05964_, _05953_);
  and (_05966_, _05160_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_05967_, _05160_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_05968_, _05967_, _05966_);
  and (_05969_, _05968_, _04608_);
  nor (_05970_, _05968_, _04608_);
  or (_05971_, _05970_, _05969_);
  or (_05972_, _05971_, _05965_);
  nor (_05973_, _05917_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_05974_, _05973_, _05943_);
  nor (_05975_, _05974_, _01144_);
  and (_05976_, _05974_, _01144_);
  or (_05977_, _05976_, _05975_);
  or (_05978_, _05977_, _05972_);
  nor (_05979_, _05946_, _01227_);
  nor (_05980_, _05939_, _00687_);
  or (_05981_, _05980_, _05979_);
  or (_05982_, _05981_, _05978_);
  or (_05983_, _05982_, _05950_);
  or (_05984_, _05983_, _05935_);
  and (_05985_, _05937_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_05986_, _05985_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_05987_, _05985_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_05988_, _05987_, _05986_);
  nand (_05989_, _05988_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_05990_, _05988_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_05991_, _05990_, _05989_);
  nor (_05992_, _05937_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_05993_, _05992_, _05985_);
  and (_05994_, _05993_, _01686_);
  nor (_05995_, _05993_, _01686_);
  nor (_05996_, _05966_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_05997_, _05996_, _05926_);
  nor (_05998_, _05997_, _01192_);
  and (_05999_, _05997_, _01192_);
  or (_06000_, _05999_, _05998_);
  nor (_06001_, _05927_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_06002_, _06001_, _05917_);
  nor (_06003_, _06002_, _01149_);
  and (_06004_, _06002_, _01149_);
  or (_06005_, _06004_, _06003_);
  or (_06006_, _06005_, _06000_);
  or (_06007_, _06006_, _05995_);
  or (_06008_, _06007_, _05994_);
  or (_06009_, _06008_, _05991_);
  and (_06010_, _05986_, _00655_);
  nor (_06011_, _05986_, _00655_);
  or (_06012_, _06011_, _06010_);
  nor (_06013_, _06012_, _00619_);
  and (_06014_, _06012_, _00619_);
  or (_06015_, _06014_, _06013_);
  or (_06016_, _06015_, _06009_);
  or (_06017_, _06016_, _05984_);
  and (_06018_, _06017_, _05230_);
  and (property_invalid_pcp3, _06018_, _05916_);
  or (_06019_, _05658_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_06020_, _05658_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_06021_, _06020_, _06019_);
  or (_06022_, _05668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_06023_, _05668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_06024_, _06023_, _06022_);
  and (_06025_, _05671_, _01149_);
  nor (_06026_, _05671_, _01149_);
  or (_06027_, _06026_, _06025_);
  nor (_06028_, _05675_, _01188_);
  and (_06029_, _05675_, _01188_);
  or (_06030_, _06029_, _06028_);
  nor (_06031_, _05682_, _01192_);
  and (_06032_, _05682_, _01192_);
  or (_06033_, _06032_, _06031_);
  and (_06034_, _05407_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_06035_, _05407_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_06036_, _06035_, _06034_);
  and (_06037_, _05692_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand (_06038_, _05956_, _05800_);
  nor (_06039_, _05692_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_06040_, _06039_, _06038_);
  or (_06041_, _06040_, _06037_);
  or (_06042_, _06041_, _06036_);
  nor (_06043_, _05688_, _04608_);
  and (_06044_, _05688_, _04608_);
  or (_06045_, _06044_, _06043_);
  or (_06046_, _06045_, _06042_);
  or (_06047_, _06046_, _06033_);
  or (_06048_, _06047_, _06030_);
  or (_06049_, _06048_, _06027_);
  or (_06050_, _06049_, _06024_);
  or (_06051_, _06050_, _05825_);
  or (_06052_, _06051_, _06021_);
  or (_06053_, _06052_, _04946_);
  or (_06054_, _06053_, _04778_);
  and (_06055_, _04931_, _05642_);
  and (_06056_, _06055_, _05644_);
  or (_06057_, _05900_, _05895_);
  or (_06058_, _06057_, _06056_);
  and (_06059_, _05871_, _05314_);
  and (_06060_, _05873_, _05904_);
  and (_06061_, _06060_, _05897_);
  or (_06062_, _06061_, _06059_);
  and (_06063_, _06062_, _05851_);
  or (_06064_, _06063_, _05646_);
  or (_06065_, _06064_, _06058_);
  and (_06066_, _05643_, _05272_);
  and (_06067_, _06066_, _05873_);
  and (_06068_, _06067_, _04879_);
  not (_06069_, _05358_);
  and (_06070_, _05897_, _06069_);
  or (_06071_, _06070_, _05645_);
  or (_06072_, _06071_, _06068_);
  and (_06073_, _06072_, _04931_);
  and (_06074_, _05898_, _05642_);
  and (_06075_, _05899_, _05314_);
  and (_06076_, _06075_, _05872_);
  or (_06077_, _06076_, _04992_);
  or (_06078_, _06077_, _06074_);
  or (_06079_, _06078_, _06073_);
  and (_06080_, _06079_, _06065_);
  and (_06081_, _06066_, _05911_);
  and (_06082_, _05644_, _04878_);
  or (_06083_, _06082_, _06081_);
  and (_06084_, _06083_, _05852_);
  and (_06085_, _05912_, _04931_);
  and (_06086_, _05897_, _04879_);
  and (_06087_, _06086_, _05641_);
  or (_06088_, _06087_, _06085_);
  or (_06089_, _06088_, _06084_);
  or (_06090_, _06089_, _06080_);
  and (_06091_, _06090_, _05230_);
  and (property_invalid_pcp2, _06091_, _06054_);
  and (_06092_, _03503_, _09009_);
  and (_06093_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_06094_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_06095_, _06094_, _06093_);
  nor (_06096_, _06095_, _13986_);
  and (_06097_, _04006_, _11821_);
  or (_06098_, _06097_, _06096_);
  or (_06099_, _06098_, _06092_);
  and (_04843_, _06099_, _06989_);
  and (_06100_, _05875_, _05895_);
  or (_06101_, _06100_, _06070_);
  and (_06102_, _06101_, _05874_);
  and (_06103_, _06069_, _05272_);
  nor (_06104_, _04992_, _04878_);
  and (_06105_, _06104_, _06103_);
  and (_06106_, _05314_, _05904_);
  and (_06107_, _06106_, _05873_);
  or (_06108_, _06107_, _05903_);
  or (_06109_, _06108_, _06105_);
  or (_06110_, _06109_, _06102_);
  and (_06111_, _06110_, _05851_);
  and (_06112_, _06067_, _05642_);
  or (_06113_, _06103_, _05902_);
  and (_06114_, _04991_, _04931_);
  and (_06115_, _06114_, _06113_);
  nor (_06116_, _06115_, _06112_);
  nor (_06117_, _06116_, _05314_);
  and (_06118_, _06069_, _04878_);
  and (_06119_, _06118_, _04992_);
  or (_06120_, _06119_, _06059_);
  or (_06121_, _06120_, _06081_);
  and (_06122_, _06121_, _04931_);
  or (_06123_, _06106_, _04991_);
  or (_06124_, _06075_, _04989_);
  and (_06125_, _06124_, _06123_);
  or (_06126_, _06066_, _05314_);
  and (_06127_, _06126_, _05641_);
  and (_06128_, _05871_, _04878_);
  and (_06129_, _06128_, _05897_);
  and (_06130_, _06129_, _05852_);
  or (_06131_, _06130_, _06127_);
  or (_06132_, _06131_, _06125_);
  or (_06133_, _06132_, _06122_);
  or (_06134_, _06133_, _06117_);
  or (_06135_, _06134_, _06111_);
  not (_06136_, _04756_);
  nand (_06137_, _04737_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_06138_, _06137_, _06136_);
  and (_06139_, _06138_, _04744_);
  and (_06140_, _06139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_06141_, _06140_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_06142_, _06141_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_06143_, _06142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_06144_, _06142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_06145_, _06144_, _06143_);
  and (_06146_, _06145_, _00619_);
  nor (_06147_, _06141_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_06148_, _06147_, _06142_);
  nand (_06149_, _06148_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or (_06150_, _06148_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and (_06151_, _06150_, _06149_);
  nor (_06152_, _06145_, _00619_);
  or (_06153_, _06152_, _06151_);
  or (_06154_, _06153_, _06146_);
  and (_06155_, _04740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_06156_, _06155_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_06157_, _06155_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_06158_, _06157_, _06156_);
  and (_06159_, _06158_, _01149_);
  nor (_06160_, _06158_, _01149_);
  and (_06161_, _06138_, _04742_);
  nor (_06162_, _06161_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_06163_, _06161_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_06164_, _06163_, _06162_);
  nor (_06165_, _06164_, _01220_);
  and (_06166_, _06164_, _01220_);
  or (_06167_, _06166_, _06165_);
  nor (_06168_, _06139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_06169_, _06168_, _06140_);
  nor (_06170_, _06169_, _00687_);
  and (_06171_, _06169_, _00687_);
  or (_06172_, _06171_, _06170_);
  or (_06173_, _06172_, _06167_);
  or (_06174_, _06173_, _06160_);
  or (_06175_, _06174_, _06159_);
  nor (_06176_, _06140_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_06177_, _06176_, _06141_);
  nor (_06178_, _06177_, _01686_);
  and (_06179_, _04739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_06180_, _06179_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_06181_, _06180_, _06155_);
  and (_06182_, _06181_, _01188_);
  nor (_06183_, _06181_, _01188_);
  or (_06184_, _06183_, _06182_);
  or (_06185_, _06184_, _06178_);
  and (_06186_, _06138_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_06187_, _06138_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_06188_, _06187_, _06186_);
  nor (_06189_, _06188_, _01144_);
  and (_06190_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _04608_);
  nor (_06191_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_06192_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_06193_, _06192_, _06191_);
  nor (_06194_, _06193_, _06137_);
  nor (_06195_, _06194_, _06190_);
  and (_06196_, _01346_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor (_06197_, _06196_, _06193_);
  or (_06198_, _06197_, _06137_);
  or (_06199_, _06198_, _06195_);
  nand (_06200_, _06197_, _06195_);
  and (_06201_, _06200_, _06199_);
  and (_06202_, _06188_, _01144_);
  or (_06203_, _06202_, _06201_);
  or (_06204_, _06203_, _06189_);
  or (_06205_, _06163_, _05922_);
  nand (_06206_, _06163_, _05922_);
  and (_06207_, _06206_, _06205_);
  nor (_06208_, _04316_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_06209_, _04316_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_06210_, _06209_, _06208_);
  or (_06211_, _05959_, _05800_);
  nor (_06212_, _04312_, _04503_);
  and (_06213_, _04312_, _04503_);
  or (_06214_, _06213_, _06212_);
  or (_06215_, _06214_, _06211_);
  or (_06216_, _06215_, _06210_);
  or (_06217_, _06216_, _06207_);
  or (_06218_, _06217_, _06204_);
  and (_06219_, _06177_, _01686_);
  and (_06220_, _06186_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_06221_, _06186_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_06222_, _06221_, _06220_);
  or (_06223_, _06222_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_06224_, _06222_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_06225_, _06224_, _06223_);
  or (_06226_, _06225_, _06219_);
  or (_06227_, _06226_, _06218_);
  or (_06228_, _06227_, _06185_);
  or (_06229_, _06228_, _06175_);
  or (_06230_, _06229_, _06154_);
  and (_06231_, _06230_, _05230_);
  and (property_invalid_pcp1, _06231_, _06135_);
  and (_06232_, _03503_, _09599_);
  and (_06233_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_06234_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_06235_, _06234_, _06233_);
  nor (_06236_, _06235_, _13986_);
  and (_06237_, _04006_, _09009_);
  or (_06238_, _06237_, _06236_);
  or (_06239_, _06238_, _06232_);
  and (_04848_, _06239_, _06989_);
  and (_06240_, _05223_, first_instr);
  or (_00000_, _06240_, rst);
  or (_06241_, _13959_, _13969_);
  nor (_06242_, _06241_, _00918_);
  and (_06243_, _00918_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_06244_, _06243_, _06242_);
  and (_06245_, _13968_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_06246_, _06245_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_06247_, _06246_, _13959_);
  nor (_06248_, _06247_, _06244_);
  nor (_06249_, _06248_, _13986_);
  and (_06250_, _04181_, _09599_);
  or (_06251_, _06250_, _06249_);
  and (_04872_, _06251_, _06989_);
  nor (_06252_, _10970_, _04286_);
  nor (_06253_, _07145_, _03252_);
  and (_06254_, _06253_, _09580_);
  nand (_06255_, _07071_, _07056_);
  and (_06256_, _06255_, _03245_);
  nor (_06257_, _06256_, _09575_);
  or (_06258_, _06257_, _07077_);
  or (_06259_, _06258_, _06254_);
  and (_06260_, _07077_, _03252_);
  nor (_06261_, _06260_, _07046_);
  and (_06262_, _06261_, _06259_);
  or (_06263_, _06262_, _07050_);
  or (_06264_, _06263_, _06252_);
  nand (_06265_, _07050_, _03245_);
  and (_06266_, _06265_, _06989_);
  and (_04889_, _06266_, _06264_);
  and (_06267_, _07077_, _03256_);
  nor (_06268_, _07145_, _03256_);
  and (_06269_, _06268_, _09580_);
  not (_06270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand (_06271_, _02808_, _06270_);
  and (_06272_, _06271_, _06255_);
  or (_06273_, _06272_, _07077_);
  nor (_06274_, _06273_, _06269_);
  or (_06275_, _06274_, _06267_);
  nand (_06276_, _06275_, _04286_);
  nand (_06277_, _07118_, _07046_);
  and (_06278_, _06277_, _06276_);
  or (_06279_, _06278_, _07050_);
  nand (_06280_, _07050_, _06270_);
  and (_06281_, _06280_, _06989_);
  and (_04896_, _06281_, _06279_);
  and (_06282_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_06283_, _06282_, _09580_);
  and (_06284_, _07071_, _07062_);
  nor (_06285_, _06284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_06286_, _06285_, _04293_);
  or (_06287_, _06286_, _07077_);
  or (_06288_, _06287_, _06283_);
  nor (_06289_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_06290_, _06289_, _07046_);
  and (_06291_, _06290_, _06288_);
  and (_06292_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_06293_, _06292_, _07050_);
  or (_06294_, _06293_, _06291_);
  nand (_06295_, _07260_, _07050_);
  and (_06296_, _06295_, _06989_);
  and (_04909_, _06296_, _06294_);
  and (_06297_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_06298_, _06297_, _09580_);
  nand (_06299_, _07071_, _07061_);
  and (_06300_, _06299_, _03049_);
  nor (_06301_, _06300_, _06284_);
  or (_06302_, _06301_, _07077_);
  or (_06303_, _06302_, _06298_);
  nor (_06304_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_06305_, _06304_, _07046_);
  and (_06306_, _06305_, _06303_);
  and (_06307_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_06308_, _06307_, _07050_);
  or (_06309_, _06308_, _06306_);
  nand (_06310_, _07317_, _07050_);
  and (_06311_, _06310_, _06989_);
  and (_04916_, _06311_, _06309_);
  and (_06312_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_06313_, _06312_, _09580_);
  and (_06314_, _07071_, _07060_);
  or (_06315_, _06314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_06316_, _06315_, _06299_);
  or (_06317_, _06316_, _07077_);
  or (_06318_, _06317_, _06313_);
  nor (_06319_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_06320_, _06319_, _07046_);
  and (_06321_, _06320_, _06318_);
  and (_06322_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_06323_, _06322_, _07050_);
  or (_06324_, _06323_, _06321_);
  nand (_06325_, _11529_, _07050_);
  and (_06326_, _06325_, _06989_);
  and (_04920_, _06326_, _06324_);
  nor (_06327_, _10970_, _14146_);
  and (_06328_, _08999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_06329_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and (_06330_, _06329_, _09002_);
  or (_06331_, _06330_, _06328_);
  or (_06332_, _06331_, _06327_);
  and (_04922_, _06332_, _06989_);
  and (_06333_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_06334_, _06333_, _09580_);
  and (_06335_, _07071_, _07059_);
  nor (_06336_, _06335_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_06337_, _06336_, _06314_);
  or (_06338_, _06337_, _07077_);
  or (_06339_, _06338_, _06334_);
  nor (_06340_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_06341_, _06340_, _07046_);
  and (_06342_, _06341_, _06339_);
  and (_06343_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_06344_, _06343_, _07050_);
  or (_06345_, _06344_, _06342_);
  nand (_06346_, _09008_, _07050_);
  and (_06347_, _06346_, _06989_);
  and (_04924_, _06347_, _06345_);
  and (_06348_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_06349_, _08139_, _04608_);
  or (_06350_, _06349_, _06348_);
  and (_04941_, _06350_, _06989_);
  and (_06351_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_06352_, _08139_, _05001_);
  or (_06353_, _06352_, _06351_);
  and (_04943_, _06353_, _06989_);
  and (_06354_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_06355_, _06354_, _09580_);
  and (_06356_, _09577_, _03143_);
  nor (_06357_, _06356_, _06335_);
  or (_06358_, _06357_, _07077_);
  or (_06359_, _06358_, _06355_);
  nor (_06360_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_06361_, _06360_, _07046_);
  and (_06362_, _06361_, _06359_);
  and (_06363_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_06364_, _06363_, _07050_);
  or (_06365_, _06364_, _06362_);
  nand (_06366_, _09598_, _07050_);
  and (_06367_, _06366_, _06989_);
  and (_04945_, _06367_, _06365_);
  nand (_06368_, _05880_, _07089_);
  nor (_06369_, _06368_, _06968_);
  or (_06370_, _05885_, _07472_);
  or (_06371_, _06370_, _05884_);
  nand (_06372_, _06371_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand (_06373_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_06374_, _06373_, _06368_);
  or (_06375_, _06374_, _07459_);
  or (_06376_, _06375_, _06369_);
  nand (_06377_, _09008_, _07459_);
  and (_06378_, _06377_, _06989_);
  and (_04978_, _06378_, _06376_);
  and (_06379_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_06380_, _08139_, _04503_);
  or (_06381_, _06380_, _06379_);
  and (_04990_, _06381_, _06989_);
  nor (_06382_, _01811_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  or (_06383_, _05887_, _07468_);
  and (_06384_, _06383_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_06385_, _06384_, _06382_);
  and (_06386_, _05880_, _07048_);
  or (_06387_, _06386_, _06385_);
  nand (_06388_, _06386_, _06968_);
  and (_06389_, _06388_, _06387_);
  or (_06390_, _06389_, _07459_);
  nand (_06391_, _07459_, _07118_);
  and (_06392_, _06391_, _06989_);
  and (_05002_, _06392_, _06390_);
  and (_06393_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_06394_, _08139_, _05013_);
  or (_06395_, _06394_, _06393_);
  and (_05018_, _06395_, _06989_);
  and (_06396_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_06397_, _08139_, _04416_);
  or (_06398_, _06397_, _06396_);
  and (_05033_, _06398_, _06989_);
  dff (first_instr, _00000_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _14649_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _14650_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _14651_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _14652_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _14653_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _14654_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _09711_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _14655_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _14707_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _09612_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _09617_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _09622_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _14708_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _14709_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _14710_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _09635_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _09522_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _14702_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _09526_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _14703_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _14704_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _14705_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _09540_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _14706_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _14694_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _14695_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _14696_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _14697_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _14698_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _14699_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _14700_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _14701_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _09328_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _14691_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _09335_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _14692_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _14693_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _09346_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _09351_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _09354_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _09235_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _09238_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _14690_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _09243_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _09247_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _09251_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _09254_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _09257_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _08840_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _14666_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _14667_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _14668_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _14669_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _14670_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _14671_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _14672_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _14642_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _14643_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _14644_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _14645_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _08749_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _14646_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _14647_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _14648_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _14680_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _14681_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _14682_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _14683_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _14684_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _14685_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _14686_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _09047_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _14673_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _14674_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _14675_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _14676_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _14677_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _08962_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _14678_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _14679_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _09135_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _09137_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _09141_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _14687_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _14688_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _14689_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _09152_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _09154_);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _07214_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _07241_);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _07280_);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _07329_);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _07388_);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _07451_);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _07503_);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _07599_);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _07673_);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _07773_);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _07869_);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _07980_);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _08081_);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _08217_);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _08347_);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _07163_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _10126_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _10131_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _10133_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _10135_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _10137_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _10139_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _10144_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _07192_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _14665_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _09956_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _09961_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _09963_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _09967_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _09971_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _09973_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _09978_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _10042_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _10047_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _10049_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _10051_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _10053_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _10055_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _10058_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _10062_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _09864_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _09867_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _09869_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _09874_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _09877_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _09880_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _14664_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _09885_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _14656_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _14657_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _14658_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _14659_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _14660_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _14661_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _14662_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _14663_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _13463_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _13118_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _13114_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _12965_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _04086_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _04206_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _04099_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _04196_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03313_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _11967_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _12000_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _11997_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _04104_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _12133_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _12387_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _04199_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11307_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _12373_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _11323_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _11318_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _11487_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _11384_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _11362_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11357_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _11434_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _08135_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _11200_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _11228_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _11222_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _11633_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _11268_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _11259_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _06825_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _06827_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _06829_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _06831_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _06833_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _06836_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _06838_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _06671_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _04487_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _06674_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _09999_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _03758_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _00258_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _03795_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _03766_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _03634_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _03693_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _03715_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _03636_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _03721_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _03638_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _03829_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _03833_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _03835_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _03837_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _03839_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _03841_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _03854_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _03641_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _03643_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _03518_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _03645_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _03541_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _03648_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _03557_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _03566_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _03655_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _03579_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _03598_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _03657_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _03719_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _03659_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _03815_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _03869_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _03879_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _03662_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _03995_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _03664_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _03666_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _03764_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _14572_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _11893_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _09305_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _13146_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _09122_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _04117_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _14014_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _01250_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _04211_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _13157_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _04214_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _02297_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _04524_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _04216_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _04034_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _03072_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _00442_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _10877_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _00494_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _03327_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _12693_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _12672_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _02737_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _03345_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _03364_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _13272_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _01662_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _00529_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _03439_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _01770_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _03992_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _08521_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _08660_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _04112_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _01526_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _12548_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _12655_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _03447_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _01800_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _11031_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _07336_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _03957_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _12976_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _03354_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _04003_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _04922_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _04207_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _02650_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _13446_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _01208_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _09596_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _13225_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _12039_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _09662_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _12810_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _01240_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _12941_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _11005_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _13597_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _08073_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _06571_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _02294_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _13343_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _08194_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _08111_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _07933_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _08088_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _03549_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _05033_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _05018_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _04990_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _04943_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _04941_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _00638_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _04566_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _02965_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _02962_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _02922_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _00667_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _02100_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _01835_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _02058_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _02001_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _14123_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _11677_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _10989_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _00681_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _01629_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _01627_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _00588_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _00575_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _00457_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _00445_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _00679_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _00663_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _06580_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _14585_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _14583_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _14403_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _14264_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _04306_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _04532_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _04360_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _10020_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _09691_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _09812_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _03712_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _03706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _10029_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _04068_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _04061_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _04059_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _10025_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _03150_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _00705_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _02578_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _01817_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _01721_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _10036_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _03489_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _03521_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _03512_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _10033_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _09687_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _14024_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _13822_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _13954_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _13872_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _10045_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _00387_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _00055_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _14019_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _14216_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _10056_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _09677_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _09795_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _14142_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _14393_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _01178_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _09919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _03539_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _09922_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _09747_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _00596_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _09929_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _10114_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _09651_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _09936_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _09733_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _04007_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _03810_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _03808_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _00250_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _03755_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _10079_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _04585_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _04582_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _04572_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _04568_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _10074_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _09791_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _04137_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _04134_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _04130_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _04122_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _04114_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _10092_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _04236_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _04233_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _03742_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _03399_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _03374_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _03372_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _10101_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _03831_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _03723_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _03682_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _03651_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _10098_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _09669_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _02056_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _01860_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _02024_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _01870_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _01865_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03726_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _14022_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _03331_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _03350_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _01023_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _01000_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _10112_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _01734_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _01732_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _01697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _01695_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _03329_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _09655_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _00647_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _03315_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _03444_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _10129_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _00160_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _00121_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _00148_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _00136_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _00130_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _00128_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03428_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _03420_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _03413_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _14255_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _14227_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _14225_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _00256_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _13207_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _13154_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _13137_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _13103_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _10142_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _09628_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _12121_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _12104_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _12057_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _10446_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _12478_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _12405_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _12475_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _12445_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _12441_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _12423_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _12414_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _10400_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _09624_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _09779_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11592_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _11544_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _10452_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _11826_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _11854_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _11847_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _11831_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _10449_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _09620_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _08105_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _03985_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _02597_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _03156_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _03146_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _03135_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01762_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01711_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01669_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _00261_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _04227_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _01821_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _14087_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _14082_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _04224_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _04219_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _04570_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _01825_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _13592_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _13580_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _13573_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _01823_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _01187_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _13423_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _04355_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _04353_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _06542_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _06536_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _03047_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _06641_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _06638_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _06626_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _02542_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _09804_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _03687_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _02805_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _02759_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _02563_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _02622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _01201_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _02756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _04485_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _07834_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _07829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _07820_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _07806_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _07785_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _07767_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _07764_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _13651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _07578_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _07635_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _07620_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _07616_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _07592_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _07584_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _07581_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _13649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _02576_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00348_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00327_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00325_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00321_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00318_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00310_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _12565_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00289_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _12832_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _12851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00275_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00272_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _03486_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00254_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00252_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _13415_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00228_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00222_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _04835_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _04978_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _05002_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _01362_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00181_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00179_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _04527_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00138_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00123_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00111_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00117_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00113_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _04529_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00050_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00048_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00031_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00028_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00026_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00024_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00009_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _04539_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _02937_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _02911_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _03081_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _02939_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _03079_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _02909_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _03077_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _00018_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _02935_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _03087_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _02907_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _03083_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _03055_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _03053_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _02933_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _14607_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _03091_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _02903_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _03089_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _03058_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _03057_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _02905_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _03085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _07448_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _02928_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _02899_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _03098_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _02930_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _03095_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _02900_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _03093_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _00502_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _03873_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _03864_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _03825_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _03793_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _03127_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _03561_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _03209_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _03456_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _04799_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _04801_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _04805_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _04813_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _04815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _04817_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _04819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _03475_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _02689_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _02698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _14456_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _14121_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _14115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _14118_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _14111_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _14105_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _14108_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _02695_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _14127_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _14085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _14090_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _14072_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _14075_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _14064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _14059_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _02692_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _02684_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _02683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _14006_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _14009_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _13910_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _13907_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _13908_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _13802_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _13798_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _02680_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _13788_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _13817_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _13809_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _13815_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _13812_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _13766_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _13768_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _02671_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _02677_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _13745_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _13710_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _13707_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _13729_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _13735_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _13919_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _13914_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _02668_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _09976_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _08250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _08297_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _08321_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _03971_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _03966_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _03942_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _03917_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _03929_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _03926_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _03920_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _08181_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _03862_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _03791_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _03821_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _03805_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _03802_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _03799_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _03761_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _08108_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _08266_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _03698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _03679_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _03675_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _03672_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _03669_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _04896_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _04889_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _08330_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _04945_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _04924_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _04920_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _04916_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _04909_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _04594_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _04592_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _10680_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _13884_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _04555_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _04550_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _04547_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _04544_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _03622_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _03619_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _03617_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _11486_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _08094_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _07997_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _07969_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _07992_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _07989_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _07976_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _07973_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _07959_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _08054_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _08100_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _08097_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _13093_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _12170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _12160_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00213_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _12208_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _12229_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _12220_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _02284_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _12214_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _02225_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _08809_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _03479_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _12211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _00465_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _00453_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _14139_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _13758_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _12863_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _12440_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _11465_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00188_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _12085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _12082_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _12075_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _12060_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01896_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _03422_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _00794_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _12052_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _04872_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _04848_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _04843_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _04563_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _04560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _04557_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _04339_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _04334_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _04282_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _04187_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00230_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _02723_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _02705_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _02703_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _02300_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _02286_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _02185_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _02212_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _12115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01673_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _00219_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _00639_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _00570_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _00334_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _13365_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _12128_);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
endmodule
