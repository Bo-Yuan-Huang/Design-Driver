
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_pcp1, property_invalid_pcp2, property_invalid_pcp3, property_invalid_sjmp, property_invalid_ljmp, property_invalid_ajmp, ABINPUT);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  wire _14608_;
  wire _14609_;
  wire _14610_;
  wire _14611_;
  wire _14612_;
  wire _14613_;
  wire _14614_;
  wire _14615_;
  wire _14616_;
  wire _14617_;
  wire _14618_;
  wire _14619_;
  wire _14620_;
  wire _14621_;
  wire _14622_;
  wire _14623_;
  wire _14624_;
  wire _14625_;
  wire _14626_;
  wire _14627_;
  wire _14628_;
  wire _14629_;
  wire _14630_;
  wire _14631_;
  wire _14632_;
  wire _14633_;
  wire _14634_;
  wire _14635_;
  wire _14636_;
  wire _14637_;
  wire _14638_;
  wire _14639_;
  wire _14640_;
  wire _14641_;
  wire _14642_;
  wire _14643_;
  wire _14644_;
  wire _14645_;
  wire _14646_;
  wire _14647_;
  wire _14648_;
  wire _14649_;
  wire _14650_;
  wire _14651_;
  wire _14652_;
  wire _14653_;
  wire _14654_;
  wire _14655_;
  wire _14656_;
  wire _14657_;
  wire _14658_;
  wire _14659_;
  wire _14660_;
  wire _14661_;
  wire _14662_;
  wire _14663_;
  wire _14664_;
  wire _14665_;
  wire _14666_;
  wire _14667_;
  wire _14668_;
  wire _14669_;
  wire _14670_;
  wire _14671_;
  wire _14672_;
  wire _14673_;
  wire _14674_;
  wire _14675_;
  wire _14676_;
  wire _14677_;
  wire _14678_;
  wire _14679_;
  wire _14680_;
  wire _14681_;
  wire _14682_;
  wire _14683_;
  wire _14684_;
  wire _14685_;
  wire _14686_;
  wire _14687_;
  wire _14688_;
  wire _14689_;
  wire _14690_;
  wire _14691_;
  wire _14692_;
  wire _14693_;
  wire _14694_;
  wire _14695_;
  wire _14696_;
  wire _14697_;
  wire _14698_;
  wire _14699_;
  wire _14700_;
  wire _14701_;
  wire _14702_;
  wire _14703_;
  wire _14704_;
  wire _14705_;
  wire _14706_;
  wire _14707_;
  wire _14708_;
  wire _14709_;
  wire _14710_;
  input [8:0] ABINPUT;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid_ajmp;
  output property_invalid_ljmp;
  output property_invalid_pcp1;
  output property_invalid_pcp2;
  output property_invalid_pcp3;
  output property_invalid_sjmp;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  or _14711_ (_06399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _14712_ (_06400_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _14713_ (_06401_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _14714_ (_06402_, _06401_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and _14715_ (_06403_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not _14716_ (_06404_, _06403_);
  not _14717_ (_06405_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not _14718_ (_06406_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _14719_ (_06407_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _06406_);
  and _14720_ (_06408_, _06407_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and _14721_ (_06409_, _06408_, _06405_);
  not _14722_ (_06410_, _06409_);
  nor _14723_ (_06411_, _06402_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _14724_ (_06412_, _06411_, _06410_);
  and _14725_ (_06413_, _06412_, _06404_);
  not _14726_ (_06414_, _06413_);
  not _14727_ (_06415_, _06407_);
  and _14728_ (_06416_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _06406_);
  and _14729_ (_06417_, _06416_, _06415_);
  and _14730_ (_06418_, _06417_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _14731_ (_06419_, _06418_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  and _14732_ (_06420_, _06408_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and _14733_ (_06421_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _06406_);
  nor _14734_ (_06422_, _06421_, _06416_);
  and _14735_ (_06423_, _06422_, _06407_);
  and _14736_ (_06424_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  or _14737_ (_06425_, _06424_, _06420_);
  nor _14738_ (_06426_, _06425_, _06419_);
  and _14739_ (_06427_, _06417_, _06405_);
  and _14740_ (_06428_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nand _14741_ (_06429_, _06422_, _06415_);
  not _14742_ (_06430_, _06429_);
  and _14743_ (_06431_, _06430_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor _14744_ (_06432_, _06431_, _06428_);
  and _14745_ (_06433_, _06432_, _06426_);
  and _14746_ (_06434_, _06433_, _06414_);
  not _14747_ (_06435_, _06402_);
  nor _14748_ (_06436_, _06401_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _14749_ (_06437_, _06436_, _06410_);
  and _14750_ (_06438_, _06437_, _06435_);
  not _14751_ (_06439_, _06438_);
  and _14752_ (_06440_, _06430_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  and _14753_ (_06441_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  nor _14754_ (_06442_, _06441_, _06440_);
  and _14755_ (_06443_, _06418_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _14756_ (_06444_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor _14757_ (_06445_, _06444_, _06443_);
  and _14758_ (_06446_, _06445_, _06442_);
  and _14759_ (_06447_, _06446_, _06439_);
  not _14760_ (_06448_, _06447_);
  and _14761_ (_06449_, _06448_, _06434_);
  and _14762_ (_06450_, _06403_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and _14763_ (_06451_, _06450_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not _14764_ (_06452_, _06451_);
  nor _14765_ (_06453_, _06450_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _14766_ (_06454_, _06453_, _06410_);
  and _14767_ (_06455_, _06454_, _06452_);
  not _14768_ (_06456_, _06455_);
  and _14769_ (_06457_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and _14770_ (_06458_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  and _14771_ (_06459_, _06418_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or _14772_ (_06460_, _06459_, _06458_);
  or _14773_ (_06461_, _06460_, _06420_);
  nor _14774_ (_06462_, _06461_, _06457_);
  and _14775_ (_06463_, _06462_, _06456_);
  not _14776_ (_06464_, _06450_);
  nor _14777_ (_06465_, _06403_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _14778_ (_06466_, _06465_, _06410_);
  and _14779_ (_06467_, _06466_, _06464_);
  not _14780_ (_06468_, _06467_);
  and _14781_ (_06469_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  not _14782_ (_06470_, _06469_);
  and _14783_ (_06471_, _06418_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  not _14784_ (_06472_, _06471_);
  and _14785_ (_06473_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  nor _14786_ (_06474_, _06473_, _06420_);
  and _14787_ (_06475_, _06474_, _06472_);
  and _14788_ (_06476_, _06475_, _06470_);
  and _14789_ (_06477_, _06476_, _06468_);
  not _14790_ (_06478_, _06477_);
  nor _14791_ (_06479_, _06478_, _06463_);
  and _14792_ (_06480_, _06479_, _06449_);
  and _14793_ (_06481_, \oc8051_top_1.oc8051_decoder1.wr , _06406_);
  not _14794_ (_06482_, _06481_);
  and _14795_ (_06483_, _06407_, _06405_);
  nor _14796_ (_06484_, _06483_, _06482_);
  and _14797_ (_06485_, _06484_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not _14798_ (_06486_, _06485_);
  not _14799_ (_06487_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor _14800_ (_06488_, _06451_, _06487_);
  and _14801_ (_06489_, _06451_, _06487_);
  nor _14802_ (_06490_, _06489_, _06488_);
  nor _14803_ (_06491_, _06490_, _06410_);
  not _14804_ (_06492_, _06491_);
  and _14805_ (_06493_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  and _14806_ (_06494_, _06427_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and _14807_ (_06495_, _06418_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  or _14808_ (_06496_, _06495_, _06494_);
  or _14809_ (_06497_, _06496_, _06420_);
  nor _14810_ (_06498_, _06497_, _06493_);
  and _14811_ (_06499_, _06498_, _06492_);
  nor _14812_ (_06500_, _06499_, _06486_);
  and _14813_ (_06501_, _06500_, _06480_);
  or _14814_ (_06502_, _06501_, _06399_);
  and _14815_ (_06503_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and _14816_ (_06504_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor _14817_ (_06505_, _06504_, _06503_);
  and _14818_ (_06506_, _06418_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  not _14819_ (_06507_, _06506_);
  not _14820_ (_06508_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and _14821_ (_06509_, _06409_, _06508_);
  and _14822_ (_06510_, _06430_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor _14823_ (_06511_, _06510_, _06509_);
  and _14824_ (_06512_, _06511_, _06507_);
  and _14825_ (_06513_, _06512_, _06505_);
  not _14826_ (_06514_, _06513_);
  nor _14827_ (_06515_, _06400_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor _14828_ (_06516_, _06515_, _06401_);
  and _14829_ (_06517_, _06516_, _06409_);
  and _14830_ (_06518_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor _14831_ (_06519_, _06518_, _06517_);
  and _14832_ (_06520_, _06418_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _14833_ (_06521_, _06427_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and _14834_ (_06522_, _06430_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or _14835_ (_06523_, _06522_, _06521_);
  nor _14836_ (_06524_, _06523_, _06520_);
  and _14837_ (_06525_, _06524_, _06519_);
  nor _14838_ (_06526_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor _14839_ (_06527_, _06526_, _06400_);
  and _14840_ (_06528_, _06527_, _06409_);
  and _14841_ (_06529_, _06423_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor _14842_ (_06530_, _06529_, _06528_);
  and _14843_ (_06531_, _06418_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and _14844_ (_06532_, _06427_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and _14845_ (_06533_, _06430_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or _14846_ (_06534_, _06533_, _06532_);
  nor _14847_ (_06535_, _06534_, _06531_);
  and _14848_ (_06537_, _06535_, _06530_);
  nor _14849_ (_06538_, _06537_, _06525_);
  and _14850_ (_06539_, _06538_, _06514_);
  not _14851_ (_06540_, _06539_);
  not _14852_ (_06541_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and _14853_ (_06543_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _06406_);
  and _14854_ (_06544_, _06543_, _06541_);
  and _14855_ (_06545_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _06406_);
  and _14856_ (_06546_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _06406_);
  nor _14857_ (_06547_, _06546_, _06545_);
  and _14858_ (_06548_, _06547_, _06544_);
  not _14859_ (_06549_, _06548_);
  not _14860_ (_06550_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not _14861_ (_06551_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand _14862_ (_06552_, _06551_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _14863_ (_06553_, _06552_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _14864_ (_06554_, _06553_, _06550_);
  nor _14865_ (_06555_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _14866_ (_06556_, _06555_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  nand _14867_ (_06557_, _06556_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and _14868_ (_06558_, _06557_, _06554_);
  not _14869_ (_06559_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  or _14870_ (_06560_, _06552_, _06559_);
  not _14871_ (_06561_, _06560_);
  nand _14872_ (_06562_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _14873_ (_06563_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _14874_ (_06564_, _06563_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _14875_ (_06565_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _14876_ (_06566_, _06565_, _06562_);
  and _14877_ (_06567_, _06566_, _06558_);
  and _14878_ (_06568_, _06555_, _06551_);
  not _14879_ (_06569_, _06568_);
  not _14880_ (_06570_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and _14881_ (_06572_, _06570_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or _14882_ (_06573_, _06572_, ABINPUT[8]);
  nand _14883_ (_06574_, _06570_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  or _14884_ (_06575_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand _14885_ (_06576_, _06575_, _06573_);
  or _14886_ (_06577_, _06576_, _06569_);
  and _14887_ (_06578_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and _14888_ (_06579_, _06578_, _06559_);
  nand _14889_ (_06581_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _14890_ (_06582_, _06578_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand _14891_ (_06583_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and _14892_ (_06584_, _06583_, _06581_);
  and _14893_ (_06585_, _06584_, _06577_);
  and _14894_ (_06586_, _06585_, _06567_);
  nor _14895_ (_06587_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not _14896_ (_06588_, _06587_);
  or _14897_ (_06589_, _06588_, _06576_);
  nand _14898_ (_06590_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _14899_ (_06591_, _06590_, _06550_);
  not _14900_ (_06592_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  not _14901_ (_06593_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand _14902_ (_06594_, _06593_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or _14903_ (_06595_, _06594_, _06592_);
  and _14904_ (_06596_, _06595_, _06591_);
  and _14905_ (_06597_, _06596_, _06589_);
  nor _14906_ (_06598_, _06597_, _06586_);
  not _14907_ (_06599_, _06598_);
  not _14908_ (_06600_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  or _14909_ (_06601_, _06553_, _06600_);
  nand _14910_ (_06602_, _06556_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  and _14911_ (_06603_, _06602_, _06601_);
  nand _14912_ (_06604_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nand _14913_ (_06605_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _14914_ (_06606_, _06605_, _06604_);
  and _14915_ (_06607_, _06606_, _06603_);
  or _14916_ (_06608_, _06572_, ABINPUT[6]);
  or _14917_ (_06609_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand _14918_ (_06610_, _06609_, _06608_);
  or _14919_ (_06611_, _06610_, _06569_);
  nand _14920_ (_06612_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  nand _14921_ (_06613_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _14922_ (_06614_, _06613_, _06612_);
  and _14923_ (_06615_, _06614_, _06611_);
  nand _14924_ (_06616_, _06615_, _06607_);
  or _14925_ (_06617_, _06610_, _06588_);
  or _14926_ (_06618_, _06590_, _06600_);
  not _14927_ (_06619_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or _14928_ (_06620_, _06594_, _06619_);
  and _14929_ (_06621_, _06620_, _06618_);
  and _14930_ (_06622_, _06621_, _06617_);
  not _14931_ (_06623_, _06622_);
  and _14932_ (_06624_, _06623_, _06616_);
  nor _14933_ (_06625_, _06623_, _06616_);
  nor _14934_ (_06627_, _06625_, _06624_);
  not _14935_ (_06628_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  or _14936_ (_06629_, _06553_, _06628_);
  nand _14937_ (_06630_, _06556_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  and _14938_ (_06631_, _06630_, _06629_);
  nand _14939_ (_06632_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nand _14940_ (_06633_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _14941_ (_06634_, _06633_, _06632_);
  and _14942_ (_06635_, _06634_, _06631_);
  or _14943_ (_06636_, _06572_, ABINPUT[5]);
  or _14944_ (_06637_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand _14945_ (_06639_, _06637_, _06636_);
  or _14946_ (_06640_, _06639_, _06569_);
  nand _14947_ (_06642_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _14948_ (_06643_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  and _14949_ (_06644_, _06643_, _06642_);
  and _14950_ (_06645_, _06644_, _06640_);
  and _14951_ (_06646_, _06645_, _06635_);
  or _14952_ (_06647_, _06639_, _06588_);
  or _14953_ (_06648_, _06590_, _06628_);
  not _14954_ (_06649_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or _14955_ (_06650_, _06594_, _06649_);
  and _14956_ (_06651_, _06650_, _06648_);
  and _14957_ (_06652_, _06651_, _06647_);
  nor _14958_ (_06653_, _06652_, _06646_);
  and _14959_ (_06654_, _06652_, _06646_);
  nor _14960_ (_06655_, _06654_, _06653_);
  nand _14961_ (_06656_, _06556_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  not _14962_ (_06657_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  or _14963_ (_06658_, _06553_, _06657_);
  and _14964_ (_06659_, _06658_, _06656_);
  nand _14965_ (_06660_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nand _14966_ (_06661_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _14967_ (_06662_, _06661_, _06660_);
  and _14968_ (_06663_, _06662_, _06659_);
  or _14969_ (_06664_, _06572_, ABINPUT[4]);
  or _14970_ (_06665_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand _14971_ (_06666_, _06665_, _06664_);
  or _14972_ (_06667_, _06666_, _06569_);
  nand _14973_ (_06668_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand _14974_ (_06669_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and _14975_ (_06670_, _06669_, _06668_);
  and _14976_ (_06672_, _06670_, _06667_);
  and _14977_ (_06673_, _06672_, _06663_);
  or _14978_ (_06675_, _06666_, _06588_);
  or _14979_ (_06676_, _06590_, _06657_);
  not _14980_ (_06677_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _14981_ (_06678_, _06594_, _06677_);
  and _14982_ (_06679_, _06678_, _06676_);
  and _14983_ (_06680_, _06679_, _06675_);
  nor _14984_ (_06681_, _06680_, _06673_);
  and _14985_ (_06682_, _06680_, _06673_);
  nor _14986_ (_06683_, _06682_, _06681_);
  nand _14987_ (_06684_, _06556_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  not _14988_ (_06685_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or _14989_ (_06686_, _06553_, _06685_);
  and _14990_ (_06687_, _06686_, _06684_);
  nand _14991_ (_06688_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  nand _14992_ (_06689_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _14993_ (_06690_, _06689_, _06688_);
  and _14994_ (_06691_, _06690_, _06687_);
  nand _14995_ (_06692_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand _14996_ (_06693_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _14997_ (_06694_, _06693_, _06692_);
  or _14998_ (_06695_, _06572_, ABINPUT[3]);
  or _14999_ (_06696_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand _15000_ (_06697_, _06696_, _06695_);
  or _15001_ (_06698_, _06697_, _06569_);
  and _15002_ (_06699_, _06698_, _06694_);
  nand _15003_ (_06700_, _06699_, _06691_);
  or _15004_ (_06701_, _06697_, _06588_);
  or _15005_ (_06702_, _06590_, _06685_);
  not _15006_ (_06703_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _15007_ (_06704_, _06594_, _06703_);
  and _15008_ (_06705_, _06704_, _06702_);
  nand _15009_ (_06706_, _06705_, _06701_);
  and _15010_ (_06707_, _06706_, _06700_);
  nor _15011_ (_06708_, _06706_, _06700_);
  nor _15012_ (_06709_, _06708_, _06707_);
  not _15013_ (_06710_, _06709_);
  nand _15014_ (_06711_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  nand _15015_ (_06712_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and _15016_ (_06713_, _06712_, _06711_);
  not _15017_ (_06714_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or _15018_ (_06715_, _06560_, _06714_);
  not _15019_ (_06716_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or _15020_ (_06717_, _06553_, _06716_);
  and _15021_ (_06718_, _06717_, _06715_);
  and _15022_ (_06719_, _06718_, _06713_);
  or _15023_ (_06720_, _06572_, ABINPUT[2]);
  or _15024_ (_06721_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand _15025_ (_06722_, _06721_, _06720_);
  or _15026_ (_06723_, _06722_, _06569_);
  nand _15027_ (_06724_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _15028_ (_06725_, _06556_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and _15029_ (_06726_, _06725_, _06724_);
  and _15030_ (_06727_, _06726_, _06723_);
  and _15031_ (_06728_, _06727_, _06719_);
  or _15032_ (_06729_, _06722_, _06588_);
  or _15033_ (_06730_, _06590_, _06716_);
  not _15034_ (_06731_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _15035_ (_06732_, _06594_, _06731_);
  and _15036_ (_06733_, _06732_, _06730_);
  nand _15037_ (_06734_, _06733_, _06729_);
  not _15038_ (_06735_, _06734_);
  nor _15039_ (_06736_, _06735_, _06728_);
  not _15040_ (_06737_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor _15041_ (_06738_, _06553_, _06737_);
  and _15042_ (_06739_, _06556_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nor _15043_ (_06740_, _06739_, _06738_);
  and _15044_ (_06741_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _15045_ (_06742_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor _15046_ (_06743_, _06742_, _06741_);
  and _15047_ (_06744_, _06743_, _06740_);
  or _15048_ (_06745_, _06572_, ABINPUT[1]);
  or _15049_ (_06746_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and _15050_ (_06747_, _06746_, _06745_);
  and _15051_ (_06748_, _06747_, _06568_);
  not _15052_ (_06749_, _06748_);
  and _15053_ (_06750_, _06561_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _15054_ (_06751_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  nor _15055_ (_06752_, _06751_, _06750_);
  and _15056_ (_06753_, _06752_, _06749_);
  and _15057_ (_06754_, _06753_, _06744_);
  nand _15058_ (_06755_, _06747_, _06587_);
  or _15059_ (_06756_, _06590_, _06737_);
  not _15060_ (_06757_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _15061_ (_06758_, _06594_, _06757_);
  and _15062_ (_06759_, _06758_, _06756_);
  nand _15063_ (_06760_, _06759_, _06755_);
  not _15064_ (_06761_, _06760_);
  nor _15065_ (_06762_, _06761_, _06754_);
  and _15066_ (_06763_, _06735_, _06728_);
  nor _15067_ (_06764_, _06763_, _06736_);
  and _15068_ (_06765_, _06764_, _06762_);
  nor _15069_ (_06766_, _06765_, _06736_);
  nor _15070_ (_06767_, _06766_, _06710_);
  nor _15071_ (_06768_, _06767_, _06707_);
  nor _15072_ (_06769_, _06768_, _06683_);
  and _15073_ (_06770_, _06768_, _06683_);
  nor _15074_ (_06771_, _06770_, _06769_);
  and _15075_ (_06772_, \oc8051_top_1.oc8051_decoder1.cy_sel [0], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _15076_ (_06773_, _06772_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nor _15077_ (_06774_, _06572_, ABINPUT[0]);
  nor _15078_ (_06775_, _06574_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _15079_ (_06776_, _06775_, _06774_);
  nor _15080_ (_06777_, _06776_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor _15081_ (_06778_, _06777_, _06773_);
  and _15082_ (_06779_, _06761_, _06754_);
  nor _15083_ (_06780_, _06779_, _06762_);
  and _15084_ (_06781_, _06780_, _06778_);
  and _15085_ (_06782_, _06781_, _06764_);
  and _15086_ (_06783_, _06766_, _06710_);
  nor _15087_ (_06784_, _06783_, _06767_);
  and _15088_ (_06785_, _06784_, _06782_);
  not _15089_ (_06786_, _06785_);
  nor _15090_ (_06787_, _06786_, _06771_);
  nor _15091_ (_06788_, _06768_, _06682_);
  or _15092_ (_06789_, _06788_, _06681_);
  or _15093_ (_06790_, _06789_, _06787_);
  and _15094_ (_06791_, _06790_, _06655_);
  and _15095_ (_06792_, _06791_, _06627_);
  nand _15096_ (_06793_, _06556_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not _15097_ (_06794_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  or _15098_ (_06795_, _06553_, _06794_);
  and _15099_ (_06796_, _06795_, _06793_);
  nand _15100_ (_06797_, _06564_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not _15101_ (_06798_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _15102_ (_06799_, _06560_, _06798_);
  and _15103_ (_06800_, _06799_, _06797_);
  and _15104_ (_06801_, _06800_, _06796_);
  or _15105_ (_06802_, _06572_, ABINPUT[7]);
  or _15106_ (_06803_, _06574_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand _15107_ (_06804_, _06803_, _06802_);
  or _15108_ (_06805_, _06804_, _06569_);
  nand _15109_ (_06806_, _06579_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand _15110_ (_06807_, _06582_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and _15111_ (_06808_, _06807_, _06806_);
  and _15112_ (_06809_, _06808_, _06805_);
  and _15113_ (_06810_, _06809_, _06801_);
  or _15114_ (_06811_, _06804_, _06588_);
  or _15115_ (_06812_, _06590_, _06794_);
  not _15116_ (_06813_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or _15117_ (_06814_, _06594_, _06813_);
  and _15118_ (_06815_, _06814_, _06812_);
  and _15119_ (_06816_, _06815_, _06811_);
  nor _15120_ (_06817_, _06816_, _06810_);
  and _15121_ (_06818_, _06816_, _06810_);
  nor _15122_ (_06819_, _06818_, _06817_);
  not _15123_ (_06820_, _06819_);
  and _15124_ (_06821_, _06653_, _06627_);
  nor _15125_ (_06822_, _06821_, _06624_);
  nor _15126_ (_06823_, _06822_, _06820_);
  and _15127_ (_06824_, _06822_, _06820_);
  nor _15128_ (_06826_, _06824_, _06823_);
  and _15129_ (_06828_, _06826_, _06792_);
  nor _15130_ (_06830_, _06823_, _06817_);
  not _15131_ (_06832_, _06830_);
  nor _15132_ (_06834_, _06832_, _06828_);
  and _15133_ (_06835_, _06597_, _06586_);
  or _15134_ (_06837_, _06835_, _06834_);
  and _15135_ (_06839_, _06837_, _06599_);
  nor _15136_ (_06840_, _06839_, _06549_);
  not _15137_ (_06841_, _06840_);
  not _15138_ (_06842_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _15139_ (_06843_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _06406_);
  and _15140_ (_06844_, _06843_, _06842_);
  and _15141_ (_06845_, _06844_, _06547_);
  not _15142_ (_06846_, _06845_);
  not _15143_ (_06847_, _06597_);
  and _15144_ (_06848_, _06847_, _06586_);
  nor _15145_ (_06849_, _06835_, _06598_);
  not _15146_ (_06850_, _06816_);
  nor _15147_ (_06851_, _06850_, _06810_);
  and _15148_ (_06852_, _06622_, _06616_);
  nand _15149_ (_06853_, _06651_, _06647_);
  and _15150_ (_06854_, _06853_, _06646_);
  nor _15151_ (_06855_, _06854_, _06627_);
  nor _15152_ (_06856_, _06855_, _06852_);
  nor _15153_ (_06857_, _06856_, _06819_);
  nor _15154_ (_06858_, _06857_, _06851_);
  and _15155_ (_06859_, _06856_, _06819_);
  nor _15156_ (_06860_, _06859_, _06857_);
  not _15157_ (_06861_, _06860_);
  and _15158_ (_06862_, _06854_, _06627_);
  nor _15159_ (_06863_, _06862_, _06855_);
  not _15160_ (_06864_, _06863_);
  not _15161_ (_06865_, _06655_);
  and _15162_ (_06866_, _06760_, _06754_);
  nor _15163_ (_06867_, _06866_, _06764_);
  nor _15164_ (_06868_, _06734_, _06728_);
  nor _15165_ (_06869_, _06868_, _06867_);
  nor _15166_ (_06870_, _06869_, _06709_);
  and _15167_ (_06871_, _06705_, _06701_);
  and _15168_ (_06872_, _06871_, _06700_);
  nor _15169_ (_06873_, _06872_, _06870_);
  nor _15170_ (_06874_, _06873_, _06683_);
  and _15171_ (_06875_, _06873_, _06683_);
  nor _15172_ (_06876_, _06875_, _06874_);
  and _15173_ (_06877_, _06869_, _06709_);
  nor _15174_ (_06878_, _06877_, _06870_);
  not _15175_ (_06879_, _06878_);
  and _15176_ (_06880_, _06866_, _06764_);
  nor _15177_ (_06881_, _06880_, _06867_);
  not _15178_ (_06882_, _06881_);
  not _15179_ (_06883_, _06778_);
  nor _15180_ (_06884_, _06780_, _06883_);
  and _15181_ (_06885_, _06884_, _06882_);
  and _15182_ (_06886_, _06885_, _06879_);
  not _15183_ (_06887_, _06886_);
  nor _15184_ (_06888_, _06887_, _06876_);
  not _15185_ (_06889_, _06680_);
  or _15186_ (_06890_, _06889_, _06673_);
  and _15187_ (_06891_, _06889_, _06673_);
  or _15188_ (_06892_, _06873_, _06891_);
  and _15189_ (_06893_, _06892_, _06890_);
  or _15190_ (_06894_, _06893_, _06888_);
  and _15191_ (_06895_, _06894_, _06865_);
  and _15192_ (_06896_, _06895_, _06864_);
  and _15193_ (_06897_, _06896_, _06861_);
  nor _15194_ (_06898_, _06897_, _06858_);
  nor _15195_ (_06899_, _06898_, _06849_);
  nor _15196_ (_06900_, _06899_, _06848_);
  nor _15197_ (_06901_, _06900_, _06846_);
  not _15198_ (_06902_, _06810_);
  nor _15199_ (_06903_, _06902_, _06616_);
  not _15200_ (_06904_, _06903_);
  not _15201_ (_06905_, _06646_);
  not _15202_ (_06906_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and _15203_ (_06907_, _06545_, _06906_);
  and _15204_ (_06908_, _06907_, _06544_);
  not _15205_ (_06909_, _06728_);
  nor _15206_ (_06910_, _06909_, _06700_);
  nor _15207_ (_06911_, _06910_, _06673_);
  and _15208_ (_06912_, _06911_, _06908_);
  and _15209_ (_06913_, _06912_, _06905_);
  nor _15210_ (_06914_, _06913_, _06904_);
  nor _15211_ (_06915_, _06914_, _06586_);
  nor _15212_ (_06916_, _06915_, _06778_);
  not _15213_ (_06917_, _06916_);
  not _15214_ (_06918_, _06908_);
  nor _15215_ (_06919_, _06883_, _06586_);
  not _15216_ (_06920_, _06919_);
  nor _15217_ (_06921_, _06920_, _06914_);
  nor _15218_ (_06922_, _06921_, _06918_);
  and _15219_ (_06923_, _06922_, _06917_);
  not _15220_ (_06924_, _06754_);
  and _15221_ (_06925_, _06546_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _15222_ (_06926_, _06925_, _06544_);
  and _15223_ (_06927_, _06926_, _06924_);
  and _15224_ (_06928_, _06776_, _06773_);
  not _15225_ (_06929_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and _15226_ (_06930_, _06546_, _06929_);
  and _15227_ (_06931_, _06930_, _06844_);
  and _15228_ (_06932_, _06843_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and _15229_ (_06933_, _06932_, _06907_);
  and _15230_ (_06934_, _06933_, _06776_);
  nor _15231_ (_06935_, _06934_, _06931_);
  nor _15232_ (_06936_, _06935_, _06928_);
  nor _15233_ (_06937_, _06936_, _06927_);
  not _15234_ (_06938_, _06912_);
  nor _15235_ (_06939_, _06778_, _06776_);
  and _15236_ (_06940_, _06930_, _06544_);
  nor _15237_ (_06941_, _06843_, _06543_);
  and _15238_ (_06942_, _06930_, _06941_);
  not _15239_ (_06943_, _06942_);
  not _15240_ (_06944_, _06776_);
  nor _15241_ (_06945_, _06944_, _06773_);
  nor _15242_ (_06946_, _06945_, _06943_);
  nor _15243_ (_06947_, _06946_, _06940_);
  nor _15244_ (_06948_, _06947_, _06939_);
  and _15245_ (_06949_, _06941_, _06925_);
  and _15246_ (_06950_, _06949_, _06944_);
  and _15247_ (_06951_, _06941_, _06547_);
  nor _15248_ (_06952_, _06951_, _06950_);
  and _15249_ (_06953_, _06952_, _06778_);
  and _15250_ (_06954_, _06907_, _06844_);
  nor _15251_ (_06955_, _06954_, _06778_);
  nor _15252_ (_06956_, _06955_, _06953_);
  not _15253_ (_06957_, _06586_);
  and _15254_ (_06958_, _06930_, _06932_);
  and _15255_ (_06959_, _06958_, _06957_);
  or _15256_ (_06960_, _06959_, _06956_);
  nor _15257_ (_06961_, _06960_, _06948_);
  and _15258_ (_06962_, _06961_, _06938_);
  and _15259_ (_06963_, _06962_, _06937_);
  not _15260_ (_06964_, _06963_);
  nor _15261_ (_06965_, _06964_, _06923_);
  not _15262_ (_06966_, _06965_);
  nor _15263_ (_06967_, _06966_, _06901_);
  and _15264_ (_06968_, _06967_, _06841_);
  nor _15265_ (_06969_, _06968_, _06540_);
  not _15266_ (_06970_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or _15267_ (_06971_, _06539_, _06970_);
  nand _15268_ (_06972_, _06971_, _06501_);
  or _15269_ (_06973_, _06972_, _06969_);
  and _15270_ (_06974_, _06973_, _06502_);
  and _15271_ (_06975_, _06477_, _06434_);
  nor _15272_ (_06976_, _06499_, _06463_);
  and _15273_ (_06977_, _06976_, _06975_);
  and _15274_ (_06978_, _06537_, _06513_);
  and _15275_ (_06979_, _06978_, _06525_);
  not _15276_ (_06980_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _15277_ (_06981_, _06481_, _06980_);
  not _15278_ (_06982_, _06981_);
  nor _15279_ (_06983_, _06982_, _06483_);
  not _15280_ (_06984_, _06983_);
  nor _15281_ (_06985_, _06984_, _06447_);
  and _15282_ (_06986_, _06985_, _06979_);
  and _15283_ (_06987_, _06986_, _06977_);
  or _15284_ (_06988_, _06987_, _06974_);
  not _15285_ (_06989_, rst);
  and _15286_ (_06990_, _06883_, _06586_);
  and _15287_ (_06991_, _06932_, _06925_);
  not _15288_ (_06992_, _06991_);
  and _15289_ (_06993_, _06778_, _06597_);
  nor _15290_ (_06994_, _06993_, _06992_);
  not _15291_ (_06995_, _06994_);
  nor _15292_ (_06996_, _06995_, _06990_);
  and _15293_ (_06997_, _06925_, _06844_);
  and _15294_ (_06998_, _06910_, _06754_);
  and _15295_ (_06999_, _06998_, _06673_);
  and _15296_ (_07000_, _06999_, _06646_);
  and _15297_ (_07001_, _07000_, _06903_);
  nor _15298_ (_07002_, _07001_, _06883_);
  not _15299_ (_07003_, _06673_);
  nor _15300_ (_07004_, _06754_, _06728_);
  and _15301_ (_07005_, _07004_, _06700_);
  and _15302_ (_07006_, _07005_, _07003_);
  and _15303_ (_07007_, _07006_, _06905_);
  and _15304_ (_07008_, _07007_, _06616_);
  and _15305_ (_07009_, _07008_, _06902_);
  nor _15306_ (_07010_, _07009_, _06778_);
  or _15307_ (_07011_, _07010_, _07002_);
  and _15308_ (_07012_, _07011_, _06586_);
  nor _15309_ (_07013_, _07011_, _06586_);
  nor _15310_ (_07014_, _07013_, _07012_);
  and _15311_ (_07015_, _07014_, _06997_);
  nor _15312_ (_07016_, _07015_, _06996_);
  not _15313_ (_07017_, _06940_);
  nor _15314_ (_07018_, _07017_, _06835_);
  and _15315_ (_07019_, _06942_, _06849_);
  nor _15316_ (_07020_, _07019_, _07018_);
  and _15317_ (_07021_, _06933_, _06598_);
  and _15318_ (_07022_, _06954_, _06586_);
  nor _15319_ (_07023_, _07022_, _07021_);
  and _15320_ (_07024_, _06941_, _06907_);
  not _15321_ (_07025_, _07024_);
  and _15322_ (_07026_, _06544_, _06906_);
  and _15323_ (_07027_, _06932_, _06547_);
  nor _15324_ (_07028_, _07027_, _07026_);
  and _15325_ (_07029_, _07028_, _07025_);
  and _15326_ (_07030_, _06925_, _06541_);
  not _15327_ (_07031_, _07030_);
  and _15328_ (_07032_, _06930_, _06843_);
  nor _15329_ (_07033_, _07032_, _06951_);
  and _15330_ (_07034_, _07033_, _07031_);
  and _15331_ (_07035_, _07034_, _07029_);
  nor _15332_ (_07036_, _07035_, _06586_);
  not _15333_ (_07037_, _07036_);
  and _15334_ (_07038_, _07037_, _07023_);
  and _15335_ (_07039_, _07038_, _07020_);
  and _15336_ (_07040_, _07039_, _07016_);
  nand _15337_ (_07041_, _07040_, _06987_);
  and _15338_ (_07042_, _07041_, _06989_);
  and _15339_ (_11486_, _07042_, _06988_);
  not _15340_ (_07043_, _06525_);
  and _15341_ (_07044_, _06978_, _07043_);
  and _15342_ (_07045_, _06985_, _07044_);
  and _15343_ (_07046_, _07045_, _06977_);
  and _15344_ (_07047_, _06537_, _06514_);
  and _15345_ (_07048_, _07047_, _07043_);
  and _15346_ (_07049_, _06985_, _07048_);
  and _15347_ (_07050_, _07049_, _06977_);
  nor _15348_ (_07051_, _07050_, _07046_);
  and _15349_ (_07052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _15350_ (_07053_, _07052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _15351_ (_07054_, _07053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and _15352_ (_07055_, _07054_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and _15353_ (_07056_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and _15354_ (_07057_, _07056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and _15355_ (_07058_, _07057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _15356_ (_07059_, _07058_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and _15357_ (_07060_, _07059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _15358_ (_07061_, _07060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _15359_ (_07062_, _07061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and _15360_ (_07063_, _07062_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _15361_ (_07064_, _07063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _15362_ (_07065_, _07064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _15363_ (_07066_, _07065_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _15364_ (_07067_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not _15365_ (_07068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _15366_ (_07069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _07068_);
  and _15367_ (_07070_, _07069_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _15368_ (_07071_, _07070_, _07067_);
  nor _15369_ (_07072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not _15370_ (_07073_, _07072_);
  not _15371_ (_07074_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _15372_ (_07075_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _15373_ (_07076_, _07075_, _07072_);
  and _15374_ (_07077_, _07076_, _07074_);
  nor _15375_ (_07078_, _07077_, _07073_);
  and _15376_ (_07079_, _07078_, _07071_);
  nand _15377_ (_07080_, _07079_, _07066_);
  nand _15378_ (_07081_, _07080_, _07051_);
  or _15379_ (_07082_, _07051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _15380_ (_07083_, _07082_, _06989_);
  and _15381_ (_13884_, _07083_, _07081_);
  not _15382_ (_07084_, _06434_);
  and _15383_ (_07085_, _06477_, _07084_);
  and _15384_ (_07086_, _06499_, _06463_);
  and _15385_ (_07087_, _07086_, _07085_);
  and _15386_ (_07088_, _06537_, _06525_);
  and _15387_ (_07089_, _07088_, _06514_);
  and _15388_ (_07090_, _07089_, _06448_);
  and _15389_ (_07091_, _07090_, _07087_);
  and _15390_ (_07092_, _06778_, _06623_);
  and _15391_ (_07093_, _06883_, _06616_);
  or _15392_ (_07094_, _07093_, _07092_);
  and _15393_ (_07095_, _07094_, _06991_);
  not _15394_ (_07096_, _06616_);
  and _15395_ (_07097_, _07007_, _06883_);
  and _15396_ (_07098_, _07000_, _06778_);
  nor _15397_ (_07099_, _07098_, _07097_);
  and _15398_ (_07100_, _07099_, _07096_);
  not _15399_ (_07101_, _06997_);
  nor _15400_ (_07102_, _07099_, _07096_);
  or _15401_ (_07103_, _07102_, _07101_);
  nor _15402_ (_07104_, _07103_, _07100_);
  nor _15403_ (_07105_, _07104_, _07095_);
  not _15404_ (_07106_, _07035_);
  and _15405_ (_07107_, _07106_, _06616_);
  not _15406_ (_07108_, _07107_);
  and _15407_ (_07109_, _06942_, _06627_);
  nor _15408_ (_07110_, _07017_, _06625_);
  not _15409_ (_07111_, _07110_);
  and _15410_ (_07112_, _06933_, _06624_);
  and _15411_ (_07113_, _06954_, _07096_);
  nor _15412_ (_07114_, _07113_, _07112_);
  nand _15413_ (_07115_, _07114_, _07111_);
  nor _15414_ (_07116_, _07115_, _07109_);
  and _15415_ (_07117_, _07116_, _07108_);
  and _15416_ (_07118_, _07117_, _07105_);
  not _15417_ (_07119_, _07118_);
  and _15418_ (_07120_, _07119_, _07091_);
  not _15419_ (_07121_, _07087_);
  nand _15420_ (_07122_, _07089_, _06447_);
  nor _15421_ (_07123_, _07122_, _07121_);
  and _15422_ (_07124_, _06525_, _06447_);
  and _15423_ (_07125_, _07124_, _06978_);
  and _15424_ (_07126_, _07125_, _07087_);
  nor _15425_ (_07127_, _07126_, _07123_);
  and _15426_ (_07128_, _06979_, _06448_);
  and _15427_ (_07129_, _07087_, _07128_);
  not _15428_ (_07130_, _07129_);
  and _15429_ (_07131_, _07130_, _07127_);
  not _15430_ (_07132_, _07131_);
  and _15431_ (_07133_, _06981_, _07088_);
  nand _15432_ (_07134_, _07133_, _07087_);
  or _15433_ (_07135_, _07134_, _07132_);
  and _15434_ (_07136_, _07135_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  or _15435_ (_07137_, _07136_, _07120_);
  or _15436_ (_07138_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and _15437_ (_07139_, _07138_, _06989_);
  and _15438_ (_06571_, _07139_, _07137_);
  and _15439_ (_07140_, _07071_, _07064_);
  and _15440_ (_07141_, _07140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _15441_ (_07142_, _07141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand _15442_ (_07143_, _07141_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _15443_ (_07144_, _07143_, _07142_);
  and _15444_ (_07145_, _07072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not _15445_ (_07146_, _07145_);
  and _15446_ (_07147_, _07146_, _07071_);
  and _15447_ (_07148_, _07147_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _15448_ (_07149_, _07148_, _07066_);
  or _15449_ (_07150_, _07149_, _07077_);
  or _15450_ (_07151_, _07150_, _07144_);
  not _15451_ (_07152_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _15452_ (_07153_, _07077_, _07152_);
  nor _15453_ (_07154_, _07153_, _07046_);
  and _15454_ (_07155_, _07154_, _07151_);
  and _15455_ (_07156_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _15456_ (_07157_, _07156_, _07050_);
  or _15457_ (_07158_, _07157_, _07155_);
  nand _15458_ (_07159_, _07050_, _07040_);
  and _15459_ (_07160_, _07159_, _06989_);
  and _15460_ (_10680_, _07160_, _07158_);
  and _15461_ (_07161_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and _15462_ (_07162_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _15463_ (_12565_, _07162_, _07161_);
  not _15464_ (_07164_, _07161_);
  not _15465_ (_07165_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not _15466_ (_07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _15467_ (_07167_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _07166_);
  and _15468_ (_07168_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _15469_ (_07169_, _07168_, _07167_);
  and _15470_ (_07170_, _07169_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor _15471_ (_07171_, _07170_, _07165_);
  not _15472_ (_07172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor _15473_ (_07173_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor _15474_ (_07174_, _07173_, _07172_);
  and _15475_ (_07175_, _07174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not _15476_ (_07176_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor _15477_ (_07177_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor _15478_ (_07178_, _07177_, _07176_);
  and _15479_ (_07179_, _07178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  nor _15480_ (_07180_, _07179_, _07175_);
  and _15481_ (_07181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _15482_ (_07182_, _07181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not _15483_ (_07183_, _07182_);
  and _15484_ (_07184_, _07183_, _07180_);
  and _15485_ (_07185_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _15486_ (_07186_, _07185_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not _15487_ (_07187_, _07186_);
  and _15488_ (_07188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and _15489_ (_07189_, _07188_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _15490_ (_07190_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _15491_ (_07191_, _07190_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor _15492_ (_07193_, _07191_, _07189_);
  and _15493_ (_07194_, _07193_, _07187_);
  and _15494_ (_07195_, _07194_, _07184_);
  nor _15495_ (_07196_, _07195_, _07171_);
  not _15496_ (_07197_, _07196_);
  and _15497_ (_07198_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _07165_);
  not _15498_ (_07199_, _07198_);
  not _15499_ (_07200_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _15500_ (_07201_, _07185_, _07200_);
  not _15501_ (_07202_, _07201_);
  not _15502_ (_07203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _15503_ (_07204_, _07188_, _07203_);
  not _15504_ (_07205_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _15505_ (_07206_, _07190_, _07205_);
  nor _15506_ (_07207_, _07206_, _07204_);
  and _15507_ (_07208_, _07207_, _07202_);
  nor _15508_ (_07209_, _07208_, _07199_);
  not _15509_ (_07210_, _07209_);
  not _15510_ (_07211_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _15511_ (_07212_, _07174_, _07211_);
  not _15512_ (_07213_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _15513_ (_07215_, _07178_, _07213_);
  nor _15514_ (_07216_, _07215_, _07212_);
  not _15515_ (_07217_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and _15516_ (_07218_, _07181_, _07217_);
  not _15517_ (_07219_, _07218_);
  and _15518_ (_07220_, _07219_, _07216_);
  or _15519_ (_07221_, _07220_, _07199_);
  and _15520_ (_07222_, _07221_, _07210_);
  and _15521_ (_07223_, _07222_, _07197_);
  and _15522_ (_07224_, _07223_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _15523_ (_07225_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and _15524_ (_07226_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor _15525_ (_07227_, _07226_, _07225_);
  nor _15526_ (_07228_, _07227_, _07197_);
  or _15527_ (_07229_, _07228_, _07224_);
  and _15528_ (_07230_, _07229_, _07164_);
  and _15529_ (_07231_, _07227_, _07161_);
  or _15530_ (_07232_, _07231_, _07230_);
  and _15531_ (_12832_, _07232_, _06989_);
  and _15532_ (_07233_, _07195_, _07165_);
  nand _15533_ (_07234_, _07233_, _07222_);
  nand _15534_ (_07235_, _07225_, _07161_);
  and _15535_ (_07236_, _07235_, _06989_);
  and _15536_ (_12851_, _07236_, _07234_);
  nor _15537_ (_07237_, _06778_, _06646_);
  and _15538_ (_07238_, _06778_, _06853_);
  or _15539_ (_07239_, _07238_, _07237_);
  and _15540_ (_07240_, _07239_, _06991_);
  nor _15541_ (_07242_, _07006_, _06778_);
  nor _15542_ (_07243_, _06999_, _06883_);
  nor _15543_ (_07244_, _07243_, _07242_);
  nor _15544_ (_07245_, _07244_, _06905_);
  and _15545_ (_07246_, _07244_, _06905_);
  nor _15546_ (_07247_, _07246_, _07245_);
  and _15547_ (_07248_, _07247_, _06997_);
  nor _15548_ (_07249_, _07248_, _07240_);
  and _15549_ (_07250_, _06942_, _06655_);
  and _15550_ (_07251_, _06933_, _06653_);
  nor _15551_ (_07252_, _07017_, _06654_);
  and _15552_ (_07253_, _06954_, _06646_);
  or _15553_ (_07254_, _07253_, _07252_);
  or _15554_ (_07255_, _07254_, _07251_);
  nor _15555_ (_07256_, _07255_, _07250_);
  nor _15556_ (_07257_, _07035_, _06646_);
  not _15557_ (_07258_, _07257_);
  and _15558_ (_07259_, _07258_, _07256_);
  and _15559_ (_07260_, _07259_, _07249_);
  and _15560_ (_07261_, _07129_, _06981_);
  not _15561_ (_07262_, _07261_);
  nor _15562_ (_07263_, _07262_, _07260_);
  and _15563_ (_07264_, _07262_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  or _15564_ (_07265_, _07264_, _07263_);
  and _15565_ (_13225_, _07265_, _06989_);
  and _15566_ (_07266_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  not _15567_ (_07267_, _07184_);
  or _15568_ (_07268_, _07194_, _07171_);
  or _15569_ (_07269_, _07268_, _07267_);
  and _15570_ (_07270_, _07269_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand _15571_ (_07271_, _07221_, _07197_);
  and _15572_ (_07272_, _07271_, _07270_);
  or _15573_ (_07273_, _07272_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor _15574_ (_07274_, _07222_, _07196_);
  nor _15575_ (_07275_, _07208_, _07166_);
  nand _15576_ (_07276_, _07275_, _07274_);
  nor _15577_ (_07277_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and _15578_ (_07278_, _07268_, _07164_);
  or _15579_ (_07279_, _07278_, _07277_);
  and _15580_ (_07281_, _07279_, _07276_);
  and _15581_ (_07282_, _07281_, _07273_);
  or _15582_ (_07283_, _07282_, _07266_);
  and _15583_ (_13415_, _07283_, _06989_);
  and _15584_ (_07284_, _07125_, _06983_);
  and _15585_ (_07285_, _07284_, _06976_);
  and _15586_ (_07286_, _06434_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _15587_ (_07287_, _07085_, _06976_);
  and _15588_ (_07288_, _07287_, _07284_);
  not _15589_ (_07289_, _07288_);
  and _15590_ (_07290_, _07289_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _15591_ (_07291_, _07285_, _07085_);
  not _15592_ (_07292_, _07291_);
  nor _15593_ (_07293_, _07292_, _07260_);
  nor _15594_ (_07294_, _07293_, _07290_);
  and _15595_ (_07295_, _07294_, _07084_);
  nor _15596_ (_07296_, _07295_, _07286_);
  and _15597_ (_07297_, _07289_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor _15598_ (_07298_, _06998_, _06883_);
  nor _15599_ (_07299_, _07005_, _06778_);
  nor _15600_ (_07300_, _07299_, _07298_);
  nor _15601_ (_07301_, _07300_, _07003_);
  not _15602_ (_07302_, _07301_);
  and _15603_ (_07303_, _07300_, _07003_);
  nor _15604_ (_07304_, _07303_, _07101_);
  and _15605_ (_07305_, _07304_, _07302_);
  nor _15606_ (_07306_, _06992_, _06680_);
  nor _15607_ (_07307_, _07306_, _07305_);
  and _15608_ (_07308_, _06933_, _06681_);
  and _15609_ (_07309_, _06954_, _06673_);
  nor _15610_ (_07310_, _07309_, _07308_);
  nor _15611_ (_07311_, _07035_, _06673_);
  and _15612_ (_07312_, _06942_, _06683_);
  nor _15613_ (_07313_, _07017_, _06682_);
  or _15614_ (_07314_, _07313_, _07312_);
  nor _15615_ (_07315_, _07314_, _07311_);
  and _15616_ (_07316_, _07315_, _07310_);
  and _15617_ (_07317_, _07316_, _07307_);
  nor _15618_ (_07318_, _07317_, _07292_);
  nor _15619_ (_07319_, _07318_, _07297_);
  and _15620_ (_07320_, _07319_, _06448_);
  not _15621_ (_07321_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor _15622_ (_07322_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _15623_ (_07323_, _07322_, _07321_);
  nor _15624_ (_07324_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  and _15625_ (_07325_, _07324_, _06406_);
  and _15626_ (_07326_, _07325_, _07323_);
  not _15627_ (_07327_, _07326_);
  not _15628_ (_07328_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _15629_ (_07330_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not _15630_ (_07331_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _15631_ (_07332_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _15632_ (_07333_, _07332_, _07331_);
  and _15633_ (_07334_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not _15634_ (_07335_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _15635_ (_07337_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], _07335_);
  and _15636_ (_07338_, _07337_, _07331_);
  and _15637_ (_07339_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _15638_ (_07340_, _07339_, _07334_);
  nor _15639_ (_07341_, _07332_, _07331_);
  nand _15640_ (_07342_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _15641_ (_07343_, _07332_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _15642_ (_07344_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _15643_ (_07345_, _07344_, _07342_);
  and _15644_ (_07346_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _15645_ (_07347_, _07346_, _07331_);
  nand _15646_ (_07348_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  not _15647_ (_07349_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _15648_ (_07350_, _07349_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _15649_ (_07351_, _07350_, _07331_);
  nand _15650_ (_07352_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and _15651_ (_07353_, _07352_, _07348_);
  and _15652_ (_07354_, _07353_, _07345_);
  nand _15653_ (_07355_, _07354_, _07340_);
  nand _15654_ (_07356_, _07355_, _07330_);
  nand _15655_ (_07357_, _07356_, _07328_);
  nor _15656_ (_07358_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _07328_);
  not _15657_ (_07359_, _07358_);
  and _15658_ (_07360_, _07359_, _07357_);
  or _15659_ (_07361_, _07360_, _07327_);
  not _15660_ (_07362_, _07323_);
  nor _15661_ (_07363_, _07325_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor _15662_ (_07364_, _07363_, _07362_);
  and _15663_ (_07365_, _07364_, _07361_);
  nor _15664_ (_07366_, _07365_, _06513_);
  not _15665_ (_07367_, _07366_);
  nand _15666_ (_07368_, _07367_, _07086_);
  nor _15667_ (_07369_, _07368_, _07320_);
  nor _15668_ (_07370_, _07319_, _06448_);
  and _15669_ (_07371_, _07365_, _06513_);
  nand _15670_ (_07372_, _06981_, _06525_);
  nand _15671_ (_07373_, _06537_, _06477_);
  or _15672_ (_07374_, _07373_, _07372_);
  or _15673_ (_07375_, _07374_, _07371_);
  nor _15674_ (_07376_, _07375_, _07370_);
  and _15675_ (_07377_, _07376_, _07369_);
  and _15676_ (_07378_, _07377_, _07296_);
  nor _15677_ (_07379_, _07365_, _07319_);
  and _15678_ (_07380_, _07379_, _07294_);
  and _15679_ (_07381_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  not _15680_ (_07382_, _07294_);
  not _15681_ (_07383_, _07365_);
  nor _15682_ (_07384_, _07383_, _07319_);
  and _15683_ (_07385_, _07384_, _07382_);
  and _15684_ (_07386_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _15685_ (_07387_, _07386_, _07381_);
  and _15686_ (_07389_, _07379_, _07382_);
  and _15687_ (_07390_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and _15688_ (_07391_, _07383_, _07319_);
  and _15689_ (_07392_, _07391_, _07382_);
  and _15690_ (_07393_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor _15691_ (_07394_, _07393_, _07390_);
  and _15692_ (_07395_, _07394_, _07387_);
  and _15693_ (_07396_, _07391_, _07294_);
  and _15694_ (_07397_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _15695_ (_07398_, _07384_, _07294_);
  and _15696_ (_07399_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor _15697_ (_07400_, _07399_, _07397_);
  and _15698_ (_07401_, _07365_, _07319_);
  and _15699_ (_07402_, _07401_, _07382_);
  and _15700_ (_07403_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  and _15701_ (_07404_, _07401_, _07294_);
  and _15702_ (_07405_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor _15703_ (_07406_, _07405_, _07403_);
  and _15704_ (_07407_, _07406_, _07400_);
  and _15705_ (_07408_, _07407_, _07395_);
  nor _15706_ (_07409_, _07408_, _07378_);
  not _15707_ (_07410_, _07317_);
  and _15708_ (_07411_, _07378_, _07410_);
  nor _15709_ (_07412_, _07411_, _07409_);
  nor _15710_ (_14142_, _07412_, rst);
  and _15711_ (_07413_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and _15712_ (_07414_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor _15713_ (_07415_, _07414_, _07413_);
  and _15714_ (_07416_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and _15715_ (_07417_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor _15716_ (_07418_, _07417_, _07416_);
  and _15717_ (_07419_, _07418_, _07415_);
  and _15718_ (_07420_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _15719_ (_07421_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor _15720_ (_07422_, _07421_, _07420_);
  and _15721_ (_07423_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and _15722_ (_07424_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor _15723_ (_07425_, _07424_, _07423_);
  and _15724_ (_07426_, _07425_, _07422_);
  and _15725_ (_07427_, _07426_, _07419_);
  nor _15726_ (_07428_, _07427_, _07378_);
  not _15727_ (_07429_, _07260_);
  and _15728_ (_07430_, _07378_, _07429_);
  nor _15729_ (_07431_, _07430_, _07428_);
  nor _15730_ (_14393_, _07431_, rst);
  and _15731_ (_07432_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _15732_ (_07433_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor _15733_ (_07434_, _07433_, _07432_);
  and _15734_ (_07435_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and _15735_ (_07436_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor _15736_ (_07437_, _07436_, _07435_);
  and _15737_ (_07438_, _07437_, _07434_);
  and _15738_ (_07439_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and _15739_ (_07440_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  nor _15740_ (_07441_, _07440_, _07439_);
  and _15741_ (_07442_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and _15742_ (_07443_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nor _15743_ (_07444_, _07443_, _07442_);
  and _15744_ (_07445_, _07444_, _07441_);
  and _15745_ (_07446_, _07445_, _07438_);
  nor _15746_ (_07447_, _07446_, _07378_);
  and _15747_ (_07449_, _07378_, _07119_);
  nor _15748_ (_07450_, _07449_, _07447_);
  nor _15749_ (_01178_, _07450_, rst);
  not _15750_ (_07452_, _06463_);
  nor _15751_ (_07453_, _06499_, _07452_);
  and _15752_ (_07454_, _07453_, _06975_);
  nor _15753_ (_07455_, _06486_, _06447_);
  and _15754_ (_07456_, _07455_, _06539_);
  and _15755_ (_07457_, _07456_, _07454_);
  nand _15756_ (_07458_, _07457_, _06968_);
  and _15757_ (_07459_, _07454_, _06986_);
  not _15758_ (_07460_, _07459_);
  nor _15759_ (_07461_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _15760_ (_07462_, _07461_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  not _15761_ (_07463_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and _15762_ (_07464_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and _15763_ (_07465_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor _15764_ (_07466_, _07465_, _07464_);
  nor _15765_ (_07467_, _07466_, _07165_);
  or _15766_ (_07468_, _07467_, _07463_);
  nor _15767_ (_07469_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _15768_ (_07470_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or _15769_ (_07471_, _07470_, _07165_);
  nor _15770_ (_07472_, _07471_, _07469_);
  and _15771_ (_07473_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _15772_ (_07474_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor _15773_ (_07475_, _07474_, _07473_);
  nand _15774_ (_07476_, _07475_, _07472_);
  or _15775_ (_07477_, _07476_, _07468_);
  and _15776_ (_07478_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or _15777_ (_07479_, _07478_, _07462_);
  or _15778_ (_07480_, _07479_, _07457_);
  and _15779_ (_07481_, _07480_, _07460_);
  and _15780_ (_07482_, _07481_, _07458_);
  nor _15781_ (_07483_, _07460_, _07040_);
  or _15782_ (_07484_, _07483_, _07482_);
  and _15783_ (_01362_, _07484_, _06989_);
  and _15784_ (_07485_, _07126_, _06981_);
  not _15785_ (_07486_, _07485_);
  nor _15786_ (_07487_, _07486_, _07317_);
  and _15787_ (_07488_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or _15788_ (_07489_, _07488_, _07487_);
  and _15789_ (_01526_, _07489_, _06989_);
  not _15790_ (_07490_, _07325_);
  nor _15791_ (_07491_, _07346_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor _15792_ (_07492_, _07491_, _07490_);
  nor _15793_ (_07493_, _07492_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and _15794_ (_07494_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  not _15795_ (_07495_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor _15796_ (_07496_, _07493_, _07495_);
  or _15797_ (_07497_, _07496_, _07494_);
  and _15798_ (_03985_, _07497_, _06989_);
  and _15799_ (_07498_, _06951_, _06734_);
  and _15800_ (_07499_, _06958_, _06616_);
  and _15801_ (_07500_, _07001_, _06586_);
  and _15802_ (_07501_, _07500_, _06761_);
  and _15803_ (_07502_, _07501_, _06778_);
  nor _15804_ (_07504_, _06761_, _06586_);
  and _15805_ (_07505_, _07504_, _07009_);
  and _15806_ (_07506_, _07505_, _06883_);
  nor _15807_ (_07507_, _07506_, _07502_);
  nor _15808_ (_07508_, _07507_, _06734_);
  and _15809_ (_07509_, _07507_, _06734_);
  nor _15810_ (_07510_, _07509_, _07508_);
  nor _15811_ (_07511_, _07510_, _07101_);
  nor _15812_ (_07512_, _06992_, _06728_);
  or _15813_ (_07513_, _07512_, _07511_);
  or _15814_ (_07514_, _07513_, _07499_);
  nor _15815_ (_07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _15816_ (_07516_, _07515_, _06586_);
  nor _15817_ (_07517_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not _15818_ (_07518_, _07517_);
  and _15819_ (_07519_, _07518_, _07516_);
  not _15820_ (_07520_, _07519_);
  or _15821_ (_07521_, _06760_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  not _15822_ (_07522_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15823_ (_07523_, _06706_, _07522_);
  and _15824_ (_07524_, _07523_, _07521_);
  or _15825_ (_07525_, _07524_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15826_ (_07526_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _15827_ (_07527_, _06853_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _15828_ (_07528_, _06816_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _15829_ (_07529_, _07528_, _07527_);
  or _15830_ (_07530_, _07529_, _07526_);
  and _15831_ (_07531_, _07530_, _07525_);
  or _15832_ (_07532_, _07531_, _07520_);
  not _15833_ (_07533_, _07531_);
  or _15834_ (_07534_, _07533_, _07519_);
  not _15835_ (_07535_, _07534_);
  nand _15836_ (_07536_, _07515_, _06810_);
  nor _15837_ (_07537_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not _15838_ (_07538_, _07537_);
  and _15839_ (_07539_, _07538_, _07536_);
  not _15840_ (_07540_, _07539_);
  and _15841_ (_07541_, _06734_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15842_ (_07542_, _07541_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand _15843_ (_07543_, _06680_, _07522_);
  nand _15844_ (_07544_, _06622_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _15845_ (_07545_, _07544_, _07543_);
  or _15846_ (_07546_, _07545_, _07526_);
  and _15847_ (_07547_, _07546_, _07542_);
  or _15848_ (_07548_, _07547_, _07540_);
  or _15849_ (_07549_, _07548_, _07535_);
  and _15850_ (_07550_, _07549_, _07532_);
  and _15851_ (_07551_, _07534_, _07532_);
  nand _15852_ (_07552_, _07547_, _07540_);
  and _15853_ (_07553_, _07552_, _07548_);
  and _15854_ (_07554_, _07553_, _07551_);
  not _15855_ (_07555_, _07515_);
  or _15856_ (_07556_, _07555_, _06616_);
  nor _15857_ (_07557_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not _15858_ (_07558_, _07557_);
  nand _15859_ (_07559_, _07558_, _07556_);
  and _15860_ (_07560_, _06760_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15861_ (_07561_, _07560_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  or _15862_ (_07562_, _06706_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _15863_ (_07563_, _06853_, _07522_);
  and _15864_ (_07564_, _07563_, _07562_);
  or _15865_ (_07565_, _07564_, _07526_);
  and _15866_ (_07566_, _07565_, _07561_);
  nor _15867_ (_07567_, _07566_, _07559_);
  or _15868_ (_07568_, _06734_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _15869_ (_07569_, _06680_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and _15870_ (_07570_, _07569_, _07568_);
  and _15871_ (_07571_, _07570_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15872_ (_07572_, _07571_);
  nand _15873_ (_07573_, _07515_, _06646_);
  nor _15874_ (_07574_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not _15875_ (_07575_, _07574_);
  and _15876_ (_07576_, _07575_, _07573_);
  and _15877_ (_07577_, _07576_, _07572_);
  and _15878_ (_07579_, _07566_, _07559_);
  or _15879_ (_07580_, _07579_, _07567_);
  not _15880_ (_07582_, _07580_);
  and _15881_ (_07583_, _07582_, _07577_);
  or _15882_ (_07585_, _07583_, _07567_);
  nand _15883_ (_07586_, _07585_, _07554_);
  and _15884_ (_07587_, _07586_, _07550_);
  and _15885_ (_07588_, _07524_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15886_ (_07589_, _07588_);
  nand _15887_ (_07590_, _07515_, _06673_);
  nor _15888_ (_07591_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not _15889_ (_07593_, _07591_);
  and _15890_ (_07594_, _07593_, _07590_);
  nand _15891_ (_07595_, _07594_, _07589_);
  or _15892_ (_07596_, _07594_, _07589_);
  nand _15893_ (_07597_, _07596_, _07595_);
  and _15894_ (_07598_, _07541_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15895_ (_07600_, _07598_);
  or _15896_ (_07601_, _07555_, _06700_);
  nor _15897_ (_07602_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not _15898_ (_07603_, _07602_);
  and _15899_ (_07604_, _07603_, _07601_);
  nand _15900_ (_07605_, _07604_, _07600_);
  and _15901_ (_07606_, _07560_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not _15902_ (_07607_, _07606_);
  nand _15903_ (_07608_, _07515_, _06728_);
  nor _15904_ (_07609_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not _15905_ (_07610_, _07609_);
  and _15906_ (_07611_, _07610_, _07608_);
  nor _15907_ (_07612_, _07611_, _07607_);
  or _15908_ (_07613_, _07604_, _07600_);
  nand _15909_ (_07614_, _07613_, _07605_);
  or _15910_ (_07615_, _07614_, _07612_);
  and _15911_ (_07617_, _07615_, _07605_);
  or _15912_ (_07618_, _07617_, _07597_);
  nand _15913_ (_07619_, _07618_, _07595_);
  nor _15914_ (_07621_, _07576_, _07572_);
  nor _15915_ (_07622_, _07621_, _07577_);
  and _15916_ (_07623_, _07582_, _07622_);
  and _15917_ (_07624_, _07623_, _07554_);
  nand _15918_ (_07625_, _07624_, _07619_);
  nand _15919_ (_07626_, _07625_, _07587_);
  nor _15920_ (_07627_, _07570_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and _15921_ (_07628_, _06622_, _07522_);
  and _15922_ (_07629_, _06597_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _15923_ (_07630_, _07629_, _07628_);
  nor _15924_ (_07631_, _07630_, _07526_);
  nor _15925_ (_07632_, _07631_, _07627_);
  not _15926_ (_07633_, _07632_);
  and _15927_ (_07634_, _06816_, _06597_);
  nor _15928_ (_07636_, _07634_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor _15929_ (_07637_, _07545_, _07529_);
  nor _15930_ (_07638_, _07630_, _07564_);
  and _15931_ (_07639_, _07638_, _07637_);
  nor _15932_ (_07640_, _07639_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor _15933_ (_07641_, _07640_, _07636_);
  and _15934_ (_07642_, _07641_, _07633_);
  and _15935_ (_07643_, _07642_, _07626_);
  and _15936_ (_07644_, _07643_, _07024_);
  nor _15937_ (_07645_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not _15938_ (_07646_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _15939_ (_07647_, _07646_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _15940_ (_07648_, _07647_, _07645_);
  not _15941_ (_07649_, _07648_);
  nor _15942_ (_07650_, _07649_, _06839_);
  nor _15943_ (_07651_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not _15944_ (_07652_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _15945_ (_07653_, _07652_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _15946_ (_07654_, _07653_, _07651_);
  nor _15947_ (_07655_, _07654_, _07650_);
  not _15948_ (_07656_, _07655_);
  and _15949_ (_07657_, _07654_, _07650_);
  nor _15950_ (_07658_, _07657_, _06549_);
  and _15951_ (_07659_, _07658_, _07656_);
  nor _15952_ (_07660_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  nand _15953_ (_07661_, _07660_, _06597_);
  not _15954_ (_07662_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  or _15955_ (_07663_, _07662_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  or _15956_ (_07664_, _07663_, _06622_);
  not _15957_ (_07665_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  or _15958_ (_07666_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _07665_);
  or _15959_ (_07667_, _07666_, _06680_);
  and _15960_ (_07668_, _07667_, _07664_);
  and _15961_ (_07669_, _07666_, _07663_);
  or _15962_ (_07670_, _06734_, _07665_);
  nand _15963_ (_07671_, _07670_, _07669_);
  nand _15964_ (_07672_, _07671_, _07668_);
  and _15965_ (_07674_, _07672_, _07661_);
  and _15966_ (_07675_, _07674_, _06909_);
  nand _15967_ (_07676_, _07660_, _06816_);
  or _15968_ (_07677_, _07663_, _06652_);
  or _15969_ (_07678_, _07666_, _06871_);
  and _15970_ (_07679_, _07678_, _07677_);
  or _15971_ (_07680_, _06760_, _07665_);
  nand _15972_ (_07681_, _07680_, _07669_);
  nand _15973_ (_07682_, _07681_, _07679_);
  and _15974_ (_07683_, _07682_, _07676_);
  and _15975_ (_07684_, _07683_, _06924_);
  and _15976_ (_07685_, _07684_, _07675_);
  and _15977_ (_07686_, _07674_, _06924_);
  not _15978_ (_07687_, _07686_);
  nand _15979_ (_07688_, _07682_, _07676_);
  or _15980_ (_07689_, _07688_, _06728_);
  and _15981_ (_07690_, _07689_, _07687_);
  nor _15982_ (_07691_, _07690_, _07685_);
  and _15983_ (_07692_, _07691_, _07027_);
  or _15984_ (_07693_, _07692_, _07659_);
  or _15985_ (_07694_, _07693_, _07644_);
  or _15986_ (_07695_, _07694_, _07514_);
  nor _15987_ (_07696_, _07695_, _07498_);
  not _15988_ (_07697_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and _15989_ (_07698_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _06406_);
  and _15990_ (_07699_, _07698_, _07697_);
  not _15991_ (_07700_, _07699_);
  nor _15992_ (_07701_, _07700_, _07696_);
  not _15993_ (_07702_, _07701_);
  not _15994_ (_07703_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _15995_ (_07704_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _06406_);
  and _15996_ (_07705_, _07704_, _07703_);
  nor _15997_ (_07706_, _06477_, _07084_);
  and _15998_ (_07707_, _07706_, _06976_);
  and _15999_ (_07708_, _07707_, _07125_);
  and _16000_ (_07709_, _07708_, _06983_);
  nor _16001_ (_07710_, _07709_, _07705_);
  nand _16002_ (_07711_, _07642_, _07626_);
  not _16003_ (_07712_, _07553_);
  and _16004_ (_07713_, _07622_, _07619_);
  nor _16005_ (_07714_, _07713_, _07577_);
  nor _16006_ (_07715_, _07714_, _07579_);
  nor _16007_ (_07716_, _07715_, _07567_);
  nor _16008_ (_07717_, _07716_, _07712_);
  and _16009_ (_07718_, _07716_, _07712_);
  nor _16010_ (_07719_, _07718_, _07717_);
  nor _16011_ (_07720_, _07719_, _07711_);
  and _16012_ (_07721_, _07711_, _07540_);
  nor _16013_ (_07722_, _07721_, _07720_);
  and _16014_ (_07723_, _07722_, _07533_);
  nor _16015_ (_07724_, _07722_, _07533_);
  nor _16016_ (_07725_, _07724_, _07723_);
  not _16017_ (_07726_, _07547_);
  and _16018_ (_07727_, _07580_, _07714_);
  nor _16019_ (_07728_, _07580_, _07714_);
  nor _16020_ (_07729_, _07728_, _07727_);
  nor _16021_ (_07730_, _07729_, _07711_);
  and _16022_ (_07731_, _07711_, _07559_);
  nor _16023_ (_07732_, _07731_, _07730_);
  and _16024_ (_07733_, _07732_, _07726_);
  nand _16025_ (_07734_, _07565_, _07561_);
  nor _16026_ (_07735_, _07622_, _07619_);
  or _16027_ (_07736_, _07735_, _07713_);
  and _16028_ (_07737_, _07736_, _07643_);
  nor _16029_ (_07738_, _07643_, _07576_);
  nor _16030_ (_07739_, _07738_, _07737_);
  and _16031_ (_07740_, _07739_, _07734_);
  not _16032_ (_07741_, _07740_);
  nor _16033_ (_07742_, _07732_, _07726_);
  or _16034_ (_07743_, _07733_, _07742_);
  nor _16035_ (_07744_, _07743_, _07741_);
  nor _16036_ (_07745_, _07744_, _07733_);
  not _16037_ (_07746_, _07745_);
  and _16038_ (_07747_, _07617_, _07597_);
  not _16039_ (_07748_, _07747_);
  and _16040_ (_07749_, _07748_, _07618_);
  nor _16041_ (_07750_, _07749_, _07711_);
  nor _16042_ (_07751_, _07643_, _07594_);
  nor _16043_ (_07752_, _07751_, _07750_);
  nor _16044_ (_07753_, _07752_, _07572_);
  not _16045_ (_07754_, _07753_);
  not _16046_ (_07755_, _07611_);
  or _16047_ (_07756_, _07711_, _07607_);
  nand _16048_ (_07757_, _07756_, _07755_);
  or _16049_ (_07758_, _07756_, _07755_);
  and _16050_ (_07759_, _07758_, _07757_);
  nand _16051_ (_07760_, _07759_, _07600_);
  or _16052_ (_07761_, _07759_, _07600_);
  and _16053_ (_07762_, _07761_, _07760_);
  and _16054_ (_07763_, _07515_, _06754_);
  nor _16055_ (_07765_, _07515_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  nor _16056_ (_07766_, _07765_, _07763_);
  nor _16057_ (_07768_, _07766_, _07607_);
  not _16058_ (_07769_, _07768_);
  nand _16059_ (_07770_, _07769_, _07762_);
  and _16060_ (_07771_, _07770_, _07760_);
  and _16061_ (_07772_, _07614_, _07612_);
  not _16062_ (_07774_, _07772_);
  and _16063_ (_07775_, _07774_, _07615_);
  or _16064_ (_07776_, _07775_, _07711_);
  or _16065_ (_07777_, _07643_, _07604_);
  and _16066_ (_07778_, _07777_, _07776_);
  and _16067_ (_07779_, _07778_, _07589_);
  nor _16068_ (_07780_, _07778_, _07589_);
  or _16069_ (_07781_, _07780_, _07779_);
  or _16070_ (_07782_, _07781_, _07771_);
  and _16071_ (_07783_, _07752_, _07572_);
  nor _16072_ (_07784_, _07783_, _07779_);
  nand _16073_ (_07786_, _07784_, _07782_);
  and _16074_ (_07787_, _07786_, _07754_);
  nor _16075_ (_07788_, _07739_, _07734_);
  nor _16076_ (_07789_, _07788_, _07740_);
  not _16077_ (_07790_, _07743_);
  and _16078_ (_07791_, _07790_, _07789_);
  and _16079_ (_07792_, _07791_, _07787_);
  or _16080_ (_07793_, _07792_, _07746_);
  and _16081_ (_07794_, _07793_, _07725_);
  and _16082_ (_07795_, _07711_, _07519_);
  not _16083_ (_07796_, _07717_);
  and _16084_ (_07797_, _07796_, _07548_);
  and _16085_ (_07798_, _07797_, _07551_);
  nor _16086_ (_07799_, _07797_, _07551_);
  or _16087_ (_07800_, _07799_, _07798_);
  and _16088_ (_07801_, _07800_, _07643_);
  or _16089_ (_07802_, _07801_, _07795_);
  and _16090_ (_07803_, _07802_, _07633_);
  or _16091_ (_07804_, _07803_, _07723_);
  or _16092_ (_07805_, _07804_, _07794_);
  not _16093_ (_07807_, _07641_);
  nor _16094_ (_07808_, _07802_, _07633_);
  nor _16095_ (_07809_, _07808_, _07807_);
  nand _16096_ (_07810_, _07809_, _07805_);
  or _16097_ (_07811_, _07769_, _07762_);
  and _16098_ (_07812_, _07811_, _07770_);
  or _16099_ (_07813_, _07812_, _07810_);
  and _16100_ (_07814_, _07809_, _07805_);
  or _16101_ (_07815_, _07814_, _07759_);
  and _16102_ (_07816_, _07815_, _07813_);
  nand _16103_ (_07817_, _07816_, _07024_);
  not _16104_ (_07818_, _07660_);
  and _16105_ (_07819_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and _16106_ (_07821_, _07674_, _06905_);
  and _16107_ (_07822_, _07683_, _07003_);
  and _16108_ (_07823_, _07822_, _07821_);
  and _16109_ (_07824_, _07683_, _06905_);
  and _16110_ (_07825_, _07674_, _06616_);
  nand _16111_ (_07826_, _07825_, _07824_);
  and _16112_ (_07827_, _07683_, _06616_);
  or _16113_ (_07828_, _07827_, _07821_);
  and _16114_ (_07830_, _07828_, _07826_);
  and _16115_ (_07831_, _07830_, _07823_);
  or _16116_ (_07832_, _07826_, _06810_);
  and _16117_ (_07833_, _07683_, _06902_);
  not _16118_ (_07835_, _07833_);
  nand _16119_ (_07836_, _07835_, _07826_);
  and _16120_ (_07837_, _07836_, _07832_);
  nand _16121_ (_07838_, _07837_, _07825_);
  or _16122_ (_07839_, _07833_, _07825_);
  and _16123_ (_07840_, _07839_, _07838_);
  nand _16124_ (_07841_, _07840_, _07831_);
  not _16125_ (_07842_, _07841_);
  not _16126_ (_07843_, _07832_);
  or _16127_ (_07844_, _07688_, _06586_);
  nand _16128_ (_07845_, _07672_, _07661_);
  or _16129_ (_07846_, _07845_, _06810_);
  or _16130_ (_07847_, _07846_, _07844_);
  nand _16131_ (_07848_, _07846_, _07844_);
  and _16132_ (_07849_, _07848_, _07847_);
  and _16133_ (_07850_, _07849_, _07843_);
  not _16134_ (_07851_, _07850_);
  and _16135_ (_07852_, _07837_, _07825_);
  nand _16136_ (_07853_, _07849_, _07852_);
  or _16137_ (_07854_, _07849_, _07852_);
  nand _16138_ (_07855_, _07854_, _07853_);
  nand _16139_ (_07856_, _07855_, _07832_);
  and _16140_ (_07857_, _07856_, _07851_);
  nand _16141_ (_07858_, _07857_, _07842_);
  or _16142_ (_07859_, _07857_, _07842_);
  nand _16143_ (_07860_, _07859_, _07858_);
  not _16144_ (_07861_, _07860_);
  and _16145_ (_07862_, _07683_, _06700_);
  nand _16146_ (_07863_, _07862_, _07675_);
  and _16147_ (_07864_, _07674_, _06700_);
  and _16148_ (_07865_, _07864_, _07689_);
  nand _16149_ (_07866_, _07865_, _07822_);
  nand _16150_ (_07867_, _07866_, _07863_);
  not _16151_ (_07868_, _07823_);
  and _16152_ (_07870_, _07674_, _07003_);
  or _16153_ (_07871_, _07870_, _07824_);
  and _16154_ (_07872_, _07871_, _07868_);
  nand _16155_ (_07873_, _07872_, _07867_);
  not _16156_ (_07874_, _07873_);
  not _16157_ (_07875_, _07831_);
  or _16158_ (_07876_, _07830_, _07823_);
  and _16159_ (_07877_, _07876_, _07875_);
  and _16160_ (_07878_, _07877_, _07874_);
  or _16161_ (_07879_, _07840_, _07831_);
  and _16162_ (_07880_, _07879_, _07841_);
  nand _16163_ (_07881_, _07880_, _07878_);
  or _16164_ (_07882_, _07862_, _07675_);
  and _16165_ (_07883_, _07882_, _07863_);
  and _16166_ (_07884_, _07883_, _07685_);
  or _16167_ (_07885_, _07865_, _07822_);
  and _16168_ (_07886_, _07885_, _07866_);
  nand _16169_ (_07887_, _07886_, _07884_);
  not _16170_ (_07888_, _07887_);
  or _16171_ (_07889_, _07872_, _07867_);
  and _16172_ (_07890_, _07889_, _07873_);
  nand _16173_ (_07891_, _07890_, _07888_);
  not _16174_ (_07892_, _07891_);
  nand _16175_ (_07893_, _07877_, _07874_);
  or _16176_ (_07894_, _07877_, _07874_);
  and _16177_ (_07895_, _07894_, _07893_);
  nand _16178_ (_07896_, _07895_, _07892_);
  not _16179_ (_07897_, _07896_);
  or _16180_ (_07898_, _07880_, _07878_);
  and _16181_ (_07899_, _07898_, _07881_);
  nand _16182_ (_07900_, _07899_, _07897_);
  nand _16183_ (_07901_, _07900_, _07881_);
  nand _16184_ (_07902_, _07901_, _07861_);
  nand _16185_ (_07903_, _07902_, _07858_);
  and _16186_ (_07904_, _07674_, _06957_);
  and _16187_ (_07905_, _07904_, _07835_);
  not _16188_ (_07906_, _07905_);
  and _16189_ (_07907_, _07851_, _07853_);
  nor _16190_ (_07908_, _07907_, _07906_);
  and _16191_ (_07909_, _07907_, _07906_);
  nor _16192_ (_07910_, _07909_, _07908_);
  nand _16193_ (_07911_, _07910_, _07903_);
  or _16194_ (_07912_, _07910_, _07903_);
  and _16195_ (_07913_, _07912_, _07911_);
  nand _16196_ (_07914_, _07913_, _07819_);
  and _16197_ (_07915_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  or _16198_ (_07916_, _07901_, _07861_);
  and _16199_ (_07917_, _07916_, _07902_);
  nand _16200_ (_07918_, _07917_, _07915_);
  or _16201_ (_07919_, _07917_, _07915_);
  nand _16202_ (_07920_, _07919_, _07918_);
  and _16203_ (_07921_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or _16204_ (_07922_, _07899_, _07897_);
  and _16205_ (_07923_, _07922_, _07900_);
  nand _16206_ (_07924_, _07923_, _07921_);
  or _16207_ (_07925_, _07923_, _07921_);
  nand _16208_ (_07926_, _07925_, _07924_);
  and _16209_ (_07927_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  or _16210_ (_07928_, _07895_, _07892_);
  and _16211_ (_07929_, _07928_, _07896_);
  nand _16212_ (_07930_, _07929_, _07927_);
  or _16213_ (_07931_, _07929_, _07927_);
  nand _16214_ (_07932_, _07931_, _07930_);
  and _16215_ (_07934_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or _16216_ (_07935_, _07890_, _07888_);
  and _16217_ (_07936_, _07935_, _07891_);
  nand _16218_ (_07937_, _07936_, _07934_);
  and _16219_ (_07938_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or _16220_ (_07939_, _07886_, _07884_);
  and _16221_ (_07940_, _07939_, _07887_);
  nand _16222_ (_07941_, _07940_, _07938_);
  and _16223_ (_07942_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  not _16224_ (_07943_, _07942_);
  nor _16225_ (_07944_, _07883_, _07685_);
  or _16226_ (_07945_, _07944_, _07884_);
  or _16227_ (_07946_, _07945_, _07943_);
  or _16228_ (_07947_, _07940_, _07938_);
  nand _16229_ (_07948_, _07947_, _07941_);
  or _16230_ (_07949_, _07948_, _07946_);
  and _16231_ (_07950_, _07949_, _07941_);
  or _16232_ (_07951_, _07936_, _07934_);
  nand _16233_ (_07952_, _07951_, _07937_);
  or _16234_ (_07953_, _07952_, _07950_);
  and _16235_ (_07954_, _07953_, _07937_);
  or _16236_ (_07955_, _07954_, _07932_);
  and _16237_ (_07956_, _07955_, _07930_);
  or _16238_ (_07957_, _07956_, _07926_);
  and _16239_ (_07958_, _07957_, _07924_);
  or _16240_ (_07960_, _07958_, _07920_);
  and _16241_ (_07961_, _07960_, _07918_);
  or _16242_ (_07962_, _07913_, _07819_);
  nand _16243_ (_07963_, _07962_, _07914_);
  or _16244_ (_07964_, _07963_, _07961_);
  and _16245_ (_07965_, _07964_, _07914_);
  and _16246_ (_07966_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  not _16247_ (_07967_, _07908_);
  and _16248_ (_07968_, _07967_, _07847_);
  nand _16249_ (_07970_, _07968_, _07911_);
  nand _16250_ (_07971_, _07970_, _07966_);
  or _16251_ (_07972_, _07970_, _07966_);
  nand _16252_ (_07974_, _07972_, _07971_);
  or _16253_ (_07975_, _07974_, _07965_);
  nand _16254_ (_07977_, _07974_, _07965_);
  and _16255_ (_07978_, _07977_, _07975_);
  nand _16256_ (_07979_, _07978_, _07027_);
  nor _16257_ (_07981_, _06884_, _06882_);
  nor _16258_ (_07982_, _07981_, _06885_);
  nor _16259_ (_07983_, _07982_, _06846_);
  not _16260_ (_07984_, _07983_);
  nor _16261_ (_07985_, _06911_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and _16262_ (_07986_, _07985_, _06909_);
  nor _16263_ (_07987_, _07985_, _06909_);
  nor _16264_ (_07988_, _07987_, _07986_);
  nor _16265_ (_07990_, _07988_, _06918_);
  and _16266_ (_07991_, _06942_, _06764_);
  nor _16267_ (_07993_, _07017_, _06763_);
  not _16268_ (_07994_, _07993_);
  and _16269_ (_07995_, _06933_, _06736_);
  and _16270_ (_07996_, _06954_, _06728_);
  nor _16271_ (_07998_, _07996_, _07995_);
  nand _16272_ (_07999_, _07998_, _07994_);
  nor _16273_ (_08000_, _07999_, _07991_);
  not _16274_ (_08001_, _07032_);
  nor _16275_ (_08002_, _08001_, _06754_);
  not _16276_ (_08003_, _08002_);
  and _16277_ (_08004_, _06951_, _06909_);
  and _16278_ (_08005_, _07030_, _06700_);
  nor _16279_ (_08006_, _08005_, _08004_);
  and _16280_ (_08007_, _08006_, _08003_);
  and _16281_ (_08008_, _08007_, _08000_);
  not _16282_ (_08009_, _08008_);
  nor _16283_ (_08010_, _08009_, _07990_);
  and _16284_ (_08011_, _06991_, _06734_);
  and _16285_ (_08012_, _06754_, _06728_);
  nor _16286_ (_08013_, _08012_, _07004_);
  nor _16287_ (_08014_, _08013_, _06778_);
  and _16288_ (_08015_, _08013_, _06778_);
  nor _16289_ (_08016_, _08015_, _08014_);
  and _16290_ (_08017_, _08016_, _06997_);
  nor _16291_ (_08018_, _08017_, _08011_);
  not _16292_ (_08019_, _08018_);
  nor _16293_ (_08020_, _06764_, _06762_);
  or _16294_ (_08021_, _08020_, _06765_);
  and _16295_ (_08022_, _08021_, _06781_);
  nor _16296_ (_08023_, _08021_, _06781_);
  or _16297_ (_08024_, _08023_, _08022_);
  and _16298_ (_08025_, _08024_, _06548_);
  nor _16299_ (_08026_, _08025_, _08019_);
  and _16300_ (_08027_, _08026_, _08010_);
  and _16301_ (_08028_, _08027_, _07984_);
  and _16302_ (_08029_, _08028_, _07979_);
  nand _16303_ (_08030_, _08029_, _07817_);
  or _16304_ (_08031_, _08030_, _07710_);
  not _16305_ (_08032_, _07089_);
  nor _16306_ (_08033_, _06968_, _08032_);
  nor _16307_ (_08034_, _07089_, _06731_);
  nor _16308_ (_08035_, _08034_, _08033_);
  nor _16309_ (_08036_, _06499_, _06448_);
  and _16310_ (_08037_, _08036_, _06434_);
  nor _16311_ (_08038_, _06477_, _06463_);
  and _16312_ (_08039_, _08038_, _06485_);
  and _16313_ (_08040_, _08039_, _08037_);
  and _16314_ (_08041_, _07710_, _07700_);
  and _16315_ (_08042_, _08041_, _08040_);
  not _16316_ (_08043_, _08042_);
  nor _16317_ (_08044_, _08043_, _08035_);
  not _16318_ (_08045_, _07710_);
  nor _16319_ (_08046_, _08040_, _06731_);
  nor _16320_ (_08047_, _08046_, _08045_);
  not _16321_ (_08048_, _08047_);
  nor _16322_ (_08049_, _08048_, _08044_);
  nor _16323_ (_08050_, _08049_, _07699_);
  nand _16324_ (_08051_, _08050_, _08031_);
  nand _16325_ (_08052_, _08051_, _07702_);
  and _16326_ (_06536_, _08052_, _06989_);
  and _16327_ (_08053_, _06951_, _06760_);
  and _16328_ (_08055_, _06958_, _06905_);
  nor _16329_ (_08056_, _06990_, _06919_);
  not _16330_ (_08057_, _08056_);
  nor _16331_ (_08058_, _08057_, _07011_);
  nor _16332_ (_08059_, _08058_, _06760_);
  and _16333_ (_08060_, _08058_, _06760_);
  nor _16334_ (_08061_, _08060_, _08059_);
  and _16335_ (_08062_, _08061_, _06997_);
  nor _16336_ (_08063_, _06992_, _06754_);
  or _16337_ (_08064_, _08063_, _08062_);
  or _16338_ (_08065_, _08064_, _08055_);
  and _16339_ (_08066_, _07814_, _07024_);
  and _16340_ (_08067_, _07649_, _06839_);
  nor _16341_ (_08068_, _08067_, _07650_);
  and _16342_ (_08069_, _08068_, _06548_);
  and _16343_ (_08070_, _07684_, _07027_);
  or _16344_ (_08071_, _08070_, _08069_);
  or _16345_ (_08072_, _08071_, _08066_);
  or _16346_ (_08074_, _08072_, _08065_);
  or _16347_ (_08075_, _08074_, _08053_);
  nand _16348_ (_08076_, _08075_, _07699_);
  nand _16349_ (_08077_, _07814_, _07606_);
  and _16350_ (_08078_, _08077_, _07766_);
  nor _16351_ (_08079_, _08077_, _07766_);
  or _16352_ (_08080_, _08079_, _08078_);
  nand _16353_ (_08082_, _08080_, _07024_);
  not _16354_ (_08083_, _07964_);
  and _16355_ (_08084_, _07963_, _07961_);
  nor _16356_ (_08085_, _08084_, _08083_);
  and _16357_ (_08086_, _08085_, _07027_);
  nor _16358_ (_08087_, _06780_, _06778_);
  nor _16359_ (_08089_, _08087_, _06781_);
  nor _16360_ (_08090_, _06845_, _06548_);
  not _16361_ (_08091_, _08090_);
  and _16362_ (_08092_, _08091_, _08089_);
  not _16363_ (_08093_, _08092_);
  nor _16364_ (_08095_, _06943_, _06762_);
  nor _16365_ (_08096_, _08095_, _06940_);
  or _16366_ (_08098_, _08096_, _06779_);
  and _16367_ (_08099_, _06997_, _06754_);
  and _16368_ (_08101_, _06991_, _06760_);
  nor _16369_ (_08102_, _08101_, _08099_);
  and _16370_ (_08103_, _06933_, _06762_);
  and _16371_ (_08104_, _06954_, _06754_);
  nor _16372_ (_08106_, _08104_, _08103_);
  and _16373_ (_08107_, _08106_, _08102_);
  and _16374_ (_08109_, _06958_, _06778_);
  nor _16375_ (_08110_, _06951_, _06908_);
  nor _16376_ (_08112_, _08110_, _06754_);
  nor _16377_ (_08113_, _08112_, _08109_);
  and _16378_ (_08114_, _06931_, _06957_);
  nor _16379_ (_08115_, _07031_, _06728_);
  nor _16380_ (_08116_, _08115_, _08114_);
  and _16381_ (_08117_, _08116_, _08113_);
  and _16382_ (_08118_, _08117_, _08107_);
  and _16383_ (_08119_, _08118_, _08098_);
  and _16384_ (_08120_, _08119_, _08093_);
  not _16385_ (_08121_, _08120_);
  nor _16386_ (_08122_, _08121_, _08086_);
  nand _16387_ (_08123_, _08122_, _08082_);
  or _16388_ (_08124_, _08123_, _07710_);
  not _16389_ (_08125_, _08040_);
  not _16390_ (_08126_, _06968_);
  and _16391_ (_08127_, _08126_, _06979_);
  nor _16392_ (_08128_, _06979_, _06757_);
  nor _16393_ (_08129_, _08128_, _08127_);
  nor _16394_ (_08130_, _08129_, _08125_);
  nor _16395_ (_08131_, _08040_, _06757_);
  nor _16396_ (_08132_, _08131_, _08045_);
  not _16397_ (_08133_, _08132_);
  nor _16398_ (_08134_, _08133_, _08130_);
  nor _16399_ (_08136_, _08134_, _07699_);
  nand _16400_ (_08137_, _08136_, _08124_);
  nand _16401_ (_08138_, _08137_, _08076_);
  and _16402_ (_06542_, _08138_, _06989_);
  and _16403_ (_08139_, _07326_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and _16404_ (_08140_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not _16405_ (_08141_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _16406_ (_08142_, _08139_, _08141_);
  or _16407_ (_08143_, _08142_, _08140_);
  and _16408_ (_06580_, _08143_, _06989_);
  and _16409_ (_08144_, _06951_, _06623_);
  and _16410_ (_08145_, _06958_, _06909_);
  and _16411_ (_08146_, _07505_, _06734_);
  and _16412_ (_08147_, _08146_, _06706_);
  and _16413_ (_08148_, _08147_, _06889_);
  nor _16414_ (_08149_, _08148_, _06778_);
  nor _16415_ (_08150_, _06760_, _06734_);
  and _16416_ (_08151_, _06871_, _06680_);
  and _16417_ (_08152_, _08151_, _08150_);
  and _16418_ (_08153_, _08152_, _07500_);
  and _16419_ (_08154_, _08153_, _06652_);
  nor _16420_ (_08155_, _08154_, _06883_);
  nor _16421_ (_08156_, _06778_, _06853_);
  or _16422_ (_08157_, _08156_, _08155_);
  nor _16423_ (_08158_, _08157_, _08149_);
  and _16424_ (_08159_, _08158_, _06622_);
  nor _16425_ (_08160_, _08158_, _06622_);
  nor _16426_ (_08161_, _08160_, _08159_);
  nor _16427_ (_08162_, _08161_, _07101_);
  nor _16428_ (_08163_, _06778_, _06622_);
  and _16429_ (_08164_, _06778_, _06616_);
  or _16430_ (_08165_, _08164_, _08163_);
  and _16431_ (_08166_, _08165_, _06991_);
  or _16432_ (_08167_, _08166_, _08162_);
  or _16433_ (_08168_, _08167_, _08145_);
  and _16434_ (_08169_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _16435_ (_08170_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not _16436_ (_08171_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _16437_ (_08172_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08171_);
  nor _16438_ (_08173_, _08172_, _08170_);
  nor _16439_ (_08174_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not _16440_ (_08175_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _16441_ (_08176_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08175_);
  nor _16442_ (_08177_, _08176_, _08174_);
  and _16443_ (_08178_, _08177_, _07657_);
  and _16444_ (_08179_, _08178_, _08173_);
  nor _16445_ (_08180_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not _16446_ (_08182_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _16447_ (_08183_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08182_);
  nor _16448_ (_08184_, _08183_, _08180_);
  and _16449_ (_08185_, _08184_, _08179_);
  nor _16450_ (_08186_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not _16451_ (_08187_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _16452_ (_08188_, _08187_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _16453_ (_08189_, _08188_, _08186_);
  nor _16454_ (_08190_, _08189_, _08185_);
  and _16455_ (_08191_, _08189_, _08185_);
  nor _16456_ (_08192_, _08191_, _08190_);
  and _16457_ (_08193_, _08192_, _06548_);
  and _16458_ (_08195_, _07954_, _07932_);
  not _16459_ (_08196_, _08195_);
  and _16460_ (_08197_, _08196_, _07955_);
  and _16461_ (_08198_, _08197_, _07027_);
  or _16462_ (_08199_, _08198_, _08193_);
  or _16463_ (_08200_, _08199_, _08169_);
  or _16464_ (_08201_, _08200_, _08168_);
  nor _16465_ (_08202_, _08201_, _08144_);
  nor _16466_ (_08203_, _08202_, _07700_);
  not _16467_ (_08204_, _08203_);
  nand _16468_ (_08205_, _07810_, _07732_);
  nand _16469_ (_08206_, _07789_, _07787_);
  and _16470_ (_08207_, _08206_, _07741_);
  nand _16471_ (_08208_, _08207_, _07790_);
  or _16472_ (_08209_, _08207_, _07790_);
  nand _16473_ (_08210_, _08209_, _08208_);
  nand _16474_ (_08211_, _08210_, _07814_);
  nand _16475_ (_08212_, _08211_, _08205_);
  nand _16476_ (_08213_, _08212_, _07024_);
  or _16477_ (_08214_, _07974_, _07914_);
  nand _16478_ (_08215_, _08214_, _07971_);
  and _16479_ (_08216_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and _16480_ (_08218_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and _16481_ (_08219_, _08218_, _08216_);
  and _16482_ (_08220_, _08219_, _08215_);
  nor _16483_ (_08221_, _07974_, _07963_);
  nand _16484_ (_08222_, _08219_, _08221_);
  nor _16485_ (_08223_, _08222_, _07961_);
  or _16486_ (_08224_, _08223_, _08220_);
  and _16487_ (_08225_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and _16488_ (_08226_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and _16489_ (_08227_, _08226_, _08225_);
  nand _16490_ (_08228_, _08227_, _08224_);
  and _16491_ (_08229_, _08224_, _08225_);
  or _16492_ (_08230_, _08226_, _08229_);
  and _16493_ (_08231_, _08230_, _08228_);
  nand _16494_ (_08232_, _08231_, _07027_);
  nor _16495_ (_08233_, _06895_, _06864_);
  nor _16496_ (_08234_, _08233_, _06896_);
  nor _16497_ (_08235_, _08234_, _06846_);
  not _16498_ (_08236_, _08235_);
  nor _16499_ (_08237_, _06653_, _06627_);
  nor _16500_ (_08238_, _08237_, _06821_);
  nor _16501_ (_08239_, _08238_, _06791_);
  not _16502_ (_08240_, _08239_);
  nor _16503_ (_08241_, _06792_, _06549_);
  and _16504_ (_08242_, _08241_, _08240_);
  nor _16505_ (_08243_, _06903_, _06586_);
  nor _16506_ (_08244_, _08243_, _06778_);
  and _16507_ (_08245_, _08244_, _06938_);
  nor _16508_ (_08246_, _08245_, _06913_);
  and _16509_ (_08247_, _08246_, _07096_);
  nor _16510_ (_08248_, _08246_, _07096_);
  nor _16511_ (_08249_, _08248_, _08247_);
  nor _16512_ (_08251_, _08249_, _06918_);
  nor _16513_ (_08252_, _07031_, _06810_);
  not _16514_ (_08253_, _08252_);
  and _16515_ (_08254_, _06951_, _06616_);
  not _16516_ (_08255_, _08254_);
  or _16517_ (_08256_, _08001_, _06646_);
  and _16518_ (_08257_, _08256_, _08255_);
  and _16519_ (_08258_, _08257_, _08253_);
  and _16520_ (_08259_, _08258_, _07116_);
  not _16521_ (_08260_, _08259_);
  nor _16522_ (_08261_, _08260_, _08251_);
  and _16523_ (_08262_, _08261_, _07105_);
  not _16524_ (_08263_, _08262_);
  nor _16525_ (_08264_, _08263_, _08242_);
  and _16526_ (_08265_, _08264_, _08236_);
  and _16527_ (_08267_, _08265_, _08232_);
  nand _16528_ (_08268_, _08267_, _08213_);
  or _16529_ (_08269_, _08268_, _07710_);
  nor _16530_ (_08270_, _08040_, _06619_);
  nor _16531_ (_08271_, _08270_, _08045_);
  and _16532_ (_08272_, _06968_, _07048_);
  or _16533_ (_08273_, _07048_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand _16534_ (_08274_, _08273_, _08040_);
  or _16535_ (_08275_, _08274_, _08272_);
  and _16536_ (_08276_, _08275_, _08271_);
  nor _16537_ (_08277_, _08276_, _07699_);
  nand _16538_ (_08278_, _08277_, _08269_);
  nand _16539_ (_08279_, _08278_, _08204_);
  and _16540_ (_06626_, _08279_, _06989_);
  and _16541_ (_08280_, _06951_, _06853_);
  and _16542_ (_08281_, _06958_, _06924_);
  nor _16543_ (_08282_, _08153_, _06883_);
  nor _16544_ (_08283_, _08282_, _08149_);
  nor _16545_ (_08284_, _08283_, _06853_);
  and _16546_ (_08285_, _08283_, _06853_);
  nor _16547_ (_08286_, _08285_, _08284_);
  and _16548_ (_08287_, _08286_, _06997_);
  and _16549_ (_08288_, _06778_, _06646_);
  nor _16550_ (_08289_, _08156_, _06992_);
  not _16551_ (_08290_, _08289_);
  nor _16552_ (_08291_, _08290_, _08288_);
  or _16553_ (_08292_, _08291_, _08287_);
  or _16554_ (_08293_, _08292_, _08281_);
  and _16555_ (_08294_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  nor _16556_ (_08295_, _08184_, _08179_);
  not _16557_ (_08296_, _08295_);
  nor _16558_ (_08298_, _08185_, _06549_);
  and _16559_ (_08299_, _08298_, _08296_);
  and _16560_ (_08300_, _07952_, _07950_);
  not _16561_ (_08301_, _08300_);
  and _16562_ (_08302_, _08301_, _07953_);
  and _16563_ (_08303_, _08302_, _07027_);
  or _16564_ (_08304_, _08303_, _08299_);
  or _16565_ (_08305_, _08304_, _08294_);
  or _16566_ (_08306_, _08305_, _08293_);
  nor _16567_ (_08307_, _08306_, _08280_);
  nor _16568_ (_08308_, _08307_, _07700_);
  not _16569_ (_08309_, _08308_);
  or _16570_ (_08310_, _07789_, _07787_);
  and _16571_ (_08311_, _08310_, _08206_);
  and _16572_ (_08312_, _08311_, _07814_);
  and _16573_ (_08313_, _07810_, _07739_);
  or _16574_ (_08314_, _08313_, _08312_);
  nand _16575_ (_08315_, _08314_, _07024_);
  nor _16576_ (_08316_, _08224_, _08225_);
  nor _16577_ (_08317_, _08316_, _08229_);
  nand _16578_ (_08318_, _08317_, _07027_);
  nor _16579_ (_08319_, _06894_, _06655_);
  and _16580_ (_08320_, _06894_, _06655_);
  nor _16581_ (_08322_, _08320_, _08319_);
  and _16582_ (_08323_, _08322_, _06845_);
  not _16583_ (_08324_, _08323_);
  nor _16584_ (_08325_, _06790_, _06655_);
  nor _16585_ (_08326_, _08325_, _06791_);
  and _16586_ (_08327_, _08326_, _06548_);
  nor _16587_ (_08328_, _06912_, _06905_);
  or _16588_ (_08329_, _08328_, _06918_);
  nor _16589_ (_08331_, _08329_, _06913_);
  not _16590_ (_08332_, _08331_);
  or _16591_ (_08333_, _08001_, _06673_);
  nand _16592_ (_08334_, _07030_, _06616_);
  not _16593_ (_08335_, _08334_);
  and _16594_ (_08336_, _06951_, _06905_);
  nor _16595_ (_08337_, _08336_, _08335_);
  and _16596_ (_08338_, _08337_, _08333_);
  and _16597_ (_08339_, _08338_, _07256_);
  and _16598_ (_08340_, _08339_, _08332_);
  and _16599_ (_08341_, _08340_, _07249_);
  not _16600_ (_08342_, _08341_);
  nor _16601_ (_08343_, _08342_, _08327_);
  and _16602_ (_08344_, _08343_, _08324_);
  and _16603_ (_08345_, _08344_, _08318_);
  nand _16604_ (_08346_, _08345_, _08315_);
  or _16605_ (_08348_, _08346_, _07710_);
  and _16606_ (_08349_, _08126_, _07044_);
  nor _16607_ (_08350_, _07044_, _06649_);
  nor _16608_ (_08351_, _08350_, _08349_);
  nor _16609_ (_08352_, _08351_, _08043_);
  nor _16610_ (_08353_, _08040_, _06649_);
  nor _16611_ (_08354_, _08353_, _08045_);
  not _16612_ (_08355_, _08354_);
  nor _16613_ (_08356_, _08355_, _08352_);
  nor _16614_ (_08357_, _08356_, _07699_);
  nand _16615_ (_08358_, _08357_, _08348_);
  nand _16616_ (_08359_, _08358_, _08309_);
  and _16617_ (_06638_, _08359_, _06989_);
  and _16618_ (_08360_, _06951_, _06889_);
  and _16619_ (_08361_, _08150_, _07500_);
  and _16620_ (_08362_, _08361_, _06871_);
  nor _16621_ (_08363_, _08362_, _06883_);
  nor _16622_ (_08364_, _08147_, _06778_);
  nor _16623_ (_08365_, _08364_, _08363_);
  and _16624_ (_08366_, _08365_, _06889_);
  not _16625_ (_08367_, _08366_);
  nor _16626_ (_08368_, _08365_, _06889_);
  nor _16627_ (_08369_, _08368_, _07101_);
  and _16628_ (_08370_, _08369_, _08367_);
  nor _16629_ (_08371_, _06992_, _06673_);
  or _16630_ (_08372_, _08371_, _08370_);
  or _16631_ (_08373_, _08372_, _06959_);
  and _16632_ (_08374_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  nor _16633_ (_08375_, _08178_, _08173_);
  nor _16634_ (_08376_, _08375_, _08179_);
  and _16635_ (_08377_, _08376_, _06548_);
  and _16636_ (_08378_, _07948_, _07946_);
  not _16637_ (_08379_, _08378_);
  and _16638_ (_08380_, _08379_, _07949_);
  and _16639_ (_08381_, _08380_, _07027_);
  or _16640_ (_08382_, _08381_, _08377_);
  or _16641_ (_08383_, _08382_, _08374_);
  or _16642_ (_08384_, _08383_, _08373_);
  nor _16643_ (_08385_, _08384_, _08360_);
  nor _16644_ (_08386_, _08385_, _07700_);
  not _16645_ (_08387_, _08386_);
  nand _16646_ (_08388_, _07810_, _07752_);
  or _16647_ (_08389_, _07783_, _07753_);
  not _16648_ (_08390_, _07779_);
  and _16649_ (_08391_, _07782_, _08390_);
  and _16650_ (_08392_, _08391_, _08389_);
  nor _16651_ (_08393_, _08391_, _08389_);
  or _16652_ (_08394_, _08393_, _08392_);
  or _16653_ (_08395_, _08394_, _07810_);
  nand _16654_ (_08396_, _08395_, _08388_);
  nand _16655_ (_08397_, _08396_, _07024_);
  nand _16656_ (_08398_, _07975_, _07971_);
  nand _16657_ (_08399_, _08398_, _08216_);
  not _16658_ (_08400_, _08218_);
  and _16659_ (_08401_, _08400_, _08399_);
  nor _16660_ (_08402_, _08401_, _08224_);
  nand _16661_ (_08403_, _08402_, _07027_);
  and _16662_ (_08404_, _06887_, _06876_);
  nor _16663_ (_08405_, _08404_, _06888_);
  nor _16664_ (_08406_, _08405_, _06846_);
  not _16665_ (_08407_, _08406_);
  and _16666_ (_08408_, _06786_, _06771_);
  or _16667_ (_08409_, _08408_, _06549_);
  nor _16668_ (_08410_, _08409_, _06787_);
  not _16669_ (_08411_, _08410_);
  not _16670_ (_08412_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _16671_ (_08413_, _06910_, _08412_);
  nor _16672_ (_08414_, _08413_, _07003_);
  not _16673_ (_08415_, _08414_);
  nor _16674_ (_08416_, _06911_, _06918_);
  and _16675_ (_08417_, _08416_, _08415_);
  not _16676_ (_08418_, _08417_);
  and _16677_ (_08419_, _06951_, _07003_);
  not _16678_ (_08420_, _08419_);
  and _16679_ (_08421_, _08420_, _07310_);
  or _16680_ (_08422_, _07031_, _06646_);
  and _16681_ (_08423_, _07032_, _06700_);
  not _16682_ (_08424_, _08423_);
  nand _16683_ (_08425_, _08424_, _08422_);
  nor _16684_ (_08426_, _08425_, _07314_);
  and _16685_ (_08427_, _08426_, _08421_);
  and _16686_ (_08428_, _08427_, _07307_);
  and _16687_ (_08429_, _08428_, _08418_);
  and _16688_ (_08430_, _08429_, _08411_);
  and _16689_ (_08431_, _08430_, _08407_);
  and _16690_ (_08432_, _08431_, _08403_);
  nand _16691_ (_08433_, _08432_, _08397_);
  or _16692_ (_08434_, _08433_, _07710_);
  nor _16693_ (_08435_, _06537_, _06513_);
  and _16694_ (_08436_, _08435_, _06525_);
  and _16695_ (_08437_, _08126_, _08436_);
  nor _16696_ (_08438_, _08436_, _06677_);
  nor _16697_ (_08439_, _08438_, _08437_);
  nor _16698_ (_08440_, _08439_, _08125_);
  nor _16699_ (_08441_, _08040_, _06677_);
  nor _16700_ (_08442_, _08441_, _08045_);
  not _16701_ (_08443_, _08442_);
  nor _16702_ (_08444_, _08443_, _08440_);
  nor _16703_ (_08445_, _08444_, _07699_);
  nand _16704_ (_08446_, _08445_, _08434_);
  nand _16705_ (_08447_, _08446_, _08387_);
  and _16706_ (_06641_, _08447_, _06989_);
  nand _16707_ (_08448_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nand _16708_ (_08449_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and _16709_ (_08450_, _08449_, _08448_);
  nand _16710_ (_08451_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand _16711_ (_08452_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _16712_ (_08453_, _08452_, _08451_);
  nand _16713_ (_08454_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand _16714_ (_08455_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and _16715_ (_08456_, _08455_, _08454_);
  and _16716_ (_08457_, _08456_, _08453_);
  nand _16717_ (_08458_, _08457_, _08450_);
  nand _16718_ (_08459_, _08458_, _07330_);
  nand _16719_ (_08460_, _08459_, _07328_);
  nor _16720_ (_08461_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _07328_);
  not _16721_ (_08462_, _08461_);
  and _16722_ (_08463_, _08462_, _08460_);
  and _16723_ (_06671_, _08463_, _06989_);
  nor _16724_ (_08464_, _07325_, _06550_);
  and _16725_ (_08465_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and _16726_ (_08466_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _16727_ (_08467_, _08466_, _08465_);
  and _16728_ (_08468_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _16729_ (_08469_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor _16730_ (_08470_, _08469_, _08468_);
  and _16731_ (_08471_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and _16732_ (_08472_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _16733_ (_08473_, _08472_, _08471_);
  and _16734_ (_08474_, _08473_, _08470_);
  and _16735_ (_08475_, _08474_, _08467_);
  and _16736_ (_08476_, _07325_, _07330_);
  not _16737_ (_08477_, _08476_);
  nor _16738_ (_08478_, _08477_, _08475_);
  nor _16739_ (_08479_, _08478_, _08464_);
  nor _16740_ (_06674_, _08479_, rst);
  and _16741_ (_06825_, _07360_, _06989_);
  and _16742_ (_08480_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and _16743_ (_08481_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _16744_ (_08482_, _08481_, _08480_);
  nand _16745_ (_08483_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and _16746_ (_08484_, _08483_, _07330_);
  and _16747_ (_08485_, _08484_, _08482_);
  and _16748_ (_08486_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not _16749_ (_08487_, _08486_);
  and _16750_ (_08488_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _16751_ (_08489_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor _16752_ (_08490_, _08489_, _08488_);
  and _16753_ (_08491_, _08490_, _08487_);
  nand _16754_ (_08492_, _08491_, _08485_);
  or _16755_ (_08493_, _08492_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _16756_ (_08494_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _07328_);
  not _16757_ (_08495_, _08494_);
  and _16758_ (_08496_, _08495_, _08493_);
  and _16759_ (_06827_, _08496_, _06989_);
  and _16760_ (_08497_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _16761_ (_08498_, _08497_);
  nand _16762_ (_08499_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand _16763_ (_08500_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _16764_ (_08501_, _08500_, _08499_);
  nand _16765_ (_08502_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nand _16766_ (_08503_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and _16767_ (_08504_, _08503_, _08502_);
  and _16768_ (_08505_, _08504_, _08501_);
  and _16769_ (_08506_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _16770_ (_08507_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor _16771_ (_08508_, _08507_, _08506_);
  and _16772_ (_08509_, _08508_, _08505_);
  or _16773_ (_08510_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or _16774_ (_08511_, _08510_, _08509_);
  and _16775_ (_08512_, _08511_, _08498_);
  nor _16776_ (_06829_, _08512_, rst);
  nand _16777_ (_08513_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nand _16778_ (_08514_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and _16779_ (_08515_, _08514_, _08513_);
  nand _16780_ (_08516_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand _16781_ (_08517_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _16782_ (_08518_, _08517_, _08516_);
  nand _16783_ (_08519_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand _16784_ (_08520_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and _16785_ (_08522_, _08520_, _08519_);
  and _16786_ (_08523_, _08522_, _08518_);
  nand _16787_ (_08524_, _08523_, _08515_);
  nand _16788_ (_08525_, _08524_, _07330_);
  nand _16789_ (_08526_, _08525_, _07328_);
  nor _16790_ (_08527_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _07328_);
  not _16791_ (_08528_, _08527_);
  and _16792_ (_08529_, _08528_, _08526_);
  and _16793_ (_06831_, _08529_, _06989_);
  and _16794_ (_08530_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _16795_ (_08531_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _16796_ (_08532_, _08531_, _08530_);
  and _16797_ (_08533_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  not _16798_ (_08534_, _08533_);
  and _16799_ (_08535_, _08534_, _08532_);
  and _16800_ (_08536_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _16801_ (_08537_, _08536_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _16802_ (_08538_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _16803_ (_08539_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor _16804_ (_08540_, _08539_, _08538_);
  and _16805_ (_08541_, _08540_, _08537_);
  and _16806_ (_08542_, _08541_, _08535_);
  and _16807_ (_08543_, _08542_, _07328_);
  nor _16808_ (_08544_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _07328_);
  nor _16809_ (_08545_, _08544_, _08543_);
  and _16810_ (_06833_, _08545_, _06989_);
  nand _16811_ (_08546_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nand _16812_ (_08547_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and _16813_ (_08548_, _08547_, _08546_);
  nand _16814_ (_08549_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand _16815_ (_08550_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _16816_ (_08551_, _08550_, _08549_);
  nand _16817_ (_08552_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand _16818_ (_08553_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  and _16819_ (_08554_, _08553_, _08552_);
  and _16820_ (_08555_, _08554_, _08551_);
  nand _16821_ (_08556_, _08555_, _08548_);
  and _16822_ (_08557_, _08556_, _07330_);
  or _16823_ (_08558_, _08557_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor _16824_ (_08559_, _07328_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  not _16825_ (_08560_, _08559_);
  and _16826_ (_08561_, _08560_, _08558_);
  and _16827_ (_06836_, _08561_, _06989_);
  nand _16828_ (_08562_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nand _16829_ (_08563_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and _16830_ (_08564_, _08563_, _08562_);
  nand _16831_ (_08565_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand _16832_ (_08566_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _16833_ (_08567_, _08566_, _08565_);
  nand _16834_ (_08568_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand _16835_ (_08569_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _16836_ (_08570_, _08569_, _08568_);
  and _16837_ (_08571_, _08570_, _08567_);
  and _16838_ (_08572_, _08571_, _08564_);
  or _16839_ (_08573_, _08572_, _08510_);
  and _16840_ (_08574_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not _16841_ (_08575_, _08574_);
  and _16842_ (_08576_, _08575_, _08573_);
  nor _16843_ (_06838_, _08576_, rst);
  nor _16844_ (_08577_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not _16845_ (_08578_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16846_ (_08579_, _08578_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor _16847_ (_08580_, _08579_, _08577_);
  nor _16848_ (_08581_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _16849_ (_08582_, _08578_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nor _16850_ (_08583_, _08582_, _08581_);
  not _16851_ (_08584_, _08583_);
  not _16852_ (_08585_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _16853_ (_08586_, _07493_, _08585_);
  and _16854_ (_08587_, _07493_, _08585_);
  nor _16855_ (_08588_, _08587_, _08586_);
  nor _16856_ (_08589_, _08588_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16857_ (_08590_, _08578_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor _16858_ (_08591_, _08590_, _08589_);
  and _16859_ (_08592_, _08591_, _08584_);
  not _16860_ (_08593_, \oc8051_symbolic_cxrom1.regvalid [13]);
  nor _16861_ (_08594_, _08586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _16862_ (_08595_, _08586_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _16863_ (_08596_, _08595_, _08594_);
  nor _16864_ (_08597_, _08596_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor _16865_ (_08598_, _08578_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor _16866_ (_08599_, _08598_, _08597_);
  and _16867_ (_08600_, _08599_, _08593_);
  nor _16868_ (_08601_, _08599_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _16869_ (_08602_, _08601_, _08600_);
  not _16870_ (_08603_, _08602_);
  nand _16871_ (_08604_, _08603_, _08592_);
  and _16872_ (_08605_, _08604_, _08580_);
  nor _16873_ (_08606_, _08591_, _08584_);
  not _16874_ (_08607_, _08606_);
  not _16875_ (_08608_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _16876_ (_08609_, _08599_, _08608_);
  and _16877_ (_08610_, _08599_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _16878_ (_08611_, _08610_, _08609_);
  nor _16879_ (_08612_, _08611_, _08607_);
  and _16880_ (_08613_, _08591_, _08583_);
  not _16881_ (_08614_, _08613_);
  not _16882_ (_08615_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _16883_ (_08616_, _08599_, _08615_);
  and _16884_ (_08617_, _08599_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _16885_ (_08618_, _08617_, _08616_);
  nor _16886_ (_08619_, _08618_, _08614_);
  nor _16887_ (_08620_, _08619_, _08612_);
  not _16888_ (_08621_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _16889_ (_08622_, _08599_, _08621_);
  nor _16890_ (_08623_, _08591_, _08583_);
  nor _16891_ (_08624_, _08599_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not _16892_ (_08625_, _08624_);
  nand _16893_ (_08626_, _08625_, _08623_);
  or _16894_ (_08627_, _08626_, _08622_);
  and _16895_ (_08628_, _08627_, _08620_);
  and _16896_ (_08629_, _08628_, _08605_);
  and _16897_ (_08630_, _08599_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _16898_ (_08631_, _08630_, _08606_);
  not _16899_ (_08632_, _08599_);
  and _16900_ (_08633_, _08606_, _08632_);
  and _16901_ (_08634_, _08633_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _16902_ (_08635_, _08634_, _08580_);
  or _16903_ (_08636_, _08635_, _08631_);
  not _16904_ (_08637_, _08623_);
  and _16905_ (_08638_, _08599_, \oc8051_symbolic_cxrom1.regvalid [8]);
  not _16906_ (_08639_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _16907_ (_08640_, _08599_, _08639_);
  nor _16908_ (_08641_, _08640_, _08638_);
  nor _16909_ (_08642_, _08641_, _08637_);
  and _16910_ (_08643_, _08632_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _16911_ (_08644_, _08599_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _16912_ (_08645_, _08644_, _08643_);
  nor _16913_ (_08646_, _08645_, _08614_);
  not _16914_ (_08647_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _16915_ (_08648_, _08599_, _08647_);
  nor _16916_ (_08649_, _08599_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or _16917_ (_08650_, _08649_, _08648_);
  not _16918_ (_08651_, _08650_);
  and _16919_ (_08652_, _08651_, _08592_);
  or _16920_ (_08653_, _08652_, _08646_);
  or _16921_ (_08654_, _08653_, _08642_);
  nor _16922_ (_08655_, _08654_, _08636_);
  nor _16923_ (_08656_, _08655_, _08629_);
  not _16924_ (_08657_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand _16925_ (_08658_, _08580_, _08657_);
  or _16926_ (_08659_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _16927_ (_08661_, _08659_, _08658_);
  and _16928_ (_08662_, _08661_, _08613_);
  not _16929_ (_08663_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand _16930_ (_08664_, _08580_, _08663_);
  or _16931_ (_08665_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _16932_ (_08666_, _08665_, _08664_);
  and _16933_ (_08667_, _08666_, _08606_);
  or _16934_ (_08668_, _08667_, _08662_);
  not _16935_ (_08669_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand _16936_ (_08670_, _08580_, _08669_);
  or _16937_ (_08671_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _16938_ (_08672_, _08671_, _08670_);
  and _16939_ (_08673_, _08672_, _08592_);
  not _16940_ (_08674_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand _16941_ (_08675_, _08580_, _08674_);
  or _16942_ (_08676_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _16943_ (_08677_, _08676_, _08675_);
  and _16944_ (_08678_, _08677_, _08623_);
  or _16945_ (_08679_, _08678_, _08673_);
  or _16946_ (_08680_, _08679_, _08668_);
  and _16947_ (_08681_, _08680_, _08599_);
  not _16948_ (_08682_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand _16949_ (_08683_, _08580_, _08682_);
  or _16950_ (_08684_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _16951_ (_08685_, _08684_, _08683_);
  and _16952_ (_08686_, _08685_, _08606_);
  not _16953_ (_08687_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand _16954_ (_08688_, _08580_, _08687_);
  or _16955_ (_08689_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _16956_ (_08690_, _08689_, _08688_);
  and _16957_ (_08691_, _08690_, _08613_);
  or _16958_ (_08692_, _08691_, _08686_);
  not _16959_ (_08693_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand _16960_ (_08694_, _08580_, _08693_);
  or _16961_ (_08695_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _16962_ (_08696_, _08695_, _08694_);
  and _16963_ (_08697_, _08696_, _08592_);
  not _16964_ (_08698_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand _16965_ (_08699_, _08580_, _08698_);
  or _16966_ (_08700_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _16967_ (_08701_, _08700_, _08699_);
  and _16968_ (_08702_, _08701_, _08623_);
  or _16969_ (_08703_, _08702_, _08697_);
  or _16970_ (_08704_, _08703_, _08692_);
  and _16971_ (_08705_, _08704_, _08632_);
  or _16972_ (_08706_, _08705_, _08681_);
  and _16973_ (_08707_, _08706_, _08656_);
  not _16974_ (_08708_, _08656_);
  and _16975_ (_08709_, _08708_, word_in[7]);
  or _16976_ (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _08709_, _08707_);
  not _16977_ (_08710_, _08580_);
  and _16978_ (_08711_, _08583_, _08710_);
  not _16979_ (_08712_, _08711_);
  and _16980_ (_08713_, _08583_, _08580_);
  and _16981_ (_08714_, _08713_, _08591_);
  nor _16982_ (_08715_, _08713_, _08591_);
  nor _16983_ (_08716_, _08715_, _08714_);
  not _16984_ (_08717_, _08716_);
  nor _16985_ (_08718_, _08717_, _08618_);
  nor _16986_ (_08719_, _08714_, _08632_);
  not _16987_ (_08720_, _08591_);
  nor _16988_ (_08721_, _08599_, _08720_);
  and _16989_ (_08722_, _08713_, _08721_);
  nor _16990_ (_08723_, _08722_, _08719_);
  and _16991_ (_08724_, _08723_, _08717_);
  and _16992_ (_08725_, _08724_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _16993_ (_08726_, _08723_, _08716_);
  and _16994_ (_08727_, _08726_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _16995_ (_08728_, _08727_, _08725_);
  nor _16996_ (_08729_, _08728_, _08718_);
  nor _16997_ (_08730_, _08729_, _08712_);
  nor _16998_ (_08731_, _08583_, _08580_);
  not _16999_ (_08732_, _08731_);
  nor _17000_ (_08733_, _08717_, _08602_);
  and _17001_ (_08734_, _08724_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _17002_ (_08735_, _08726_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _17003_ (_08736_, _08735_, _08734_);
  nor _17004_ (_08737_, _08736_, _08733_);
  nor _17005_ (_08738_, _08737_, _08732_);
  nor _17006_ (_08739_, _08738_, _08730_);
  and _17007_ (_08740_, _08584_, _08580_);
  not _17008_ (_08741_, _08740_);
  nor _17009_ (_08742_, _08717_, _08645_);
  and _17010_ (_08743_, _08724_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _17011_ (_08744_, _08726_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17012_ (_08745_, _08744_, _08743_);
  nor _17013_ (_08746_, _08745_, _08742_);
  nor _17014_ (_08747_, _08746_, _08741_);
  not _17015_ (_08748_, _08713_);
  nor _17016_ (_08750_, _08717_, _08650_);
  and _17017_ (_08751_, _08724_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _17018_ (_08752_, _08726_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _17019_ (_08753_, _08752_, _08751_);
  nor _17020_ (_08754_, _08753_, _08750_);
  nor _17021_ (_08755_, _08754_, _08748_);
  nor _17022_ (_08756_, _08755_, _08747_);
  and _17023_ (_08757_, _08756_, _08739_);
  or _17024_ (_08758_, _08713_, _08731_);
  not _17025_ (_08759_, _08758_);
  not _17026_ (_08760_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand _17027_ (_08761_, _08580_, _08760_);
  or _17028_ (_08762_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and _17029_ (_08763_, _08762_, _08761_);
  and _17030_ (_08764_, _08763_, _08759_);
  not _17031_ (_08765_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand _17032_ (_08766_, _08580_, _08765_);
  or _17033_ (_08767_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _17034_ (_08768_, _08767_, _08766_);
  and _17035_ (_08769_, _08768_, _08758_);
  or _17036_ (_08770_, _08769_, _08764_);
  and _17037_ (_08771_, _08770_, _08726_);
  not _17038_ (_08772_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand _17039_ (_08773_, _08580_, _08772_);
  or _17040_ (_08774_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _17041_ (_08775_, _08774_, _08773_);
  and _17042_ (_08776_, _08775_, _08759_);
  not _17043_ (_08777_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand _17044_ (_08778_, _08580_, _08777_);
  or _17045_ (_08779_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and _17046_ (_08780_, _08779_, _08778_);
  and _17047_ (_08781_, _08780_, _08758_);
  or _17048_ (_08782_, _08781_, _08776_);
  and _17049_ (_08783_, _08782_, _08724_);
  and _17050_ (_08784_, _08716_, _08632_);
  not _17051_ (_08785_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand _17052_ (_08786_, _08580_, _08785_);
  or _17053_ (_08787_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _17054_ (_08788_, _08787_, _08786_);
  and _17055_ (_08789_, _08788_, _08759_);
  not _17056_ (_08790_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand _17057_ (_08791_, _08580_, _08790_);
  or _17058_ (_08792_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and _17059_ (_08793_, _08792_, _08791_);
  and _17060_ (_08794_, _08793_, _08758_);
  or _17061_ (_08795_, _08794_, _08789_);
  and _17062_ (_08796_, _08795_, _08784_);
  and _17063_ (_08797_, _08716_, _08599_);
  not _17064_ (_08798_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand _17065_ (_08799_, _08580_, _08798_);
  or _17066_ (_08800_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _17067_ (_08801_, _08800_, _08799_);
  and _17068_ (_08802_, _08801_, _08759_);
  not _17069_ (_08803_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand _17070_ (_08804_, _08580_, _08803_);
  or _17071_ (_08805_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and _17072_ (_08806_, _08805_, _08804_);
  and _17073_ (_08807_, _08806_, _08758_);
  or _17074_ (_08808_, _08807_, _08802_);
  and _17075_ (_08810_, _08808_, _08797_);
  or _17076_ (_08811_, _08810_, _08796_);
  or _17077_ (_08812_, _08811_, _08783_);
  nor _17078_ (_08813_, _08812_, _08771_);
  nor _17079_ (_08814_, _08813_, _08757_);
  and _17080_ (_08815_, _08757_, word_in[15]);
  or _17081_ (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _08815_, _08814_);
  nor _17082_ (_08816_, _08613_, _08623_);
  not _17083_ (_08817_, _08816_);
  nor _17084_ (_08818_, _08817_, _08602_);
  and _17085_ (_08819_, _08613_, _08599_);
  nor _17086_ (_08820_, _08613_, _08599_);
  nor _17087_ (_08821_, _08820_, _08819_);
  and _17088_ (_08822_, _08821_, _08817_);
  and _17089_ (_08823_, _08822_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _17090_ (_08824_, _08821_, _08816_);
  and _17091_ (_08825_, _08824_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or _17092_ (_08826_, _08825_, _08823_);
  nor _17093_ (_08827_, _08826_, _08818_);
  nor _17094_ (_08828_, _08827_, _08748_);
  nor _17095_ (_08829_, _08817_, _08618_);
  and _17096_ (_08830_, _08824_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _17097_ (_08831_, _08822_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _17098_ (_08832_, _08831_, _08830_);
  nor _17099_ (_08833_, _08832_, _08829_);
  nor _17100_ (_08834_, _08833_, _08741_);
  nor _17101_ (_08835_, _08834_, _08828_);
  nor _17102_ (_08836_, _08817_, _08645_);
  and _17103_ (_08837_, _08824_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and _17104_ (_08838_, _08822_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17105_ (_08839_, _08838_, _08837_);
  nor _17106_ (_08841_, _08839_, _08836_);
  nor _17107_ (_08842_, _08841_, _08732_);
  nor _17108_ (_08843_, _08817_, _08650_);
  and _17109_ (_08844_, _08822_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and _17110_ (_08845_, _08824_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _17111_ (_08846_, _08845_, _08844_);
  nor _17112_ (_08847_, _08846_, _08843_);
  nor _17113_ (_08848_, _08847_, _08712_);
  nor _17114_ (_08849_, _08848_, _08842_);
  and _17115_ (_08850_, _08849_, _08835_);
  and _17116_ (_08851_, _08850_, word_in[23]);
  and _17117_ (_08852_, _08696_, _08606_);
  and _17118_ (_08853_, _08685_, _08623_);
  or _17119_ (_08854_, _08853_, _08852_);
  and _17120_ (_08855_, _08690_, _08592_);
  and _17121_ (_08856_, _08701_, _08613_);
  or _17122_ (_08857_, _08856_, _08855_);
  or _17123_ (_08858_, _08857_, _08854_);
  or _17124_ (_08859_, _08858_, _08821_);
  not _17125_ (_08860_, _08821_);
  and _17126_ (_08861_, _08672_, _08606_);
  and _17127_ (_08862_, _08677_, _08632_);
  or _17128_ (_08863_, _08862_, _08861_);
  and _17129_ (_08864_, _08661_, _08592_);
  and _17130_ (_08865_, _08666_, _08623_);
  or _17131_ (_08866_, _08865_, _08864_);
  or _17132_ (_08867_, _08866_, _08863_);
  or _17133_ (_08868_, _08867_, _08860_);
  nand _17134_ (_08869_, _08868_, _08859_);
  nor _17135_ (_08870_, _08869_, _08850_);
  or _17136_ (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _08870_, _08851_);
  nand _17137_ (_08871_, _08732_, _08591_);
  nor _17138_ (_08872_, _08732_, _08591_);
  not _17139_ (_08873_, _08872_);
  and _17140_ (_08874_, _08873_, _08871_);
  not _17141_ (_08875_, _08874_);
  nor _17142_ (_08876_, _08875_, _08618_);
  nor _17143_ (_08877_, _08871_, _08599_);
  and _17144_ (_08878_, _08871_, _08599_);
  nor _17145_ (_08879_, _08878_, _08877_);
  nor _17146_ (_08880_, _08879_, _08874_);
  and _17147_ (_08881_, _08880_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _17148_ (_08882_, _08881_, _08876_);
  nor _17149_ (_08883_, _08882_, _08732_);
  nor _17150_ (_08884_, _08650_, _08875_);
  and _17151_ (_08885_, _08879_, _08875_);
  and _17152_ (_08886_, _08885_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _17153_ (_08887_, _08886_, _08884_);
  and _17154_ (_08888_, _08887_, _08740_);
  and _17155_ (_08889_, _08872_, _08609_);
  and _17156_ (_08890_, _08740_, _08721_);
  and _17157_ (_08891_, _08890_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or _17158_ (_08892_, _08891_, _08889_);
  or _17159_ (_08893_, _08892_, _08888_);
  or _17160_ (_08894_, _08893_, _08883_);
  nor _17161_ (_08895_, _08645_, _08875_);
  and _17162_ (_08896_, _08880_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17163_ (_08897_, _08885_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _17164_ (_08898_, _08897_, _08896_);
  nor _17165_ (_08899_, _08898_, _08895_);
  nor _17166_ (_08900_, _08899_, _08748_);
  nor _17167_ (_08901_, _08875_, _08602_);
  and _17168_ (_08902_, _08885_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _17169_ (_08903_, _08880_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or _17170_ (_08904_, _08903_, _08902_);
  nor _17171_ (_08905_, _08904_, _08901_);
  nor _17172_ (_08906_, _08905_, _08712_);
  or _17173_ (_08907_, _08906_, _08900_);
  nor _17174_ (_08908_, _08907_, _08894_);
  and _17175_ (_08909_, _08768_, _08759_);
  and _17176_ (_08910_, _08763_, _08758_);
  or _17177_ (_08911_, _08910_, _08909_);
  and _17178_ (_08912_, _08911_, _08880_);
  and _17179_ (_08913_, _08780_, _08759_);
  and _17180_ (_08914_, _08775_, _08758_);
  or _17181_ (_08915_, _08914_, _08913_);
  and _17182_ (_08916_, _08915_, _08885_);
  and _17183_ (_08917_, _08874_, _08632_);
  and _17184_ (_08918_, _08793_, _08759_);
  and _17185_ (_08919_, _08788_, _08758_);
  or _17186_ (_08920_, _08919_, _08918_);
  and _17187_ (_08921_, _08920_, _08917_);
  and _17188_ (_08922_, _08806_, _08759_);
  and _17189_ (_08923_, _08801_, _08758_);
  or _17190_ (_08924_, _08923_, _08922_);
  and _17191_ (_08925_, _08878_, _08873_);
  and _17192_ (_08926_, _08925_, _08924_);
  or _17193_ (_08927_, _08926_, _08921_);
  or _17194_ (_08928_, _08927_, _08916_);
  nor _17195_ (_08929_, _08928_, _08912_);
  nor _17196_ (_08930_, _08929_, _08908_);
  and _17197_ (_08931_, _08908_, word_in[31]);
  or _17198_ (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08931_, _08930_);
  and _17199_ (_08932_, _08599_, _08591_);
  or _17200_ (_08933_, _08932_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _17201_ (_07163_, _08933_, _06989_);
  and _17202_ (_08934_, _08932_, _08731_);
  and _17203_ (_08935_, _08908_, _06989_);
  and _17204_ (_08936_, _08935_, _08934_);
  and _17205_ (_08937_, _08850_, _06989_);
  and _17206_ (_08938_, _08937_, _08816_);
  and _17207_ (_08939_, _08938_, _08821_);
  and _17208_ (_08940_, _08939_, _08740_);
  not _17209_ (_08941_, _08940_);
  and _17210_ (_08942_, _08937_, word_in[23]);
  or _17211_ (_08943_, _08942_, _08941_);
  and _17212_ (_08944_, _08757_, _06989_);
  and _17213_ (_08945_, _08944_, _08711_);
  and _17214_ (_08946_, _08945_, _08797_);
  and _17215_ (_08947_, _08629_, _06989_);
  and _17216_ (_08948_, _08947_, _08583_);
  nor _17217_ (_08949_, _08656_, rst);
  and _17218_ (_08950_, _08949_, _08932_);
  and _17219_ (_08951_, _08950_, _08948_);
  nor _17220_ (_08952_, _08951_, _08657_);
  and _17221_ (_08953_, _08949_, word_in[7]);
  and _17222_ (_08954_, _08953_, _08951_);
  or _17223_ (_08955_, _08954_, _08952_);
  or _17224_ (_08956_, _08955_, _08946_);
  not _17225_ (_08957_, _08946_);
  or _17226_ (_08958_, _08957_, word_in[15]);
  and _17227_ (_08959_, _08958_, _08956_);
  or _17228_ (_08960_, _08959_, _08940_);
  and _17229_ (_08961_, _08960_, _08943_);
  or _17230_ (_08963_, _08961_, _08936_);
  not _17231_ (_08964_, _08936_);
  or _17232_ (_08965_, _08964_, word_in[31]);
  and _17233_ (_07192_, _08965_, _08963_);
  or _17234_ (_08966_, _08885_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _17235_ (_07214_, _08966_, _06989_);
  not _17236_ (_08967_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand _17237_ (_08968_, _08623_, _08632_);
  nand _17238_ (_08969_, _08968_, _08967_);
  or _17239_ (_08970_, _08969_, _08819_);
  and _17240_ (_07241_, _08970_, _06989_);
  and _17241_ (_08971_, _08714_, _08599_);
  not _17242_ (_08972_, _08971_);
  and _17243_ (_08973_, _08968_, _08972_);
  not _17244_ (_08974_, _08973_);
  and _17245_ (_08975_, _08740_, _08917_);
  and _17246_ (_08976_, _08711_, _08917_);
  nor _17247_ (_08977_, _08976_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _17248_ (_08978_, _08977_, _08975_);
  or _17249_ (_08979_, _08978_, _08974_);
  and _17250_ (_07280_, _08979_, _06989_);
  not _17251_ (_08980_, _08724_);
  and _17252_ (_08981_, _08713_, _08917_);
  or _17253_ (_08982_, _08981_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _17254_ (_08983_, _08982_, _08980_);
  and _17255_ (_08984_, _08609_, _08623_);
  or _17256_ (_08985_, _08984_, _08976_);
  or _17257_ (_08986_, _08985_, _08983_);
  and _17258_ (_08987_, _08986_, _08973_);
  not _17259_ (_08988_, _08968_);
  and _17260_ (_08989_, _08982_, _08971_);
  or _17261_ (_08990_, _08989_, _08988_);
  or _17262_ (_08991_, _08990_, _08987_);
  and _17263_ (_07329_, _08991_, _06989_);
  not _17264_ (_08992_, _07090_);
  nand _17265_ (_08993_, _07086_, _06975_);
  nor _17266_ (_08994_, _08993_, _08992_);
  not _17267_ (_08995_, _07128_);
  nor _17268_ (_08996_, _08993_, _08995_);
  nor _17269_ (_08997_, _08996_, _08994_);
  and _17270_ (_08998_, _08997_, _07127_);
  or _17271_ (_08999_, _08998_, _06982_);
  and _17272_ (_09000_, _08999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  not _17273_ (_09001_, _07126_);
  nand _17274_ (_09002_, _08997_, _09001_);
  and _17275_ (_09003_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and _17276_ (_09004_, _09003_, _09002_);
  nor _17277_ (_09005_, _07035_, _06728_);
  not _17278_ (_09006_, _09005_);
  and _17279_ (_09007_, _09006_, _08000_);
  and _17280_ (_09008_, _09007_, _08018_);
  not _17281_ (_09009_, _09008_);
  and _17282_ (_09010_, _07123_, _06981_);
  and _17283_ (_09011_, _09010_, _09009_);
  or _17284_ (_09012_, _09011_, _09004_);
  or _17285_ (_09013_, _09012_, _09000_);
  and _17286_ (_07336_, _09013_, _06989_);
  or _17287_ (_09014_, _08975_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _17288_ (_09015_, _09014_, _08974_);
  and _17289_ (_09016_, _08721_, _08731_);
  or _17290_ (_09017_, _09016_, _08981_);
  or _17291_ (_09018_, _09017_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _17292_ (_09019_, _09018_, _08980_);
  or _17293_ (_09020_, _09019_, _09015_);
  or _17294_ (_09021_, _09020_, _08976_);
  and _17295_ (_07388_, _09021_, _06989_);
  and _17296_ (_09022_, _06478_, _06463_);
  and _17297_ (_09023_, _09022_, _08037_);
  and _17298_ (_09024_, _09023_, _06539_);
  nand _17299_ (_09025_, _09024_, _06968_);
  or _17300_ (_09026_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and _17301_ (_09027_, _09026_, _06485_);
  and _17302_ (_09028_, _09027_, _09025_);
  and _17303_ (_09029_, _07706_, _07453_);
  and _17304_ (_09030_, _09029_, _07125_);
  not _17305_ (_09031_, _09030_);
  nor _17306_ (_09032_, _09031_, _07040_);
  not _17307_ (_09033_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  nor _17308_ (_09034_, _09030_, _09033_);
  or _17309_ (_09035_, _09034_, _09032_);
  and _17310_ (_09036_, _09035_, _06983_);
  nor _17311_ (_09037_, _06484_, _09033_);
  or _17312_ (_09038_, _09037_, rst);
  or _17313_ (_09039_, _09038_, _09036_);
  or _17314_ (_07448_, _09039_, _09028_);
  and _17315_ (_09040_, _08872_, _08632_);
  nor _17316_ (_09041_, _09040_, _08917_);
  not _17317_ (_09042_, _08820_);
  or _17318_ (_09043_, _09042_, _09017_);
  and _17319_ (_09044_, _09043_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and _17320_ (_09045_, _08976_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _17321_ (_09046_, _09045_, _08890_);
  or _17322_ (_09048_, _09046_, _09044_);
  and _17323_ (_09049_, _09048_, _09041_);
  and _17324_ (_09050_, _08988_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or _17325_ (_09051_, _09050_, _08976_);
  or _17326_ (_09052_, _09051_, _09016_);
  or _17327_ (_09053_, _09052_, _08981_);
  or _17328_ (_09054_, _09053_, _09049_);
  and _17329_ (_07451_, _09054_, _06989_);
  or _17330_ (_09055_, _08719_, _08877_);
  and _17331_ (_09056_, _08932_, _08711_);
  or _17332_ (_09057_, _08821_, _09056_);
  and _17333_ (_09058_, _08711_, _08721_);
  or _17334_ (_09059_, _09058_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and _17335_ (_09060_, _09059_, _09057_);
  and _17336_ (_09061_, _09017_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _17337_ (_09062_, _09061_, _08890_);
  or _17338_ (_09063_, _09062_, _09060_);
  and _17339_ (_09064_, _09063_, _09055_);
  and _17340_ (_09065_, _09059_, _08971_);
  and _17341_ (_09066_, _08715_, _08643_);
  or _17342_ (_09067_, _09066_, _08981_);
  or _17343_ (_09068_, _09067_, _09016_);
  or _17344_ (_09069_, _09068_, _09065_);
  or _17345_ (_09070_, _09069_, _09064_);
  and _17346_ (_07503_, _09070_, _06989_);
  and _17347_ (_09071_, _07704_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and _17348_ (_09072_, _06983_, _06447_);
  nor _17349_ (_09073_, _06537_, _06514_);
  and _17350_ (_09074_, _09073_, _06525_);
  and _17351_ (_09075_, _07454_, _09074_);
  and _17352_ (_09076_, _09075_, _09072_);
  nor _17353_ (_09077_, _09076_, _09071_);
  or _17354_ (_09078_, _09077_, _08123_);
  not _17355_ (_09079_, _09077_);
  or _17356_ (_09080_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and _17357_ (_09081_, _09080_, _06989_);
  and _17358_ (_07578_, _09081_, _09078_);
  nor _17359_ (_09082_, _07793_, _07725_);
  or _17360_ (_09083_, _09082_, _07794_);
  nand _17361_ (_09084_, _09083_, _07814_);
  or _17362_ (_09085_, _07814_, _07722_);
  and _17363_ (_09086_, _09085_, _09084_);
  nand _17364_ (_09087_, _09086_, _07024_);
  and _17365_ (_09088_, _08227_, _08224_);
  and _17366_ (_09089_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  nand _17367_ (_09090_, _09089_, _09088_);
  or _17368_ (_09091_, _09089_, _09088_);
  and _17369_ (_09092_, _09091_, _09090_);
  nand _17370_ (_09093_, _09092_, _07027_);
  nor _17371_ (_09094_, _06826_, _06792_);
  not _17372_ (_09095_, _09094_);
  nor _17373_ (_09096_, _06828_, _06549_);
  and _17374_ (_09097_, _09096_, _09095_);
  not _17375_ (_09098_, _09097_);
  nor _17376_ (_09099_, _06896_, _06861_);
  nor _17377_ (_09100_, _09099_, _06897_);
  nor _17378_ (_09101_, _09100_, _06846_);
  and _17379_ (_09102_, _06810_, _06883_);
  not _17380_ (_09103_, _09102_);
  and _17381_ (_09104_, _06816_, _06778_);
  nor _17382_ (_09105_, _09104_, _06992_);
  and _17383_ (_09106_, _09105_, _09103_);
  or _17384_ (_09107_, _07008_, _06902_);
  and _17385_ (_09108_, _09107_, _07010_);
  and _17386_ (_09109_, _07000_, _07096_);
  nor _17387_ (_09110_, _09109_, _06810_);
  or _17388_ (_09111_, _09110_, _07001_);
  and _17389_ (_09112_, _09111_, _06778_);
  or _17390_ (_09113_, _09112_, _09108_);
  and _17391_ (_09114_, _09113_, _06997_);
  nor _17392_ (_09115_, _09114_, _09106_);
  nor _17393_ (_09116_, _08247_, _06810_);
  and _17394_ (_09117_, _08247_, _06810_);
  nor _17395_ (_09118_, _09117_, _09116_);
  nor _17396_ (_09119_, _09118_, _06918_);
  and _17397_ (_09120_, _06951_, _06902_);
  not _17398_ (_09121_, _09120_);
  or _17399_ (_09123_, _07031_, _06586_);
  nand _17400_ (_09124_, _07032_, _06616_);
  and _17401_ (_09125_, _09124_, _09123_);
  and _17402_ (_09126_, _09125_, _09121_);
  and _17403_ (_09127_, _06942_, _06819_);
  and _17404_ (_09128_, _06933_, _06817_);
  nor _17405_ (_09129_, _07017_, _06818_);
  and _17406_ (_09130_, _06954_, _06810_);
  or _17407_ (_09131_, _09130_, _09129_);
  or _17408_ (_09132_, _09131_, _09128_);
  nor _17409_ (_09133_, _09132_, _09127_);
  and _17410_ (_09134_, _09133_, _09126_);
  not _17411_ (_09136_, _09134_);
  nor _17412_ (_09138_, _09136_, _09119_);
  and _17413_ (_09139_, _09138_, _09115_);
  not _17414_ (_09140_, _09139_);
  nor _17415_ (_09142_, _09140_, _09101_);
  and _17416_ (_09143_, _09142_, _09098_);
  and _17417_ (_09144_, _09143_, _09093_);
  and _17418_ (_09145_, _09144_, _09087_);
  nand _17419_ (_09146_, _09145_, _09079_);
  or _17420_ (_09147_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _17421_ (_09148_, _09147_, _06989_);
  and _17422_ (_07581_, _09148_, _09146_);
  or _17423_ (_09149_, _09077_, _08268_);
  or _17424_ (_09150_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and _17425_ (_09151_, _09150_, _06989_);
  and _17426_ (_07584_, _09151_, _09149_);
  or _17427_ (_09153_, _09077_, _08346_);
  or _17428_ (_09155_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and _17429_ (_09156_, _09155_, _06989_);
  and _17430_ (_07592_, _09156_, _09153_);
  or _17431_ (_09157_, _08714_, _08599_);
  nor _17432_ (_09158_, _08599_, _08710_);
  or _17433_ (_09159_, _09158_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and _17434_ (_09160_, _09159_, _09042_);
  and _17435_ (_09161_, _08616_, _08614_);
  or _17436_ (_09162_, _09161_, _09160_);
  and _17437_ (_09163_, _09162_, _09157_);
  and _17438_ (_09164_, _08874_, _08616_);
  and _17439_ (_09165_, _09040_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or _17440_ (_09166_, _09165_, _09016_);
  or _17441_ (_09167_, _09166_, _09164_);
  or _17442_ (_09168_, _09167_, _08890_);
  or _17443_ (_09169_, _09168_, _09058_);
  or _17444_ (_09170_, _09169_, _09163_);
  and _17445_ (_07599_, _09170_, _06989_);
  or _17446_ (_09171_, _09077_, _08433_);
  or _17447_ (_09172_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _17448_ (_09173_, _09172_, _06989_);
  and _17449_ (_07616_, _09173_, _09171_);
  and _17450_ (_09174_, _07781_, _07771_);
  not _17451_ (_09175_, _09174_);
  and _17452_ (_09176_, _09175_, _07782_);
  or _17453_ (_09177_, _09176_, _07810_);
  or _17454_ (_09178_, _07814_, _07778_);
  and _17455_ (_09179_, _09178_, _09177_);
  nand _17456_ (_09180_, _09179_, _07024_);
  or _17457_ (_09181_, _08398_, _08216_);
  and _17458_ (_09182_, _09181_, _08399_);
  nand _17459_ (_09183_, _09182_, _07027_);
  nor _17460_ (_09184_, _06784_, _06782_);
  not _17461_ (_09185_, _09184_);
  nor _17462_ (_09186_, _06785_, _06549_);
  and _17463_ (_09187_, _09186_, _09185_);
  not _17464_ (_09188_, _09187_);
  nor _17465_ (_09189_, _06885_, _06879_);
  nor _17466_ (_09190_, _09189_, _06886_);
  nor _17467_ (_09191_, _09190_, _06846_);
  not _17468_ (_09192_, _09191_);
  and _17469_ (_09193_, _06991_, _06706_);
  nor _17470_ (_09194_, _07004_, _06778_);
  nor _17471_ (_09195_, _08012_, _06883_);
  nor _17472_ (_09196_, _09195_, _09194_);
  and _17473_ (_09197_, _09196_, _06700_);
  not _17474_ (_09198_, _09197_);
  nor _17475_ (_09199_, _09196_, _06700_);
  nor _17476_ (_09200_, _09199_, _07101_);
  and _17477_ (_09201_, _09200_, _09198_);
  nor _17478_ (_09202_, _09201_, _09193_);
  and _17479_ (_09203_, _06910_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  not _17480_ (_09204_, _06700_);
  nor _17481_ (_09205_, _07987_, _09204_);
  nor _17482_ (_09206_, _09205_, _09203_);
  nor _17483_ (_09207_, _09206_, _06918_);
  nor _17484_ (_09208_, _07017_, _06708_);
  and _17485_ (_09209_, _06942_, _06709_);
  nor _17486_ (_09210_, _09209_, _09208_);
  and _17487_ (_09211_, _06933_, _06707_);
  and _17488_ (_09212_, _06954_, _09204_);
  nor _17489_ (_09213_, _09212_, _09211_);
  or _17490_ (_09214_, _07031_, _06673_);
  nor _17491_ (_09215_, _08001_, _06728_);
  and _17492_ (_09216_, _06951_, _06700_);
  nor _17493_ (_09217_, _09216_, _09215_);
  and _17494_ (_09218_, _09217_, _09214_);
  and _17495_ (_09219_, _09218_, _09213_);
  and _17496_ (_09220_, _09219_, _09210_);
  not _17497_ (_09221_, _09220_);
  nor _17498_ (_09222_, _09221_, _09207_);
  and _17499_ (_09223_, _09222_, _09202_);
  and _17500_ (_09224_, _09223_, _09192_);
  and _17501_ (_09225_, _09224_, _09188_);
  and _17502_ (_09226_, _09225_, _09183_);
  and _17503_ (_09227_, _09226_, _09180_);
  nand _17504_ (_09228_, _09227_, _09079_);
  or _17505_ (_09229_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and _17506_ (_09230_, _09229_, _06989_);
  and _17507_ (_07620_, _09230_, _09228_);
  or _17508_ (_09231_, _09077_, _08030_);
  or _17509_ (_09232_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _17510_ (_09233_, _09232_, _06989_);
  and _17511_ (_07635_, _09233_, _09231_);
  not _17512_ (_09234_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _17513_ (_09236_, _08877_, _09234_);
  or _17514_ (_09237_, _09236_, _08880_);
  and _17515_ (_07673_, _09237_, _06989_);
  and _17516_ (_09239_, _07454_, _09072_);
  nand _17517_ (_09240_, _09239_, _08436_);
  nor _17518_ (_09241_, _09240_, _09145_);
  and _17519_ (_09242_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _17520_ (_09244_, _09242_, _09071_);
  or _17521_ (_09245_, _09244_, _09241_);
  and _17522_ (_09246_, _06951_, _06850_);
  and _17523_ (_09248_, _06958_, _06700_);
  and _17524_ (_09249_, _08148_, _06853_);
  and _17525_ (_09250_, _09249_, _06623_);
  or _17526_ (_09252_, _09250_, _06778_);
  and _17527_ (_09253_, _08154_, _06622_);
  or _17528_ (_09255_, _09253_, _06883_);
  and _17529_ (_09256_, _09255_, _09252_);
  and _17530_ (_09258_, _09256_, _06816_);
  nor _17531_ (_09259_, _09256_, _06816_);
  or _17532_ (_09260_, _09259_, _09258_);
  and _17533_ (_09261_, _09260_, _06997_);
  nor _17534_ (_09262_, _06816_, _06778_);
  nor _17535_ (_09263_, _06810_, _06883_);
  or _17536_ (_09264_, _09263_, _09262_);
  and _17537_ (_09265_, _09264_, _06991_);
  or _17538_ (_09266_, _09265_, _09261_);
  or _17539_ (_09267_, _09266_, _09248_);
  and _17540_ (_09268_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor _17541_ (_09269_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not _17542_ (_09270_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _17543_ (_09271_, _09270_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor _17544_ (_09272_, _09271_, _09269_);
  nor _17545_ (_09273_, _09272_, _08191_);
  not _17546_ (_09274_, _09273_);
  and _17547_ (_09275_, _09272_, _08191_);
  nor _17548_ (_09276_, _09275_, _06549_);
  and _17549_ (_09277_, _09276_, _09274_);
  and _17550_ (_09278_, _07956_, _07926_);
  not _17551_ (_09279_, _09278_);
  and _17552_ (_09280_, _09279_, _07957_);
  and _17553_ (_09281_, _09280_, _07027_);
  or _17554_ (_09282_, _09281_, _09277_);
  or _17555_ (_09283_, _09282_, _09268_);
  or _17556_ (_09284_, _09283_, _09267_);
  nor _17557_ (_09285_, _09284_, _09246_);
  nand _17558_ (_09286_, _09285_, _09071_);
  and _17559_ (_09287_, _09286_, _06989_);
  and _17560_ (_07764_, _09287_, _09245_);
  and _17561_ (_09288_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _17562_ (_09289_, _07124_, _08435_);
  and _17563_ (_09290_, _09289_, _07454_);
  and _17564_ (_09291_, _09290_, _06484_);
  and _17565_ (_09292_, _09291_, _06980_);
  and _17566_ (_09293_, _09292_, _08268_);
  or _17567_ (_09294_, _09293_, _09288_);
  or _17568_ (_09295_, _09294_, _09071_);
  nand _17569_ (_09296_, _09071_, _08202_);
  and _17570_ (_09297_, _09296_, _06989_);
  and _17571_ (_07767_, _09297_, _09295_);
  and _17572_ (_09298_, _08820_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _17573_ (_09299_, _08872_, _08599_);
  and _17574_ (_09300_, _08719_, _08873_);
  and _17575_ (_09301_, _08925_, _08740_);
  nor _17576_ (_09302_, _08820_, _08621_);
  or _17577_ (_09303_, _09302_, _09301_);
  and _17578_ (_09304_, _09303_, _09300_);
  or _17579_ (_09306_, _09304_, _09299_);
  and _17580_ (_09307_, _09303_, _08971_);
  or _17581_ (_09308_, _09307_, _09058_);
  or _17582_ (_09309_, _09308_, _08722_);
  or _17583_ (_09310_, _09309_, _09306_);
  or _17584_ (_09311_, _09310_, _09298_);
  and _17585_ (_07773_, _09311_, _06989_);
  and _17586_ (_09312_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _17587_ (_09313_, _09292_, _08346_);
  or _17588_ (_09314_, _09313_, _09312_);
  or _17589_ (_09315_, _09314_, _09071_);
  nand _17590_ (_09316_, _09071_, _08307_);
  and _17591_ (_09317_, _09316_, _06989_);
  and _17592_ (_07785_, _09317_, _09315_);
  and _17593_ (_09318_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  and _17594_ (_09319_, _09292_, _08433_);
  or _17595_ (_09320_, _09319_, _09318_);
  or _17596_ (_09321_, _09320_, _09071_);
  nand _17597_ (_09322_, _09071_, _08385_);
  and _17598_ (_09323_, _09322_, _06989_);
  and _17599_ (_07806_, _09323_, _09321_);
  nor _17600_ (_09324_, _09240_, _09227_);
  and _17601_ (_09325_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or _17602_ (_09326_, _09325_, _09071_);
  or _17603_ (_09327_, _09326_, _09324_);
  and _17604_ (_09329_, _06951_, _06706_);
  and _17605_ (_09330_, _06958_, _06902_);
  nor _17606_ (_09331_, _08146_, _06778_);
  nor _17607_ (_09332_, _08361_, _06883_);
  nor _17608_ (_09333_, _09332_, _09331_);
  nor _17609_ (_09334_, _09333_, _06706_);
  and _17610_ (_09336_, _09333_, _06706_);
  nor _17611_ (_09337_, _09336_, _09334_);
  and _17612_ (_09338_, _09337_, _06997_);
  and _17613_ (_09339_, _06991_, _06700_);
  or _17614_ (_09340_, _09339_, _09338_);
  or _17615_ (_09341_, _09340_, _09330_);
  and _17616_ (_09342_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor _17617_ (_09343_, _08177_, _07657_);
  nor _17618_ (_09344_, _09343_, _08178_);
  and _17619_ (_09345_, _09344_, _06548_);
  and _17620_ (_09347_, _07945_, _07943_);
  not _17621_ (_09348_, _09347_);
  and _17622_ (_09349_, _09348_, _07946_);
  and _17623_ (_09350_, _09349_, _07027_);
  or _17624_ (_09352_, _09350_, _09345_);
  or _17625_ (_09353_, _09352_, _09342_);
  or _17626_ (_09355_, _09353_, _09341_);
  nor _17627_ (_09356_, _09355_, _09329_);
  nand _17628_ (_09357_, _09356_, _09071_);
  and _17629_ (_09358_, _09357_, _06989_);
  and _17630_ (_07820_, _09358_, _09327_);
  and _17631_ (_09359_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  and _17632_ (_09360_, _09292_, _08030_);
  or _17633_ (_09361_, _09360_, _09359_);
  or _17634_ (_09362_, _09361_, _09071_);
  nand _17635_ (_09363_, _09071_, _07696_);
  and _17636_ (_09364_, _09363_, _06989_);
  and _17637_ (_07829_, _09364_, _09362_);
  and _17638_ (_09365_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _17639_ (_09366_, _09292_, _08123_);
  or _17640_ (_09367_, _09366_, _09365_);
  or _17641_ (_09368_, _09367_, _09071_);
  not _17642_ (_09369_, _09071_);
  or _17643_ (_09370_, _09369_, _08075_);
  and _17644_ (_09371_, _09370_, _06989_);
  and _17645_ (_07834_, _09371_, _09368_);
  and _17646_ (_09372_, _08711_, _08878_);
  not _17647_ (_09373_, _08715_);
  and _17648_ (_09374_, _09373_, _08630_);
  or _17649_ (_09375_, _09374_, _09372_);
  or _17650_ (_09376_, _09058_, _08988_);
  and _17651_ (_09377_, _09376_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _17652_ (_09378_, _08816_, _08632_);
  and _17653_ (_09379_, _09378_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _17654_ (_09380_, _09379_, _08722_);
  or _17655_ (_09381_, _09380_, _09377_);
  or _17656_ (_09382_, _09381_, _09301_);
  or _17657_ (_09383_, _09382_, _09299_);
  or _17658_ (_09384_, _09383_, _09375_);
  and _17659_ (_07869_, _09384_, _06989_);
  nand _17660_ (_09385_, _08512_, _07326_);
  nor _17661_ (_09386_, _07325_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor _17662_ (_09387_, _09386_, _07362_);
  and _17663_ (_09388_, _09387_, _09385_);
  and _17664_ (_07933_, _09388_, _06989_);
  not _17665_ (_09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _17666_ (_09390_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _17667_ (_09391_, _09390_, _06989_);
  nor _17668_ (_09392_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not _17669_ (_09393_, _09392_);
  and _17670_ (_09394_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _17671_ (_09395_, _09394_, _09393_);
  not _17672_ (_09396_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor _17673_ (_09397_, _09396_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not _17674_ (_09398_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor _17675_ (_09399_, _09398_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _17676_ (_09400_, _09399_, _09397_);
  not _17677_ (_09401_, _09400_);
  and _17678_ (_09402_, _09401_, _09395_);
  and _17679_ (_09403_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and _17680_ (_09404_, _09403_, _09393_);
  not _17681_ (_09405_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor _17682_ (_09406_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _09405_);
  not _17683_ (_09407_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and _17684_ (_09408_, _09392_, _09407_);
  and _17685_ (_09409_, _09408_, _09406_);
  nor _17686_ (_09410_, _09409_, _09395_);
  not _17687_ (_09411_, _09410_);
  nor _17688_ (_09412_, _09411_, _09404_);
  nor _17689_ (_09413_, _09412_, _09402_);
  and _17690_ (_09414_, _09392_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and _17691_ (_09415_, _09414_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or _17692_ (_09416_, _09415_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or _17693_ (_09417_, _09416_, _09413_);
  and _17694_ (_09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _06989_);
  and _17695_ (_09419_, _09400_, _09395_);
  nor _17696_ (_09420_, _09419_, _09415_);
  or _17697_ (_09421_, _09420_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _17698_ (_09422_, _09421_, _09418_);
  and _17699_ (_09423_, _09422_, _09417_);
  or _17700_ (_07959_, _09423_, _09391_);
  not _17701_ (_09424_, _09420_);
  nor _17702_ (_09425_, _09409_, _09404_);
  nor _17703_ (_09426_, _09425_, _09395_);
  nor _17704_ (_09427_, _09426_, _09424_);
  nor _17705_ (_09428_, _09427_, _09389_);
  or _17706_ (_09429_, _09428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _17707_ (_09430_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or _17708_ (_09431_, _09430_, _09420_);
  and _17709_ (_09432_, _09431_, _06989_);
  and _17710_ (_07969_, _09432_, _09429_);
  and _17711_ (_09433_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and _17712_ (_09434_, _09433_, _06989_);
  or _17713_ (_09435_, _09426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _17714_ (_09436_, _09435_, _09424_);
  or _17715_ (_09437_, _09420_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and _17716_ (_09438_, _09437_, _09418_);
  and _17717_ (_09439_, _09438_, _09436_);
  or _17718_ (_07973_, _09439_, _09434_);
  and _17719_ (_09440_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _17720_ (_09441_, _09440_, _06989_);
  or _17721_ (_09442_, _09426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and _17722_ (_09443_, _09442_, _09420_);
  and _17723_ (_09444_, _09424_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or _17724_ (_09445_, _09444_, _09443_);
  and _17725_ (_09446_, _09445_, _09418_);
  or _17726_ (_07976_, _09446_, _09441_);
  and _17727_ (_09447_, _08713_, _08878_);
  and _17728_ (_09448_, _08932_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _17729_ (_09449_, _09448_, _09447_);
  or _17730_ (_09450_, _08599_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and _17731_ (_09451_, _09450_, _08872_);
  or _17732_ (_09452_, _09451_, _09301_);
  or _17733_ (_09453_, _09452_, _09449_);
  nor _17734_ (_09454_, _08872_, _08599_);
  and _17735_ (_09455_, _09454_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _17736_ (_09456_, _09455_, _09372_);
  or _17737_ (_09457_, _09456_, _09453_);
  and _17738_ (_07980_, _09457_, _06989_);
  and _17739_ (_09458_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _17740_ (_09459_, _09458_, _06989_);
  or _17741_ (_09460_, _09426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and _17742_ (_09461_, _09460_, _09420_);
  and _17743_ (_09462_, _09424_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or _17744_ (_09463_, _09462_, _09461_);
  and _17745_ (_09464_, _09463_, _09418_);
  or _17746_ (_07989_, _09464_, _09459_);
  and _17747_ (_09465_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _17748_ (_09466_, _09465_, _06989_);
  or _17749_ (_09467_, _09426_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and _17750_ (_09468_, _09467_, _09420_);
  and _17751_ (_09469_, _09424_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or _17752_ (_09470_, _09469_, _09468_);
  and _17753_ (_09471_, _09470_, _09418_);
  or _17754_ (_07992_, _09471_, _09466_);
  or _17755_ (_09472_, _09428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _17756_ (_09473_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or _17757_ (_09474_, _09473_, _09420_);
  and _17758_ (_09475_, _09474_, _06989_);
  and _17759_ (_07997_, _09475_, _09472_);
  and _17760_ (_09476_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _17761_ (_09477_, _09476_, _06989_);
  and _17762_ (_09478_, _09424_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _17763_ (_09479_, _09402_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or _17764_ (_09480_, _09479_, _09410_);
  not _17765_ (_09481_, _09415_);
  or _17766_ (_09482_, _09404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and _17767_ (_09483_, _09482_, _09481_);
  and _17768_ (_09484_, _09483_, _09480_);
  or _17769_ (_09485_, _09484_, _09478_);
  and _17770_ (_09486_, _09485_, _09418_);
  or _17771_ (_08054_, _09486_, _09477_);
  and _17772_ (_09487_, _07135_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and _17773_ (_09488_, _07091_, _06981_);
  not _17774_ (_09489_, _09488_);
  nor _17775_ (_09490_, _09489_, _07260_);
  or _17776_ (_09491_, _09490_, _09487_);
  and _17777_ (_08073_, _09491_, _06989_);
  and _17778_ (_09492_, _08932_, _08732_);
  and _17779_ (_09493_, _09492_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _17780_ (_09494_, _08721_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and _17781_ (_09495_, _08633_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _17782_ (_09496_, _09495_, _08925_);
  or _17783_ (_09497_, _08975_, _08872_);
  and _17784_ (_09498_, _09497_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _17785_ (_09499_, _09498_, _09496_);
  or _17786_ (_09500_, _09499_, _09494_);
  or _17787_ (_09501_, _09500_, _09493_);
  and _17788_ (_08081_, _09501_, _06989_);
  nor _17789_ (_08088_, _07319_, rst);
  or _17790_ (_09502_, _09428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _17791_ (_09503_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or _17792_ (_09504_, _09503_, _09420_);
  and _17793_ (_09505_, _09504_, _06989_);
  and _17794_ (_08094_, _09505_, _09502_);
  and _17795_ (_09506_, _09400_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _17796_ (_09507_, _09506_, _09425_);
  or _17797_ (_09508_, _09507_, _09427_);
  and _17798_ (_09509_, _09508_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _17799_ (_09510_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nand _17800_ (_09511_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor _17801_ (_09512_, _09511_, _09420_);
  or _17802_ (_09513_, _09512_, _09510_);
  or _17803_ (_09514_, _09513_, _09509_);
  and _17804_ (_08097_, _09514_, _06989_);
  not _17805_ (_09515_, _09428_);
  and _17806_ (_09516_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and _17807_ (_09517_, _09516_, _09515_);
  and _17808_ (_09518_, _09400_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nand _17809_ (_09519_, _09518_, _09425_);
  nand _17810_ (_09520_, _09519_, _09420_);
  and _17811_ (_09521_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and _17812_ (_09523_, _09521_, _09520_);
  or _17813_ (_08100_, _09523_, _09517_);
  and _17814_ (_09524_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  not _17815_ (_09525_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nor _17816_ (_09527_, _07493_, _09525_);
  or _17817_ (_09528_, _09527_, _09524_);
  and _17818_ (_08105_, _09528_, _06989_);
  and _17819_ (_09529_, _08436_, _06448_);
  and _17820_ (_09530_, _09529_, _06983_);
  and _17821_ (_09531_, _09530_, _06977_);
  nand _17822_ (_09532_, _09531_, _07040_);
  and _17823_ (_09533_, _07145_, _07075_);
  not _17824_ (_09534_, _09533_);
  and _17825_ (_09535_, _06985_, _09074_);
  and _17826_ (_09536_, _09535_, _06977_);
  nor _17827_ (_09537_, _09536_, _09534_);
  nor _17828_ (_09538_, _09537_, _07152_);
  and _17829_ (_09539_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or _17830_ (_09541_, _09539_, _09538_);
  or _17831_ (_09542_, _09531_, _09541_);
  and _17832_ (_09543_, _09542_, _06989_);
  and _17833_ (_08108_, _09543_, _09532_);
  or _17834_ (_09544_, _08496_, _07327_);
  nor _17835_ (_09545_, _07325_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor _17836_ (_09546_, _09545_, _07362_);
  and _17837_ (_09547_, _09546_, _09544_);
  and _17838_ (_08111_, _09547_, _06989_);
  and _17839_ (_09548_, _07958_, _07920_);
  not _17840_ (_09549_, _09548_);
  and _17841_ (_09550_, _09549_, _07960_);
  and _17842_ (_08135_, _09550_, _06989_);
  nand _17843_ (_09551_, _09536_, _07040_);
  not _17844_ (_09552_, _09531_);
  not _17845_ (_09553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor _17846_ (_09554_, _09533_, _09553_);
  and _17847_ (_09555_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or _17848_ (_09556_, _09555_, _09554_);
  or _17849_ (_09557_, _09556_, _09536_);
  and _17850_ (_09558_, _09557_, _09552_);
  and _17851_ (_09559_, _09558_, _09551_);
  and _17852_ (_09560_, _06985_, _08436_);
  and _17853_ (_09561_, _09560_, _06977_);
  and _17854_ (_09562_, _09561_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _17855_ (_09563_, _09562_, _09559_);
  and _17856_ (_08181_, _09563_, _06989_);
  and _17857_ (_08194_, _07365_, _06989_);
  and _17858_ (_09564_, _08821_, _08816_);
  or _17859_ (_09565_, _09564_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _17860_ (_08217_, _09565_, _06989_);
  nor _17861_ (_09566_, t2_i, rst);
  and _17862_ (_08250_, _09566_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  not _17863_ (_09567_, _07066_);
  and _17864_ (_09568_, _07073_, _07071_);
  and _17865_ (_09569_, _09568_, _07051_);
  nand _17866_ (_09570_, _09569_, _09567_);
  or _17867_ (_09571_, _09569_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and _17868_ (_09572_, _09571_, _06989_);
  and _17869_ (_08266_, _09572_, _09570_);
  nand _17870_ (_09573_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _06989_);
  nor _17871_ (_08297_, _09573_, t2ex_i);
  and _17872_ (_08321_, t2ex_i, _06989_);
  not _17873_ (_09574_, _07077_);
  and _17874_ (_09575_, _07071_, _07057_);
  or _17875_ (_09576_, _09575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand _17876_ (_09577_, _07071_, _07058_);
  and _17877_ (_09578_, _09577_, _09576_);
  nor _17878_ (_09579_, _07145_, _09553_);
  and _17879_ (_09580_, _07071_, _07066_);
  and _17880_ (_09581_, _09580_, _09579_);
  or _17881_ (_09582_, _09581_, _09578_);
  and _17882_ (_09583_, _09582_, _09574_);
  and _17883_ (_09584_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or _17884_ (_09585_, _09584_, _07046_);
  or _17885_ (_09586_, _09585_, _09583_);
  nand _17886_ (_09587_, _07046_, _07040_);
  and _17887_ (_09588_, _09587_, _09586_);
  or _17888_ (_09589_, _09588_, _07050_);
  not _17889_ (_09590_, _07050_);
  or _17890_ (_09591_, _09590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _17891_ (_09592_, _09591_, _06989_);
  and _17892_ (_08330_, _09592_, _09589_);
  or _17893_ (_09593_, _08797_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and _17894_ (_08347_, _09593_, _06989_);
  nor _17895_ (_09594_, _07035_, _06754_);
  not _17896_ (_09595_, _09594_);
  and _17897_ (_09597_, _09595_, _08107_);
  and _17898_ (_09598_, _09597_, _08098_);
  not _17899_ (_09599_, _09598_);
  and _17900_ (_09600_, _09599_, _07485_);
  and _17901_ (_09601_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  or _17902_ (_09602_, _09601_, _09600_);
  and _17903_ (_08521_, _09602_, _06989_);
  not _17904_ (_09603_, _07125_);
  nor _17905_ (_09604_, _08993_, _09603_);
  nor _17906_ (_09605_, _08993_, _07122_);
  nor _17907_ (_09606_, _09604_, _09605_);
  and _17908_ (_09607_, _09606_, _08997_);
  and _17909_ (_09608_, _09607_, _09001_);
  or _17910_ (_09609_, _09608_, _06982_);
  or _17911_ (_09610_, _09609_, _09604_);
  and _17912_ (_09611_, _09610_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _17913_ (_09613_, _09009_, _07485_);
  not _17914_ (_09614_, _09605_);
  nand _17915_ (_09615_, _09614_, _08997_);
  and _17916_ (_09616_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _17917_ (_09618_, _09616_, _09615_);
  or _17918_ (_09619_, _09618_, _09613_);
  or _17919_ (_09621_, _09619_, _09611_);
  and _17920_ (_08660_, _09621_, _06989_);
  and _17921_ (_09623_, _08944_, _08971_);
  not _17922_ (_09625_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _17923_ (_09626_, _08949_, _08583_);
  nor _17924_ (_09627_, _09626_, _08947_);
  and _17925_ (_09629_, _08949_, _08591_);
  and _17926_ (_09630_, _08949_, _08599_);
  nor _17927_ (_09631_, _09630_, _09629_);
  and _17928_ (_09632_, _09631_, _08949_);
  and _17929_ (_09633_, _09632_, _09627_);
  nor _17930_ (_09634_, _09633_, _09625_);
  and _17931_ (_09636_, _08949_, word_in[0]);
  and _17932_ (_09637_, _09636_, _09633_);
  or _17933_ (_09638_, _09637_, _09634_);
  or _17934_ (_09639_, _09638_, _09623_);
  and _17935_ (_09640_, _08937_, _09056_);
  not _17936_ (_09641_, _09640_);
  not _17937_ (_09642_, _09623_);
  or _17938_ (_09643_, _09642_, word_in[8]);
  and _17939_ (_09644_, _09643_, _09641_);
  and _17940_ (_09645_, _09644_, _09639_);
  and _17941_ (_09646_, _08740_, _08932_);
  and _17942_ (_09647_, _08935_, _09646_);
  and _17943_ (_09648_, _08937_, word_in[16]);
  and _17944_ (_09649_, _09648_, _09056_);
  or _17945_ (_09650_, _09649_, _09647_);
  or _17946_ (_09652_, _09650_, _09645_);
  not _17947_ (_09653_, _09647_);
  or _17948_ (_09654_, _09653_, word_in[24]);
  and _17949_ (_14642_, _09654_, _09652_);
  and _17950_ (_09656_, _08935_, word_in[25]);
  and _17951_ (_09657_, _09656_, _09647_);
  not _17952_ (_09658_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _17953_ (_09659_, _09633_, _09658_);
  and _17954_ (_09660_, _08949_, word_in[1]);
  and _17955_ (_09661_, _09660_, _09633_);
  or _17956_ (_09663_, _09661_, _09659_);
  or _17957_ (_09664_, _09663_, _09623_);
  or _17958_ (_09665_, _09642_, word_in[9]);
  and _17959_ (_09666_, _09665_, _09664_);
  or _17960_ (_09667_, _09666_, _09640_);
  nor _17961_ (_09668_, _09641_, word_in[17]);
  nor _17962_ (_09670_, _09668_, _09647_);
  and _17963_ (_09671_, _09670_, _09667_);
  or _17964_ (_14643_, _09671_, _09657_);
  not _17965_ (_09672_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _17966_ (_09673_, _09633_, _09672_);
  and _17967_ (_09674_, _08949_, word_in[2]);
  and _17968_ (_09675_, _09674_, _09633_);
  or _17969_ (_09676_, _09675_, _09673_);
  and _17970_ (_09678_, _09676_, _09642_);
  and _17971_ (_09679_, _09623_, word_in[10]);
  or _17972_ (_09680_, _09679_, _09678_);
  or _17973_ (_09681_, _09680_, _09640_);
  or _17974_ (_09682_, _09641_, word_in[18]);
  and _17975_ (_09683_, _09682_, _09653_);
  and _17976_ (_09684_, _09683_, _09681_);
  and _17977_ (_09685_, _08935_, word_in[26]);
  and _17978_ (_09686_, _09685_, _09647_);
  or _17979_ (_14644_, _09686_, _09684_);
  not _17980_ (_09688_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _17981_ (_09689_, _09633_, _09688_);
  and _17982_ (_09690_, _08949_, word_in[3]);
  and _17983_ (_09692_, _09690_, _09633_);
  or _17984_ (_09693_, _09692_, _09689_);
  or _17985_ (_09694_, _09693_, _09623_);
  or _17986_ (_09695_, _09642_, word_in[11]);
  and _17987_ (_09696_, _09695_, _09694_);
  or _17988_ (_09697_, _09696_, _09640_);
  or _17989_ (_09698_, _09641_, word_in[19]);
  and _17990_ (_09699_, _09698_, _09653_);
  and _17991_ (_09700_, _09699_, _09697_);
  and _17992_ (_09701_, _08935_, word_in[27]);
  and _17993_ (_09702_, _09701_, _09647_);
  or _17994_ (_14645_, _09702_, _09700_);
  and _17995_ (_09703_, _08935_, word_in[28]);
  and _17996_ (_09704_, _09703_, _09647_);
  not _17997_ (_09705_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _17998_ (_09706_, _09633_, _09705_);
  and _17999_ (_09707_, _08949_, word_in[4]);
  and _18000_ (_09708_, _09707_, _09633_);
  or _18001_ (_09709_, _09708_, _09706_);
  and _18002_ (_09710_, _09709_, _09642_);
  and _18003_ (_09712_, _09623_, word_in[12]);
  or _18004_ (_09713_, _09712_, _09710_);
  or _18005_ (_09714_, _09713_, _09640_);
  nor _18006_ (_09715_, _09641_, word_in[20]);
  nor _18007_ (_09716_, _09715_, _09647_);
  and _18008_ (_09717_, _09716_, _09714_);
  or _18009_ (_08749_, _09717_, _09704_);
  and _18010_ (_09718_, _08935_, word_in[29]);
  and _18011_ (_09719_, _09718_, _09647_);
  not _18012_ (_09720_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _18013_ (_09721_, _09633_, _09720_);
  and _18014_ (_09722_, _08949_, word_in[5]);
  and _18015_ (_09723_, _09722_, _09633_);
  or _18016_ (_09724_, _09723_, _09721_);
  or _18017_ (_09725_, _09724_, _09623_);
  or _18018_ (_09726_, _09642_, word_in[13]);
  and _18019_ (_09727_, _09726_, _09725_);
  or _18020_ (_09728_, _09727_, _09640_);
  nor _18021_ (_09729_, _09641_, word_in[21]);
  nor _18022_ (_09730_, _09729_, _09647_);
  and _18023_ (_09731_, _09730_, _09728_);
  or _18024_ (_14646_, _09731_, _09719_);
  not _18025_ (_09732_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _18026_ (_09734_, _09633_, _09732_);
  and _18027_ (_09735_, _08949_, word_in[6]);
  and _18028_ (_09736_, _09735_, _09633_);
  or _18029_ (_09737_, _09736_, _09734_);
  or _18030_ (_09738_, _09737_, _09623_);
  or _18031_ (_09739_, _09642_, word_in[14]);
  and _18032_ (_09740_, _09739_, _09738_);
  or _18033_ (_09741_, _09740_, _09640_);
  nor _18034_ (_09742_, _09641_, word_in[22]);
  nor _18035_ (_09743_, _09742_, _09647_);
  and _18036_ (_09744_, _09743_, _09741_);
  and _18037_ (_09745_, _08935_, word_in[30]);
  and _18038_ (_09746_, _09745_, _09647_);
  or _18039_ (_14647_, _09746_, _09744_);
  nor _18040_ (_09748_, _09633_, _08777_);
  and _18041_ (_09749_, _09633_, _08953_);
  or _18042_ (_09750_, _09749_, _09748_);
  and _18043_ (_09751_, _09750_, _09642_);
  and _18044_ (_09752_, _09623_, word_in[15]);
  or _18045_ (_09753_, _09752_, _09751_);
  or _18046_ (_09754_, _09753_, _09640_);
  or _18047_ (_09755_, _09641_, word_in[23]);
  and _18048_ (_09756_, _09755_, _09653_);
  and _18049_ (_09757_, _09756_, _09754_);
  and _18050_ (_09758_, _09647_, word_in[31]);
  or _18051_ (_14648_, _09758_, _09757_);
  nor _18052_ (_09759_, _09404_, _09395_);
  or _18053_ (_09760_, _09759_, _09389_);
  and _18054_ (_09761_, _09760_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and _18055_ (_09762_, _09395_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _18056_ (_09763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _18057_ (_09764_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor _18058_ (_09765_, _09764_, _09763_);
  and _18059_ (_09766_, _09765_, _09762_);
  or _18060_ (_09767_, _09766_, _09761_);
  and _18061_ (_08809_, _09767_, _06989_);
  and _18062_ (_09768_, _08944_, _08731_);
  and _18063_ (_09769_, _09768_, _08724_);
  not _18064_ (_09770_, _09769_);
  not _18065_ (_09771_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _18066_ (_09772_, _08947_, _08584_);
  and _18067_ (_09773_, _09772_, _09631_);
  nor _18068_ (_09774_, _09773_, _09771_);
  and _18069_ (_09775_, _09773_, _09636_);
  or _18070_ (_09776_, _09775_, _09774_);
  and _18071_ (_09777_, _09776_, _09770_);
  and _18072_ (_09778_, _08937_, _08713_);
  and _18073_ (_09780_, _09778_, _08824_);
  and _18074_ (_09781_, _09769_, word_in[8]);
  or _18075_ (_09782_, _09781_, _09780_);
  or _18076_ (_09783_, _09782_, _09777_);
  and _18077_ (_09784_, _08935_, _09056_);
  not _18078_ (_09785_, _09784_);
  not _18079_ (_09786_, _09780_);
  or _18080_ (_09787_, _09786_, _09648_);
  and _18081_ (_09788_, _09787_, _09785_);
  and _18082_ (_09789_, _09788_, _09783_);
  and _18083_ (_09790_, _09784_, word_in[24]);
  or _18084_ (_08840_, _09790_, _09789_);
  not _18085_ (_09792_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _18086_ (_09793_, _09773_, _09792_);
  and _18087_ (_09794_, _09773_, _09660_);
  or _18088_ (_09796_, _09794_, _09793_);
  and _18089_ (_09797_, _09796_, _09770_);
  and _18090_ (_09798_, _09769_, word_in[9]);
  or _18091_ (_09799_, _09798_, _09780_);
  or _18092_ (_09800_, _09799_, _09797_);
  and _18093_ (_09801_, _08937_, word_in[17]);
  or _18094_ (_09802_, _09786_, _09801_);
  and _18095_ (_09803_, _09802_, _09785_);
  and _18096_ (_09805_, _09803_, _09800_);
  and _18097_ (_09806_, _09784_, word_in[25]);
  or _18098_ (_14666_, _09806_, _09805_);
  not _18099_ (_09807_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _18100_ (_09808_, _09773_, _09807_);
  and _18101_ (_09809_, _09773_, _09674_);
  or _18102_ (_09810_, _09809_, _09808_);
  and _18103_ (_09811_, _09810_, _09770_);
  and _18104_ (_09813_, _09769_, word_in[10]);
  or _18105_ (_09814_, _09813_, _09780_);
  or _18106_ (_09815_, _09814_, _09811_);
  and _18107_ (_09816_, _08937_, word_in[18]);
  or _18108_ (_09817_, _09786_, _09816_);
  and _18109_ (_09818_, _09817_, _09785_);
  and _18110_ (_09819_, _09818_, _09815_);
  and _18111_ (_09820_, _09784_, word_in[26]);
  or _18112_ (_14667_, _09820_, _09819_);
  not _18113_ (_09821_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _18114_ (_09822_, _09773_, _09821_);
  and _18115_ (_09823_, _09773_, _09690_);
  or _18116_ (_09824_, _09823_, _09822_);
  and _18117_ (_09825_, _09824_, _09770_);
  and _18118_ (_09826_, _09769_, word_in[11]);
  or _18119_ (_09827_, _09826_, _09780_);
  or _18120_ (_09828_, _09827_, _09825_);
  and _18121_ (_09829_, _08937_, word_in[19]);
  or _18122_ (_09830_, _09786_, _09829_);
  and _18123_ (_09831_, _09830_, _09785_);
  and _18124_ (_09832_, _09831_, _09828_);
  and _18125_ (_09833_, _09784_, word_in[27]);
  or _18126_ (_14668_, _09833_, _09832_);
  not _18127_ (_09834_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor _18128_ (_09835_, _09773_, _09834_);
  and _18129_ (_09836_, _09773_, _09707_);
  or _18130_ (_09837_, _09836_, _09835_);
  and _18131_ (_09838_, _09837_, _09770_);
  and _18132_ (_09839_, _09769_, word_in[12]);
  or _18133_ (_09840_, _09839_, _09780_);
  or _18134_ (_09841_, _09840_, _09838_);
  and _18135_ (_09842_, _08937_, word_in[20]);
  or _18136_ (_09843_, _09786_, _09842_);
  and _18137_ (_09844_, _09843_, _09785_);
  and _18138_ (_09845_, _09844_, _09841_);
  and _18139_ (_09846_, _09784_, word_in[28]);
  or _18140_ (_14669_, _09846_, _09845_);
  not _18141_ (_09847_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor _18142_ (_09848_, _09773_, _09847_);
  and _18143_ (_09849_, _09773_, _09722_);
  or _18144_ (_09850_, _09849_, _09848_);
  and _18145_ (_09851_, _09850_, _09770_);
  and _18146_ (_09852_, _09769_, word_in[13]);
  or _18147_ (_09853_, _09852_, _09780_);
  or _18148_ (_09854_, _09853_, _09851_);
  and _18149_ (_09855_, _08937_, word_in[21]);
  or _18150_ (_09856_, _09786_, _09855_);
  and _18151_ (_09857_, _09856_, _09785_);
  and _18152_ (_09858_, _09857_, _09854_);
  and _18153_ (_09859_, _09784_, word_in[29]);
  or _18154_ (_14670_, _09859_, _09858_);
  not _18155_ (_09860_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor _18156_ (_09861_, _09773_, _09860_);
  and _18157_ (_09862_, _09773_, _09735_);
  or _18158_ (_09863_, _09862_, _09861_);
  and _18159_ (_09865_, _09863_, _09770_);
  and _18160_ (_09866_, _09769_, word_in[14]);
  or _18161_ (_09868_, _09866_, _09780_);
  or _18162_ (_09870_, _09868_, _09865_);
  and _18163_ (_09871_, _08937_, word_in[22]);
  or _18164_ (_09872_, _09786_, _09871_);
  and _18165_ (_09873_, _09872_, _09785_);
  and _18166_ (_09875_, _09873_, _09870_);
  and _18167_ (_09876_, _09784_, word_in[30]);
  or _18168_ (_14671_, _09876_, _09875_);
  nor _18169_ (_09878_, _09773_, _08698_);
  and _18170_ (_09879_, _09773_, _08953_);
  or _18171_ (_09881_, _09879_, _09878_);
  and _18172_ (_09882_, _09881_, _09770_);
  and _18173_ (_09883_, _09769_, word_in[15]);
  or _18174_ (_09884_, _09883_, _09780_);
  or _18175_ (_09886_, _09884_, _09882_);
  or _18176_ (_09887_, _09786_, _08942_);
  and _18177_ (_09888_, _09887_, _09785_);
  and _18178_ (_09889_, _09888_, _09886_);
  and _18179_ (_09890_, _09784_, word_in[31]);
  or _18180_ (_14672_, _09890_, _09889_);
  and _18181_ (_09891_, _08935_, _08713_);
  and _18182_ (_09892_, _09891_, _08885_);
  and _18183_ (_09893_, _08937_, _08731_);
  and _18184_ (_09894_, _09893_, _08824_);
  not _18185_ (_09895_, _09894_);
  or _18186_ (_09896_, _09895_, _09648_);
  and _18187_ (_09897_, _08944_, _08740_);
  and _18188_ (_09898_, _09897_, _08724_);
  not _18189_ (_09899_, _09898_);
  not _18190_ (_09900_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  not _18191_ (_09901_, _08947_);
  and _18192_ (_09902_, _09626_, _09901_);
  and _18193_ (_09903_, _09902_, _09631_);
  nor _18194_ (_09904_, _09903_, _09900_);
  and _18195_ (_09905_, _09903_, _09636_);
  or _18196_ (_09906_, _09905_, _09904_);
  and _18197_ (_09907_, _09906_, _09899_);
  and _18198_ (_09908_, _09898_, word_in[8]);
  or _18199_ (_09909_, _09908_, _09894_);
  or _18200_ (_09910_, _09909_, _09907_);
  and _18201_ (_09911_, _09910_, _09896_);
  or _18202_ (_09912_, _09911_, _09892_);
  not _18203_ (_09913_, _09892_);
  or _18204_ (_09914_, _09913_, word_in[24]);
  and _18205_ (_14673_, _09914_, _09912_);
  or _18206_ (_09915_, _09895_, _09801_);
  not _18207_ (_09916_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor _18208_ (_09917_, _09903_, _09916_);
  and _18209_ (_09918_, _09903_, _09660_);
  or _18210_ (_09920_, _09918_, _09917_);
  and _18211_ (_09921_, _09920_, _09899_);
  and _18212_ (_09923_, _09898_, word_in[9]);
  or _18213_ (_09924_, _09923_, _09894_);
  or _18214_ (_09925_, _09924_, _09921_);
  and _18215_ (_09926_, _09925_, _09915_);
  or _18216_ (_09927_, _09926_, _09892_);
  or _18217_ (_09928_, _09913_, word_in[25]);
  and _18218_ (_14674_, _09928_, _09927_);
  or _18219_ (_09930_, _09895_, _09816_);
  not _18220_ (_09931_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor _18221_ (_09932_, _09903_, _09931_);
  and _18222_ (_09933_, _09903_, _09674_);
  or _18223_ (_09934_, _09933_, _09932_);
  and _18224_ (_09935_, _09934_, _09899_);
  and _18225_ (_09937_, _09898_, word_in[10]);
  or _18226_ (_09938_, _09937_, _09894_);
  or _18227_ (_09939_, _09938_, _09935_);
  and _18228_ (_09940_, _09939_, _09930_);
  or _18229_ (_09941_, _09940_, _09892_);
  or _18230_ (_09942_, _09913_, word_in[26]);
  and _18231_ (_14675_, _09942_, _09941_);
  or _18232_ (_09943_, _09895_, _09829_);
  not _18233_ (_09944_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor _18234_ (_09945_, _09903_, _09944_);
  and _18235_ (_09946_, _09903_, _09690_);
  or _18236_ (_09947_, _09946_, _09945_);
  and _18237_ (_09948_, _09947_, _09899_);
  and _18238_ (_09949_, _09898_, word_in[11]);
  or _18239_ (_09950_, _09949_, _09894_);
  or _18240_ (_09951_, _09950_, _09948_);
  and _18241_ (_09952_, _09951_, _09943_);
  or _18242_ (_09953_, _09952_, _09892_);
  or _18243_ (_09954_, _09913_, word_in[27]);
  and _18244_ (_14676_, _09954_, _09953_);
  or _18245_ (_09955_, _09895_, _09842_);
  not _18246_ (_09957_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor _18247_ (_09958_, _09903_, _09957_);
  and _18248_ (_09959_, _09903_, _09707_);
  or _18249_ (_09960_, _09959_, _09958_);
  and _18250_ (_09962_, _09960_, _09899_);
  and _18251_ (_09964_, _09898_, word_in[12]);
  or _18252_ (_09965_, _09964_, _09894_);
  or _18253_ (_09966_, _09965_, _09962_);
  and _18254_ (_09968_, _09966_, _09955_);
  or _18255_ (_09969_, _09968_, _09892_);
  or _18256_ (_09970_, _09913_, word_in[28]);
  and _18257_ (_14677_, _09970_, _09969_);
  or _18258_ (_09972_, _09895_, _09855_);
  not _18259_ (_09974_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _18260_ (_09975_, _09903_, _09974_);
  and _18261_ (_09977_, _09903_, _09722_);
  or _18262_ (_09979_, _09977_, _09975_);
  and _18263_ (_09980_, _09979_, _09899_);
  and _18264_ (_09981_, _09898_, word_in[13]);
  or _18265_ (_09982_, _09981_, _09894_);
  or _18266_ (_09983_, _09982_, _09980_);
  and _18267_ (_09984_, _09983_, _09972_);
  and _18268_ (_09985_, _09984_, _09913_);
  and _18269_ (_09986_, _09892_, word_in[29]);
  or _18270_ (_08962_, _09986_, _09985_);
  or _18271_ (_09987_, _09895_, _09871_);
  not _18272_ (_09988_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _18273_ (_09989_, _09903_, _09988_);
  and _18274_ (_09990_, _09903_, _09735_);
  or _18275_ (_09991_, _09990_, _09989_);
  and _18276_ (_09992_, _09991_, _09899_);
  and _18277_ (_09993_, _09898_, word_in[14]);
  or _18278_ (_09994_, _09993_, _09894_);
  or _18279_ (_09995_, _09994_, _09992_);
  and _18280_ (_09996_, _09995_, _09987_);
  and _18281_ (_09997_, _09996_, _09913_);
  and _18282_ (_09998_, _09892_, word_in[30]);
  or _18283_ (_14678_, _09998_, _09997_);
  or _18284_ (_10000_, _09895_, _08942_);
  nor _18285_ (_10001_, _09903_, _08772_);
  and _18286_ (_10002_, _09903_, _08953_);
  or _18287_ (_10003_, _10002_, _10001_);
  and _18288_ (_10004_, _10003_, _09899_);
  and _18289_ (_10005_, _09898_, word_in[15]);
  or _18290_ (_10006_, _10005_, _09894_);
  or _18291_ (_10007_, _10006_, _10004_);
  and _18292_ (_10008_, _10007_, _10000_);
  and _18293_ (_10009_, _10008_, _09913_);
  and _18294_ (_10010_, _09892_, word_in[31]);
  or _18295_ (_14679_, _10010_, _10009_);
  and _18296_ (_10011_, _08935_, _08731_);
  and _18297_ (_10012_, _10011_, _08885_);
  not _18298_ (_10013_, _10012_);
  and _18299_ (_10014_, _08945_, _08724_);
  not _18300_ (_10015_, _10014_);
  not _18301_ (_10016_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _18302_ (_10017_, _09631_, _08948_);
  nor _18303_ (_10018_, _10017_, _10016_);
  and _18304_ (_10019_, _10017_, _09636_);
  or _18305_ (_10021_, _10019_, _10018_);
  and _18306_ (_10022_, _10021_, _10015_);
  and _18307_ (_10023_, _08937_, _08740_);
  and _18308_ (_10024_, _10023_, _08824_);
  and _18309_ (_10026_, _10014_, word_in[8]);
  or _18310_ (_10027_, _10026_, _10024_);
  or _18311_ (_10028_, _10027_, _10022_);
  not _18312_ (_10030_, _10024_);
  or _18313_ (_10031_, _10030_, _09648_);
  and _18314_ (_10032_, _10031_, _10028_);
  and _18315_ (_10034_, _10032_, _10013_);
  and _18316_ (_10035_, _10012_, word_in[24]);
  or _18317_ (_14680_, _10035_, _10034_);
  not _18318_ (_10037_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor _18319_ (_10038_, _10017_, _10037_);
  and _18320_ (_10039_, _10017_, _09660_);
  or _18321_ (_10040_, _10039_, _10038_);
  and _18322_ (_10041_, _10040_, _10015_);
  and _18323_ (_10043_, _10014_, word_in[9]);
  or _18324_ (_10044_, _10043_, _10024_);
  or _18325_ (_10046_, _10044_, _10041_);
  or _18326_ (_10048_, _10030_, _09801_);
  and _18327_ (_10050_, _10048_, _10046_);
  or _18328_ (_10052_, _10050_, _10012_);
  or _18329_ (_10054_, _10013_, word_in[25]);
  and _18330_ (_14681_, _10054_, _10052_);
  not _18331_ (_10057_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor _18332_ (_10059_, _10017_, _10057_);
  and _18333_ (_10060_, _10017_, _09674_);
  or _18334_ (_10061_, _10060_, _10059_);
  and _18335_ (_10063_, _10061_, _10015_);
  and _18336_ (_10064_, _10014_, word_in[10]);
  or _18337_ (_10065_, _10064_, _10024_);
  or _18338_ (_10066_, _10065_, _10063_);
  or _18339_ (_10067_, _10030_, _09816_);
  and _18340_ (_10068_, _10067_, _10066_);
  or _18341_ (_10069_, _10068_, _10012_);
  or _18342_ (_10070_, _10013_, word_in[26]);
  and _18343_ (_14682_, _10070_, _10069_);
  and _18344_ (_10071_, _10017_, _09690_);
  not _18345_ (_10072_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor _18346_ (_10073_, _10017_, _10072_);
  or _18347_ (_10075_, _10073_, _10071_);
  and _18348_ (_10076_, _10075_, _10015_);
  and _18349_ (_10077_, _10014_, word_in[11]);
  or _18350_ (_10078_, _10077_, _10024_);
  or _18351_ (_10080_, _10078_, _10076_);
  or _18352_ (_10081_, _10030_, _09829_);
  and _18353_ (_10082_, _10081_, _10080_);
  and _18354_ (_10083_, _10082_, _10013_);
  and _18355_ (_10084_, _10012_, word_in[27]);
  or _18356_ (_14683_, _10084_, _10083_);
  and _18357_ (_10085_, _10017_, _09707_);
  not _18358_ (_10086_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _18359_ (_10087_, _10017_, _10086_);
  or _18360_ (_10088_, _10087_, _10085_);
  and _18361_ (_10089_, _10088_, _10015_);
  and _18362_ (_10090_, _10014_, word_in[12]);
  or _18363_ (_10091_, _10090_, _10024_);
  or _18364_ (_10093_, _10091_, _10089_);
  or _18365_ (_10094_, _10030_, _09842_);
  and _18366_ (_10095_, _10094_, _10093_);
  and _18367_ (_10096_, _10095_, _10013_);
  and _18368_ (_10097_, _10012_, word_in[28]);
  or _18369_ (_14684_, _10097_, _10096_);
  or _18370_ (_10099_, _10030_, _09855_);
  not _18371_ (_10100_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor _18372_ (_10102_, _10017_, _10100_);
  and _18373_ (_10103_, _10017_, _09722_);
  or _18374_ (_10104_, _10103_, _10102_);
  and _18375_ (_10105_, _10104_, _10015_);
  and _18376_ (_10106_, _10014_, word_in[13]);
  or _18377_ (_10107_, _10106_, _10024_);
  or _18378_ (_10108_, _10107_, _10105_);
  and _18379_ (_10109_, _10108_, _10099_);
  or _18380_ (_10110_, _10109_, _10012_);
  or _18381_ (_10111_, _10013_, word_in[29]);
  and _18382_ (_14685_, _10111_, _10110_);
  not _18383_ (_10113_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor _18384_ (_10115_, _10017_, _10113_);
  and _18385_ (_10116_, _10017_, _09735_);
  or _18386_ (_10117_, _10116_, _10115_);
  and _18387_ (_10118_, _10117_, _10015_);
  and _18388_ (_10119_, _10014_, word_in[14]);
  or _18389_ (_10120_, _10119_, _10024_);
  or _18390_ (_10121_, _10120_, _10118_);
  or _18391_ (_10122_, _10030_, _09871_);
  and _18392_ (_10123_, _10122_, _10121_);
  and _18393_ (_10124_, _10123_, _10013_);
  and _18394_ (_10125_, _10012_, word_in[30]);
  or _18395_ (_14686_, _10125_, _10124_);
  and _18396_ (_10127_, _10017_, _08953_);
  nor _18397_ (_10128_, _10017_, _08682_);
  or _18398_ (_10130_, _10128_, _10127_);
  and _18399_ (_10132_, _10130_, _10015_);
  and _18400_ (_10134_, _10014_, word_in[15]);
  or _18401_ (_10136_, _10134_, _10024_);
  or _18402_ (_10138_, _10136_, _10132_);
  or _18403_ (_10140_, _10030_, _08942_);
  and _18404_ (_10141_, _10140_, _10138_);
  and _18405_ (_10143_, _10141_, _10013_);
  and _18406_ (_10145_, _10012_, word_in[31]);
  or _18407_ (_09047_, _10145_, _10143_);
  and _18408_ (_10146_, _09604_, _06981_);
  nand _18409_ (_10147_, _10146_, _07118_);
  or _18410_ (_10148_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and _18411_ (_10149_, _10148_, _06989_);
  and _18412_ (_09122_, _10149_, _10147_);
  and _18413_ (_10150_, _08935_, _08874_);
  and _18414_ (_10151_, _10150_, _08879_);
  and _18415_ (_10152_, _10151_, _08740_);
  and _18416_ (_10153_, _08938_, _08860_);
  and _18417_ (_10154_, _10153_, _08711_);
  not _18418_ (_10155_, _10154_);
  or _18419_ (_10156_, _10155_, _09648_);
  and _18420_ (_10157_, _08944_, _08981_);
  not _18421_ (_10158_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _18422_ (_10159_, _08949_, _08721_);
  and _18423_ (_10160_, _10159_, _09627_);
  nor _18424_ (_10161_, _10160_, _10158_);
  and _18425_ (_10162_, _10160_, _09636_);
  or _18426_ (_10163_, _10162_, _10161_);
  or _18427_ (_10164_, _10163_, _10157_);
  not _18428_ (_10165_, _10157_);
  or _18429_ (_10166_, _10165_, word_in[8]);
  and _18430_ (_10167_, _10166_, _10164_);
  or _18431_ (_10168_, _10167_, _10154_);
  and _18432_ (_10169_, _10168_, _10156_);
  or _18433_ (_10170_, _10169_, _10152_);
  and _18434_ (_10171_, _08935_, word_in[24]);
  not _18435_ (_10172_, _10152_);
  or _18436_ (_10173_, _10172_, _10171_);
  and _18437_ (_09135_, _10173_, _10170_);
  or _18438_ (_10174_, _10155_, _09801_);
  not _18439_ (_10175_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _18440_ (_10176_, _10160_, _10175_);
  and _18441_ (_10177_, _10160_, _09660_);
  or _18442_ (_10178_, _10177_, _10176_);
  or _18443_ (_10179_, _10178_, _10157_);
  or _18444_ (_10180_, _10165_, word_in[9]);
  and _18445_ (_10181_, _10180_, _10179_);
  or _18446_ (_10182_, _10181_, _10154_);
  and _18447_ (_10183_, _10182_, _10174_);
  or _18448_ (_10184_, _10183_, _10152_);
  or _18449_ (_10185_, _10172_, _09656_);
  and _18450_ (_09137_, _10185_, _10184_);
  or _18451_ (_10186_, _10155_, _09816_);
  not _18452_ (_10187_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _18453_ (_10188_, _10160_, _10187_);
  and _18454_ (_10189_, _10160_, _09674_);
  or _18455_ (_10190_, _10189_, _10188_);
  or _18456_ (_10191_, _10190_, _10157_);
  or _18457_ (_10192_, _10165_, word_in[10]);
  and _18458_ (_10193_, _10192_, _10191_);
  or _18459_ (_10194_, _10193_, _10154_);
  and _18460_ (_10195_, _10194_, _10186_);
  or _18461_ (_10196_, _10195_, _10152_);
  or _18462_ (_10197_, _10172_, _09685_);
  and _18463_ (_09141_, _10197_, _10196_);
  or _18464_ (_10198_, _10155_, _09829_);
  not _18465_ (_10199_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _18466_ (_10200_, _10160_, _10199_);
  and _18467_ (_10201_, _10160_, _09690_);
  or _18468_ (_10202_, _10201_, _10200_);
  or _18469_ (_10203_, _10202_, _10157_);
  or _18470_ (_10204_, _10165_, word_in[11]);
  and _18471_ (_10205_, _10204_, _10203_);
  or _18472_ (_10206_, _10205_, _10154_);
  and _18473_ (_10207_, _10206_, _10198_);
  or _18474_ (_10208_, _10207_, _10152_);
  or _18475_ (_10209_, _10172_, _09701_);
  and _18476_ (_14687_, _10209_, _10208_);
  and _18477_ (_10210_, _10154_, _09842_);
  and _18478_ (_10211_, _10160_, word_in[4]);
  not _18479_ (_10212_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _18480_ (_10213_, _10160_, _10212_);
  or _18481_ (_10214_, _10213_, _10211_);
  and _18482_ (_10215_, _10214_, _10165_);
  and _18483_ (_10216_, _10157_, word_in[12]);
  or _18484_ (_10217_, _10216_, _10215_);
  and _18485_ (_10218_, _10217_, _10155_);
  or _18486_ (_10219_, _10218_, _10210_);
  and _18487_ (_10220_, _10219_, _10172_);
  and _18488_ (_10221_, _10152_, _09703_);
  or _18489_ (_14688_, _10221_, _10220_);
  or _18490_ (_10222_, _10155_, _09855_);
  not _18491_ (_10223_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _18492_ (_10224_, _10160_, _10223_);
  and _18493_ (_10225_, _10160_, _09722_);
  or _18494_ (_10226_, _10225_, _10224_);
  or _18495_ (_10227_, _10226_, _10157_);
  or _18496_ (_10228_, _10165_, word_in[13]);
  and _18497_ (_10229_, _10228_, _10227_);
  or _18498_ (_10230_, _10229_, _10154_);
  and _18499_ (_10231_, _10230_, _10222_);
  or _18500_ (_10232_, _10231_, _10152_);
  or _18501_ (_10233_, _10172_, _09718_);
  and _18502_ (_14689_, _10233_, _10232_);
  and _18503_ (_10234_, _10160_, word_in[6]);
  not _18504_ (_10235_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _18505_ (_10236_, _10160_, _10235_);
  or _18506_ (_10237_, _10236_, _10234_);
  or _18507_ (_10238_, _10237_, _10157_);
  or _18508_ (_10239_, _10165_, word_in[14]);
  and _18509_ (_10240_, _10239_, _10155_);
  and _18510_ (_10241_, _10240_, _10238_);
  and _18511_ (_10242_, _10154_, _09871_);
  or _18512_ (_10243_, _10242_, _10152_);
  or _18513_ (_10244_, _10243_, _10241_);
  or _18514_ (_10245_, _10172_, _09745_);
  and _18515_ (_09152_, _10245_, _10244_);
  and _18516_ (_10246_, _10154_, _08942_);
  and _18517_ (_10247_, _10160_, word_in[7]);
  nor _18518_ (_10248_, _10160_, _08790_);
  or _18519_ (_10249_, _10248_, _10247_);
  and _18520_ (_10250_, _10249_, _10165_);
  and _18521_ (_10251_, _10157_, word_in[15]);
  or _18522_ (_10252_, _10251_, _10250_);
  and _18523_ (_10253_, _10252_, _10155_);
  or _18524_ (_10254_, _10253_, _10246_);
  and _18525_ (_10255_, _10254_, _10172_);
  and _18526_ (_10256_, _08935_, word_in[31]);
  and _18527_ (_10257_, _10152_, _10256_);
  or _18528_ (_09154_, _10257_, _10255_);
  and _18529_ (_10258_, _10153_, _08713_);
  not _18530_ (_10259_, _10258_);
  and _18531_ (_10260_, _09768_, _08784_);
  and _18532_ (_10261_, _10159_, _09772_);
  and _18533_ (_10262_, _10261_, _09636_);
  not _18534_ (_10263_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _18535_ (_10264_, _10261_, _10263_);
  nor _18536_ (_10265_, _10264_, _10262_);
  nor _18537_ (_10266_, _10265_, _10260_);
  and _18538_ (_10267_, _10260_, word_in[8]);
  or _18539_ (_10268_, _10267_, _10266_);
  and _18540_ (_10269_, _10268_, _10259_);
  and _18541_ (_10270_, _10151_, _08711_);
  and _18542_ (_10271_, _10258_, _09648_);
  or _18543_ (_10272_, _10271_, _10270_);
  or _18544_ (_10273_, _10272_, _10269_);
  not _18545_ (_10274_, _10270_);
  or _18546_ (_10275_, _10274_, word_in[24]);
  and _18547_ (_09235_, _10275_, _10273_);
  not _18548_ (_10276_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _18549_ (_10277_, _10261_, _10276_);
  and _18550_ (_10278_, _10261_, _09660_);
  nor _18551_ (_10279_, _10278_, _10277_);
  nor _18552_ (_10280_, _10279_, _10260_);
  and _18553_ (_10281_, _10260_, word_in[9]);
  or _18554_ (_10282_, _10281_, _10280_);
  and _18555_ (_10283_, _10282_, _10259_);
  and _18556_ (_10284_, _10258_, _09801_);
  or _18557_ (_10285_, _10284_, _10270_);
  or _18558_ (_10286_, _10285_, _10283_);
  or _18559_ (_10287_, _10274_, word_in[25]);
  and _18560_ (_09238_, _10287_, _10286_);
  not _18561_ (_10288_, _10260_);
  or _18562_ (_10289_, _10288_, word_in[10]);
  not _18563_ (_10290_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _18564_ (_10291_, _10261_, _10290_);
  and _18565_ (_10292_, _10261_, _09674_);
  or _18566_ (_10293_, _10292_, _10291_);
  or _18567_ (_10294_, _10293_, _10260_);
  and _18568_ (_10295_, _10294_, _10259_);
  and _18569_ (_10296_, _10295_, _10289_);
  and _18570_ (_10297_, _10258_, _09816_);
  or _18571_ (_10298_, _10297_, _10270_);
  or _18572_ (_10299_, _10298_, _10296_);
  or _18573_ (_10300_, _10274_, word_in[26]);
  and _18574_ (_14690_, _10300_, _10299_);
  not _18575_ (_10301_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _18576_ (_10302_, _10261_, _10301_);
  and _18577_ (_10303_, _10261_, _09690_);
  or _18578_ (_10304_, _10303_, _10302_);
  or _18579_ (_10305_, _10304_, _10260_);
  or _18580_ (_10306_, _10288_, word_in[11]);
  and _18581_ (_10307_, _10306_, _10305_);
  or _18582_ (_10308_, _10307_, _10258_);
  or _18583_ (_10309_, _10259_, _09829_);
  and _18584_ (_10310_, _10309_, _10308_);
  or _18585_ (_10311_, _10310_, _10270_);
  or _18586_ (_10312_, _10274_, word_in[27]);
  and _18587_ (_09243_, _10312_, _10311_);
  and _18588_ (_10313_, _10258_, _09842_);
  and _18589_ (_10314_, _10261_, _09707_);
  not _18590_ (_10315_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _18591_ (_10316_, _10261_, _10315_);
  nor _18592_ (_10317_, _10316_, _10314_);
  nor _18593_ (_10318_, _10317_, _10260_);
  and _18594_ (_10319_, _10260_, word_in[12]);
  or _18595_ (_10320_, _10319_, _10318_);
  and _18596_ (_10321_, _10320_, _10259_);
  or _18597_ (_10322_, _10321_, _10313_);
  and _18598_ (_10323_, _10322_, _10274_);
  and _18599_ (_10324_, _10270_, word_in[28]);
  or _18600_ (_09247_, _10324_, _10323_);
  not _18601_ (_10325_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _18602_ (_10326_, _10261_, _10325_);
  and _18603_ (_10327_, _10261_, _09722_);
  or _18604_ (_10328_, _10327_, _10326_);
  or _18605_ (_10329_, _10328_, _10260_);
  or _18606_ (_10330_, _10288_, word_in[13]);
  and _18607_ (_10331_, _10330_, _10329_);
  or _18608_ (_10332_, _10331_, _10258_);
  or _18609_ (_10333_, _10259_, _09855_);
  and _18610_ (_10334_, _10333_, _10332_);
  or _18611_ (_10335_, _10334_, _10270_);
  or _18612_ (_10336_, _10274_, word_in[29]);
  and _18613_ (_09251_, _10336_, _10335_);
  or _18614_ (_10337_, _10288_, word_in[14]);
  not _18615_ (_10338_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _18616_ (_10339_, _10261_, _10338_);
  and _18617_ (_10340_, _10261_, _09735_);
  or _18618_ (_10341_, _10340_, _10339_);
  or _18619_ (_10342_, _10341_, _10260_);
  and _18620_ (_10343_, _10342_, _10259_);
  and _18621_ (_10344_, _10343_, _10337_);
  and _18622_ (_10345_, _10258_, _09871_);
  or _18623_ (_10346_, _10345_, _10270_);
  or _18624_ (_10347_, _10346_, _10344_);
  or _18625_ (_10348_, _10274_, word_in[30]);
  and _18626_ (_09254_, _10348_, _10347_);
  nor _18627_ (_10349_, _10261_, _08693_);
  and _18628_ (_10350_, _10261_, _08953_);
  or _18629_ (_10351_, _10350_, _10349_);
  or _18630_ (_10352_, _10351_, _10260_);
  or _18631_ (_10353_, _10288_, word_in[15]);
  and _18632_ (_10354_, _10353_, _10352_);
  or _18633_ (_10355_, _10354_, _10258_);
  or _18634_ (_10356_, _10259_, _08942_);
  and _18635_ (_10357_, _10356_, _10355_);
  or _18636_ (_10358_, _10357_, _10270_);
  or _18637_ (_10359_, _10274_, word_in[31]);
  and _18638_ (_09257_, _10359_, _10358_);
  nand _18639_ (_10360_, _10146_, _07317_);
  or _18640_ (_10361_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and _18641_ (_10362_, _10361_, _06989_);
  and _18642_ (_09305_, _10362_, _10360_);
  and _18643_ (_10363_, _10151_, _08713_);
  and _18644_ (_10364_, _10153_, _08731_);
  not _18645_ (_10365_, _10364_);
  or _18646_ (_10366_, _10365_, _09648_);
  and _18647_ (_10367_, _09897_, _08784_);
  not _18648_ (_10368_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _18649_ (_10369_, _09902_, _08721_);
  nor _18650_ (_10370_, _10369_, _10368_);
  and _18651_ (_10371_, _10369_, _09636_);
  or _18652_ (_10372_, _10371_, _10370_);
  or _18653_ (_10373_, _10372_, _10367_);
  not _18654_ (_10374_, _10367_);
  or _18655_ (_10375_, _10374_, word_in[8]);
  and _18656_ (_10376_, _10375_, _10373_);
  or _18657_ (_10377_, _10376_, _10364_);
  and _18658_ (_10378_, _10377_, _10366_);
  or _18659_ (_10379_, _10378_, _10363_);
  not _18660_ (_10380_, _10363_);
  or _18661_ (_10381_, _10380_, word_in[24]);
  and _18662_ (_09328_, _10381_, _10379_);
  not _18663_ (_10382_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor _18664_ (_10383_, _10369_, _10382_);
  and _18665_ (_10384_, _10369_, _09660_);
  or _18666_ (_10385_, _10384_, _10383_);
  and _18667_ (_10386_, _10385_, _10374_);
  and _18668_ (_10387_, _10367_, word_in[9]);
  or _18669_ (_10388_, _10387_, _10364_);
  or _18670_ (_10389_, _10388_, _10386_);
  or _18671_ (_10390_, _10365_, _09801_);
  and _18672_ (_10391_, _10390_, _10389_);
  or _18673_ (_10392_, _10391_, _10363_);
  or _18674_ (_10393_, _10380_, word_in[25]);
  and _18675_ (_14691_, _10393_, _10392_);
  or _18676_ (_10394_, _10365_, _09816_);
  not _18677_ (_10395_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor _18678_ (_10396_, _10369_, _10395_);
  and _18679_ (_10397_, _10369_, _09674_);
  or _18680_ (_10398_, _10397_, _10396_);
  and _18681_ (_10399_, _10398_, _10374_);
  and _18682_ (_10401_, _10367_, word_in[10]);
  or _18683_ (_10402_, _10401_, _10364_);
  or _18684_ (_10403_, _10402_, _10399_);
  and _18685_ (_10404_, _10403_, _10394_);
  or _18686_ (_10405_, _10404_, _10363_);
  or _18687_ (_10406_, _10380_, word_in[26]);
  and _18688_ (_09335_, _10406_, _10405_);
  not _18689_ (_10407_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor _18690_ (_10408_, _10369_, _10407_);
  and _18691_ (_10409_, _10369_, _09690_);
  or _18692_ (_10410_, _10409_, _10408_);
  or _18693_ (_10411_, _10410_, _10367_);
  or _18694_ (_10412_, _10374_, word_in[11]);
  and _18695_ (_10413_, _10412_, _10411_);
  or _18696_ (_10414_, _10413_, _10364_);
  or _18697_ (_10415_, _10365_, _09829_);
  and _18698_ (_10416_, _10415_, _10414_);
  and _18699_ (_10417_, _10416_, _10380_);
  and _18700_ (_10418_, _10363_, word_in[27]);
  or _18701_ (_14692_, _10418_, _10417_);
  or _18702_ (_10419_, _10365_, _09842_);
  not _18703_ (_10420_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor _18704_ (_10421_, _10369_, _10420_);
  and _18705_ (_10422_, _10369_, _09707_);
  or _18706_ (_10423_, _10422_, _10421_);
  and _18707_ (_10424_, _10423_, _10374_);
  and _18708_ (_10425_, _10367_, word_in[12]);
  or _18709_ (_10426_, _10425_, _10364_);
  or _18710_ (_10427_, _10426_, _10424_);
  and _18711_ (_10428_, _10427_, _10419_);
  or _18712_ (_10429_, _10428_, _10363_);
  or _18713_ (_10430_, _10380_, word_in[28]);
  and _18714_ (_14693_, _10430_, _10429_);
  not _18715_ (_10431_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor _18716_ (_10432_, _10369_, _10431_);
  and _18717_ (_10433_, _10369_, _09722_);
  or _18718_ (_10434_, _10433_, _10432_);
  or _18719_ (_10435_, _10434_, _10367_);
  or _18720_ (_10436_, _10374_, word_in[13]);
  and _18721_ (_10437_, _10436_, _10435_);
  or _18722_ (_10438_, _10437_, _10364_);
  or _18723_ (_10439_, _10365_, _09855_);
  and _18724_ (_10440_, _10439_, _10438_);
  and _18725_ (_10441_, _10440_, _10380_);
  and _18726_ (_10442_, _10363_, word_in[29]);
  or _18727_ (_09346_, _10442_, _10441_);
  or _18728_ (_10443_, _10365_, _09871_);
  not _18729_ (_10444_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor _18730_ (_10445_, _10369_, _10444_);
  and _18731_ (_10447_, _10369_, _09735_);
  or _18732_ (_10448_, _10447_, _10445_);
  and _18733_ (_10450_, _10448_, _10374_);
  and _18734_ (_10451_, _10367_, word_in[14]);
  or _18735_ (_10453_, _10451_, _10364_);
  or _18736_ (_10454_, _10453_, _10450_);
  and _18737_ (_10455_, _10454_, _10443_);
  or _18738_ (_10456_, _10455_, _10363_);
  or _18739_ (_10457_, _10380_, word_in[30]);
  and _18740_ (_09351_, _10457_, _10456_);
  or _18741_ (_10458_, _10365_, _08942_);
  nor _18742_ (_10459_, _10369_, _08785_);
  and _18743_ (_10460_, _10369_, _08953_);
  or _18744_ (_10461_, _10460_, _10459_);
  and _18745_ (_10462_, _10461_, _10374_);
  and _18746_ (_10463_, _10367_, word_in[15]);
  or _18747_ (_10464_, _10463_, _10364_);
  or _18748_ (_10465_, _10464_, _10462_);
  and _18749_ (_10466_, _10465_, _10458_);
  or _18750_ (_10467_, _10466_, _10363_);
  or _18751_ (_10468_, _10380_, word_in[31]);
  and _18752_ (_09354_, _10468_, _10467_);
  and _18753_ (_10469_, _08935_, _09016_);
  and _18754_ (_10470_, _10153_, _08740_);
  not _18755_ (_10471_, _10470_);
  or _18756_ (_10472_, _10471_, _09648_);
  and _18757_ (_10473_, _08945_, _08784_);
  not _18758_ (_10474_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _18759_ (_10475_, _10159_, _08948_);
  nor _18760_ (_10476_, _10475_, _10474_);
  and _18761_ (_10477_, _10475_, _09636_);
  or _18762_ (_10478_, _10477_, _10476_);
  or _18763_ (_10479_, _10478_, _10473_);
  not _18764_ (_10480_, _10473_);
  or _18765_ (_10481_, _10480_, word_in[8]);
  and _18766_ (_10482_, _10481_, _10479_);
  or _18767_ (_10483_, _10482_, _10470_);
  and _18768_ (_10484_, _10483_, _10472_);
  or _18769_ (_10485_, _10484_, _10469_);
  not _18770_ (_10486_, _10469_);
  or _18771_ (_10487_, _10486_, word_in[24]);
  and _18772_ (_14694_, _10487_, _10485_);
  or _18773_ (_10488_, _10480_, word_in[9]);
  not _18774_ (_10489_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor _18775_ (_10490_, _10475_, _10489_);
  and _18776_ (_10491_, _10475_, _09660_);
  or _18777_ (_10492_, _10491_, _10490_);
  or _18778_ (_10493_, _10492_, _10473_);
  and _18779_ (_10494_, _10493_, _10471_);
  and _18780_ (_10495_, _10494_, _10488_);
  and _18781_ (_10496_, _10470_, _09801_);
  or _18782_ (_10497_, _10496_, _10469_);
  or _18783_ (_10498_, _10497_, _10495_);
  or _18784_ (_10499_, _10486_, word_in[25]);
  and _18785_ (_14695_, _10499_, _10498_);
  or _18786_ (_10500_, _10471_, _09816_);
  not _18787_ (_10501_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor _18788_ (_10502_, _10475_, _10501_);
  and _18789_ (_10503_, _10475_, _09674_);
  or _18790_ (_10504_, _10503_, _10502_);
  or _18791_ (_10505_, _10504_, _10473_);
  or _18792_ (_10506_, _10480_, word_in[10]);
  and _18793_ (_10507_, _10506_, _10505_);
  or _18794_ (_10508_, _10507_, _10470_);
  and _18795_ (_10509_, _10508_, _10500_);
  and _18796_ (_10510_, _10509_, _10486_);
  and _18797_ (_10511_, _10469_, word_in[26]);
  or _18798_ (_14696_, _10511_, _10510_);
  not _18799_ (_10512_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor _18800_ (_10513_, _10475_, _10512_);
  and _18801_ (_10514_, _10475_, _09690_);
  nor _18802_ (_10515_, _10514_, _10513_);
  nor _18803_ (_10516_, _10515_, _10473_);
  and _18804_ (_10517_, _10473_, word_in[11]);
  or _18805_ (_10518_, _10517_, _10516_);
  and _18806_ (_10519_, _10518_, _10471_);
  and _18807_ (_10520_, _10470_, _09829_);
  or _18808_ (_10521_, _10520_, _10469_);
  or _18809_ (_10522_, _10521_, _10519_);
  or _18810_ (_10523_, _10486_, word_in[27]);
  and _18811_ (_14697_, _10523_, _10522_);
  or _18812_ (_10524_, _10480_, word_in[12]);
  not _18813_ (_10525_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor _18814_ (_10526_, _10475_, _10525_);
  and _18815_ (_10527_, _10475_, _09707_);
  or _18816_ (_10528_, _10527_, _10526_);
  or _18817_ (_10529_, _10528_, _10473_);
  and _18818_ (_10530_, _10529_, _10471_);
  and _18819_ (_10531_, _10530_, _10524_);
  and _18820_ (_10532_, _10470_, _09842_);
  or _18821_ (_10533_, _10532_, _10469_);
  or _18822_ (_10534_, _10533_, _10531_);
  or _18823_ (_10535_, _10486_, word_in[28]);
  and _18824_ (_14698_, _10535_, _10534_);
  or _18825_ (_10536_, _10471_, _09855_);
  not _18826_ (_10537_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor _18827_ (_10538_, _10475_, _10537_);
  and _18828_ (_10539_, _10475_, _09722_);
  or _18829_ (_10540_, _10539_, _10538_);
  or _18830_ (_10541_, _10540_, _10473_);
  or _18831_ (_10542_, _10480_, word_in[13]);
  and _18832_ (_10543_, _10542_, _10541_);
  or _18833_ (_10544_, _10543_, _10470_);
  and _18834_ (_10545_, _10544_, _10536_);
  or _18835_ (_10546_, _10545_, _10469_);
  or _18836_ (_10547_, _10486_, word_in[29]);
  and _18837_ (_14699_, _10547_, _10546_);
  not _18838_ (_10548_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor _18839_ (_10549_, _10475_, _10548_);
  and _18840_ (_10550_, _10475_, _09735_);
  nor _18841_ (_10551_, _10550_, _10549_);
  nor _18842_ (_10552_, _10551_, _10473_);
  and _18843_ (_10553_, _10473_, word_in[14]);
  or _18844_ (_10554_, _10553_, _10552_);
  and _18845_ (_10555_, _10554_, _10471_);
  and _18846_ (_10556_, _10470_, _09871_);
  or _18847_ (_10557_, _10556_, _10469_);
  or _18848_ (_10558_, _10557_, _10555_);
  or _18849_ (_10559_, _10486_, word_in[30]);
  and _18850_ (_14700_, _10559_, _10558_);
  or _18851_ (_10560_, _10471_, _08942_);
  nor _18852_ (_10561_, _10475_, _08687_);
  and _18853_ (_10562_, _10475_, _08953_);
  or _18854_ (_10563_, _10562_, _10561_);
  or _18855_ (_10564_, _10563_, _10473_);
  or _18856_ (_10565_, _10480_, word_in[15]);
  and _18857_ (_10566_, _10565_, _10564_);
  or _18858_ (_10567_, _10566_, _10470_);
  and _18859_ (_10568_, _10567_, _10560_);
  or _18860_ (_10569_, _10568_, _10469_);
  or _18861_ (_10570_, _10486_, word_in[31]);
  and _18862_ (_14701_, _10570_, _10569_);
  and _18863_ (_10571_, _08937_, _09058_);
  and _18864_ (_10572_, _08944_, _08722_);
  not _18865_ (_10573_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _18866_ (_10574_, _09630_, _08720_);
  and _18867_ (_10575_, _10574_, _09627_);
  nor _18868_ (_10576_, _10575_, _10573_);
  and _18869_ (_10577_, _10575_, _09636_);
  or _18870_ (_10578_, _10577_, _10576_);
  or _18871_ (_10579_, _10578_, _10572_);
  not _18872_ (_10580_, _10572_);
  or _18873_ (_10581_, _10580_, word_in[8]);
  and _18874_ (_10582_, _10581_, _10579_);
  or _18875_ (_10583_, _10582_, _10571_);
  and _18876_ (_10584_, _08935_, _08890_);
  not _18877_ (_10585_, _10584_);
  not _18878_ (_10586_, _10571_);
  or _18879_ (_10587_, _10586_, word_in[16]);
  and _18880_ (_10588_, _10587_, _10585_);
  and _18881_ (_10589_, _10588_, _10583_);
  and _18882_ (_10590_, _10584_, word_in[24]);
  or _18883_ (_09522_, _10590_, _10589_);
  not _18884_ (_10591_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _18885_ (_10592_, _10575_, _10591_);
  and _18886_ (_10593_, _10575_, _09660_);
  or _18887_ (_10594_, _10593_, _10592_);
  or _18888_ (_10595_, _10594_, _10572_);
  or _18889_ (_10596_, _10580_, word_in[9]);
  and _18890_ (_10597_, _10596_, _10595_);
  or _18891_ (_10598_, _10597_, _10571_);
  or _18892_ (_10599_, _10586_, word_in[17]);
  and _18893_ (_10600_, _10599_, _10585_);
  and _18894_ (_10601_, _10600_, _10598_);
  and _18895_ (_10602_, _10584_, word_in[25]);
  or _18896_ (_14702_, _10602_, _10601_);
  not _18897_ (_10603_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _18898_ (_10604_, _10575_, _10603_);
  and _18899_ (_10605_, _10575_, _09674_);
  or _18900_ (_10606_, _10605_, _10604_);
  or _18901_ (_10607_, _10606_, _10572_);
  or _18902_ (_10608_, _10580_, word_in[10]);
  and _18903_ (_10609_, _10608_, _10607_);
  or _18904_ (_10610_, _10609_, _10571_);
  or _18905_ (_10611_, _10586_, word_in[18]);
  and _18906_ (_10612_, _10611_, _10585_);
  and _18907_ (_10613_, _10612_, _10610_);
  and _18908_ (_10614_, _10584_, word_in[26]);
  or _18909_ (_09526_, _10614_, _10613_);
  not _18910_ (_10615_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _18911_ (_10616_, _10575_, _10615_);
  and _18912_ (_10617_, _10575_, _09690_);
  or _18913_ (_10618_, _10617_, _10616_);
  or _18914_ (_10619_, _10618_, _10572_);
  or _18915_ (_10620_, _10580_, word_in[11]);
  and _18916_ (_10621_, _10620_, _10619_);
  or _18917_ (_10622_, _10621_, _10571_);
  or _18918_ (_10623_, _10586_, word_in[19]);
  and _18919_ (_10624_, _10623_, _10585_);
  and _18920_ (_10625_, _10624_, _10622_);
  and _18921_ (_10626_, _10584_, word_in[27]);
  or _18922_ (_14703_, _10626_, _10625_);
  not _18923_ (_10627_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _18924_ (_10628_, _10575_, _10627_);
  and _18925_ (_10629_, _10575_, _09707_);
  or _18926_ (_10630_, _10629_, _10628_);
  or _18927_ (_10631_, _10630_, _10572_);
  or _18928_ (_10632_, _10580_, word_in[12]);
  and _18929_ (_10633_, _10632_, _10631_);
  or _18930_ (_10634_, _10633_, _10571_);
  or _18931_ (_10635_, _10586_, word_in[20]);
  and _18932_ (_10636_, _10635_, _10585_);
  and _18933_ (_10637_, _10636_, _10634_);
  and _18934_ (_10638_, _10584_, word_in[28]);
  or _18935_ (_14704_, _10638_, _10637_);
  not _18936_ (_10639_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _18937_ (_10640_, _10575_, _10639_);
  and _18938_ (_10641_, _10575_, _09722_);
  or _18939_ (_10642_, _10641_, _10640_);
  or _18940_ (_10643_, _10642_, _10572_);
  or _18941_ (_10644_, _10580_, word_in[13]);
  and _18942_ (_10645_, _10644_, _10643_);
  or _18943_ (_10646_, _10645_, _10571_);
  or _18944_ (_10647_, _10586_, word_in[21]);
  and _18945_ (_10648_, _10647_, _10585_);
  and _18946_ (_10649_, _10648_, _10646_);
  and _18947_ (_10650_, _10584_, word_in[29]);
  or _18948_ (_14705_, _10650_, _10649_);
  and _18949_ (_10651_, _10584_, word_in[30]);
  not _18950_ (_10652_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _18951_ (_10653_, _10575_, _10652_);
  and _18952_ (_10654_, _10575_, _09735_);
  or _18953_ (_10655_, _10654_, _10653_);
  and _18954_ (_10656_, _10655_, _10580_);
  and _18955_ (_10657_, _10572_, word_in[14]);
  or _18956_ (_10658_, _10657_, _10656_);
  or _18957_ (_10659_, _10658_, _10571_);
  nor _18958_ (_10660_, _10586_, word_in[22]);
  nor _18959_ (_10661_, _10660_, _10584_);
  and _18960_ (_10662_, _10661_, _10659_);
  or _18961_ (_09540_, _10662_, _10651_);
  nor _18962_ (_10663_, _10575_, _08765_);
  and _18963_ (_10664_, _10575_, _08953_);
  or _18964_ (_10665_, _10664_, _10663_);
  or _18965_ (_10666_, _10665_, _10572_);
  or _18966_ (_10667_, _10580_, word_in[15]);
  and _18967_ (_10668_, _10667_, _10666_);
  or _18968_ (_10669_, _10668_, _10571_);
  or _18969_ (_10670_, _10586_, word_in[23]);
  and _18970_ (_10671_, _10670_, _10585_);
  and _18971_ (_10672_, _10671_, _10669_);
  and _18972_ (_10673_, _10584_, word_in[31]);
  or _18973_ (_14706_, _10673_, _10672_);
  and _18974_ (_10674_, _07262_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nor _18975_ (_10675_, _07317_, _07262_);
  or _18976_ (_10676_, _10675_, _10674_);
  and _18977_ (_09596_, _10676_, _06989_);
  and _18978_ (_10677_, _08935_, _08711_);
  and _18979_ (_10678_, _10677_, _08880_);
  and _18980_ (_10679_, _09778_, _08822_);
  not _18981_ (_10681_, _10679_);
  or _18982_ (_10682_, _10681_, _09648_);
  and _18983_ (_10683_, _09768_, _08726_);
  not _18984_ (_10684_, _10683_);
  not _18985_ (_10685_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _18986_ (_10686_, _10574_, _09772_);
  nor _18987_ (_10687_, _10686_, _10685_);
  and _18988_ (_10688_, _10686_, _09636_);
  or _18989_ (_10689_, _10688_, _10687_);
  and _18990_ (_10690_, _10689_, _10684_);
  and _18991_ (_10691_, _10683_, word_in[8]);
  or _18992_ (_10692_, _10691_, _10679_);
  or _18993_ (_10693_, _10692_, _10690_);
  and _18994_ (_10694_, _10693_, _10682_);
  or _18995_ (_10695_, _10694_, _10678_);
  not _18996_ (_10696_, _10678_);
  or _18997_ (_10697_, _10696_, word_in[24]);
  and _18998_ (_14707_, _10697_, _10695_);
  or _18999_ (_10698_, _10681_, _09801_);
  not _19000_ (_10699_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _19001_ (_10700_, _10686_, _10699_);
  and _19002_ (_10701_, _10686_, _09660_);
  or _19003_ (_10702_, _10701_, _10700_);
  and _19004_ (_10703_, _10702_, _10684_);
  and _19005_ (_10704_, _10683_, word_in[9]);
  or _19006_ (_10705_, _10704_, _10679_);
  or _19007_ (_10706_, _10705_, _10703_);
  and _19008_ (_10707_, _10706_, _10698_);
  or _19009_ (_10708_, _10707_, _10678_);
  or _19010_ (_10709_, _10696_, word_in[25]);
  and _19011_ (_09612_, _10709_, _10708_);
  not _19012_ (_10710_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _19013_ (_10711_, _10686_, _10710_);
  and _19014_ (_10712_, _10686_, _09674_);
  or _19015_ (_10713_, _10712_, _10711_);
  and _19016_ (_10714_, _10713_, _10684_);
  and _19017_ (_10715_, _10683_, word_in[10]);
  or _19018_ (_10716_, _10715_, _10679_);
  or _19019_ (_10717_, _10716_, _10714_);
  or _19020_ (_10718_, _10681_, _09816_);
  and _19021_ (_10719_, _10718_, _10717_);
  or _19022_ (_10720_, _10719_, _10678_);
  or _19023_ (_10721_, _10696_, word_in[26]);
  and _19024_ (_09617_, _10721_, _10720_);
  and _19025_ (_10722_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  not _19026_ (_10723_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor _19027_ (_10724_, _07493_, _10723_);
  or _19028_ (_10725_, _10724_, _10722_);
  and _19029_ (_09620_, _10725_, _06989_);
  or _19030_ (_10726_, _10681_, _09829_);
  not _19031_ (_10727_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _19032_ (_10728_, _10686_, _10727_);
  and _19033_ (_10729_, _10686_, _09690_);
  or _19034_ (_10730_, _10729_, _10728_);
  and _19035_ (_10731_, _10730_, _10684_);
  and _19036_ (_10732_, _10683_, word_in[11]);
  or _19037_ (_10733_, _10732_, _10679_);
  or _19038_ (_10734_, _10733_, _10731_);
  and _19039_ (_10735_, _10734_, _10726_);
  or _19040_ (_10736_, _10735_, _10678_);
  or _19041_ (_10737_, _10696_, word_in[27]);
  and _19042_ (_09622_, _10737_, _10736_);
  and _19043_ (_10738_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  not _19044_ (_10739_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor _19045_ (_10740_, _07493_, _10739_);
  or _19046_ (_10741_, _10740_, _10738_);
  and _19047_ (_09624_, _10741_, _06989_);
  or _19048_ (_10742_, _10681_, _09842_);
  not _19049_ (_10743_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor _19050_ (_10744_, _10686_, _10743_);
  and _19051_ (_10745_, _10686_, _09707_);
  or _19052_ (_10746_, _10745_, _10744_);
  and _19053_ (_10747_, _10746_, _10684_);
  and _19054_ (_10748_, _10683_, word_in[12]);
  or _19055_ (_10749_, _10748_, _10679_);
  or _19056_ (_10750_, _10749_, _10747_);
  and _19057_ (_10751_, _10750_, _10742_);
  or _19058_ (_10752_, _10751_, _10678_);
  or _19059_ (_10753_, _10696_, word_in[28]);
  and _19060_ (_14708_, _10753_, _10752_);
  and _19061_ (_10754_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not _19062_ (_10755_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _19063_ (_10756_, _07493_, _10755_);
  or _19064_ (_10757_, _10756_, _10754_);
  and _19065_ (_09628_, _10757_, _06989_);
  or _19066_ (_10758_, _10681_, _09855_);
  not _19067_ (_10759_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _19068_ (_10760_, _10686_, _10759_);
  and _19069_ (_10761_, _10686_, _09722_);
  or _19070_ (_10762_, _10761_, _10760_);
  and _19071_ (_10763_, _10762_, _10684_);
  and _19072_ (_10764_, _10683_, word_in[13]);
  or _19073_ (_10765_, _10764_, _10679_);
  or _19074_ (_10766_, _10765_, _10763_);
  and _19075_ (_10767_, _10766_, _10758_);
  or _19076_ (_10768_, _10767_, _10678_);
  or _19077_ (_10769_, _10696_, word_in[29]);
  and _19078_ (_14709_, _10769_, _10768_);
  or _19079_ (_10770_, _10681_, _09871_);
  not _19080_ (_10771_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _19081_ (_10772_, _10686_, _10771_);
  and _19082_ (_10773_, _10686_, _09735_);
  or _19083_ (_10774_, _10773_, _10772_);
  and _19084_ (_10775_, _10774_, _10684_);
  and _19085_ (_10776_, _10683_, word_in[14]);
  or _19086_ (_10777_, _10776_, _10679_);
  or _19087_ (_10778_, _10777_, _10775_);
  and _19088_ (_10779_, _10778_, _10770_);
  or _19089_ (_10780_, _10779_, _10678_);
  or _19090_ (_10781_, _10696_, word_in[30]);
  and _19091_ (_14710_, _10781_, _10780_);
  or _19092_ (_10782_, _10681_, _08942_);
  nor _19093_ (_10783_, _10686_, _08674_);
  and _19094_ (_10784_, _10686_, _08953_);
  or _19095_ (_10785_, _10784_, _10783_);
  and _19096_ (_10786_, _10785_, _10684_);
  and _19097_ (_10787_, _10683_, word_in[15]);
  or _19098_ (_10788_, _10787_, _10679_);
  or _19099_ (_10789_, _10788_, _10786_);
  and _19100_ (_10790_, _10789_, _10782_);
  or _19101_ (_10791_, _10790_, _10678_);
  or _19102_ (_10792_, _10696_, word_in[31]);
  and _19103_ (_09635_, _10792_, _10791_);
  nor _19104_ (_10793_, _07325_, _06794_);
  and _19105_ (_10794_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and _19106_ (_10795_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor _19107_ (_10796_, _10795_, _10794_);
  and _19108_ (_10797_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _19109_ (_10798_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _19110_ (_10799_, _10798_, _10797_);
  and _19111_ (_10800_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and _19112_ (_10801_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _19113_ (_10802_, _10801_, _10800_);
  and _19114_ (_10803_, _10802_, _10799_);
  and _19115_ (_10804_, _10803_, _10796_);
  nor _19116_ (_10805_, _10804_, _08477_);
  nor _19117_ (_10806_, _10805_, _10793_);
  nor _19118_ (_09651_, _10806_, rst);
  not _19119_ (_10807_, _07360_);
  not _19120_ (_10808_, _08496_);
  not _19121_ (_10809_, _08529_);
  and _19122_ (_10810_, _10809_, _08512_);
  and _19123_ (_10811_, _10810_, _10808_);
  and _19124_ (_10812_, _10811_, _10807_);
  nor _19125_ (_10813_, _08576_, _08463_);
  nor _19126_ (_10814_, _08561_, _08545_);
  and _19127_ (_10815_, _10814_, _10813_);
  and _19128_ (_10816_, _10815_, _10812_);
  and _19129_ (_10817_, _08561_, _08545_);
  and _19130_ (_10818_, _10817_, _10813_);
  not _19131_ (_10819_, _08512_);
  and _19132_ (_10820_, _10819_, _08496_);
  and _19133_ (_10821_, _10820_, _10809_);
  and _19134_ (_10822_, _10821_, _10818_);
  nor _19135_ (_10823_, _10822_, _10816_);
  and _19136_ (_10824_, _08576_, _08463_);
  and _19137_ (_10825_, _10824_, _10817_);
  and _19138_ (_10826_, _10825_, _10812_);
  and _19139_ (_10827_, _10813_, _08561_);
  and _19140_ (_10828_, _10827_, _10812_);
  nor _19141_ (_10829_, _10828_, _10826_);
  and _19142_ (_10830_, _10829_, _10823_);
  and _19143_ (_10831_, _10811_, _07360_);
  nor _19144_ (_10832_, _08512_, _08496_);
  and _19145_ (_10833_, _10832_, _10809_);
  and _19146_ (_10834_, _10833_, _10807_);
  not _19147_ (_10835_, _08576_);
  nor _19148_ (_10836_, _10835_, _08463_);
  and _19149_ (_10837_, _10836_, _08561_);
  and _19150_ (_10838_, _10837_, _10834_);
  nor _19151_ (_10839_, _10838_, _10831_);
  not _19152_ (_10840_, _08545_);
  and _19153_ (_10841_, _10824_, _10840_);
  and _19154_ (_10842_, _10841_, _10821_);
  and _19155_ (_10843_, _10821_, _08545_);
  and _19156_ (_10844_, _10824_, _08561_);
  and _19157_ (_10845_, _10844_, _10843_);
  nor _19158_ (_10846_, _10845_, _10842_);
  and _19159_ (_10847_, _10846_, _10839_);
  and _19160_ (_10848_, _10847_, _10830_);
  and _19161_ (_10849_, _10833_, _07360_);
  and _19162_ (_10850_, _10835_, _08463_);
  and _19163_ (_10851_, _10850_, _08561_);
  and _19164_ (_10852_, _10851_, _10849_);
  not _19165_ (_10853_, _10852_);
  not _19166_ (_10854_, _08561_);
  and _19167_ (_10855_, _10854_, _08463_);
  and _19168_ (_10856_, _10855_, _10835_);
  and _19169_ (_10857_, _10856_, _10812_);
  not _19170_ (_10858_, _10857_);
  and _19171_ (_10859_, _10824_, _10814_);
  and _19172_ (_10860_, _10859_, _10812_);
  and _19173_ (_10861_, _10825_, _08529_);
  nor _19174_ (_10862_, _10861_, _10860_);
  and _19175_ (_10863_, _10862_, _10858_);
  and _19176_ (_10864_, _10863_, _10853_);
  and _19177_ (_10865_, _10864_, _10848_);
  nor _19178_ (_10866_, _10854_, _08545_);
  and _19179_ (_10867_, _10866_, _10824_);
  not _19180_ (_10868_, _10867_);
  and _19181_ (_10869_, _08512_, _08496_);
  and _19182_ (_10870_, _10869_, _10809_);
  and _19183_ (_10871_, _10870_, _10807_);
  nor _19184_ (_10872_, _10871_, _10812_);
  nor _19185_ (_10873_, _10872_, _10868_);
  not _19186_ (_10874_, _10873_);
  and _19187_ (_10875_, _10854_, _08545_);
  and _19188_ (_10876_, _10875_, _10850_);
  and _19189_ (_10878_, _10876_, _08529_);
  and _19190_ (_10879_, _10875_, _10813_);
  not _19191_ (_10880_, _10879_);
  nor _19192_ (_10881_, _10871_, _10833_);
  nor _19193_ (_10882_, _10881_, _10880_);
  nor _19194_ (_10883_, _10882_, _10878_);
  and _19195_ (_10884_, _10883_, _10874_);
  not _19196_ (_10885_, _10815_);
  nor _19197_ (_10886_, _10881_, _10885_);
  and _19198_ (_10887_, _10849_, _10836_);
  nor _19199_ (_10888_, _10887_, _10886_);
  and _19200_ (_10889_, _10866_, _10813_);
  nor _19201_ (_10890_, _10869_, _10832_);
  nor _19202_ (_10891_, _10890_, _08529_);
  and _19203_ (_10892_, _10891_, _10889_);
  not _19204_ (_10893_, _10859_);
  nor _19205_ (_10894_, _10871_, _08529_);
  nor _19206_ (_10895_, _10894_, _10893_);
  nor _19207_ (_10896_, _10895_, _10892_);
  and _19208_ (_10897_, _10896_, _10888_);
  and _19209_ (_10898_, _10897_, _10884_);
  and _19210_ (_10899_, _10898_, _10865_);
  nor _19211_ (_10900_, _10859_, _10818_);
  not _19212_ (_10901_, _10900_);
  and _19213_ (_10902_, _10901_, _10849_);
  and _19214_ (_10903_, _10836_, _10854_);
  and _19215_ (_10904_, _10903_, _10871_);
  nor _19216_ (_10905_, _10904_, _10902_);
  and _19217_ (_10906_, _10876_, _10849_);
  not _19218_ (_10907_, _10817_);
  not _19219_ (_10908_, _10814_);
  and _19220_ (_10909_, _10836_, _10908_);
  and _19221_ (_10910_, _10909_, _10907_);
  and _19222_ (_10911_, _10910_, _10812_);
  and _19223_ (_10912_, _10833_, _10825_);
  and _19224_ (_10913_, _10912_, _10807_);
  or _19225_ (_10914_, _10913_, _10911_);
  nor _19226_ (_10915_, _10914_, _10906_);
  and _19227_ (_10916_, _10915_, _10905_);
  and _19228_ (_10917_, _10870_, _07360_);
  and _19229_ (_10918_, _10917_, _10815_);
  and _19230_ (_10919_, _10875_, _10824_);
  and _19231_ (_10920_, _10919_, _10812_);
  nor _19232_ (_10921_, _10920_, _10918_);
  nor _19233_ (_10922_, _10867_, _10818_);
  nor _19234_ (_10923_, _10922_, _10809_);
  not _19235_ (_10924_, _10871_);
  not _19236_ (_10925_, _10876_);
  nor _19237_ (_10926_, _10825_, _10818_);
  and _19238_ (_10927_, _10926_, _10925_);
  nor _19239_ (_10928_, _10927_, _10924_);
  nor _19240_ (_10929_, _10928_, _10923_);
  and _19241_ (_10930_, _10929_, _10921_);
  and _19242_ (_10931_, _10849_, _10825_);
  and _19243_ (_10932_, _10917_, _10879_);
  or _19244_ (_10933_, _10932_, _10931_);
  and _19245_ (_10934_, _10850_, _10814_);
  nor _19246_ (_10935_, _10934_, _10919_);
  nor _19247_ (_10936_, _10871_, _10849_);
  nor _19248_ (_10937_, _10936_, _10935_);
  nor _19249_ (_10938_, _10937_, _10933_);
  and _19250_ (_10939_, _10836_, _10817_);
  or _19251_ (_10940_, _10939_, _10879_);
  nand _19252_ (_10941_, _10940_, _10812_);
  not _19253_ (_10942_, _10834_);
  nor _19254_ (_10943_, _10919_, _10818_);
  nor _19255_ (_10944_, _10943_, _10942_);
  not _19256_ (_10945_, _10944_);
  and _19257_ (_10946_, _10945_, _10941_);
  and _19258_ (_10947_, _10946_, _10938_);
  and _19259_ (_10948_, _10947_, _10930_);
  and _19260_ (_10949_, _10948_, _10916_);
  and _19261_ (_10950_, _10949_, _10899_);
  nor _19262_ (_10951_, _10861_, _10845_);
  and _19263_ (_10952_, _10917_, _10889_);
  and _19264_ (_10953_, _10939_, _10812_);
  nor _19265_ (_10954_, _10953_, _10952_);
  and _19266_ (_10955_, _10954_, _10951_);
  not _19267_ (_10956_, _10933_);
  and _19268_ (_10957_, _10956_, _10921_);
  and _19269_ (_10958_, _10957_, _10955_);
  and _19270_ (_10959_, _10958_, _10916_);
  not _19271_ (_10960_, _10959_);
  nor _19272_ (_10961_, _10960_, _10950_);
  nor _19273_ (_10962_, _10961_, _07490_);
  nand _19274_ (_10963_, _10962_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _19275_ (_10964_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  or _19276_ (_10965_, _10962_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and _19277_ (_10966_, _10965_, _10964_);
  and _19278_ (_09655_, _10966_, _10963_);
  nor _19279_ (_10967_, _07035_, _06810_);
  not _19280_ (_10968_, _10967_);
  and _19281_ (_10969_, _10968_, _09133_);
  and _19282_ (_10970_, _10969_, _09115_);
  nor _19283_ (_10971_, _10970_, _07262_);
  nor _19284_ (_10972_, _08994_, _06982_);
  nand _19285_ (_10973_, _10972_, _07127_);
  or _19286_ (_10974_, _10973_, _07131_);
  and _19287_ (_10975_, _10974_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or _19288_ (_10976_, _10975_, _10971_);
  and _19289_ (_09662_, _10976_, _06989_);
  and _19290_ (_10977_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _06989_);
  and _19291_ (_10978_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not _19292_ (_10979_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _19293_ (_10980_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _19294_ (_10981_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _19295_ (_10982_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _19296_ (_10983_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor _19297_ (_10984_, _10983_, _10981_);
  and _19298_ (_10985_, _10984_, _10982_);
  nor _19299_ (_10986_, _10985_, _10981_);
  nor _19300_ (_10987_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _19301_ (_10988_, _10987_, _10980_);
  not _19302_ (_10990_, _10988_);
  nor _19303_ (_10991_, _10990_, _10986_);
  nor _19304_ (_10992_, _10991_, _10980_);
  not _19305_ (_10993_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not _19306_ (_10994_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  not _19307_ (_10995_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not _19308_ (_10996_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _19309_ (_10997_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _19310_ (_10998_, _10997_, _10996_);
  and _19311_ (_10999_, _10998_, _10995_);
  and _19312_ (_11000_, _10999_, _10994_);
  and _19313_ (_11001_, _11000_, _10993_);
  and _19314_ (_11002_, _11001_, _10992_);
  nor _19315_ (_11003_, _11002_, _10979_);
  and _19316_ (_11004_, _11002_, _10979_);
  nor _19317_ (_11006_, _11004_, _11003_);
  not _19318_ (_11007_, _11006_);
  and _19319_ (_11008_, _10999_, _10992_);
  and _19320_ (_11009_, _11008_, _10994_);
  nor _19321_ (_11010_, _11009_, _10993_);
  nor _19322_ (_11011_, _11010_, _11002_);
  nor _19323_ (_11012_, _11008_, _10994_);
  nor _19324_ (_11013_, _11012_, _11009_);
  not _19325_ (_11014_, _11013_);
  and _19326_ (_11015_, _10998_, _10992_);
  nor _19327_ (_11016_, _11015_, _10995_);
  nor _19328_ (_11017_, _11016_, _11008_);
  not _19329_ (_11018_, _11017_);
  and _19330_ (_11019_, _10992_, _10997_);
  nor _19331_ (_11020_, _11019_, _10996_);
  nor _19332_ (_11021_, _11020_, _11015_);
  not _19333_ (_11022_, _11021_);
  nor _19334_ (_11023_, _10992_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and _19335_ (_11024_, _10992_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or _19336_ (_11025_, _11024_, _11023_);
  not _19337_ (_11026_, _11025_);
  nor _19338_ (_11027_, _10984_, _10982_);
  nor _19339_ (_11028_, _11027_, _10985_);
  not _19340_ (_11029_, _11028_);
  nor _19341_ (_11030_, _11029_, _10950_);
  not _19342_ (_11032_, _10961_);
  nor _19343_ (_11033_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor _19344_ (_11034_, _11033_, _10982_);
  and _19345_ (_11035_, _11034_, _11032_);
  and _19346_ (_11036_, _11029_, _10950_);
  nor _19347_ (_11037_, _11036_, _11030_);
  and _19348_ (_11038_, _11037_, _11035_);
  nor _19349_ (_11039_, _11038_, _11030_);
  not _19350_ (_11040_, _11039_);
  and _19351_ (_11041_, _10990_, _10986_);
  nor _19352_ (_11042_, _11041_, _10991_);
  and _19353_ (_11043_, _11042_, _11040_);
  and _19354_ (_11044_, _11043_, _11026_);
  and _19355_ (_11045_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _19356_ (_11046_, _11045_, _10997_);
  nand _19357_ (_11047_, _11046_, _11023_);
  or _19358_ (_11048_, _11046_, _11023_);
  and _19359_ (_11049_, _11048_, _11047_);
  and _19360_ (_11050_, _11049_, _11044_);
  and _19361_ (_11051_, _11050_, _11022_);
  and _19362_ (_11052_, _11051_, _11018_);
  nand _19363_ (_11053_, _11052_, _11014_);
  nor _19364_ (_11054_, _11053_, _11011_);
  and _19365_ (_11055_, _11054_, _11007_);
  nor _19366_ (_11056_, _11054_, _11007_);
  nor _19367_ (_11057_, _11056_, _11055_);
  or _19368_ (_11058_, _11057_, _08477_);
  or _19369_ (_11059_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _19370_ (_11060_, _11059_, _10964_);
  and _19371_ (_11061_, _11060_, _11058_);
  or _19372_ (_09669_, _11061_, _10978_);
  and _19373_ (_11062_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and _19374_ (_11063_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor _19375_ (_11064_, _11063_, _11062_);
  and _19376_ (_11065_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _19377_ (_11066_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor _19378_ (_11067_, _11066_, _11065_);
  and _19379_ (_11068_, _11067_, _11064_);
  and _19380_ (_11069_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _19381_ (_11070_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  nor _19382_ (_11071_, _11070_, _11069_);
  and _19383_ (_11072_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _19384_ (_11073_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor _19385_ (_11074_, _11073_, _11072_);
  and _19386_ (_11075_, _11074_, _11071_);
  and _19387_ (_11076_, _11075_, _11068_);
  nor _19388_ (_11077_, _11076_, _07378_);
  and _19389_ (_11078_, _09009_, _07378_);
  nor _19390_ (_11079_, _11078_, _11077_);
  nor _19391_ (_09677_, _11079_, rst);
  or _19392_ (_11080_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  not _19393_ (_11081_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand _19394_ (_11082_, _07493_, _11081_);
  and _19395_ (_11083_, _11082_, _06989_);
  and _19396_ (_09687_, _11083_, _11080_);
  or _19397_ (_11084_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  not _19398_ (_11085_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand _19399_ (_11086_, _07493_, _11085_);
  and _19400_ (_11087_, _11086_, _06989_);
  and _19401_ (_09691_, _11087_, _11084_);
  and _19402_ (_11088_, _09891_, _08880_);
  and _19403_ (_11089_, _09893_, _08822_);
  not _19404_ (_11090_, _11089_);
  or _19405_ (_11091_, _11090_, _09648_);
  and _19406_ (_11092_, _09897_, _08726_);
  not _19407_ (_11093_, _11092_);
  not _19408_ (_11094_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _19409_ (_11095_, _10574_, _09902_);
  nor _19410_ (_11096_, _11095_, _11094_);
  and _19411_ (_11097_, _11095_, _09636_);
  or _19412_ (_11098_, _11097_, _11096_);
  and _19413_ (_11099_, _11098_, _11093_);
  and _19414_ (_11100_, _11092_, word_in[8]);
  or _19415_ (_11101_, _11100_, _11089_);
  or _19416_ (_11102_, _11101_, _11099_);
  and _19417_ (_11103_, _11102_, _11091_);
  or _19418_ (_11104_, _11103_, _11088_);
  not _19419_ (_11105_, _11088_);
  or _19420_ (_11106_, _11105_, word_in[24]);
  and _19421_ (_14649_, _11106_, _11104_);
  or _19422_ (_11107_, _11090_, _09801_);
  not _19423_ (_11108_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor _19424_ (_11109_, _11095_, _11108_);
  and _19425_ (_11110_, _11095_, _09660_);
  or _19426_ (_11111_, _11110_, _11109_);
  and _19427_ (_11112_, _11111_, _11093_);
  and _19428_ (_11113_, _11092_, word_in[9]);
  or _19429_ (_11114_, _11113_, _11089_);
  or _19430_ (_11115_, _11114_, _11112_);
  and _19431_ (_11116_, _11115_, _11107_);
  or _19432_ (_11117_, _11116_, _11088_);
  or _19433_ (_11118_, _11105_, word_in[25]);
  and _19434_ (_14650_, _11118_, _11117_);
  or _19435_ (_11119_, _11090_, _09816_);
  not _19436_ (_11120_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor _19437_ (_11121_, _11095_, _11120_);
  and _19438_ (_11122_, _11095_, _09674_);
  or _19439_ (_11123_, _11122_, _11121_);
  and _19440_ (_11124_, _11123_, _11093_);
  and _19441_ (_11125_, _11092_, word_in[10]);
  or _19442_ (_11126_, _11125_, _11089_);
  or _19443_ (_11127_, _11126_, _11124_);
  and _19444_ (_11128_, _11127_, _11119_);
  and _19445_ (_11129_, _11128_, _11105_);
  and _19446_ (_11130_, _11088_, word_in[26]);
  or _19447_ (_14651_, _11130_, _11129_);
  or _19448_ (_11131_, _11090_, _09829_);
  not _19449_ (_11132_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor _19450_ (_11133_, _11095_, _11132_);
  and _19451_ (_11134_, _11095_, _09690_);
  or _19452_ (_11135_, _11134_, _11133_);
  and _19453_ (_11136_, _11135_, _11093_);
  and _19454_ (_11137_, _11092_, word_in[11]);
  or _19455_ (_11138_, _11137_, _11089_);
  or _19456_ (_11139_, _11138_, _11136_);
  and _19457_ (_11140_, _11139_, _11131_);
  or _19458_ (_11141_, _11140_, _11088_);
  or _19459_ (_11142_, _11105_, word_in[27]);
  and _19460_ (_14652_, _11142_, _11141_);
  or _19461_ (_11143_, _11090_, _09842_);
  not _19462_ (_11144_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor _19463_ (_11145_, _11095_, _11144_);
  and _19464_ (_11146_, _11095_, _09707_);
  or _19465_ (_11147_, _11146_, _11145_);
  and _19466_ (_11148_, _11147_, _11093_);
  and _19467_ (_11149_, _11092_, word_in[12]);
  or _19468_ (_11150_, _11149_, _11089_);
  or _19469_ (_11151_, _11150_, _11148_);
  and _19470_ (_11152_, _11151_, _11143_);
  or _19471_ (_11153_, _11152_, _11088_);
  or _19472_ (_11154_, _11105_, word_in[28]);
  and _19473_ (_14653_, _11154_, _11153_);
  or _19474_ (_11155_, _11090_, _09855_);
  not _19475_ (_11156_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor _19476_ (_11157_, _11095_, _11156_);
  and _19477_ (_11158_, _11095_, _09722_);
  or _19478_ (_11159_, _11158_, _11157_);
  and _19479_ (_11160_, _11159_, _11093_);
  and _19480_ (_11161_, _11092_, word_in[13]);
  or _19481_ (_11162_, _11161_, _11089_);
  or _19482_ (_11163_, _11162_, _11160_);
  and _19483_ (_11164_, _11163_, _11155_);
  or _19484_ (_11165_, _11164_, _11088_);
  or _19485_ (_11166_, _11105_, word_in[29]);
  and _19486_ (_14654_, _11166_, _11165_);
  or _19487_ (_11167_, _11090_, _09871_);
  not _19488_ (_11168_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor _19489_ (_11169_, _11095_, _11168_);
  and _19490_ (_11170_, _11095_, _09735_);
  or _19491_ (_11171_, _11170_, _11169_);
  and _19492_ (_11172_, _11171_, _11093_);
  and _19493_ (_11173_, _11092_, word_in[14]);
  or _19494_ (_11174_, _11173_, _11089_);
  or _19495_ (_11175_, _11174_, _11172_);
  and _19496_ (_11176_, _11175_, _11167_);
  or _19497_ (_11177_, _11176_, _11088_);
  or _19498_ (_11178_, _11105_, word_in[30]);
  and _19499_ (_09711_, _11178_, _11177_);
  or _19500_ (_11179_, _11090_, _08942_);
  nor _19501_ (_11180_, _11095_, _08760_);
  and _19502_ (_11181_, _11095_, _08953_);
  or _19503_ (_11182_, _11181_, _11180_);
  and _19504_ (_11183_, _11182_, _11093_);
  and _19505_ (_11184_, _11092_, word_in[15]);
  or _19506_ (_11185_, _11184_, _11089_);
  or _19507_ (_11186_, _11185_, _11183_);
  and _19508_ (_11187_, _11186_, _11179_);
  or _19509_ (_11188_, _11187_, _11088_);
  or _19510_ (_11189_, _11105_, word_in[31]);
  and _19511_ (_14655_, _11189_, _11188_);
  and _19512_ (_11190_, _07490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and _19513_ (_11191_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _19514_ (_11192_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _19515_ (_11193_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _19516_ (_11194_, _11193_, _11192_);
  and _19517_ (_11195_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _19518_ (_11196_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _19519_ (_11197_, _11196_, _11195_);
  and _19520_ (_11198_, _11197_, _11194_);
  and _19521_ (_11199_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _19522_ (_11201_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _19523_ (_11202_, _11201_, _11199_);
  and _19524_ (_11203_, _11202_, _11198_);
  nor _19525_ (_11204_, _11203_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _19526_ (_11205_, _11204_, _11191_);
  nor _19527_ (_11206_, _11205_, _07490_);
  nor _19528_ (_11207_, _11206_, _11190_);
  nor _19529_ (_09733_, _11207_, rst);
  nor _19530_ (_11208_, _07325_, _06716_);
  and _19531_ (_11209_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _19532_ (_11210_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _19533_ (_11211_, _11210_, _11209_);
  and _19534_ (_11212_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _19535_ (_11213_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor _19536_ (_11214_, _11213_, _11212_);
  and _19537_ (_11215_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _19538_ (_11216_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _19539_ (_11217_, _11216_, _11215_);
  and _19540_ (_11218_, _11217_, _11214_);
  and _19541_ (_11219_, _11218_, _11211_);
  nor _19542_ (_11220_, _11219_, _08477_);
  nor _19543_ (_11221_, _11220_, _11208_);
  nor _19544_ (_09747_, _11221_, rst);
  and _19545_ (_11223_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  not _19546_ (_11224_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor _19547_ (_11225_, _07493_, _11224_);
  or _19548_ (_11226_, _11225_, _11223_);
  and _19549_ (_09779_, _11226_, _06989_);
  and _19550_ (_11227_, _08945_, _08726_);
  not _19551_ (_11229_, _11227_);
  not _19552_ (_11230_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _19553_ (_11231_, _10574_, _08948_);
  nor _19554_ (_11232_, _11231_, _11230_);
  and _19555_ (_11233_, _11231_, _09636_);
  or _19556_ (_11234_, _11233_, _11232_);
  and _19557_ (_11235_, _11234_, _11229_);
  and _19558_ (_11236_, _10023_, _08822_);
  and _19559_ (_11237_, _11227_, word_in[8]);
  or _19560_ (_11238_, _11237_, _11236_);
  or _19561_ (_11239_, _11238_, _11235_);
  and _19562_ (_11240_, _08935_, _09299_);
  not _19563_ (_11241_, _11240_);
  not _19564_ (_11242_, _11236_);
  or _19565_ (_11243_, _11242_, _09648_);
  and _19566_ (_11244_, _11243_, _11241_);
  and _19567_ (_11245_, _11244_, _11239_);
  and _19568_ (_11246_, _11240_, word_in[24]);
  or _19569_ (_14656_, _11246_, _11245_);
  not _19570_ (_11247_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor _19571_ (_11248_, _11231_, _11247_);
  and _19572_ (_11249_, _11231_, _09660_);
  or _19573_ (_11250_, _11249_, _11248_);
  and _19574_ (_11251_, _11250_, _11229_);
  and _19575_ (_11252_, _11227_, word_in[9]);
  or _19576_ (_11253_, _11252_, _11236_);
  or _19577_ (_11254_, _11253_, _11251_);
  or _19578_ (_11255_, _11242_, _09801_);
  and _19579_ (_11256_, _11255_, _11241_);
  and _19580_ (_11257_, _11256_, _11254_);
  and _19581_ (_11258_, _11240_, word_in[25]);
  or _19582_ (_14657_, _11258_, _11257_);
  not _19583_ (_11260_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor _19584_ (_11261_, _11231_, _11260_);
  and _19585_ (_11262_, _11231_, _09674_);
  or _19586_ (_11263_, _11262_, _11261_);
  and _19587_ (_11264_, _11263_, _11229_);
  and _19588_ (_11265_, _11227_, word_in[10]);
  or _19589_ (_11266_, _11265_, _11236_);
  or _19590_ (_11267_, _11266_, _11264_);
  or _19591_ (_11269_, _11242_, _09816_);
  and _19592_ (_11270_, _11269_, _11241_);
  and _19593_ (_11271_, _11270_, _11267_);
  and _19594_ (_11272_, _11240_, word_in[26]);
  or _19595_ (_14658_, _11272_, _11271_);
  not _19596_ (_11273_, _07493_);
  and _19597_ (_11274_, _11045_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and _19598_ (_11275_, _11274_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and _19599_ (_11276_, _11275_, _11273_);
  and _19600_ (_11277_, _11276_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor _19601_ (_11278_, _11276_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or _19602_ (_11279_, _11278_, _11277_);
  not _19603_ (_11280_, _07412_);
  and _19604_ (_11281_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _19605_ (_11282_, _07324_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _19606_ (_11283_, _11282_);
  or _19607_ (_11284_, _08529_, _07327_);
  nor _19608_ (_11285_, _07325_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor _19609_ (_11286_, _11285_, _07362_);
  and _19610_ (_11287_, _11286_, _11284_);
  nor _19611_ (_11288_, _11287_, _09388_);
  and _19612_ (_11289_, _11288_, _09547_);
  and _19613_ (_11290_, _11289_, _07365_);
  or _19614_ (_11291_, _08561_, _07327_);
  nor _19615_ (_11292_, _07325_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor _19616_ (_11293_, _11292_, _07362_);
  and _19617_ (_11294_, _11293_, _11291_);
  not _19618_ (_11295_, _11294_);
  or _19619_ (_11296_, _08463_, _07327_);
  nor _19620_ (_11297_, _07325_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor _19621_ (_11298_, _11297_, _07362_);
  and _19622_ (_11299_, _11298_, _11296_);
  nand _19623_ (_11300_, _08576_, _07326_);
  nor _19624_ (_11301_, _07325_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor _19625_ (_11302_, _11301_, _07362_);
  and _19626_ (_11303_, _11302_, _11300_);
  not _19627_ (_11304_, _11303_);
  and _19628_ (_11305_, _11304_, _11299_);
  and _19629_ (_11306_, _11305_, _11295_);
  nor _19630_ (_11308_, _08545_, _07327_);
  not _19631_ (_11309_, _11308_);
  nor _19632_ (_11310_, _07325_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor _19633_ (_11311_, _11310_, _07362_);
  and _19634_ (_11312_, _11311_, _11309_);
  and _19635_ (_11313_, _11312_, _11306_);
  and _19636_ (_11314_, _11313_, _11290_);
  not _19637_ (_11315_, _11314_);
  not _19638_ (_11316_, _11312_);
  and _19639_ (_11317_, _11305_, _11294_);
  and _19640_ (_11319_, _11317_, _11316_);
  and _19641_ (_11320_, _11319_, _11290_);
  nor _19642_ (_11321_, _11304_, _11299_);
  and _19643_ (_11322_, _11321_, _11294_);
  and _19644_ (_11324_, _11322_, _11312_);
  and _19645_ (_11325_, _11324_, _11290_);
  nor _19646_ (_11326_, _11325_, _11320_);
  and _19647_ (_11327_, _11326_, _11315_);
  and _19648_ (_11328_, _11316_, _11306_);
  nor _19649_ (_11329_, _09547_, _07365_);
  not _19650_ (_11330_, _11287_);
  and _19651_ (_11331_, _11330_, _09388_);
  and _19652_ (_11332_, _11331_, _11329_);
  and _19653_ (_11333_, _11332_, _11328_);
  and _19654_ (_11334_, _11332_, _11319_);
  nor _19655_ (_11335_, _11334_, _11333_);
  and _19656_ (_11336_, _11335_, _11327_);
  nor _19657_ (_11337_, _11336_, _11283_);
  not _19658_ (_11338_, _11337_);
  and _19659_ (_11339_, _11329_, _11288_);
  not _19660_ (_11340_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _19661_ (_11341_, \oc8051_top_1.oc8051_decoder1.state [1], _06406_);
  and _19662_ (_11342_, _11341_, _11340_);
  and _19663_ (_11343_, _11342_, _11321_);
  and _19664_ (_11344_, _11343_, _11339_);
  not _19665_ (_11345_, _07324_);
  nor _19666_ (_11346_, _11335_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and _19667_ (_11347_, _11346_, _11345_);
  nor _19668_ (_11348_, _11347_, _11344_);
  and _19669_ (_11349_, _11348_, _11338_);
  nor _19670_ (_11350_, _11349_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _19671_ (_11351_, _11350_, _11281_);
  and _19672_ (_11352_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _19673_ (_11353_, _06406_, \oc8051_top_1.oc8051_decoder1.state [0]);
  nor _19674_ (_11354_, _11303_, _11299_);
  and _19675_ (_11355_, _11354_, _11295_);
  and _19676_ (_11356_, _11355_, _11312_);
  and _19677_ (_11358_, _11356_, _11339_);
  and _19678_ (_11359_, _11354_, _11294_);
  and _19679_ (_11360_, _11359_, _11339_);
  nor _19680_ (_11361_, _11360_, _11358_);
  not _19681_ (_11363_, _11361_);
  and _19682_ (_11364_, _11321_, _11295_);
  and _19683_ (_11365_, _11364_, _11339_);
  and _19684_ (_11366_, _11365_, _11342_);
  nor _19685_ (_11367_, _11366_, _11363_);
  nor _19686_ (_11368_, _11367_, _11353_);
  and _19687_ (_11369_, _11339_, _11321_);
  and _19688_ (_11370_, _11369_, _11342_);
  not _19689_ (_11371_, _11370_);
  nor _19690_ (_11372_, _11371_, _11368_);
  nor _19691_ (_11373_, _11304_, _11294_);
  and _19692_ (_11374_, _11373_, _11299_);
  and _19693_ (_11375_, _11374_, _11312_);
  and _19694_ (_11376_, _11375_, _11339_);
  and _19695_ (_11377_, _09547_, _09388_);
  nor _19696_ (_11378_, _11287_, _11312_);
  and _19697_ (_11379_, _11378_, _11377_);
  and _19698_ (_11380_, _11379_, _11306_);
  nor _19699_ (_11381_, _11380_, _11376_);
  and _19700_ (_11382_, _11289_, _07383_);
  and _19701_ (_11383_, _11359_, _11382_);
  and _19702_ (_11385_, _11379_, _11322_);
  nor _19703_ (_11386_, _11385_, _11383_);
  and _19704_ (_11387_, _11379_, _11364_);
  and _19705_ (_11388_, _11303_, _11294_);
  and _19706_ (_11389_, _11388_, _11299_);
  and _19707_ (_11390_, _11379_, _11389_);
  nor _19708_ (_11391_, _11390_, _11387_);
  and _19709_ (_11392_, _11391_, _11386_);
  and _19710_ (_11393_, _11392_, _11381_);
  and _19711_ (_11394_, _11377_, _11330_);
  and _19712_ (_11395_, _11394_, _11374_);
  and _19713_ (_11396_, _11394_, _11312_);
  and _19714_ (_11397_, _11396_, _11306_);
  nor _19715_ (_11398_, _11397_, _11395_);
  and _19716_ (_11399_, _11317_, _11312_);
  and _19717_ (_11400_, _11399_, _11394_);
  and _19718_ (_11401_, _11355_, _11394_);
  nor _19719_ (_11402_, _11401_, _11400_);
  and _19720_ (_11403_, _11364_, _11312_);
  and _19721_ (_11404_, _11403_, _11394_);
  and _19722_ (_11405_, _11359_, _11394_);
  nor _19723_ (_11406_, _11405_, _11404_);
  and _19724_ (_11407_, _11406_, _11402_);
  and _19725_ (_11408_, _11407_, _11398_);
  and _19726_ (_11409_, _11408_, _11393_);
  and _19727_ (_11410_, _11409_, _11327_);
  nor _19728_ (_11411_, _11410_, _11283_);
  and _19729_ (_11412_, _11341_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and _19730_ (_11413_, _11412_, _11383_);
  or _19731_ (_11414_, _11413_, _11411_);
  nor _19732_ (_11415_, _11414_, _11372_);
  nor _19733_ (_11416_, _11415_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _19734_ (_11417_, _11416_, _11352_);
  not _19735_ (_11418_, _11417_);
  and _19736_ (_11419_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _19737_ (_11420_, _09547_);
  and _19738_ (_11421_, _11420_, _07365_);
  and _19739_ (_11422_, _11421_, _11331_);
  and _19740_ (_11423_, _11422_, _11356_);
  not _19741_ (_11424_, _11423_);
  and _19742_ (_11425_, _11422_, _11375_);
  and _19743_ (_11426_, _11399_, _11339_);
  nor _19744_ (_11427_, _11426_, _11425_);
  and _19745_ (_11428_, _11427_, _11424_);
  and _19746_ (_11429_, _11382_, _11324_);
  and _19747_ (_11430_, _11364_, _11316_);
  and _19748_ (_11431_, _11430_, _11289_);
  nor _19749_ (_11432_, _11431_, _11429_);
  and _19750_ (_11433_, _11339_, _11319_);
  and _19751_ (_11435_, _11430_, _11422_);
  nor _19752_ (_11436_, _11435_, _11433_);
  and _19753_ (_11437_, _11399_, _11382_);
  and _19754_ (_11438_, _11374_, _11316_);
  and _19755_ (_11439_, _11438_, _11382_);
  nor _19756_ (_11440_, _11439_, _11437_);
  and _19757_ (_11441_, _11440_, _11436_);
  and _19758_ (_11442_, _11441_, _11432_);
  and _19759_ (_11443_, _11442_, _11428_);
  not _19760_ (_11444_, _11443_);
  nor _19761_ (_11445_, _11403_, _11359_);
  not _19762_ (_11446_, _11422_);
  nor _19763_ (_11447_, _11446_, _11445_);
  or _19764_ (_11448_, _11375_, _11313_);
  and _19765_ (_11449_, _11448_, _11382_);
  or _19766_ (_11450_, _11449_, _11447_);
  and _19767_ (_11451_, _11322_, _11316_);
  and _19768_ (_11452_, _11422_, _11451_);
  and _19769_ (_11453_, _11438_, _11422_);
  nor _19770_ (_11454_, _11453_, _11452_);
  and _19771_ (_11455_, _11382_, _11328_);
  and _19772_ (_11456_, _11403_, _11289_);
  nor _19773_ (_11457_, _11456_, _11455_);
  nand _19774_ (_11458_, _11457_, _11454_);
  or _19775_ (_11459_, _11458_, _11450_);
  and _19776_ (_11460_, _11451_, _11289_);
  and _19777_ (_11461_, _11422_, _11328_);
  and _19778_ (_11462_, _11394_, _11316_);
  and _19779_ (_11463_, _11462_, _11317_);
  or _19780_ (_11464_, _11463_, _11461_);
  or _19781_ (_11466_, _11464_, _11460_);
  and _19782_ (_11467_, _11389_, _11316_);
  and _19783_ (_11468_, _11467_, _11422_);
  and _19784_ (_11469_, _11422_, _11312_);
  and _19785_ (_11470_, _11469_, _11305_);
  or _19786_ (_11471_, _11470_, _11468_);
  and _19787_ (_11472_, _11355_, _11316_);
  and _19788_ (_11473_, _11472_, _11422_);
  and _19789_ (_11474_, _11382_, _11319_);
  or _19790_ (_11475_, _11474_, _11473_);
  or _19791_ (_11476_, _11475_, _11471_);
  and _19792_ (_11477_, _11374_, _11339_);
  nor _19793_ (_11478_, _11330_, _11312_);
  and _19794_ (_11479_, _11478_, _11305_);
  and _19795_ (_11480_, _11479_, _11294_);
  or _19796_ (_11481_, _11480_, _11477_);
  or _19797_ (_11482_, _11481_, _11383_);
  or _19798_ (_11483_, _11482_, _11363_);
  or _19799_ (_11484_, _11483_, _11476_);
  or _19800_ (_11485_, _11484_, _11466_);
  or _19801_ (_11488_, _11485_, _11459_);
  nor _19802_ (_11489_, _11488_, _11444_);
  nor _19803_ (_11490_, _11489_, _11283_);
  nor _19804_ (_11491_, _11490_, _11413_);
  and _19805_ (_11492_, _11491_, _11371_);
  nor _19806_ (_11493_, _11492_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor _19807_ (_11494_, _11493_, _11419_);
  and _19808_ (_11495_, _11494_, _11418_);
  and _19809_ (_11496_, _11495_, _11351_);
  and _19810_ (_11497_, _11496_, _11280_);
  nor _19811_ (_11498_, _11494_, _11418_);
  and _19812_ (_11499_, _11351_, _11498_);
  nor _19813_ (_11500_, _07325_, _06657_);
  and _19814_ (_11501_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and _19815_ (_11502_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _19816_ (_11503_, _11502_, _11501_);
  and _19817_ (_11504_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _19818_ (_11505_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor _19819_ (_11506_, _11505_, _11504_);
  and _19820_ (_11507_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _19821_ (_11508_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _19822_ (_11509_, _11508_, _11507_);
  and _19823_ (_11510_, _11509_, _11506_);
  and _19824_ (_11511_, _11510_, _11503_);
  nor _19825_ (_11512_, _11511_, _08477_);
  nor _19826_ (_11513_, _11512_, _11500_);
  not _19827_ (_11514_, _11513_);
  and _19828_ (_11515_, _11514_, _11499_);
  nor _19829_ (_11516_, _11515_, _11497_);
  nor _19830_ (_11517_, _11494_, _11417_);
  and _19831_ (_11518_, _11351_, _11517_);
  and _19832_ (_11519_, _09239_, _07089_);
  not _19833_ (_11520_, _11519_);
  nor _19834_ (_11521_, _11520_, _07317_);
  and _19835_ (_11522_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor _19836_ (_11523_, _11521_, _11522_);
  and _19837_ (_11524_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and _19838_ (_11525_, _07106_, _06700_);
  not _19839_ (_11526_, _11525_);
  and _19840_ (_11527_, _11526_, _09213_);
  and _19841_ (_11528_, _11527_, _09210_);
  and _19842_ (_11529_, _11528_, _09202_);
  nor _19843_ (_11530_, _11529_, _11520_);
  nor _19844_ (_11531_, _11530_, _11524_);
  and _19845_ (_11532_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and _19846_ (_11533_, _11519_, _09009_);
  nor _19847_ (_11534_, _11533_, _11532_);
  nor _19848_ (_11535_, _11519_, _06508_);
  and _19849_ (_11536_, _11519_, _09599_);
  nor _19850_ (_11537_, _11536_, _11535_);
  and _19851_ (_11538_, _11537_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and _19852_ (_11539_, _11538_, _11534_);
  and _19853_ (_11540_, _11539_, _11531_);
  and _19854_ (_11541_, _11540_, _11523_);
  nor _19855_ (_11542_, _11540_, _11523_);
  nor _19856_ (_11543_, _11542_, _11541_);
  nor _19857_ (_11545_, _11543_, _06409_);
  nor _19858_ (_11546_, _11545_, _06438_);
  nor _19859_ (_11547_, _11546_, _11519_);
  nor _19860_ (_11548_, _11547_, _11521_);
  not _19861_ (_11549_, _11548_);
  and _19862_ (_11550_, _11549_, _11518_);
  not _19863_ (_11551_, _07319_);
  and _19864_ (_11552_, _11351_, _11417_);
  and _19865_ (_11553_, _11552_, _11494_);
  and _19866_ (_11554_, _11553_, _11551_);
  nor _19867_ (_11555_, _11554_, _11550_);
  and _19868_ (_11556_, _11555_, _11516_);
  nor _19869_ (_11557_, _11556_, _06448_);
  and _19870_ (_11558_, _11556_, _06448_);
  nor _19871_ (_11559_, _11558_, _11557_);
  not _19872_ (_11560_, _06499_);
  and _19873_ (_11561_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and _19874_ (_11562_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor _19875_ (_11563_, _11562_, _11561_);
  and _19876_ (_11564_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _19877_ (_11565_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  nor _19878_ (_11566_, _11565_, _11564_);
  and _19879_ (_11567_, _11566_, _11563_);
  and _19880_ (_11568_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _19881_ (_11569_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor _19882_ (_11570_, _11569_, _11568_);
  and _19883_ (_11571_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and _19884_ (_11572_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor _19885_ (_11573_, _11572_, _11571_);
  and _19886_ (_11574_, _11573_, _11570_);
  and _19887_ (_11575_, _11574_, _11567_);
  nor _19888_ (_11576_, _11575_, _07378_);
  not _19889_ (_11577_, _07040_);
  and _19890_ (_11578_, _07378_, _11577_);
  nor _19891_ (_11579_, _11578_, _11576_);
  not _19892_ (_11580_, _11579_);
  and _19893_ (_11581_, _11496_, _11580_);
  not _19894_ (_11582_, _11581_);
  and _19895_ (_11583_, _11519_, _07040_);
  nor _19896_ (_11584_, _11520_, _07260_);
  and _19897_ (_11585_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor _19898_ (_11586_, _11585_, _11584_);
  and _19899_ (_11587_, _11586_, _11541_);
  and _19900_ (_11588_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor _19901_ (_11589_, _11520_, _07118_);
  nor _19902_ (_11590_, _11589_, _11588_);
  and _19903_ (_11591_, _11590_, _11587_);
  and _19904_ (_11593_, _11520_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor _19905_ (_11594_, _11520_, _10970_);
  nor _19906_ (_11595_, _11594_, _11593_);
  and _19907_ (_11596_, _11595_, _11591_);
  nor _19908_ (_11597_, _11519_, _06487_);
  nor _19909_ (_11598_, _11597_, _11596_);
  and _19910_ (_11599_, _11597_, _11596_);
  or _19911_ (_11600_, _11599_, _11598_);
  nor _19912_ (_11601_, _11600_, _06409_);
  nor _19913_ (_11602_, _11519_, _06491_);
  not _19914_ (_11603_, _11602_);
  nor _19915_ (_11604_, _11603_, _11601_);
  nor _19916_ (_11605_, _11604_, _11583_);
  and _19917_ (_11606_, _11605_, _11517_);
  not _19918_ (_11607_, _11606_);
  not _19919_ (_11608_, _08479_);
  and _19920_ (_11609_, _11498_, _11608_);
  not _19921_ (_11610_, _11351_);
  nor _19922_ (_11611_, _11610_, _11609_);
  and _19923_ (_11612_, _11611_, _11607_);
  and _19924_ (_11613_, _11612_, _11582_);
  nor _19925_ (_11614_, _11613_, _11560_);
  and _19926_ (_11615_, _11613_, _11560_);
  nor _19927_ (_11616_, _11615_, _11614_);
  nor _19928_ (_11617_, _11495_, _11351_);
  not _19929_ (_11618_, _10806_);
  and _19930_ (_11619_, _11499_, _11618_);
  nor _19931_ (_11620_, _11619_, _11617_);
  nor _19932_ (_11621_, _11595_, _11591_);
  nor _19933_ (_11622_, _11621_, _11596_);
  nor _19934_ (_11623_, _11622_, _06409_);
  nor _19935_ (_11624_, _11623_, _06455_);
  nor _19936_ (_11625_, _11624_, _11519_);
  nor _19937_ (_11626_, _11625_, _11594_);
  not _19938_ (_11627_, _11626_);
  and _19939_ (_11628_, _11627_, _11518_);
  and _19940_ (_11629_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and _19941_ (_11630_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor _19942_ (_11631_, _11630_, _11629_);
  and _19943_ (_11632_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _19944_ (_11634_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor _19945_ (_11635_, _11634_, _11632_);
  and _19946_ (_11636_, _11635_, _11631_);
  and _19947_ (_11637_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and _19948_ (_11638_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor _19949_ (_11639_, _11638_, _11637_);
  and _19950_ (_11640_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and _19951_ (_11641_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor _19952_ (_11642_, _11641_, _11640_);
  and _19953_ (_11643_, _11642_, _11639_);
  and _19954_ (_11644_, _11643_, _11636_);
  nor _19955_ (_11645_, _11644_, _07378_);
  not _19956_ (_11646_, _10970_);
  and _19957_ (_11647_, _11646_, _07378_);
  nor _19958_ (_11648_, _11647_, _11645_);
  not _19959_ (_11649_, _11648_);
  and _19960_ (_11650_, _11649_, _11496_);
  nor _19961_ (_11651_, _11650_, _11628_);
  and _19962_ (_11652_, _11651_, _11620_);
  nor _19963_ (_11653_, _11652_, _07452_);
  and _19964_ (_11654_, _11652_, _07452_);
  nor _19965_ (_11655_, _11654_, _11653_);
  and _19966_ (_11656_, _11655_, _11616_);
  nor _19967_ (_11657_, _07325_, _06600_);
  and _19968_ (_11658_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and _19969_ (_11659_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _19970_ (_11660_, _11659_, _11658_);
  and _19971_ (_11661_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _19972_ (_11662_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor _19973_ (_11663_, _11662_, _11661_);
  and _19974_ (_11664_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _19975_ (_11665_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _19976_ (_11666_, _11665_, _11664_);
  and _19977_ (_11667_, _11666_, _11663_);
  and _19978_ (_11668_, _11667_, _11660_);
  nor _19979_ (_11669_, _11668_, _08477_);
  nor _19980_ (_11670_, _11669_, _11657_);
  not _19981_ (_11671_, _11670_);
  and _19982_ (_11672_, _11671_, _11499_);
  not _19983_ (_11673_, _11498_);
  and _19984_ (_11674_, _11617_, _11673_);
  nor _19985_ (_11675_, _11674_, _11672_);
  nor _19986_ (_11676_, _11590_, _11587_);
  nor _19987_ (_11678_, _11676_, _11591_);
  nor _19988_ (_11679_, _11678_, _06409_);
  nor _19989_ (_11680_, _11679_, _06467_);
  nor _19990_ (_11681_, _11680_, _11519_);
  nor _19991_ (_11682_, _11681_, _11589_);
  not _19992_ (_11683_, _11682_);
  and _19993_ (_11684_, _11683_, _11518_);
  not _19994_ (_11685_, _07450_);
  and _19995_ (_11686_, _11496_, _11685_);
  nor _19996_ (_11687_, _11686_, _11684_);
  and _19997_ (_11688_, _11687_, _11675_);
  nor _19998_ (_11689_, _11688_, _06478_);
  and _19999_ (_11690_, _11688_, _06478_);
  nor _20000_ (_11691_, _11690_, _11689_);
  nor _20001_ (_11692_, _11586_, _11541_);
  nor _20002_ (_11693_, _11692_, _11587_);
  nor _20003_ (_11694_, _11693_, _06409_);
  nor _20004_ (_11695_, _11694_, _06413_);
  nor _20005_ (_11696_, _11695_, _11519_);
  nor _20006_ (_11697_, _11696_, _11584_);
  not _20007_ (_11698_, _11697_);
  and _20008_ (_11699_, _11698_, _11518_);
  and _20009_ (_11700_, _11610_, _11417_);
  nor _20010_ (_11701_, _11700_, _11699_);
  not _20011_ (_11702_, _07431_);
  and _20012_ (_11703_, _11496_, _11702_);
  nor _20013_ (_11704_, _07325_, _06628_);
  and _20014_ (_11705_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and _20015_ (_11706_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor _20016_ (_11707_, _11706_, _11705_);
  and _20017_ (_11708_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _20018_ (_11709_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor _20019_ (_11710_, _11709_, _11708_);
  and _20020_ (_11711_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _20021_ (_11712_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _20022_ (_11713_, _11712_, _11711_);
  and _20023_ (_11714_, _11713_, _11710_);
  and _20024_ (_11715_, _11714_, _11707_);
  nor _20025_ (_11716_, _11715_, _08477_);
  nor _20026_ (_11717_, _11716_, _11704_);
  not _20027_ (_11718_, _11717_);
  and _20028_ (_11719_, _11718_, _11499_);
  nor _20029_ (_11720_, _11719_, _11703_);
  and _20030_ (_11721_, _11553_, _07382_);
  not _20031_ (_11722_, _11721_);
  and _20032_ (_11723_, _11722_, _11720_);
  and _20033_ (_11724_, _11723_, _11701_);
  nor _20034_ (_11725_, _11724_, _07084_);
  and _20035_ (_11726_, _11724_, _07084_);
  nor _20036_ (_11727_, _11726_, _11725_);
  and _20037_ (_11728_, _11727_, _11691_);
  and _20038_ (_11729_, _11728_, _11656_);
  and _20039_ (_11730_, _11729_, _11559_);
  not _20040_ (_11731_, _11079_);
  and _20041_ (_11732_, _11496_, _11731_);
  and _20042_ (_11733_, _11495_, _11610_);
  nor _20043_ (_11734_, _11538_, _11534_);
  nor _20044_ (_11735_, _11734_, _11539_);
  nor _20045_ (_11736_, _11735_, _06409_);
  nor _20046_ (_11737_, _11736_, _06528_);
  nor _20047_ (_11738_, _11737_, _11519_);
  nor _20048_ (_11739_, _11738_, _11533_);
  not _20049_ (_11740_, _11739_);
  and _20050_ (_11741_, _11740_, _11518_);
  or _20051_ (_11742_, _11741_, _11733_);
  and _20052_ (_11743_, _11553_, _09547_);
  not _20053_ (_11744_, _11221_);
  and _20054_ (_11745_, _11499_, _11744_);
  or _20055_ (_11746_, _11745_, _11743_);
  or _20056_ (_11747_, _11746_, _11742_);
  nor _20057_ (_11748_, _11747_, _11732_);
  nor _20058_ (_11749_, _11748_, _06537_);
  and _20059_ (_11750_, _11748_, _06537_);
  nor _20060_ (_11751_, _11750_, _11749_);
  and _20061_ (_11752_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _20062_ (_11753_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor _20063_ (_11754_, _11753_, _11752_);
  and _20064_ (_11755_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and _20065_ (_11756_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor _20066_ (_11757_, _11756_, _11755_);
  and _20067_ (_11758_, _11757_, _11754_);
  and _20068_ (_11759_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _20069_ (_11760_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor _20070_ (_11761_, _11760_, _11759_);
  and _20071_ (_11762_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and _20072_ (_11763_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  nor _20073_ (_11764_, _11763_, _11762_);
  and _20074_ (_11765_, _11764_, _11761_);
  and _20075_ (_11766_, _11765_, _11758_);
  nor _20076_ (_11767_, _11766_, _07378_);
  and _20077_ (_11768_, _09599_, _07378_);
  nor _20078_ (_11769_, _11768_, _11767_);
  not _20079_ (_11770_, _11769_);
  and _20080_ (_11771_, _11770_, _11496_);
  nor _20081_ (_11772_, _07325_, _06737_);
  and _20082_ (_11773_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and _20083_ (_11774_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _20084_ (_11775_, _11774_, _11773_);
  and _20085_ (_11776_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _20086_ (_11777_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _20087_ (_11778_, _11777_, _11776_);
  and _20088_ (_11779_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _20089_ (_11780_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _20090_ (_11781_, _11780_, _11779_);
  and _20091_ (_11782_, _11781_, _11778_);
  and _20092_ (_11783_, _11782_, _11775_);
  nor _20093_ (_11784_, _11783_, _08477_);
  nor _20094_ (_11785_, _11784_, _11772_);
  not _20095_ (_11786_, _11785_);
  and _20096_ (_11787_, _11786_, _11499_);
  nor _20097_ (_11788_, _11787_, _11771_);
  nor _20098_ (_11789_, _11537_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor _20099_ (_11790_, _11789_, _11538_);
  nor _20100_ (_11791_, _11790_, _06409_);
  nor _20101_ (_11792_, _11791_, _06509_);
  nor _20102_ (_11793_, _11792_, _11519_);
  nor _20103_ (_11794_, _11793_, _11536_);
  not _20104_ (_11795_, _11794_);
  and _20105_ (_11796_, _11795_, _11518_);
  and _20106_ (_11797_, _11553_, _07365_);
  nor _20107_ (_11798_, _11797_, _11796_);
  and _20108_ (_11799_, _11798_, _11788_);
  nor _20109_ (_11800_, _11799_, _06514_);
  and _20110_ (_11801_, _11799_, _06514_);
  or _20111_ (_11802_, _11801_, _11800_);
  nor _20112_ (_11803_, _11802_, _11751_);
  not _20113_ (_11804_, _06484_);
  and _20114_ (_11805_, _07396_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _20115_ (_11806_, _07404_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor _20116_ (_11807_, _11806_, _11805_);
  and _20117_ (_11808_, _07398_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _20118_ (_11809_, _07402_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor _20119_ (_11810_, _11809_, _11808_);
  and _20120_ (_11811_, _11810_, _11807_);
  and _20121_ (_11812_, _07389_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  and _20122_ (_11813_, _07392_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor _20123_ (_11814_, _11813_, _11812_);
  and _20124_ (_11815_, _07380_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and _20125_ (_11816_, _07385_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _20126_ (_11817_, _11816_, _11815_);
  and _20127_ (_11818_, _11817_, _11814_);
  and _20128_ (_11819_, _11818_, _11811_);
  nor _20129_ (_11820_, _11819_, _07378_);
  not _20130_ (_11821_, _11529_);
  and _20131_ (_11822_, _11821_, _07378_);
  nor _20132_ (_11823_, _11822_, _11820_);
  not _20133_ (_11824_, _11823_);
  and _20134_ (_11825_, _11824_, _11496_);
  nor _20135_ (_11827_, _07325_, _06685_);
  and _20136_ (_11828_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and _20137_ (_11829_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor _20138_ (_11830_, _11829_, _11828_);
  and _20139_ (_11832_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and _20140_ (_11833_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor _20141_ (_11834_, _11833_, _11832_);
  and _20142_ (_11835_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _20143_ (_11836_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor _20144_ (_11837_, _11836_, _11835_);
  and _20145_ (_11838_, _11837_, _11834_);
  and _20146_ (_11839_, _11838_, _11830_);
  nor _20147_ (_11840_, _11839_, _08477_);
  nor _20148_ (_11841_, _11840_, _11827_);
  not _20149_ (_11842_, _11841_);
  and _20150_ (_11843_, _11842_, _11499_);
  nor _20151_ (_11844_, _11843_, _11825_);
  nor _20152_ (_11845_, _11539_, _11531_);
  nor _20153_ (_11846_, _11845_, _11540_);
  nor _20154_ (_11848_, _11846_, _06409_);
  nor _20155_ (_11849_, _11848_, _06517_);
  nor _20156_ (_11850_, _11849_, _11519_);
  nor _20157_ (_11851_, _11850_, _11530_);
  not _20158_ (_11852_, _11851_);
  and _20159_ (_11853_, _11852_, _11518_);
  and _20160_ (_11855_, _11553_, _09388_);
  nor _20161_ (_11856_, _11855_, _11853_);
  and _20162_ (_11857_, _11856_, _11844_);
  nor _20163_ (_11858_, _11857_, _06525_);
  and _20164_ (_11859_, _11857_, _06525_);
  nor _20165_ (_11860_, _11859_, _11858_);
  nor _20166_ (_11861_, _11860_, _11804_);
  and _20167_ (_11862_, _11861_, _11803_);
  and _20168_ (_11863_, _11862_, _11730_);
  nor _20169_ (_11864_, _06499_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _20170_ (_11865_, _11864_, _11863_);
  not _20171_ (_11866_, _11865_);
  not _20172_ (_11867_, _11344_);
  and _20173_ (_11868_, _11344_, _11295_);
  nor _20174_ (_11869_, _11868_, _11363_);
  nor _20175_ (_11870_, _11869_, _11353_);
  and _20176_ (_11871_, _11870_, _11867_);
  nor _20177_ (_11872_, _06984_, _06539_);
  and _20178_ (_11873_, _11872_, _11730_);
  and _20179_ (_11874_, _11873_, _11871_);
  not _20180_ (_11875_, _11342_);
  not _20181_ (_11876_, _06849_);
  and _20182_ (_11877_, _06898_, _11876_);
  nor _20183_ (_11878_, _06898_, _11876_);
  nor _20184_ (_11879_, _11878_, _11877_);
  not _20185_ (_11880_, _11879_);
  or _20186_ (_11881_, _08089_, _06881_);
  nor _20187_ (_11882_, _11881_, _06878_);
  and _20188_ (_11883_, _11882_, _11867_);
  and _20189_ (_11884_, _11883_, _08405_);
  nand _20190_ (_11885_, _11884_, _08234_);
  nor _20191_ (_11886_, _11885_, _11368_);
  not _20192_ (_11887_, _08322_);
  and _20193_ (_11888_, _09100_, _11887_);
  and _20194_ (_11889_, _11888_, _11886_);
  and _20195_ (_11890_, _11889_, _11880_);
  not _20196_ (_11891_, _11890_);
  and _20197_ (_11892_, _11868_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  not _20198_ (_11894_, _11892_);
  nor _20199_ (_11895_, _11870_, _11867_);
  nor _20200_ (_11896_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor _20201_ (_11897_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _20202_ (_11898_, _11897_, _11896_);
  nor _20203_ (_11899_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor _20204_ (_11900_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _20205_ (_11901_, _11900_, _11899_);
  and _20206_ (_11902_, _11901_, _11898_);
  and _20207_ (_11903_, _11902_, _11895_);
  and _20208_ (_11904_, _11871_, _06776_);
  nor _20209_ (_11905_, _11904_, _11903_);
  and _20210_ (_11906_, _11905_, _11894_);
  and _20211_ (_11907_, _11906_, _11891_);
  and _20212_ (_11908_, _11331_, _11420_);
  and _20213_ (_11909_, _11908_, _11399_);
  nor _20214_ (_11910_, _11909_, _11425_);
  and _20215_ (_11911_, _11287_, _11312_);
  and _20216_ (_11912_, _11911_, _11374_);
  and _20217_ (_11913_, _11360_, _11312_);
  nor _20218_ (_11914_, _11913_, _11912_);
  and _20219_ (_11915_, _11914_, _11910_);
  not _20220_ (_11916_, _11339_);
  nor _20221_ (_11917_, _11403_, _11324_);
  nor _20222_ (_11918_, _11917_, _11916_);
  and _20223_ (_11919_, _11911_, _11317_);
  nor _20224_ (_11920_, _11919_, _11400_);
  not _20225_ (_11921_, _11920_);
  nor _20226_ (_11922_, _11921_, _11918_);
  and _20227_ (_11923_, _11922_, _11915_);
  and _20228_ (_11924_, _11923_, _11907_);
  or _20229_ (_11925_, _11430_, _11451_);
  nand _20230_ (_11926_, _11925_, _11339_);
  and _20231_ (_11927_, _11359_, _11316_);
  and _20232_ (_11928_, _11927_, _11339_);
  or _20233_ (_11929_, _11928_, _11358_);
  nor _20234_ (_11930_, _11907_, _11929_);
  and _20235_ (_11931_, _11930_, _11926_);
  nor _20236_ (_11932_, _11931_, _11924_);
  not _20237_ (_11933_, _11932_);
  and _20238_ (_11934_, _11290_, _11312_);
  and _20239_ (_11935_, _11322_, _11934_);
  and _20240_ (_11936_, _11328_, _11339_);
  nor _20241_ (_11937_, _11936_, _11935_);
  and _20242_ (_11938_, _11937_, _11933_);
  nor _20243_ (_11939_, _11938_, _11875_);
  and _20244_ (_11940_, _11421_, _11288_);
  and _20245_ (_11941_, _11355_, _11382_);
  nor _20246_ (_11942_, _11941_, _11940_);
  nor _20247_ (_11943_, _11942_, _11283_);
  and _20248_ (_11944_, _11383_, _11341_);
  nor _20249_ (_11945_, _11944_, _11943_);
  not _20250_ (_11946_, _11945_);
  nor _20251_ (_11947_, _11946_, _11939_);
  nand _20252_ (_11948_, _08041_, _08125_);
  and _20253_ (_11949_, _11948_, _11895_);
  nor _20254_ (_11950_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not _20255_ (_11951_, _11950_);
  nor _20256_ (_11952_, _06448_, _06463_);
  and _20257_ (_11953_, _11952_, _07085_);
  and _20258_ (_11954_, _11953_, _06500_);
  or _20259_ (_11955_, _11954_, _11951_);
  nor _20260_ (_11956_, _11955_, _07291_);
  not _20261_ (_11957_, _11956_);
  and _20262_ (_11958_, _11957_, _11868_);
  nor _20263_ (_11959_, _11958_, _11949_);
  not _20264_ (_11960_, _11959_);
  nor _20265_ (_11961_, _11960_, _11947_);
  not _20266_ (_11962_, _11961_);
  nor _20267_ (_11963_, _11962_, _11874_);
  and _20268_ (_11964_, _11963_, _11866_);
  nor _20269_ (_11965_, _11964_, _11279_);
  not _20270_ (_11966_, _09145_);
  and _20271_ (_11968_, _11342_, _11325_);
  nor _20272_ (_11969_, _11968_, _11943_);
  nand _20273_ (_11970_, _11910_, _11361_);
  or _20274_ (_11971_, _11970_, _11921_);
  and _20275_ (_11972_, _11971_, _11342_);
  not _20276_ (_11973_, _11972_);
  and _20277_ (_11974_, _11941_, _11282_);
  nor _20278_ (_11975_, _11974_, _11413_);
  and _20279_ (_11976_, _11975_, _11973_);
  nor _20280_ (_11977_, _11912_, _11369_);
  and _20281_ (_11978_, _11977_, _11937_);
  nor _20282_ (_11979_, _11978_, _11875_);
  not _20283_ (_11980_, _11979_);
  nand _20284_ (_11981_, _11360_, _11282_);
  and _20285_ (_11982_, _11981_, _11973_);
  and _20286_ (_11983_, _11982_, _11980_);
  and _20287_ (_11984_, _11983_, _11976_);
  and _20288_ (_11985_, _11984_, _11969_);
  or _20289_ (_11986_, _11985_, _11968_);
  and _20290_ (_11987_, _11986_, _11966_);
  not _20291_ (_11988_, _11974_);
  not _20292_ (_11989_, _11413_);
  and _20293_ (_11990_, _11981_, _11989_);
  and _20294_ (_11991_, _11990_, _11988_);
  and _20295_ (_11992_, _11991_, _11973_);
  and _20296_ (_11993_, _11992_, _11670_);
  nand _20297_ (_11994_, _11991_, _11973_);
  and _20298_ (_11995_, _07490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  and _20299_ (_11996_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20300_ (_11998_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and _20301_ (_11999_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor _20302_ (_12001_, _11999_, _11998_);
  and _20303_ (_12002_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and _20304_ (_12003_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor _20305_ (_12004_, _12003_, _12002_);
  and _20306_ (_12005_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _20307_ (_12006_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor _20308_ (_12007_, _12006_, _12005_);
  and _20309_ (_12008_, _12007_, _12004_);
  and _20310_ (_12009_, _12008_, _12001_);
  nor _20311_ (_12010_, _12009_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20312_ (_12011_, _12010_, _11996_);
  nor _20313_ (_12012_, _12011_, _07490_);
  nor _20314_ (_12013_, _12012_, _11995_);
  and _20315_ (_12014_, _12013_, _11994_);
  nor _20316_ (_12015_, _12014_, _11993_);
  and _20317_ (_12016_, _12015_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _20318_ (_12017_, _12015_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _20319_ (_12018_, _12017_, _12016_);
  and _20320_ (_12019_, _11992_, _11717_);
  and _20321_ (_12020_, _07490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  and _20322_ (_12021_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20323_ (_12022_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _20324_ (_12023_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor _20325_ (_12024_, _12023_, _12022_);
  and _20326_ (_12025_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and _20327_ (_12026_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor _20328_ (_12027_, _12026_, _12025_);
  and _20329_ (_12028_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and _20330_ (_12029_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor _20331_ (_12030_, _12029_, _12028_);
  and _20332_ (_12031_, _12030_, _12027_);
  and _20333_ (_12032_, _12031_, _12024_);
  nor _20334_ (_12033_, _12032_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20335_ (_12034_, _12033_, _12021_);
  nor _20336_ (_12035_, _12034_, _07490_);
  nor _20337_ (_12036_, _12035_, _12020_);
  and _20338_ (_12037_, _12036_, _11994_);
  nor _20339_ (_12038_, _12037_, _12019_);
  nand _20340_ (_12040_, _12038_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _20341_ (_12041_, _11992_, _11513_);
  and _20342_ (_12042_, _07490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and _20343_ (_12043_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20344_ (_12044_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _20345_ (_12045_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor _20346_ (_12046_, _12045_, _12044_);
  and _20347_ (_12047_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and _20348_ (_12048_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor _20349_ (_12049_, _12048_, _12047_);
  and _20350_ (_12050_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and _20351_ (_12051_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor _20352_ (_12053_, _12051_, _12050_);
  and _20353_ (_12054_, _12053_, _12049_);
  and _20354_ (_12055_, _12054_, _12046_);
  nor _20355_ (_12056_, _12055_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20356_ (_12058_, _12056_, _12043_);
  nor _20357_ (_12059_, _12058_, _07490_);
  nor _20358_ (_12061_, _12059_, _12042_);
  and _20359_ (_12062_, _12061_, _11994_);
  nor _20360_ (_12063_, _12062_, _12041_);
  nor _20361_ (_12064_, _12063_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _20362_ (_12065_, _12063_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _20363_ (_12066_, _11992_, _11841_);
  and _20364_ (_12067_, _11994_, _11207_);
  nor _20365_ (_12068_, _12067_, _12066_);
  and _20366_ (_12069_, _12068_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or _20367_ (_12070_, _11994_, _11744_);
  and _20368_ (_12071_, _07490_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and _20369_ (_12072_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20370_ (_12073_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _20371_ (_12074_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor _20372_ (_12076_, _12074_, _12073_);
  and _20373_ (_12077_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _20374_ (_12078_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor _20375_ (_12079_, _12078_, _12077_);
  and _20376_ (_12080_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _20377_ (_12081_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor _20378_ (_12083_, _12081_, _12080_);
  and _20379_ (_12084_, _12083_, _12079_);
  and _20380_ (_12086_, _12084_, _12076_);
  nor _20381_ (_12087_, _12086_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20382_ (_12088_, _12087_, _12072_);
  nor _20383_ (_12089_, _12088_, _07490_);
  nor _20384_ (_12090_, _12089_, _12071_);
  not _20385_ (_12091_, _12090_);
  or _20386_ (_12092_, _12091_, _11992_);
  nand _20387_ (_12093_, _12092_, _12070_);
  or _20388_ (_12094_, _12093_, _06714_);
  or _20389_ (_12095_, _11994_, _11786_);
  and _20390_ (_12096_, _07490_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and _20391_ (_12097_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20392_ (_12098_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and _20393_ (_12099_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor _20394_ (_12100_, _12099_, _12098_);
  and _20395_ (_12101_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _20396_ (_12102_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _20397_ (_12103_, _12102_, _12101_);
  and _20398_ (_12105_, _12103_, _12100_);
  and _20399_ (_12106_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _20400_ (_12107_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor _20401_ (_12108_, _12107_, _12106_);
  and _20402_ (_12109_, _12108_, _12105_);
  nor _20403_ (_12110_, _12109_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20404_ (_12111_, _12110_, _12097_);
  nor _20405_ (_12112_, _12111_, _07490_);
  nor _20406_ (_12113_, _12112_, _12096_);
  not _20407_ (_12114_, _12113_);
  or _20408_ (_12116_, _12114_, _11992_);
  and _20409_ (_12117_, _12116_, _12095_);
  and _20410_ (_12118_, _12117_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nand _20411_ (_12119_, _12093_, _06714_);
  and _20412_ (_12120_, _12119_, _12094_);
  and _20413_ (_12122_, _12120_, _12118_);
  not _20414_ (_12123_, _12122_);
  nand _20415_ (_12124_, _12123_, _12094_);
  nor _20416_ (_12125_, _12068_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _20417_ (_12126_, _12125_, _12069_);
  and _20418_ (_12127_, _12126_, _12124_);
  or _20419_ (_12129_, _12127_, _12069_);
  nor _20420_ (_12130_, _12129_, _12065_);
  nor _20421_ (_12131_, _12130_, _12064_);
  or _20422_ (_12132_, _12038_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _20423_ (_12134_, _12132_, _12040_);
  nand _20424_ (_12135_, _12134_, _12131_);
  nand _20425_ (_12136_, _12135_, _12040_);
  and _20426_ (_12137_, _12136_, _12018_);
  or _20427_ (_12138_, _12137_, _12016_);
  and _20428_ (_12139_, _11992_, _10806_);
  and _20429_ (_12140_, _07490_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and _20430_ (_12141_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _20431_ (_12142_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _20432_ (_12143_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor _20433_ (_12144_, _12143_, _12142_);
  and _20434_ (_12145_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and _20435_ (_12146_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _20436_ (_12147_, _12146_, _12145_);
  and _20437_ (_12148_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and _20438_ (_12149_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _20439_ (_12150_, _12149_, _12148_);
  and _20440_ (_12151_, _12150_, _12147_);
  and _20441_ (_12152_, _12151_, _12144_);
  nor _20442_ (_12153_, _12152_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _20443_ (_12154_, _12153_, _12141_);
  nor _20444_ (_12155_, _12154_, _07490_);
  nor _20445_ (_12156_, _12155_, _12140_);
  and _20446_ (_12157_, _12156_, _11994_);
  nor _20447_ (_12158_, _12157_, _12139_);
  nand _20448_ (_12159_, _12158_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or _20449_ (_12161_, _12158_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and _20450_ (_12162_, _12161_, _12159_);
  nand _20451_ (_12163_, _12162_, _12138_);
  or _20452_ (_12164_, _12162_, _12138_);
  nor _20453_ (_12165_, _11979_, _11972_);
  and _20454_ (_12166_, _11981_, _12165_);
  and _20455_ (_12167_, _11342_, _11935_);
  nor _20456_ (_12168_, _12167_, _11943_);
  nor _20457_ (_12169_, _12168_, _11994_);
  nor _20458_ (_12171_, _12169_, _12166_);
  and _20459_ (_12172_, _12171_, _12164_);
  and _20460_ (_12173_, _12172_, _12163_);
  nor _20461_ (_12174_, _12156_, _11988_);
  and _20462_ (_12175_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _20463_ (_12176_, _12169_, _12165_);
  and _20464_ (_12177_, _12176_, _11618_);
  or _20465_ (_12178_, _12177_, _12175_);
  or _20466_ (_12179_, _12178_, _12174_);
  or _20467_ (_12180_, _12179_, _12173_);
  or _20468_ (_12181_, _12180_, _11987_);
  and _20469_ (_12182_, _12181_, _11964_);
  or _20470_ (_12183_, _12182_, _11965_);
  and _20471_ (_09791_, _12183_, _06989_);
  and _20472_ (_12184_, _11240_, word_in[27]);
  not _20473_ (_12185_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor _20474_ (_12186_, _11231_, _12185_);
  and _20475_ (_12187_, _11231_, _09690_);
  or _20476_ (_12188_, _12187_, _12186_);
  and _20477_ (_12189_, _12188_, _11229_);
  and _20478_ (_12190_, _11227_, word_in[11]);
  or _20479_ (_12191_, _12190_, _11236_);
  or _20480_ (_12192_, _12191_, _12189_);
  or _20481_ (_12193_, _11242_, _09829_);
  and _20482_ (_12194_, _12193_, _11241_);
  and _20483_ (_12195_, _12194_, _12192_);
  or _20484_ (_14659_, _12195_, _12184_);
  nor _20485_ (_09795_, _11823_, rst);
  not _20486_ (_12196_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _20487_ (_12197_, _11231_, _12196_);
  and _20488_ (_12198_, _11231_, _09707_);
  or _20489_ (_12199_, _12198_, _12197_);
  and _20490_ (_12200_, _12199_, _11229_);
  and _20491_ (_12201_, _11227_, word_in[12]);
  or _20492_ (_12202_, _12201_, _11236_);
  or _20493_ (_12203_, _12202_, _12200_);
  or _20494_ (_12204_, _11242_, _09842_);
  and _20495_ (_12205_, _12204_, _11241_);
  and _20496_ (_12206_, _12205_, _12203_);
  and _20497_ (_12207_, _11240_, word_in[28]);
  or _20498_ (_14660_, _12207_, _12206_);
  not _20499_ (_12209_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor _20500_ (_12210_, _11231_, _12209_);
  and _20501_ (_12212_, _11231_, _09722_);
  or _20502_ (_12213_, _12212_, _12210_);
  and _20503_ (_12215_, _12213_, _11229_);
  and _20504_ (_12216_, _11227_, word_in[13]);
  or _20505_ (_12217_, _12216_, _11236_);
  or _20506_ (_12218_, _12217_, _12215_);
  or _20507_ (_12219_, _11242_, _09855_);
  and _20508_ (_12221_, _12219_, _11241_);
  and _20509_ (_12222_, _12221_, _12218_);
  and _20510_ (_12223_, _11240_, word_in[29]);
  or _20511_ (_14661_, _12223_, _12222_);
  and _20512_ (_12224_, _11240_, word_in[30]);
  not _20513_ (_12225_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor _20514_ (_12226_, _11231_, _12225_);
  and _20515_ (_12227_, _11231_, _09735_);
  or _20516_ (_12228_, _12227_, _12226_);
  and _20517_ (_12230_, _12228_, _11229_);
  and _20518_ (_12231_, _11227_, word_in[14]);
  or _20519_ (_12232_, _12231_, _11236_);
  or _20520_ (_12233_, _12232_, _12230_);
  or _20521_ (_12234_, _11242_, _09871_);
  and _20522_ (_12235_, _12234_, _11241_);
  and _20523_ (_12236_, _12235_, _12233_);
  or _20524_ (_14662_, _12236_, _12224_);
  or _20525_ (_12237_, _07808_, _07803_);
  or _20526_ (_12238_, _07794_, _07723_);
  nand _20527_ (_12239_, _12238_, _12237_);
  or _20528_ (_12240_, _12238_, _12237_);
  nand _20529_ (_12241_, _12240_, _12239_);
  nand _20530_ (_12242_, _12241_, _07814_);
  nand _20531_ (_12243_, _07810_, _07802_);
  nand _20532_ (_12244_, _12243_, _12242_);
  nand _20533_ (_12245_, _12244_, _07024_);
  and _20534_ (_12246_, _07818_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand _20535_ (_12247_, _12246_, _09090_);
  or _20536_ (_12248_, _09090_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand _20537_ (_12249_, _12248_, _12247_);
  nand _20538_ (_12250_, _12249_, _07027_);
  and _20539_ (_12251_, _11879_, _06845_);
  not _20540_ (_12252_, _12251_);
  nor _20541_ (_12253_, _11876_, _06834_);
  and _20542_ (_12254_, _11876_, _06834_);
  or _20543_ (_12255_, _12254_, _12253_);
  nor _20544_ (_12256_, _12255_, _06549_);
  nor _20545_ (_12257_, _08245_, _06914_);
  nor _20546_ (_12258_, _12257_, _06586_);
  and _20547_ (_12259_, _12257_, _06586_);
  nor _20548_ (_12260_, _12259_, _12258_);
  nor _20549_ (_12261_, _12260_, _06918_);
  nor _20550_ (_12262_, _08001_, _06810_);
  and _20551_ (_12263_, _06926_, _06778_);
  nor _20552_ (_12264_, _12263_, _12262_);
  and _20553_ (_12265_, _06951_, _06957_);
  and _20554_ (_12266_, _06949_, _06924_);
  nor _20555_ (_12267_, _12266_, _12265_);
  and _20556_ (_12268_, _12267_, _12264_);
  and _20557_ (_12269_, _12268_, _07023_);
  and _20558_ (_12270_, _12269_, _07020_);
  not _20559_ (_12271_, _12270_);
  nor _20560_ (_12272_, _12271_, _12261_);
  and _20561_ (_12273_, _12272_, _07016_);
  not _20562_ (_12274_, _12273_);
  nor _20563_ (_12275_, _12274_, _12256_);
  and _20564_ (_12276_, _12275_, _12252_);
  and _20565_ (_12277_, _12276_, _12250_);
  nand _20566_ (_12278_, _12277_, _12245_);
  nand _20567_ (_12279_, _12278_, _08045_);
  nor _20568_ (_12280_, _06539_, _06592_);
  nor _20569_ (_12281_, _12280_, _06969_);
  nor _20570_ (_12282_, _12281_, _08043_);
  nor _20571_ (_12283_, _11948_, _06592_);
  or _20572_ (_12284_, _12283_, _07699_);
  nor _20573_ (_12285_, _12284_, _12282_);
  nand _20574_ (_12286_, _12285_, _12279_);
  and _20575_ (_12287_, _06951_, _06847_);
  and _20576_ (_12288_, _06958_, _07003_);
  nor _20577_ (_12289_, _09262_, _09104_);
  not _20578_ (_12290_, _12289_);
  and _20579_ (_12291_, _12290_, _09256_);
  nor _20580_ (_12292_, _12291_, _06847_);
  and _20581_ (_12293_, _12291_, _06847_);
  nor _20582_ (_12294_, _12293_, _12292_);
  and _20583_ (_12295_, _12294_, _06997_);
  nor _20584_ (_12296_, _06778_, _06597_);
  nor _20585_ (_12297_, _12296_, _06919_);
  nor _20586_ (_12298_, _12297_, _06992_);
  or _20587_ (_12299_, _12298_, _12295_);
  or _20588_ (_12300_, _12299_, _12288_);
  and _20589_ (_12301_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor _20590_ (_12302_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not _20591_ (_12303_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _20592_ (_12304_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _12303_);
  nor _20593_ (_12305_, _12304_, _12302_);
  nand _20594_ (_12306_, _12305_, _09275_);
  or _20595_ (_12307_, _12305_, _09275_);
  and _20596_ (_12308_, _12307_, _06548_);
  and _20597_ (_12309_, _12308_, _12306_);
  and _20598_ (_12310_, _09550_, _07027_);
  or _20599_ (_12311_, _12310_, _12309_);
  or _20600_ (_12312_, _12311_, _12301_);
  or _20601_ (_12313_, _12312_, _12300_);
  or _20602_ (_12314_, _12313_, _12287_);
  or _20603_ (_12315_, _12314_, _07700_);
  and _20604_ (_12316_, _12315_, _12286_);
  and _20605_ (_09804_, _12316_, _06989_);
  and _20606_ (_12317_, _11240_, word_in[31]);
  nor _20607_ (_12318_, _11231_, _08663_);
  and _20608_ (_12319_, _11231_, _08953_);
  or _20609_ (_12320_, _12319_, _12318_);
  and _20610_ (_12321_, _12320_, _11229_);
  and _20611_ (_12322_, _11227_, word_in[15]);
  or _20612_ (_12323_, _12322_, _11236_);
  or _20613_ (_12324_, _12323_, _12321_);
  or _20614_ (_12325_, _11242_, _08942_);
  and _20615_ (_12326_, _12325_, _11241_);
  and _20616_ (_12327_, _12326_, _12324_);
  or _20617_ (_14663_, _12327_, _12317_);
  or _20618_ (_12328_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand _20619_ (_12329_, _07493_, _10755_);
  and _20620_ (_12330_, _12329_, _06989_);
  and _20621_ (_09812_, _12330_, _12328_);
  and _20622_ (_12331_, _08939_, _08711_);
  and _20623_ (_12332_, _08944_, _09447_);
  not _20624_ (_12333_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _20625_ (_12334_, _09627_, _08950_);
  nor _20626_ (_12335_, _12334_, _12333_);
  and _20627_ (_12336_, _12334_, _09636_);
  or _20628_ (_12337_, _12336_, _12335_);
  or _20629_ (_12338_, _12337_, _12332_);
  not _20630_ (_12339_, _12332_);
  or _20631_ (_12340_, _12339_, word_in[8]);
  and _20632_ (_12341_, _12340_, _12338_);
  or _20633_ (_12342_, _12341_, _12331_);
  not _20634_ (_12343_, _08879_);
  and _20635_ (_12344_, _10150_, _12343_);
  and _20636_ (_12345_, _12344_, _08740_);
  not _20637_ (_12346_, _12345_);
  not _20638_ (_12347_, _12331_);
  or _20639_ (_12348_, _12347_, _09648_);
  and _20640_ (_12349_, _12348_, _12346_);
  and _20641_ (_12350_, _12349_, _12342_);
  and _20642_ (_12351_, _12345_, _10171_);
  or _20643_ (_09864_, _12351_, _12350_);
  not _20644_ (_12352_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _20645_ (_12353_, _12334_, _12352_);
  and _20646_ (_12354_, _12334_, word_in[1]);
  or _20647_ (_12355_, _12354_, _12353_);
  and _20648_ (_12356_, _12355_, _12339_);
  and _20649_ (_12357_, _12332_, word_in[9]);
  or _20650_ (_12358_, _12357_, _12356_);
  and _20651_ (_12359_, _12358_, _12347_);
  and _20652_ (_12360_, _12331_, _09801_);
  or _20653_ (_12361_, _12360_, _12359_);
  and _20654_ (_12362_, _12361_, _12346_);
  and _20655_ (_12363_, _12345_, _09656_);
  or _20656_ (_09867_, _12363_, _12362_);
  or _20657_ (_12364_, _12347_, _09816_);
  not _20658_ (_12365_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _20659_ (_12366_, _12334_, _12365_);
  and _20660_ (_12367_, _12334_, _09674_);
  or _20661_ (_12368_, _12367_, _12366_);
  or _20662_ (_12369_, _12368_, _12332_);
  or _20663_ (_12370_, _12339_, word_in[10]);
  and _20664_ (_12371_, _12370_, _12369_);
  or _20665_ (_12372_, _12371_, _12331_);
  and _20666_ (_12374_, _12372_, _12364_);
  or _20667_ (_12375_, _12374_, _12345_);
  or _20668_ (_12376_, _12346_, _09685_);
  and _20669_ (_09869_, _12376_, _12375_);
  or _20670_ (_12377_, _12347_, _09829_);
  not _20671_ (_12378_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _20672_ (_12379_, _12334_, _12378_);
  and _20673_ (_12380_, _12334_, _09690_);
  or _20674_ (_12381_, _12380_, _12379_);
  or _20675_ (_12382_, _12381_, _12332_);
  or _20676_ (_12383_, _12339_, word_in[11]);
  and _20677_ (_12384_, _12383_, _12382_);
  or _20678_ (_12385_, _12384_, _12331_);
  and _20679_ (_12386_, _12385_, _12377_);
  or _20680_ (_12388_, _12386_, _12345_);
  or _20681_ (_12389_, _12346_, _09701_);
  and _20682_ (_09874_, _12389_, _12388_);
  not _20683_ (_12390_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _20684_ (_12391_, _12334_, _12390_);
  and _20685_ (_12392_, _12334_, word_in[4]);
  or _20686_ (_12393_, _12392_, _12391_);
  and _20687_ (_12394_, _12393_, _12339_);
  and _20688_ (_12395_, _12332_, word_in[12]);
  or _20689_ (_12396_, _12395_, _12394_);
  or _20690_ (_12397_, _12396_, _12331_);
  nor _20691_ (_12398_, _12347_, _09842_);
  nor _20692_ (_12399_, _12398_, _12345_);
  and _20693_ (_12400_, _12399_, _12397_);
  and _20694_ (_12401_, _12345_, _09703_);
  or _20695_ (_09877_, _12401_, _12400_);
  or _20696_ (_12402_, _12347_, _09855_);
  not _20697_ (_12403_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _20698_ (_12404_, _12334_, _12403_);
  and _20699_ (_12406_, _12334_, _09722_);
  or _20700_ (_12407_, _12406_, _12404_);
  or _20701_ (_12408_, _12407_, _12332_);
  or _20702_ (_12409_, _12339_, word_in[13]);
  and _20703_ (_12410_, _12409_, _12408_);
  or _20704_ (_12411_, _12410_, _12331_);
  and _20705_ (_12412_, _12411_, _12402_);
  or _20706_ (_12413_, _12412_, _12345_);
  or _20707_ (_12415_, _12346_, _09718_);
  and _20708_ (_09880_, _12415_, _12413_);
  or _20709_ (_12416_, _12347_, _09871_);
  not _20710_ (_12417_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _20711_ (_12418_, _12334_, _12417_);
  and _20712_ (_12419_, _12334_, _09735_);
  or _20713_ (_12420_, _12419_, _12418_);
  or _20714_ (_12421_, _12420_, _12332_);
  or _20715_ (_12422_, _12339_, word_in[14]);
  and _20716_ (_12424_, _12422_, _12421_);
  or _20717_ (_12425_, _12424_, _12331_);
  and _20718_ (_12426_, _12425_, _12416_);
  or _20719_ (_12427_, _12426_, _12345_);
  or _20720_ (_12428_, _12346_, _09745_);
  and _20721_ (_14664_, _12428_, _12427_);
  nor _20722_ (_12429_, _12334_, _08803_);
  and _20723_ (_12430_, _12334_, word_in[7]);
  or _20724_ (_12431_, _12430_, _12429_);
  and _20725_ (_12432_, _12431_, _12339_);
  and _20726_ (_12433_, _12332_, word_in[15]);
  or _20727_ (_12434_, _12433_, _12432_);
  and _20728_ (_12435_, _12434_, _12347_);
  and _20729_ (_12436_, _12331_, _08942_);
  or _20730_ (_12437_, _12436_, _12435_);
  and _20731_ (_12438_, _12437_, _12346_);
  and _20732_ (_12439_, _12345_, _10256_);
  or _20733_ (_09885_, _12439_, _12438_);
  nor _20734_ (_09919_, _11648_, rst);
  nor _20735_ (_09922_, _11785_, rst);
  nor _20736_ (_09929_, _11717_, rst);
  nor _20737_ (_09936_, _12090_, rst);
  and _20738_ (_12442_, _09768_, _08797_);
  not _20739_ (_12443_, _12442_);
  or _20740_ (_12444_, _12443_, word_in[8]);
  and _20741_ (_12446_, _08939_, _08713_);
  not _20742_ (_12447_, _12446_);
  not _20743_ (_12448_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _20744_ (_12449_, _09772_, _08950_);
  nor _20745_ (_12450_, _12449_, _12448_);
  and _20746_ (_12451_, _12449_, _09636_);
  or _20747_ (_12452_, _12451_, _12450_);
  or _20748_ (_12453_, _12452_, _12442_);
  and _20749_ (_12454_, _12453_, _12447_);
  and _20750_ (_12455_, _12454_, _12444_);
  and _20751_ (_12456_, _12344_, _08711_);
  and _20752_ (_12457_, _12446_, _09648_);
  or _20753_ (_12458_, _12457_, _12456_);
  or _20754_ (_12459_, _12458_, _12455_);
  not _20755_ (_12460_, _12456_);
  or _20756_ (_12461_, _12460_, word_in[24]);
  and _20757_ (_14665_, _12461_, _12459_);
  or _20758_ (_12462_, _12443_, word_in[9]);
  not _20759_ (_12463_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _20760_ (_12464_, _12449_, _12463_);
  and _20761_ (_12465_, _12449_, _09660_);
  or _20762_ (_12466_, _12465_, _12464_);
  or _20763_ (_12467_, _12466_, _12442_);
  and _20764_ (_12468_, _12467_, _12447_);
  and _20765_ (_12469_, _12468_, _12462_);
  and _20766_ (_12470_, _12446_, _09801_);
  or _20767_ (_12471_, _12470_, _12456_);
  or _20768_ (_12472_, _12471_, _12469_);
  or _20769_ (_12473_, _12460_, word_in[25]);
  and _20770_ (_09956_, _12473_, _12472_);
  not _20771_ (_12474_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _20772_ (_12476_, _12449_, _12474_);
  and _20773_ (_12477_, _12449_, _09674_);
  nor _20774_ (_12479_, _12477_, _12476_);
  nor _20775_ (_12480_, _12479_, _12442_);
  and _20776_ (_12481_, _12442_, word_in[10]);
  or _20777_ (_12482_, _12481_, _12480_);
  and _20778_ (_12483_, _12482_, _12447_);
  and _20779_ (_12484_, _12446_, _09816_);
  or _20780_ (_12485_, _12484_, _12456_);
  or _20781_ (_12486_, _12485_, _12483_);
  or _20782_ (_12487_, _12460_, word_in[26]);
  and _20783_ (_09961_, _12487_, _12486_);
  not _20784_ (_12488_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _20785_ (_12489_, _12449_, _12488_);
  and _20786_ (_12490_, _12449_, _09690_);
  nor _20787_ (_12491_, _12490_, _12489_);
  nor _20788_ (_12492_, _12491_, _12442_);
  and _20789_ (_12493_, _12442_, word_in[11]);
  or _20790_ (_12494_, _12493_, _12492_);
  and _20791_ (_12495_, _12494_, _12447_);
  and _20792_ (_12496_, _12446_, _09829_);
  or _20793_ (_12497_, _12496_, _12456_);
  or _20794_ (_12498_, _12497_, _12495_);
  or _20795_ (_12499_, _12460_, word_in[27]);
  and _20796_ (_09963_, _12499_, _12498_);
  or _20797_ (_12500_, _12443_, word_in[12]);
  not _20798_ (_12501_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _20799_ (_12502_, _12449_, _12501_);
  and _20800_ (_12503_, _12449_, _09707_);
  or _20801_ (_12504_, _12503_, _12502_);
  or _20802_ (_12505_, _12504_, _12442_);
  and _20803_ (_12506_, _12505_, _12447_);
  and _20804_ (_12507_, _12506_, _12500_);
  and _20805_ (_12508_, _12446_, _09842_);
  or _20806_ (_12509_, _12508_, _12456_);
  or _20807_ (_12510_, _12509_, _12507_);
  or _20808_ (_12511_, _12460_, word_in[28]);
  and _20809_ (_09967_, _12511_, _12510_);
  or _20810_ (_12512_, _12443_, word_in[13]);
  not _20811_ (_12513_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _20812_ (_12514_, _12449_, _12513_);
  and _20813_ (_12515_, _12449_, _09722_);
  or _20814_ (_12516_, _12515_, _12514_);
  or _20815_ (_12517_, _12516_, _12442_);
  and _20816_ (_12518_, _12517_, _12447_);
  and _20817_ (_12519_, _12518_, _12512_);
  and _20818_ (_12520_, _12446_, _09855_);
  or _20819_ (_12521_, _12520_, _12456_);
  or _20820_ (_12522_, _12521_, _12519_);
  or _20821_ (_12523_, _12460_, word_in[29]);
  and _20822_ (_09971_, _12523_, _12522_);
  not _20823_ (_12524_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _20824_ (_12525_, _12449_, _12524_);
  and _20825_ (_12526_, _12449_, _09735_);
  nor _20826_ (_12527_, _12526_, _12525_);
  nor _20827_ (_12528_, _12527_, _12442_);
  and _20828_ (_12529_, _12442_, word_in[14]);
  or _20829_ (_12530_, _12529_, _12528_);
  and _20830_ (_12531_, _12530_, _12447_);
  and _20831_ (_12532_, _12446_, _09871_);
  or _20832_ (_12533_, _12532_, _12456_);
  or _20833_ (_12534_, _12533_, _12531_);
  or _20834_ (_12535_, _12460_, word_in[30]);
  and _20835_ (_09973_, _12535_, _12534_);
  and _20836_ (_09976_, t2_i, _06989_);
  or _20837_ (_12536_, _12443_, word_in[15]);
  nor _20838_ (_12537_, _12449_, _08669_);
  and _20839_ (_12538_, _12449_, _08953_);
  or _20840_ (_12539_, _12538_, _12537_);
  or _20841_ (_12540_, _12539_, _12442_);
  and _20842_ (_12541_, _12540_, _12447_);
  and _20843_ (_12542_, _12541_, _12536_);
  and _20844_ (_12543_, _12446_, _08942_);
  or _20845_ (_12544_, _12543_, _12456_);
  or _20846_ (_12545_, _12544_, _12542_);
  or _20847_ (_12546_, _12460_, word_in[31]);
  and _20848_ (_09978_, _12546_, _12545_);
  nor _20849_ (_09999_, _12113_, rst);
  or _20850_ (_12547_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  not _20851_ (_12549_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nand _20852_ (_12550_, _07493_, _12549_);
  and _20853_ (_12551_, _12550_, _06989_);
  and _20854_ (_10020_, _12551_, _12547_);
  and _20855_ (_12552_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and _20856_ (_12553_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  or _20857_ (_12554_, _12553_, _12552_);
  and _20858_ (_10025_, _12554_, _06989_);
  or _20859_ (_12555_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not _20860_ (_12556_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand _20861_ (_12557_, _07493_, _12556_);
  and _20862_ (_12558_, _12557_, _06989_);
  and _20863_ (_10029_, _12558_, _12555_);
  and _20864_ (_12559_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and _20865_ (_12560_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or _20866_ (_12561_, _12560_, _12559_);
  and _20867_ (_10033_, _12561_, _06989_);
  or _20868_ (_12562_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  nand _20869_ (_12563_, _07493_, _10739_);
  and _20870_ (_12564_, _12563_, _06989_);
  and _20871_ (_10036_, _12564_, _12562_);
  and _20872_ (_12566_, _12344_, _08713_);
  and _20873_ (_12567_, _08939_, _08731_);
  not _20874_ (_12568_, _12567_);
  or _20875_ (_12569_, _12568_, _09648_);
  and _20876_ (_12570_, _09897_, _08797_);
  not _20877_ (_12571_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _20878_ (_12572_, _09902_, _08932_);
  nor _20879_ (_12573_, _12572_, _12571_);
  and _20880_ (_12574_, _12572_, _09636_);
  or _20881_ (_12575_, _12574_, _12573_);
  or _20882_ (_12576_, _12575_, _12570_);
  not _20883_ (_12577_, _12570_);
  or _20884_ (_12578_, _12577_, word_in[8]);
  and _20885_ (_12579_, _12578_, _12576_);
  or _20886_ (_12580_, _12579_, _12567_);
  and _20887_ (_12581_, _12580_, _12569_);
  or _20888_ (_12582_, _12581_, _12566_);
  not _20889_ (_12583_, _12566_);
  or _20890_ (_12584_, _12583_, word_in[24]);
  and _20891_ (_10042_, _12584_, _12582_);
  or _20892_ (_12585_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  nand _20893_ (_12586_, _07493_, _10723_);
  and _20894_ (_12587_, _12586_, _06989_);
  and _20895_ (_10045_, _12587_, _12585_);
  or _20896_ (_12588_, _12568_, _09801_);
  not _20897_ (_12589_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor _20898_ (_12590_, _12572_, _12589_);
  and _20899_ (_12591_, _12572_, _09660_);
  or _20900_ (_12592_, _12591_, _12590_);
  or _20901_ (_12593_, _12592_, _12570_);
  or _20902_ (_12594_, _12577_, word_in[9]);
  and _20903_ (_12595_, _12594_, _12593_);
  or _20904_ (_12596_, _12595_, _12567_);
  and _20905_ (_12597_, _12596_, _12588_);
  or _20906_ (_12598_, _12597_, _12566_);
  or _20907_ (_12599_, _12583_, word_in[25]);
  and _20908_ (_10047_, _12599_, _12598_);
  or _20909_ (_12600_, _12568_, _09816_);
  not _20910_ (_12601_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor _20911_ (_12602_, _12572_, _12601_);
  and _20912_ (_12603_, _12572_, _09674_);
  or _20913_ (_12604_, _12603_, _12602_);
  or _20914_ (_12605_, _12604_, _12570_);
  or _20915_ (_12606_, _12577_, word_in[10]);
  and _20916_ (_12607_, _12606_, _12605_);
  or _20917_ (_12608_, _12607_, _12567_);
  and _20918_ (_12609_, _12608_, _12600_);
  or _20919_ (_12610_, _12609_, _12566_);
  or _20920_ (_12611_, _12583_, word_in[26]);
  and _20921_ (_10049_, _12611_, _12610_);
  or _20922_ (_12612_, _12568_, _09829_);
  not _20923_ (_12613_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor _20924_ (_12614_, _12572_, _12613_);
  and _20925_ (_12615_, _12572_, _09690_);
  or _20926_ (_12616_, _12615_, _12614_);
  or _20927_ (_12617_, _12616_, _12570_);
  or _20928_ (_12618_, _12577_, word_in[11]);
  and _20929_ (_12619_, _12618_, _12617_);
  or _20930_ (_12620_, _12619_, _12567_);
  and _20931_ (_12621_, _12620_, _12612_);
  and _20932_ (_12622_, _12621_, _12583_);
  and _20933_ (_12623_, _12566_, word_in[27]);
  or _20934_ (_10051_, _12623_, _12622_);
  or _20935_ (_12624_, _12568_, _09842_);
  not _20936_ (_12625_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor _20937_ (_12626_, _12572_, _12625_);
  and _20938_ (_12627_, _12572_, _09707_);
  or _20939_ (_12628_, _12627_, _12626_);
  or _20940_ (_12629_, _12628_, _12570_);
  or _20941_ (_12630_, _12577_, word_in[12]);
  and _20942_ (_12631_, _12630_, _12629_);
  or _20943_ (_12632_, _12631_, _12567_);
  and _20944_ (_12633_, _12632_, _12624_);
  or _20945_ (_12634_, _12633_, _12566_);
  or _20946_ (_12635_, _12583_, word_in[28]);
  and _20947_ (_10053_, _12635_, _12634_);
  or _20948_ (_12636_, _12568_, _09855_);
  not _20949_ (_12637_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor _20950_ (_12638_, _12572_, _12637_);
  and _20951_ (_12639_, _12572_, _09722_);
  or _20952_ (_12640_, _12639_, _12638_);
  or _20953_ (_12641_, _12640_, _12570_);
  or _20954_ (_12642_, _12577_, word_in[13]);
  and _20955_ (_12643_, _12642_, _12641_);
  or _20956_ (_12644_, _12643_, _12567_);
  and _20957_ (_12645_, _12644_, _12636_);
  and _20958_ (_12646_, _12645_, _12583_);
  and _20959_ (_12647_, _12566_, word_in[29]);
  or _20960_ (_10055_, _12647_, _12646_);
  nor _20961_ (_10056_, _11769_, rst);
  or _20962_ (_12648_, _12568_, _09871_);
  not _20963_ (_12649_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor _20964_ (_12650_, _12572_, _12649_);
  and _20965_ (_12651_, _12572_, _09735_);
  or _20966_ (_12652_, _12651_, _12650_);
  or _20967_ (_12653_, _12652_, _12570_);
  or _20968_ (_12654_, _12577_, word_in[14]);
  and _20969_ (_12656_, _12654_, _12653_);
  or _20970_ (_12657_, _12656_, _12567_);
  and _20971_ (_12658_, _12657_, _12648_);
  or _20972_ (_12659_, _12658_, _12566_);
  or _20973_ (_12660_, _12583_, word_in[30]);
  and _20974_ (_10058_, _12660_, _12659_);
  nor _20975_ (_12661_, _12572_, _08798_);
  and _20976_ (_12662_, _12572_, _08953_);
  or _20977_ (_12663_, _12662_, _12661_);
  and _20978_ (_12664_, _12663_, _12577_);
  and _20979_ (_12665_, _12570_, word_in[15]);
  or _20980_ (_12666_, _12665_, _12664_);
  or _20981_ (_12667_, _12666_, _12567_);
  or _20982_ (_12668_, _12568_, _08942_);
  and _20983_ (_12669_, _12668_, _12667_);
  and _20984_ (_12670_, _12669_, _12583_);
  and _20985_ (_12671_, _12566_, word_in[31]);
  or _20986_ (_10062_, _12671_, _12670_);
  and _20987_ (_12673_, _11045_, _08586_);
  nor _20988_ (_12674_, _12673_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _20989_ (_12675_, _12674_, _11276_);
  nor _20990_ (_12676_, _12675_, _11964_);
  and _20991_ (_12677_, _11986_, _08268_);
  or _20992_ (_12678_, _12136_, _12018_);
  not _20993_ (_12679_, _12137_);
  and _20994_ (_12680_, _12171_, _12679_);
  and _20995_ (_12681_, _12680_, _12678_);
  and _20996_ (_12682_, _12176_, _11671_);
  and _20997_ (_12683_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor _20998_ (_12684_, _12013_, _11988_);
  or _20999_ (_12685_, _12684_, _12683_);
  or _21000_ (_12686_, _12685_, _12682_);
  or _21001_ (_12687_, _12686_, _12681_);
  or _21002_ (_12688_, _12687_, _12677_);
  and _21003_ (_12689_, _12688_, _11964_);
  or _21004_ (_12690_, _12689_, _12676_);
  and _21005_ (_10074_, _12690_, _06989_);
  not _21006_ (_12691_, _11964_);
  and _21007_ (_12692_, _12691_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _21008_ (_12694_, _11986_, _08123_);
  or _21009_ (_12695_, _12117_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not _21010_ (_12696_, _12118_);
  and _21011_ (_12697_, _12171_, _12696_);
  and _21012_ (_12698_, _12697_, _12695_);
  and _21013_ (_12699_, _12114_, _11974_);
  and _21014_ (_12700_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and _21015_ (_12701_, _12176_, _11786_);
  or _21016_ (_12702_, _12701_, _12700_);
  or _21017_ (_12703_, _12702_, _12699_);
  or _21018_ (_12704_, _12703_, _12698_);
  or _21019_ (_12705_, _12704_, _12694_);
  and _21020_ (_12706_, _12705_, _11964_);
  or _21021_ (_12707_, _12706_, _12692_);
  and _21022_ (_10079_, _12707_, _06989_);
  and _21023_ (_12708_, _11275_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and _21024_ (_12709_, _12708_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _21025_ (_12710_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _21026_ (_12711_, _12710_, _12709_);
  and _21027_ (_12712_, _12711_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _21028_ (_12713_, _12712_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _21029_ (_12714_, _12713_, _11273_);
  nor _21030_ (_12715_, _12714_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _21031_ (_12716_, _12714_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor _21032_ (_12717_, _12716_, _12715_);
  or _21033_ (_12718_, _12717_, _11964_);
  and _21034_ (_12719_, _12718_, _06989_);
  nand _21035_ (_12720_, _11976_, _11981_);
  nor _21036_ (_12721_, _12720_, _11969_);
  nor _21037_ (_12722_, _12721_, _11983_);
  and _21038_ (_12723_, _11992_, _08479_);
  and _21039_ (_12724_, _07490_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and _21040_ (_12725_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and _21041_ (_12726_, _07343_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and _21042_ (_12727_, _07351_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor _21043_ (_12728_, _12727_, _12726_);
  and _21044_ (_12729_, _07341_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _21045_ (_12730_, _07338_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _21046_ (_12731_, _12730_, _12729_);
  and _21047_ (_12732_, _07333_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and _21048_ (_12733_, _07347_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _21049_ (_12734_, _12733_, _12732_);
  and _21050_ (_12735_, _12734_, _12731_);
  and _21051_ (_12736_, _12735_, _12728_);
  nor _21052_ (_12737_, _12736_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor _21053_ (_12738_, _12737_, _12725_);
  nor _21054_ (_12739_, _12738_, _07490_);
  nor _21055_ (_12740_, _12739_, _12724_);
  and _21056_ (_12741_, _12740_, _11994_);
  nor _21057_ (_12742_, _12741_, _12723_);
  nor _21058_ (_12743_, _12742_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _21059_ (_12744_, _12742_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nand _21060_ (_12745_, _12163_, _12159_);
  nor _21061_ (_12746_, _12745_, _12744_);
  nor _21062_ (_12747_, _12746_, _12743_);
  or _21063_ (_12748_, _12747_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _21064_ (_12749_, _12748_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or _21065_ (_12750_, _12749_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or _21066_ (_12751_, _12750_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand _21067_ (_12752_, _12751_, _12742_);
  not _21068_ (_12753_, _12742_);
  and _21069_ (_12754_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _21070_ (_12755_, _12754_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _21071_ (_12756_, _12755_, _12747_);
  nand _21072_ (_12757_, _12756_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand _21073_ (_12758_, _12757_, _12753_);
  and _21074_ (_12759_, _12758_, _12752_);
  or _21075_ (_12760_, _12759_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand _21076_ (_12761_, _12759_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _21077_ (_12762_, _12761_, _12760_);
  and _21078_ (_12763_, _12762_, _12722_);
  and _21079_ (_12764_, _11863_, _11560_);
  and _21080_ (_12765_, _12764_, _06980_);
  nor _21081_ (_12766_, _11936_, _11325_);
  not _21082_ (_12767_, _12766_);
  or _21083_ (_12768_, _12767_, _11383_);
  nor _21084_ (_12769_, _12768_, _11932_);
  nor _21085_ (_12770_, _11342_, _11413_);
  nor _21086_ (_12771_, _12770_, _12769_);
  nor _21087_ (_12772_, _12771_, _11943_);
  and _21088_ (_12773_, _11370_, _11368_);
  and _21089_ (_12774_, _11957_, _12773_);
  or _21090_ (_12775_, _12774_, _12772_);
  or _21091_ (_12776_, _12775_, _12765_);
  and _21092_ (_12777_, _11948_, _11372_);
  and _21093_ (_12778_, _11371_, _11368_);
  and _21094_ (_12779_, _12778_, _11873_);
  or _21095_ (_12780_, _12779_, _12777_);
  or _21096_ (_12781_, _12780_, _12776_);
  not _21097_ (_12782_, _11969_);
  and _21098_ (_12783_, _11984_, _12782_);
  and _21099_ (_12784_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _21100_ (_12785_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _21101_ (_12786_, _12785_, _12784_);
  and _21102_ (_12787_, \oc8051_top_1.oc8051_memory_interface1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _21103_ (_12788_, _12787_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _21104_ (_12789_, _12788_, _12755_);
  and _21105_ (_12790_, _12789_, _12786_);
  and _21106_ (_12791_, _12790_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _21107_ (_12792_, _12791_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _21108_ (_12793_, _12791_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _21109_ (_12794_, _12793_, _12792_);
  and _21110_ (_12795_, _12794_, _12783_);
  and _21111_ (_12796_, _11413_, _08346_);
  not _21112_ (_12797_, _11968_);
  nor _21113_ (_12798_, _12797_, _08307_);
  and _21114_ (_12799_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _21115_ (_12800_, _11974_, _11718_);
  or _21116_ (_12801_, _12800_, _12799_);
  or _21117_ (_12802_, _12801_, _12798_);
  or _21118_ (_12803_, _12802_, _12796_);
  or _21119_ (_12804_, _12803_, _12795_);
  or _21120_ (_12805_, _12804_, _12781_);
  or _21121_ (_12806_, _12805_, _12763_);
  and _21122_ (_10092_, _12806_, _12719_);
  and _21123_ (_12807_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _21124_ (_12808_, _11053_, _11011_);
  nor _21125_ (_12809_, _12808_, _11054_);
  or _21126_ (_12811_, _12809_, _08477_);
  or _21127_ (_12812_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and _21128_ (_12813_, _12812_, _10964_);
  and _21129_ (_12814_, _12813_, _12811_);
  or _21130_ (_10098_, _12814_, _12807_);
  and _21131_ (_12815_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _21132_ (_12816_, _11043_, _11026_);
  nor _21133_ (_12817_, _12816_, _11044_);
  or _21134_ (_12818_, _12817_, _08477_);
  or _21135_ (_12819_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and _21136_ (_12820_, _12819_, _10964_);
  and _21137_ (_12821_, _12820_, _12818_);
  or _21138_ (_10101_, _12821_, _12815_);
  and _21139_ (_12822_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _06989_);
  nor _21140_ (_12823_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _21141_ (_12824_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  and _21142_ (_12825_, _12824_, _12823_);
  nor _21143_ (_12826_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  nor _21144_ (_12827_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _21145_ (_12828_, _12827_, _12826_);
  and _21146_ (_12829_, _12828_, _12825_);
  and _21147_ (_12830_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _06989_);
  and _21148_ (_12831_, _12830_, _12829_);
  or _21149_ (_10112_, _12831_, _12822_);
  nor _21150_ (_10114_, _11670_, rst);
  not _21151_ (_12833_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor _21152_ (_12834_, _08951_, _12833_);
  and _21153_ (_12835_, _08951_, word_in[0]);
  nor _21154_ (_12836_, _12835_, _12834_);
  nor _21155_ (_12837_, _12836_, _08946_);
  and _21156_ (_12838_, _08946_, word_in[8]);
  or _21157_ (_12839_, _12838_, _12837_);
  and _21158_ (_12840_, _12839_, _08941_);
  and _21159_ (_12841_, _09648_, _08940_);
  or _21160_ (_12842_, _12841_, _12840_);
  and _21161_ (_12843_, _12842_, _08964_);
  and _21162_ (_12844_, _08936_, word_in[24]);
  or _21163_ (_10126_, _12844_, _12843_);
  and _21164_ (_12845_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _08578_);
  and _21165_ (_12846_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _21166_ (_12847_, _12846_, _12845_);
  and _21167_ (_10129_, _12847_, _06989_);
  not _21168_ (_12848_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor _21169_ (_12849_, _08951_, _12848_);
  and _21170_ (_12850_, _08951_, word_in[1]);
  nor _21171_ (_12852_, _12850_, _12849_);
  nor _21172_ (_12853_, _12852_, _08946_);
  and _21173_ (_12854_, _08946_, word_in[9]);
  or _21174_ (_12855_, _12854_, _12853_);
  and _21175_ (_12856_, _12855_, _08941_);
  and _21176_ (_12857_, _09801_, _08940_);
  or _21177_ (_12858_, _12857_, _12856_);
  and _21178_ (_12859_, _12858_, _08964_);
  and _21179_ (_12860_, _08936_, word_in[25]);
  or _21180_ (_10131_, _12860_, _12859_);
  not _21181_ (_12861_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor _21182_ (_12862_, _08951_, _12861_);
  and _21183_ (_12864_, _08951_, word_in[2]);
  or _21184_ (_12865_, _12864_, _12862_);
  or _21185_ (_12866_, _12865_, _08946_);
  or _21186_ (_12867_, _08957_, word_in[10]);
  and _21187_ (_12868_, _12867_, _12866_);
  or _21188_ (_12869_, _12868_, _08940_);
  or _21189_ (_12870_, _09816_, _08941_);
  and _21190_ (_12871_, _12870_, _08964_);
  and _21191_ (_12872_, _12871_, _12869_);
  and _21192_ (_12873_, _09685_, _08936_);
  or _21193_ (_10133_, _12873_, _12872_);
  not _21194_ (_12874_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor _21195_ (_12875_, _08951_, _12874_);
  and _21196_ (_12876_, _08951_, word_in[3]);
  or _21197_ (_12877_, _12876_, _12875_);
  or _21198_ (_12878_, _12877_, _08946_);
  or _21199_ (_12879_, _08957_, word_in[11]);
  and _21200_ (_12880_, _12879_, _12878_);
  or _21201_ (_12881_, _12880_, _08940_);
  or _21202_ (_12882_, _09829_, _08941_);
  and _21203_ (_12883_, _12882_, _08964_);
  and _21204_ (_12884_, _12883_, _12881_);
  and _21205_ (_12885_, _09701_, _08936_);
  or _21206_ (_10135_, _12885_, _12884_);
  and _21207_ (_12886_, _09842_, _08940_);
  not _21208_ (_12887_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor _21209_ (_12888_, _08951_, _12887_);
  and _21210_ (_12889_, _08951_, word_in[4]);
  nor _21211_ (_12890_, _12889_, _12888_);
  nor _21212_ (_12891_, _12890_, _08946_);
  and _21213_ (_12892_, _08946_, word_in[12]);
  or _21214_ (_12893_, _12892_, _12891_);
  and _21215_ (_12894_, _12893_, _08941_);
  or _21216_ (_12895_, _12894_, _12886_);
  and _21217_ (_12896_, _12895_, _08964_);
  and _21218_ (_12897_, _08936_, word_in[28]);
  or _21219_ (_10137_, _12897_, _12896_);
  and _21220_ (_12898_, _09855_, _08940_);
  not _21221_ (_12899_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor _21222_ (_12900_, _08951_, _12899_);
  and _21223_ (_12901_, _08951_, word_in[5]);
  nor _21224_ (_12902_, _12901_, _12900_);
  nor _21225_ (_12903_, _12902_, _08946_);
  and _21226_ (_12904_, _08946_, word_in[13]);
  or _21227_ (_12905_, _12904_, _12903_);
  and _21228_ (_12906_, _12905_, _08941_);
  or _21229_ (_12907_, _12906_, _12898_);
  and _21230_ (_12908_, _12907_, _08964_);
  and _21231_ (_12909_, _08936_, word_in[29]);
  or _21232_ (_10139_, _12909_, _12908_);
  and _21233_ (_12910_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor _21234_ (_12911_, _07493_, _11085_);
  or _21235_ (_12912_, _12911_, _12910_);
  and _21236_ (_10142_, _12912_, _06989_);
  and _21237_ (_12913_, _08951_, word_in[6]);
  not _21238_ (_12914_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor _21239_ (_12915_, _08951_, _12914_);
  nor _21240_ (_12916_, _12915_, _12913_);
  nor _21241_ (_12917_, _12916_, _08946_);
  and _21242_ (_12918_, _08946_, word_in[14]);
  or _21243_ (_12919_, _12918_, _12917_);
  or _21244_ (_12920_, _12919_, _08940_);
  or _21245_ (_12921_, _09871_, _08941_);
  and _21246_ (_12922_, _12921_, _08964_);
  and _21247_ (_12923_, _12922_, _12920_);
  and _21248_ (_12924_, _08936_, word_in[30]);
  or _21249_ (_10144_, _12924_, _12923_);
  or _21250_ (_12925_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  or _21251_ (_12926_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and _21252_ (_12927_, _12926_, _06989_);
  and _21253_ (_10400_, _12927_, _12925_);
  and _21254_ (_12928_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and _21255_ (_12929_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or _21256_ (_12930_, _12929_, _12928_);
  and _21257_ (_10446_, _12930_, _06989_);
  or _21258_ (_12931_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  or _21259_ (_12932_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  and _21260_ (_12933_, _12932_, _06989_);
  and _21261_ (_10449_, _12933_, _12931_);
  or _21262_ (_12934_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or _21263_ (_12935_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and _21264_ (_12936_, _12935_, _06989_);
  and _21265_ (_10452_, _12936_, _12934_);
  and _21266_ (_12937_, _08996_, _06981_);
  not _21267_ (_12938_, _12937_);
  nor _21268_ (_12939_, _12938_, _11529_);
  not _21269_ (_12940_, _08996_);
  and _21270_ (_12942_, _09606_, _12940_);
  nor _21271_ (_12943_, _12942_, _06982_);
  or _21272_ (_12944_, _09606_, _06982_);
  nand _21273_ (_12945_, _12944_, _12943_);
  and _21274_ (_12946_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  or _21275_ (_12947_, _12946_, _12939_);
  and _21276_ (_10877_, _12947_, _06989_);
  and _21277_ (_12948_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not _21278_ (_12949_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _21279_ (_12950_, _08139_, _12949_);
  or _21280_ (_12951_, _12950_, _12948_);
  and _21281_ (_10989_, _12951_, _06989_);
  and _21282_ (_12952_, _07134_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _21283_ (_12953_, _11529_, _09489_);
  or _21284_ (_12954_, _12953_, _12952_);
  nand _21285_ (_12955_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nor _21286_ (_12956_, _12955_, _07131_);
  or _21287_ (_12957_, _12956_, _12954_);
  and _21288_ (_11005_, _12957_, _06989_);
  not _21289_ (_12958_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor _21290_ (_12959_, _07123_, _12958_);
  and _21291_ (_12960_, _09599_, _07123_);
  or _21292_ (_12961_, _12960_, _06982_);
  or _21293_ (_12962_, _12961_, _12959_);
  or _21294_ (_12963_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and _21295_ (_12964_, _12963_, _06989_);
  and _21296_ (_11031_, _12964_, _12962_);
  and _21297_ (_12966_, _08708_, word_in[0]);
  nand _21298_ (_12967_, _08580_, _10685_);
  or _21299_ (_12968_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and _21300_ (_12969_, _12968_, _12967_);
  and _21301_ (_12970_, _12969_, _08623_);
  nand _21302_ (_12971_, _08580_, _11230_);
  or _21303_ (_12972_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _21304_ (_12973_, _12972_, _12971_);
  and _21305_ (_12974_, _12973_, _08606_);
  nand _21306_ (_12975_, _08580_, _12448_);
  or _21307_ (_12977_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and _21308_ (_12978_, _12977_, _12975_);
  and _21309_ (_12979_, _12978_, _08592_);
  or _21310_ (_12980_, _12979_, _12974_);
  or _21311_ (_12981_, _12980_, _12970_);
  nand _21312_ (_12982_, _08580_, _12833_);
  or _21313_ (_12983_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _21314_ (_12984_, _12983_, _12982_);
  and _21315_ (_12985_, _12984_, _08613_);
  or _21316_ (_12986_, _12985_, _08632_);
  or _21317_ (_12987_, _12986_, _12981_);
  nand _21318_ (_12988_, _08580_, _09771_);
  or _21319_ (_12989_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and _21320_ (_12990_, _12989_, _12988_);
  and _21321_ (_12991_, _12990_, _08623_);
  nand _21322_ (_12992_, _08580_, _10016_);
  or _21323_ (_12993_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _21324_ (_12994_, _12993_, _12992_);
  and _21325_ (_12995_, _12994_, _08606_);
  nand _21326_ (_12996_, _08580_, _10263_);
  or _21327_ (_12997_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and _21328_ (_12998_, _12997_, _12996_);
  and _21329_ (_12999_, _12998_, _08592_);
  or _21330_ (_13000_, _12999_, _12995_);
  or _21331_ (_13001_, _13000_, _12991_);
  nand _21332_ (_13002_, _08580_, _10474_);
  or _21333_ (_13003_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _21334_ (_13004_, _13003_, _13002_);
  and _21335_ (_13005_, _13004_, _08613_);
  or _21336_ (_13006_, _13005_, _08599_);
  or _21337_ (_13007_, _13006_, _13001_);
  and _21338_ (_13008_, _13007_, _12987_);
  and _21339_ (_13009_, _13008_, _08656_);
  or _21340_ (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _13009_, _12966_);
  and _21341_ (_13010_, _08708_, word_in[1]);
  nand _21342_ (_13011_, _08580_, _11247_);
  or _21343_ (_13012_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _21344_ (_13013_, _13012_, _13011_);
  and _21345_ (_13014_, _13013_, _08606_);
  nand _21346_ (_13015_, _08580_, _12463_);
  or _21347_ (_13016_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and _21348_ (_13017_, _13016_, _13015_);
  and _21349_ (_13018_, _13017_, _08592_);
  nand _21350_ (_13019_, _08580_, _10699_);
  or _21351_ (_13020_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and _21352_ (_13021_, _13020_, _13019_);
  and _21353_ (_13022_, _13021_, _08623_);
  or _21354_ (_13023_, _13022_, _13018_);
  or _21355_ (_13024_, _13023_, _13014_);
  nand _21356_ (_13025_, _08580_, _12848_);
  or _21357_ (_13026_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _21358_ (_13027_, _13026_, _13025_);
  and _21359_ (_13028_, _13027_, _08613_);
  or _21360_ (_13029_, _13028_, _08632_);
  or _21361_ (_13030_, _13029_, _13024_);
  nand _21362_ (_13031_, _08580_, _10037_);
  or _21363_ (_13032_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _21364_ (_13033_, _13032_, _13031_);
  and _21365_ (_13034_, _13033_, _08606_);
  nand _21366_ (_13035_, _08580_, _09792_);
  or _21367_ (_13036_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and _21368_ (_13037_, _13036_, _13035_);
  and _21369_ (_13038_, _13037_, _08623_);
  nand _21370_ (_13039_, _08580_, _10276_);
  or _21371_ (_13040_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and _21372_ (_13041_, _13040_, _13039_);
  and _21373_ (_13042_, _13041_, _08592_);
  or _21374_ (_13043_, _13042_, _13038_);
  or _21375_ (_13044_, _13043_, _13034_);
  nand _21376_ (_13045_, _08580_, _10489_);
  or _21377_ (_13046_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _21378_ (_13047_, _13046_, _13045_);
  and _21379_ (_13048_, _13047_, _08613_);
  or _21380_ (_13049_, _13048_, _08599_);
  or _21381_ (_13050_, _13049_, _13044_);
  and _21382_ (_13051_, _13050_, _13030_);
  and _21383_ (_13052_, _13051_, _08656_);
  or _21384_ (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _13052_, _13010_);
  and _21385_ (_13053_, _08708_, word_in[2]);
  nand _21386_ (_13054_, _08580_, _10710_);
  or _21387_ (_13055_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and _21388_ (_13056_, _13055_, _13054_);
  and _21389_ (_13057_, _13056_, _08623_);
  nand _21390_ (_13058_, _08580_, _11260_);
  or _21391_ (_13059_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _21392_ (_13060_, _13059_, _13058_);
  and _21393_ (_13061_, _13060_, _08606_);
  nand _21394_ (_13062_, _08580_, _12474_);
  or _21395_ (_13063_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and _21396_ (_13064_, _13063_, _13062_);
  and _21397_ (_13065_, _13064_, _08592_);
  or _21398_ (_13066_, _13065_, _13061_);
  or _21399_ (_13067_, _13066_, _13057_);
  nand _21400_ (_13068_, _08580_, _12861_);
  or _21401_ (_13069_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _21402_ (_13070_, _13069_, _13068_);
  and _21403_ (_13071_, _13070_, _08613_);
  or _21404_ (_13072_, _13071_, _08632_);
  or _21405_ (_13073_, _13072_, _13067_);
  nand _21406_ (_13074_, _08580_, _09807_);
  or _21407_ (_13075_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and _21408_ (_13076_, _13075_, _13074_);
  and _21409_ (_13077_, _13076_, _08623_);
  nand _21410_ (_13078_, _08580_, _10057_);
  or _21411_ (_13079_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _21412_ (_13080_, _13079_, _13078_);
  and _21413_ (_13081_, _13080_, _08606_);
  nand _21414_ (_13082_, _08580_, _10290_);
  or _21415_ (_13083_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and _21416_ (_13084_, _13083_, _13082_);
  and _21417_ (_13085_, _13084_, _08592_);
  or _21418_ (_13086_, _13085_, _13081_);
  or _21419_ (_13087_, _13086_, _13077_);
  nand _21420_ (_13088_, _08580_, _10501_);
  or _21421_ (_13089_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _21422_ (_13090_, _13089_, _13088_);
  and _21423_ (_13091_, _13090_, _08613_);
  or _21424_ (_13092_, _13091_, _08599_);
  or _21425_ (_13094_, _13092_, _13087_);
  and _21426_ (_13095_, _13094_, _13073_);
  and _21427_ (_13096_, _13095_, _08656_);
  or _21428_ (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _13096_, _13053_);
  and _21429_ (_13097_, _08708_, word_in[3]);
  nand _21430_ (_13098_, _08580_, _10727_);
  or _21431_ (_13099_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and _21432_ (_13100_, _13099_, _13098_);
  and _21433_ (_13101_, _13100_, _08623_);
  nand _21434_ (_13102_, _08580_, _12185_);
  or _21435_ (_13104_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _21436_ (_13105_, _13104_, _13102_);
  and _21437_ (_13106_, _13105_, _08606_);
  nand _21438_ (_13107_, _08580_, _12488_);
  or _21439_ (_13108_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and _21440_ (_13109_, _13108_, _13107_);
  and _21441_ (_13110_, _13109_, _08592_);
  or _21442_ (_13111_, _13110_, _13106_);
  or _21443_ (_13112_, _13111_, _13101_);
  nand _21444_ (_13113_, _08580_, _12874_);
  or _21445_ (_13115_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _21446_ (_13116_, _13115_, _13113_);
  and _21447_ (_13117_, _13116_, _08613_);
  or _21448_ (_13119_, _13117_, _08632_);
  or _21449_ (_13120_, _13119_, _13112_);
  nand _21450_ (_13121_, _08580_, _09821_);
  or _21451_ (_13122_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and _21452_ (_13123_, _13122_, _13121_);
  and _21453_ (_13124_, _13123_, _08623_);
  nand _21454_ (_13125_, _08580_, _10072_);
  or _21455_ (_13126_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _21456_ (_13127_, _13126_, _13125_);
  and _21457_ (_13128_, _13127_, _08606_);
  nand _21458_ (_13129_, _08580_, _10301_);
  or _21459_ (_13130_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and _21460_ (_13131_, _13130_, _13129_);
  and _21461_ (_13132_, _13131_, _08592_);
  or _21462_ (_13133_, _13132_, _13128_);
  or _21463_ (_13134_, _13133_, _13124_);
  nand _21464_ (_13135_, _08580_, _10512_);
  or _21465_ (_13136_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _21466_ (_13138_, _13136_, _13135_);
  and _21467_ (_13139_, _13138_, _08613_);
  or _21468_ (_13140_, _13139_, _08599_);
  or _21469_ (_13141_, _13140_, _13134_);
  and _21470_ (_13142_, _13141_, _13120_);
  and _21471_ (_13143_, _13142_, _08656_);
  or _21472_ (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _13143_, _13097_);
  and _21473_ (_13144_, _08708_, word_in[4]);
  nand _21474_ (_13145_, _08580_, _10743_);
  or _21475_ (_13147_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and _21476_ (_13148_, _13147_, _13145_);
  and _21477_ (_13149_, _13148_, _08623_);
  nand _21478_ (_13150_, _08580_, _12196_);
  or _21479_ (_13151_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _21480_ (_13152_, _13151_, _13150_);
  and _21481_ (_13153_, _13152_, _08606_);
  nand _21482_ (_13155_, _08580_, _12501_);
  or _21483_ (_13156_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and _21484_ (_13158_, _13156_, _13155_);
  and _21485_ (_13159_, _13158_, _08592_);
  or _21486_ (_13160_, _13159_, _13153_);
  or _21487_ (_13161_, _13160_, _13149_);
  nand _21488_ (_13162_, _08580_, _12887_);
  or _21489_ (_13163_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _21490_ (_13164_, _13163_, _13162_);
  and _21491_ (_13165_, _13164_, _08613_);
  or _21492_ (_13166_, _13165_, _08632_);
  or _21493_ (_13167_, _13166_, _13161_);
  nand _21494_ (_13168_, _08580_, _09834_);
  or _21495_ (_13169_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and _21496_ (_13170_, _13169_, _13168_);
  and _21497_ (_13171_, _13170_, _08623_);
  nand _21498_ (_13172_, _08580_, _10086_);
  or _21499_ (_13173_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _21500_ (_13174_, _13173_, _13172_);
  and _21501_ (_13175_, _13174_, _08606_);
  nand _21502_ (_13176_, _08580_, _10315_);
  or _21503_ (_13177_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and _21504_ (_13178_, _13177_, _13176_);
  and _21505_ (_13179_, _13178_, _08592_);
  or _21506_ (_13180_, _13179_, _13175_);
  or _21507_ (_13181_, _13180_, _13171_);
  nand _21508_ (_13182_, _08580_, _10525_);
  or _21509_ (_13183_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _21510_ (_13184_, _13183_, _13182_);
  and _21511_ (_13185_, _13184_, _08613_);
  or _21512_ (_13186_, _13185_, _08599_);
  or _21513_ (_13187_, _13186_, _13181_);
  and _21514_ (_13188_, _13187_, _13167_);
  and _21515_ (_13189_, _13188_, _08656_);
  or _21516_ (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _13189_, _13144_);
  and _21517_ (_13190_, _08708_, word_in[5]);
  nand _21518_ (_13191_, _08580_, _10759_);
  or _21519_ (_13192_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and _21520_ (_13193_, _13192_, _13191_);
  and _21521_ (_13194_, _13193_, _08623_);
  nand _21522_ (_13195_, _08580_, _12209_);
  or _21523_ (_13196_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _21524_ (_13197_, _13196_, _13195_);
  and _21525_ (_13198_, _13197_, _08606_);
  nand _21526_ (_13199_, _08580_, _12513_);
  or _21527_ (_13200_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and _21528_ (_13201_, _13200_, _13199_);
  and _21529_ (_13202_, _13201_, _08592_);
  or _21530_ (_13203_, _13202_, _13198_);
  or _21531_ (_13204_, _13203_, _13194_);
  nand _21532_ (_13205_, _08580_, _12899_);
  or _21533_ (_13206_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _21534_ (_13208_, _13206_, _13205_);
  and _21535_ (_13209_, _13208_, _08613_);
  or _21536_ (_13210_, _13209_, _08632_);
  or _21537_ (_13211_, _13210_, _13204_);
  nand _21538_ (_13212_, _08580_, _09847_);
  or _21539_ (_13213_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and _21540_ (_13214_, _13213_, _13212_);
  and _21541_ (_13215_, _13214_, _08623_);
  nand _21542_ (_13216_, _08580_, _10100_);
  or _21543_ (_13217_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and _21544_ (_13218_, _13217_, _13216_);
  and _21545_ (_13219_, _13218_, _08606_);
  nand _21546_ (_13220_, _08580_, _10325_);
  or _21547_ (_13221_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and _21548_ (_13222_, _13221_, _13220_);
  and _21549_ (_13223_, _13222_, _08592_);
  or _21550_ (_13224_, _13223_, _13219_);
  or _21551_ (_13226_, _13224_, _13215_);
  nand _21552_ (_13227_, _08580_, _10537_);
  or _21553_ (_13228_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _21554_ (_13229_, _13228_, _13227_);
  and _21555_ (_13230_, _13229_, _08613_);
  or _21556_ (_13231_, _13230_, _08599_);
  or _21557_ (_13232_, _13231_, _13226_);
  and _21558_ (_13233_, _13232_, _13211_);
  and _21559_ (_13234_, _13233_, _08656_);
  or _21560_ (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _13234_, _13190_);
  and _21561_ (_13235_, _08708_, word_in[6]);
  nand _21562_ (_13236_, _08580_, _10771_);
  or _21563_ (_13237_, _08580_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and _21564_ (_13238_, _13237_, _13236_);
  and _21565_ (_13239_, _13238_, _08623_);
  nand _21566_ (_13240_, _08580_, _12225_);
  or _21567_ (_13241_, _08580_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _21568_ (_13242_, _13241_, _13240_);
  and _21569_ (_13243_, _13242_, _08606_);
  nand _21570_ (_13244_, _08580_, _12524_);
  or _21571_ (_13245_, _08580_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and _21572_ (_13246_, _13245_, _13244_);
  and _21573_ (_13247_, _13246_, _08592_);
  or _21574_ (_13248_, _13247_, _13243_);
  or _21575_ (_13249_, _13248_, _13239_);
  nand _21576_ (_13250_, _08580_, _12914_);
  or _21577_ (_13251_, _08580_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _21578_ (_13252_, _13251_, _13250_);
  and _21579_ (_13253_, _13252_, _08613_);
  or _21580_ (_13254_, _13253_, _08632_);
  or _21581_ (_13255_, _13254_, _13249_);
  nand _21582_ (_13256_, _08580_, _09860_);
  or _21583_ (_13257_, _08580_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and _21584_ (_13258_, _13257_, _13256_);
  and _21585_ (_13259_, _13258_, _08623_);
  nand _21586_ (_13260_, _08580_, _10113_);
  or _21587_ (_13261_, _08580_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and _21588_ (_13262_, _13261_, _13260_);
  and _21589_ (_13263_, _13262_, _08606_);
  nand _21590_ (_13264_, _08580_, _10338_);
  or _21591_ (_13265_, _08580_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and _21592_ (_13266_, _13265_, _13264_);
  and _21593_ (_13267_, _13266_, _08592_);
  or _21594_ (_13268_, _13267_, _13263_);
  or _21595_ (_13269_, _13268_, _13259_);
  nand _21596_ (_13270_, _08580_, _10548_);
  or _21597_ (_13271_, _08580_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _21598_ (_13273_, _13271_, _13270_);
  and _21599_ (_13274_, _13273_, _08613_);
  or _21600_ (_13275_, _13274_, _08599_);
  or _21601_ (_13276_, _13275_, _13269_);
  and _21602_ (_13277_, _13276_, _13255_);
  and _21603_ (_13278_, _13277_, _08656_);
  or _21604_ (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _13278_, _13235_);
  and _21605_ (_13279_, _08757_, word_in[8]);
  nand _21606_ (_13280_, _08580_, _09900_);
  or _21607_ (_13281_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _21608_ (_13282_, _13281_, _13280_);
  and _21609_ (_13283_, _13282_, _08759_);
  nand _21610_ (_13284_, _08580_, _09625_);
  or _21611_ (_13285_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and _21612_ (_13286_, _13285_, _13284_);
  and _21613_ (_13287_, _13286_, _08758_);
  or _21614_ (_13288_, _13287_, _13283_);
  and _21615_ (_13289_, _13288_, _08724_);
  nand _21616_ (_13290_, _08580_, _11094_);
  or _21617_ (_13291_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _21618_ (_13292_, _13291_, _13290_);
  and _21619_ (_13293_, _13292_, _08759_);
  nand _21620_ (_13294_, _08580_, _10573_);
  or _21621_ (_13295_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and _21622_ (_13296_, _13295_, _13294_);
  and _21623_ (_13297_, _13296_, _08758_);
  or _21624_ (_13298_, _13297_, _13293_);
  and _21625_ (_13299_, _13298_, _08726_);
  nand _21626_ (_13300_, _08580_, _10368_);
  or _21627_ (_13301_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _21628_ (_13302_, _13301_, _13300_);
  and _21629_ (_13303_, _13302_, _08759_);
  nand _21630_ (_13304_, _08580_, _10158_);
  or _21631_ (_13305_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and _21632_ (_13306_, _13305_, _13304_);
  and _21633_ (_13307_, _13306_, _08758_);
  or _21634_ (_13308_, _13307_, _13303_);
  and _21635_ (_13309_, _13308_, _08784_);
  nand _21636_ (_13310_, _08580_, _12571_);
  or _21637_ (_13311_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _21638_ (_13312_, _13311_, _13310_);
  and _21639_ (_13313_, _13312_, _08759_);
  nand _21640_ (_13314_, _08580_, _12333_);
  or _21641_ (_13315_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and _21642_ (_13316_, _13315_, _13314_);
  and _21643_ (_13317_, _13316_, _08758_);
  or _21644_ (_13318_, _13317_, _13313_);
  and _21645_ (_13319_, _13318_, _08797_);
  or _21646_ (_13320_, _13319_, _13309_);
  or _21647_ (_13321_, _13320_, _13299_);
  nor _21648_ (_13322_, _13321_, _13289_);
  nor _21649_ (_13323_, _13322_, _08757_);
  or _21650_ (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _13323_, _13279_);
  and _21651_ (_13324_, _08757_, word_in[9]);
  nand _21652_ (_13325_, _08580_, _09916_);
  or _21653_ (_13326_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _21654_ (_13327_, _13326_, _13325_);
  and _21655_ (_13328_, _13327_, _08759_);
  nand _21656_ (_13329_, _08580_, _09658_);
  or _21657_ (_13330_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and _21658_ (_13331_, _13330_, _13329_);
  and _21659_ (_13332_, _13331_, _08758_);
  or _21660_ (_13333_, _13332_, _13328_);
  and _21661_ (_13334_, _13333_, _08724_);
  nand _21662_ (_13335_, _08580_, _11108_);
  or _21663_ (_13336_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _21664_ (_13337_, _13336_, _13335_);
  and _21665_ (_13338_, _13337_, _08759_);
  nand _21666_ (_13339_, _08580_, _10591_);
  or _21667_ (_13340_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and _21668_ (_13341_, _13340_, _13339_);
  and _21669_ (_13342_, _13341_, _08758_);
  or _21670_ (_13344_, _13342_, _13338_);
  and _21671_ (_13345_, _13344_, _08726_);
  nand _21672_ (_13346_, _08580_, _10382_);
  or _21673_ (_13347_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _21674_ (_13348_, _13347_, _13346_);
  and _21675_ (_13349_, _13348_, _08759_);
  nand _21676_ (_13350_, _08580_, _10175_);
  or _21677_ (_13351_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and _21678_ (_13352_, _13351_, _13350_);
  and _21679_ (_13353_, _13352_, _08758_);
  or _21680_ (_13354_, _13353_, _13349_);
  and _21681_ (_13355_, _13354_, _08784_);
  nand _21682_ (_13356_, _08580_, _12589_);
  or _21683_ (_13357_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _21684_ (_13358_, _13357_, _13356_);
  and _21685_ (_13359_, _13358_, _08759_);
  nand _21686_ (_13360_, _08580_, _12352_);
  or _21687_ (_13361_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and _21688_ (_13362_, _13361_, _13360_);
  and _21689_ (_13363_, _13362_, _08758_);
  or _21690_ (_13364_, _13363_, _13359_);
  and _21691_ (_13366_, _13364_, _08797_);
  or _21692_ (_13367_, _13366_, _13355_);
  or _21693_ (_13368_, _13367_, _13345_);
  nor _21694_ (_13369_, _13368_, _13334_);
  nor _21695_ (_13370_, _13369_, _08757_);
  or _21696_ (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _13370_, _13324_);
  and _21697_ (_13371_, _08757_, word_in[10]);
  nand _21698_ (_13372_, _08580_, _09931_);
  or _21699_ (_13373_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _21700_ (_13374_, _13373_, _13372_);
  and _21701_ (_13375_, _13374_, _08759_);
  nand _21702_ (_13376_, _08580_, _09672_);
  or _21703_ (_13377_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  and _21704_ (_13378_, _13377_, _13376_);
  and _21705_ (_13379_, _13378_, _08758_);
  or _21706_ (_13380_, _13379_, _13375_);
  and _21707_ (_13381_, _13380_, _08724_);
  nand _21708_ (_13382_, _08580_, _11120_);
  or _21709_ (_13383_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _21710_ (_13384_, _13383_, _13382_);
  and _21711_ (_13385_, _13384_, _08759_);
  nand _21712_ (_13386_, _08580_, _10603_);
  or _21713_ (_13387_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and _21714_ (_13388_, _13387_, _13386_);
  and _21715_ (_13389_, _13388_, _08758_);
  or _21716_ (_13390_, _13389_, _13385_);
  and _21717_ (_13391_, _13390_, _08726_);
  nand _21718_ (_13392_, _08580_, _10395_);
  or _21719_ (_13393_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _21720_ (_13394_, _13393_, _13392_);
  and _21721_ (_13395_, _13394_, _08759_);
  nand _21722_ (_13396_, _08580_, _10187_);
  or _21723_ (_13397_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and _21724_ (_13398_, _13397_, _13396_);
  and _21725_ (_13399_, _13398_, _08758_);
  or _21726_ (_13400_, _13399_, _13395_);
  and _21727_ (_13401_, _13400_, _08784_);
  nand _21728_ (_13402_, _08580_, _12601_);
  or _21729_ (_13403_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _21730_ (_13404_, _13403_, _13402_);
  and _21731_ (_13405_, _13404_, _08759_);
  nand _21732_ (_13406_, _08580_, _12365_);
  or _21733_ (_13407_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and _21734_ (_13408_, _13407_, _13406_);
  and _21735_ (_13409_, _13408_, _08758_);
  or _21736_ (_13410_, _13409_, _13405_);
  and _21737_ (_13411_, _13410_, _08797_);
  or _21738_ (_13412_, _13411_, _13401_);
  or _21739_ (_13413_, _13412_, _13391_);
  nor _21740_ (_13414_, _13413_, _13381_);
  nor _21741_ (_13416_, _13414_, _08757_);
  or _21742_ (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _13416_, _13371_);
  and _21743_ (_13417_, _08757_, word_in[11]);
  nand _21744_ (_13418_, _08580_, _09944_);
  or _21745_ (_13419_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _21746_ (_13420_, _13419_, _13418_);
  and _21747_ (_13421_, _13420_, _08759_);
  nand _21748_ (_13422_, _08580_, _09688_);
  or _21749_ (_13424_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  and _21750_ (_13425_, _13424_, _13422_);
  and _21751_ (_13426_, _13425_, _08758_);
  or _21752_ (_13427_, _13426_, _13421_);
  and _21753_ (_13428_, _13427_, _08724_);
  nand _21754_ (_13429_, _08580_, _11132_);
  or _21755_ (_13430_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _21756_ (_13431_, _13430_, _13429_);
  and _21757_ (_13432_, _13431_, _08759_);
  nand _21758_ (_13433_, _08580_, _10615_);
  or _21759_ (_13434_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and _21760_ (_13435_, _13434_, _13433_);
  and _21761_ (_13436_, _13435_, _08758_);
  or _21762_ (_13437_, _13436_, _13432_);
  and _21763_ (_13438_, _13437_, _08726_);
  nand _21764_ (_13439_, _08580_, _10407_);
  or _21765_ (_13440_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _21766_ (_13441_, _13440_, _13439_);
  and _21767_ (_13442_, _13441_, _08759_);
  nand _21768_ (_13443_, _08580_, _10199_);
  or _21769_ (_13444_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and _21770_ (_13445_, _13444_, _13443_);
  and _21771_ (_13447_, _13445_, _08758_);
  or _21772_ (_13448_, _13447_, _13442_);
  and _21773_ (_13449_, _13448_, _08784_);
  nand _21774_ (_13450_, _08580_, _12613_);
  or _21775_ (_13451_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _21776_ (_13452_, _13451_, _13450_);
  and _21777_ (_13453_, _13452_, _08759_);
  nand _21778_ (_13454_, _08580_, _12378_);
  or _21779_ (_13455_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and _21780_ (_13456_, _13455_, _13454_);
  and _21781_ (_13457_, _13456_, _08758_);
  or _21782_ (_13458_, _13457_, _13453_);
  and _21783_ (_13459_, _13458_, _08797_);
  or _21784_ (_13460_, _13459_, _13449_);
  or _21785_ (_13461_, _13460_, _13438_);
  nor _21786_ (_13462_, _13461_, _13428_);
  nor _21787_ (_13464_, _13462_, _08757_);
  or _21788_ (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _13464_, _13417_);
  and _21789_ (_13465_, _08757_, word_in[12]);
  nand _21790_ (_13466_, _08580_, _09957_);
  or _21791_ (_13467_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and _21792_ (_13468_, _13467_, _13466_);
  and _21793_ (_13469_, _13468_, _08759_);
  nand _21794_ (_13470_, _08580_, _09705_);
  or _21795_ (_13471_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _21796_ (_13472_, _13471_, _13470_);
  and _21797_ (_13473_, _13472_, _08758_);
  or _21798_ (_13474_, _13473_, _13469_);
  and _21799_ (_13475_, _13474_, _08724_);
  nand _21800_ (_13476_, _08580_, _11144_);
  or _21801_ (_13477_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and _21802_ (_13478_, _13477_, _13476_);
  and _21803_ (_13479_, _13478_, _08759_);
  nand _21804_ (_13480_, _08580_, _10627_);
  or _21805_ (_13481_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _21806_ (_13482_, _13481_, _13480_);
  and _21807_ (_13483_, _13482_, _08758_);
  or _21808_ (_13484_, _13483_, _13479_);
  and _21809_ (_13485_, _13484_, _08726_);
  nand _21810_ (_13486_, _08580_, _10420_);
  or _21811_ (_13487_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _21812_ (_13488_, _13487_, _13486_);
  and _21813_ (_13489_, _13488_, _08759_);
  nand _21814_ (_13490_, _08580_, _10212_);
  or _21815_ (_13491_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and _21816_ (_13492_, _13491_, _13490_);
  and _21817_ (_13493_, _13492_, _08758_);
  or _21818_ (_13494_, _13493_, _13489_);
  and _21819_ (_13495_, _13494_, _08784_);
  nand _21820_ (_13496_, _08580_, _12625_);
  or _21821_ (_13497_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _21822_ (_13498_, _13497_, _13496_);
  and _21823_ (_13499_, _13498_, _08759_);
  nand _21824_ (_13500_, _08580_, _12390_);
  or _21825_ (_13501_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and _21826_ (_13502_, _13501_, _13500_);
  and _21827_ (_13503_, _13502_, _08758_);
  or _21828_ (_13504_, _13503_, _13499_);
  and _21829_ (_13505_, _13504_, _08797_);
  or _21830_ (_13506_, _13505_, _13495_);
  or _21831_ (_13507_, _13506_, _13485_);
  nor _21832_ (_13508_, _13507_, _13475_);
  nor _21833_ (_13509_, _13508_, _08757_);
  or _21834_ (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _13509_, _13465_);
  and _21835_ (_13510_, _08757_, word_in[13]);
  nand _21836_ (_13511_, _08580_, _09974_);
  or _21837_ (_13512_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _21838_ (_13513_, _13512_, _13511_);
  and _21839_ (_13514_, _13513_, _08759_);
  nand _21840_ (_13515_, _08580_, _09720_);
  or _21841_ (_13516_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _21842_ (_13517_, _13516_, _13515_);
  and _21843_ (_13518_, _13517_, _08758_);
  or _21844_ (_13519_, _13518_, _13514_);
  and _21845_ (_13520_, _13519_, _08724_);
  nand _21846_ (_13521_, _08580_, _11156_);
  or _21847_ (_13522_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _21848_ (_13523_, _13522_, _13521_);
  and _21849_ (_13524_, _13523_, _08759_);
  nand _21850_ (_13525_, _08580_, _10639_);
  or _21851_ (_13526_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and _21852_ (_13527_, _13526_, _13525_);
  and _21853_ (_13528_, _13527_, _08758_);
  or _21854_ (_13529_, _13528_, _13524_);
  and _21855_ (_13530_, _13529_, _08726_);
  nand _21856_ (_13531_, _08580_, _10431_);
  or _21857_ (_13532_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _21858_ (_13533_, _13532_, _13531_);
  and _21859_ (_13534_, _13533_, _08759_);
  nand _21860_ (_13535_, _08580_, _10223_);
  or _21861_ (_13536_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and _21862_ (_13537_, _13536_, _13535_);
  and _21863_ (_13538_, _13537_, _08758_);
  or _21864_ (_13539_, _13538_, _13534_);
  and _21865_ (_13540_, _13539_, _08784_);
  nand _21866_ (_13541_, _08580_, _12637_);
  or _21867_ (_13542_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _21868_ (_13543_, _13542_, _13541_);
  and _21869_ (_13544_, _13543_, _08759_);
  nand _21870_ (_13545_, _08580_, _12403_);
  or _21871_ (_13546_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and _21872_ (_13547_, _13546_, _13545_);
  and _21873_ (_13548_, _13547_, _08758_);
  or _21874_ (_13549_, _13548_, _13544_);
  and _21875_ (_13550_, _13549_, _08797_);
  or _21876_ (_13551_, _13550_, _13540_);
  or _21877_ (_13552_, _13551_, _13530_);
  nor _21878_ (_13553_, _13552_, _13520_);
  nor _21879_ (_13554_, _13553_, _08757_);
  or _21880_ (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _13554_, _13510_);
  and _21881_ (_13555_, _08757_, word_in[14]);
  nand _21882_ (_13556_, _08580_, _09988_);
  or _21883_ (_13557_, _08580_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _21884_ (_13558_, _13557_, _13556_);
  and _21885_ (_13559_, _13558_, _08759_);
  nand _21886_ (_13560_, _08580_, _09732_);
  or _21887_ (_13561_, _08580_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _21888_ (_13562_, _13561_, _13560_);
  and _21889_ (_13563_, _13562_, _08758_);
  or _21890_ (_13564_, _13563_, _13559_);
  and _21891_ (_13565_, _13564_, _08724_);
  nand _21892_ (_13566_, _08580_, _11168_);
  or _21893_ (_13567_, _08580_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _21894_ (_13568_, _13567_, _13566_);
  and _21895_ (_13569_, _13568_, _08759_);
  nand _21896_ (_13570_, _08580_, _10652_);
  or _21897_ (_13571_, _08580_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and _21898_ (_13572_, _13571_, _13570_);
  and _21899_ (_13574_, _13572_, _08758_);
  or _21900_ (_13575_, _13574_, _13569_);
  and _21901_ (_13576_, _13575_, _08726_);
  nand _21902_ (_13577_, _08580_, _10444_);
  or _21903_ (_13578_, _08580_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _21904_ (_13579_, _13578_, _13577_);
  and _21905_ (_13581_, _13579_, _08759_);
  nand _21906_ (_13582_, _08580_, _10235_);
  or _21907_ (_13583_, _08580_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and _21908_ (_13584_, _13583_, _13582_);
  and _21909_ (_13585_, _13584_, _08758_);
  or _21910_ (_13586_, _13585_, _13581_);
  and _21911_ (_13587_, _13586_, _08784_);
  nand _21912_ (_13588_, _08580_, _12649_);
  or _21913_ (_13589_, _08580_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _21914_ (_13590_, _13589_, _13588_);
  and _21915_ (_13591_, _13590_, _08759_);
  nand _21916_ (_13593_, _08580_, _12417_);
  or _21917_ (_13594_, _08580_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and _21918_ (_13595_, _13594_, _13593_);
  and _21919_ (_13596_, _13595_, _08758_);
  or _21920_ (_13598_, _13596_, _13591_);
  and _21921_ (_13599_, _13598_, _08797_);
  or _21922_ (_13600_, _13599_, _13587_);
  or _21923_ (_13601_, _13600_, _13576_);
  nor _21924_ (_13602_, _13601_, _13565_);
  nor _21925_ (_13603_, _13602_, _08757_);
  or _21926_ (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _13603_, _13555_);
  and _21927_ (_13604_, _08850_, word_in[16]);
  and _21928_ (_13605_, _12998_, _08606_);
  and _21929_ (_13606_, _12990_, _08613_);
  or _21930_ (_13607_, _13606_, _13605_);
  and _21931_ (_13608_, _13004_, _08592_);
  and _21932_ (_13609_, _12994_, _08623_);
  or _21933_ (_13610_, _13609_, _13608_);
  or _21934_ (_13611_, _13610_, _13607_);
  or _21935_ (_13612_, _13611_, _08821_);
  and _21936_ (_13613_, _12978_, _08606_);
  and _21937_ (_13614_, _12969_, _08613_);
  or _21938_ (_13615_, _13614_, _13613_);
  and _21939_ (_13616_, _12984_, _08592_);
  and _21940_ (_13617_, _12973_, _08623_);
  or _21941_ (_13618_, _13617_, _13616_);
  or _21942_ (_13619_, _13618_, _13615_);
  or _21943_ (_13620_, _13619_, _08860_);
  nand _21944_ (_13621_, _13620_, _13612_);
  nor _21945_ (_13622_, _13621_, _08850_);
  or _21946_ (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _13622_, _13604_);
  and _21947_ (_13623_, _08850_, word_in[17]);
  and _21948_ (_13624_, _13037_, _08613_);
  and _21949_ (_13625_, _13047_, _08592_);
  or _21950_ (_13626_, _13625_, _13624_);
  and _21951_ (_13627_, _13041_, _08606_);
  and _21952_ (_13628_, _13033_, _08623_);
  or _21953_ (_13629_, _13628_, _13627_);
  or _21954_ (_13630_, _13629_, _13626_);
  or _21955_ (_13631_, _13630_, _08821_);
  and _21956_ (_13632_, _13017_, _08606_);
  and _21957_ (_13633_, _13021_, _08613_);
  or _21958_ (_13634_, _13633_, _13632_);
  and _21959_ (_13635_, _13027_, _08592_);
  and _21960_ (_13636_, _13013_, _08623_);
  or _21961_ (_13637_, _13636_, _13635_);
  or _21962_ (_13638_, _13637_, _13634_);
  or _21963_ (_13639_, _13638_, _08860_);
  nand _21964_ (_13640_, _13639_, _13631_);
  nor _21965_ (_13641_, _13640_, _08850_);
  or _21966_ (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _13641_, _13623_);
  and _21967_ (_13642_, _08850_, word_in[18]);
  and _21968_ (_13643_, _13084_, _08606_);
  and _21969_ (_13644_, _13076_, _08613_);
  or _21970_ (_13645_, _13644_, _13643_);
  and _21971_ (_13646_, _13090_, _08592_);
  and _21972_ (_13647_, _13080_, _08623_);
  or _21973_ (_13648_, _13647_, _13646_);
  or _21974_ (_13650_, _13648_, _13645_);
  or _21975_ (_13652_, _13650_, _08821_);
  and _21976_ (_13653_, _13064_, _08606_);
  and _21977_ (_13654_, _13056_, _08613_);
  or _21978_ (_13655_, _13654_, _13653_);
  and _21979_ (_13656_, _13070_, _08592_);
  and _21980_ (_13657_, _13060_, _08623_);
  or _21981_ (_13658_, _13657_, _13656_);
  or _21982_ (_13659_, _13658_, _13655_);
  or _21983_ (_13660_, _13659_, _08860_);
  nand _21984_ (_13661_, _13660_, _13652_);
  nor _21985_ (_13662_, _13661_, _08850_);
  or _21986_ (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _13662_, _13642_);
  and _21987_ (_13663_, _08850_, word_in[19]);
  and _21988_ (_13664_, _13131_, _08606_);
  and _21989_ (_13665_, _13123_, _08613_);
  or _21990_ (_13666_, _13665_, _13664_);
  and _21991_ (_13667_, _13138_, _08592_);
  and _21992_ (_13668_, _13127_, _08623_);
  or _21993_ (_13669_, _13668_, _13667_);
  or _21994_ (_13670_, _13669_, _13666_);
  or _21995_ (_13671_, _13670_, _08821_);
  and _21996_ (_13672_, _13100_, _08613_);
  and _21997_ (_13673_, _13116_, _08592_);
  or _21998_ (_13674_, _13673_, _13672_);
  and _21999_ (_13675_, _13109_, _08606_);
  and _22000_ (_13676_, _13105_, _08623_);
  or _22001_ (_13677_, _13676_, _13675_);
  or _22002_ (_13678_, _13677_, _13674_);
  or _22003_ (_13679_, _13678_, _08860_);
  nand _22004_ (_13680_, _13679_, _13671_);
  nor _22005_ (_13681_, _13680_, _08850_);
  or _22006_ (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _13681_, _13663_);
  and _22007_ (_13682_, _08850_, word_in[20]);
  and _22008_ (_13683_, _13178_, _08606_);
  and _22009_ (_13684_, _13170_, _08613_);
  or _22010_ (_13685_, _13684_, _13683_);
  and _22011_ (_13686_, _13184_, _08592_);
  and _22012_ (_13687_, _13174_, _08623_);
  or _22013_ (_13688_, _13687_, _13686_);
  or _22014_ (_13689_, _13688_, _13685_);
  or _22015_ (_13690_, _13689_, _08821_);
  and _22016_ (_13691_, _13158_, _08606_);
  and _22017_ (_13692_, _13148_, _08613_);
  or _22018_ (_13693_, _13692_, _13691_);
  and _22019_ (_13694_, _13164_, _08592_);
  and _22020_ (_13695_, _13152_, _08623_);
  or _22021_ (_13696_, _13695_, _13694_);
  or _22022_ (_13697_, _13696_, _13693_);
  or _22023_ (_13698_, _13697_, _08860_);
  nand _22024_ (_13699_, _13698_, _13690_);
  nor _22025_ (_13700_, _13699_, _08850_);
  or _22026_ (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _13700_, _13682_);
  and _22027_ (_13701_, _08850_, word_in[21]);
  and _22028_ (_13702_, _13222_, _08606_);
  and _22029_ (_13703_, _13214_, _08613_);
  or _22030_ (_13704_, _13703_, _13702_);
  and _22031_ (_13705_, _13229_, _08592_);
  and _22032_ (_13706_, _13218_, _08623_);
  or _22033_ (_13708_, _13706_, _13705_);
  or _22034_ (_13709_, _13708_, _13704_);
  or _22035_ (_13711_, _13709_, _08821_);
  and _22036_ (_13712_, _13193_, _08613_);
  and _22037_ (_13713_, _13208_, _08592_);
  or _22038_ (_13714_, _13713_, _13712_);
  and _22039_ (_13715_, _13201_, _08606_);
  and _22040_ (_13716_, _13197_, _08623_);
  or _22041_ (_13717_, _13716_, _13715_);
  or _22042_ (_13718_, _13717_, _13714_);
  or _22043_ (_13719_, _13718_, _08860_);
  nand _22044_ (_13720_, _13719_, _13711_);
  nor _22045_ (_13721_, _13720_, _08850_);
  or _22046_ (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _13721_, _13701_);
  and _22047_ (_13722_, _08850_, word_in[22]);
  and _22048_ (_13723_, _13258_, _08613_);
  and _22049_ (_13724_, _13273_, _08592_);
  or _22050_ (_13725_, _13724_, _13723_);
  and _22051_ (_13726_, _13266_, _08606_);
  and _22052_ (_13727_, _13262_, _08623_);
  or _22053_ (_13728_, _13727_, _13726_);
  or _22054_ (_13730_, _13728_, _13725_);
  or _22055_ (_13731_, _13730_, _08821_);
  and _22056_ (_13732_, _13246_, _08606_);
  and _22057_ (_13733_, _13238_, _08613_);
  or _22058_ (_13734_, _13733_, _13732_);
  and _22059_ (_13736_, _13252_, _08592_);
  and _22060_ (_13737_, _13242_, _08623_);
  or _22061_ (_13738_, _13737_, _13736_);
  or _22062_ (_13739_, _13738_, _13734_);
  or _22063_ (_13740_, _13739_, _08860_);
  nand _22064_ (_13741_, _13740_, _13731_);
  nor _22065_ (_13742_, _13741_, _08850_);
  or _22066_ (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _13742_, _13722_);
  and _22067_ (_13743_, _08908_, word_in[24]);
  and _22068_ (_13744_, _13286_, _08759_);
  and _22069_ (_13746_, _13282_, _08758_);
  or _22070_ (_13747_, _13746_, _13744_);
  and _22071_ (_13748_, _13747_, _08885_);
  and _22072_ (_13749_, _13296_, _08759_);
  and _22073_ (_13750_, _13292_, _08758_);
  or _22074_ (_13751_, _13750_, _13749_);
  and _22075_ (_13752_, _13751_, _08880_);
  and _22076_ (_13753_, _13306_, _08759_);
  and _22077_ (_13754_, _13302_, _08758_);
  or _22078_ (_13755_, _13754_, _13753_);
  and _22079_ (_13756_, _13755_, _08917_);
  and _22080_ (_13757_, _13316_, _08759_);
  and _22081_ (_13759_, _13312_, _08758_);
  or _22082_ (_13760_, _13759_, _13757_);
  and _22083_ (_13761_, _13760_, _08925_);
  or _22084_ (_13762_, _13761_, _13756_);
  or _22085_ (_13763_, _13762_, _13752_);
  nor _22086_ (_13764_, _13763_, _13748_);
  nor _22087_ (_13765_, _13764_, _08908_);
  or _22088_ (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _13765_, _13743_);
  and _22089_ (_13767_, _08908_, word_in[25]);
  and _22090_ (_13769_, _13331_, _08759_);
  and _22091_ (_13770_, _13327_, _08758_);
  or _22092_ (_13771_, _13770_, _13769_);
  and _22093_ (_13772_, _13771_, _08885_);
  and _22094_ (_13773_, _13341_, _08759_);
  and _22095_ (_13774_, _13337_, _08758_);
  or _22096_ (_13775_, _13774_, _13773_);
  and _22097_ (_13776_, _13775_, _08880_);
  and _22098_ (_13777_, _13352_, _08759_);
  and _22099_ (_13778_, _13348_, _08758_);
  or _22100_ (_13779_, _13778_, _13777_);
  and _22101_ (_13780_, _13779_, _08917_);
  and _22102_ (_13781_, _13362_, _08759_);
  and _22103_ (_13782_, _13358_, _08758_);
  or _22104_ (_13783_, _13782_, _13781_);
  and _22105_ (_13784_, _13783_, _08925_);
  or _22106_ (_13785_, _13784_, _13780_);
  or _22107_ (_13786_, _13785_, _13776_);
  nor _22108_ (_13787_, _13786_, _13772_);
  nor _22109_ (_13789_, _13787_, _08908_);
  or _22110_ (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _13789_, _13767_);
  and _22111_ (_13790_, _08908_, word_in[26]);
  and _22112_ (_13791_, _13378_, _08759_);
  and _22113_ (_13792_, _13374_, _08758_);
  or _22114_ (_13793_, _13792_, _13791_);
  and _22115_ (_13794_, _13793_, _08885_);
  and _22116_ (_13795_, _13388_, _08759_);
  and _22117_ (_13796_, _13384_, _08758_);
  or _22118_ (_13797_, _13796_, _13795_);
  and _22119_ (_13799_, _13797_, _08880_);
  and _22120_ (_13800_, _13398_, _08759_);
  and _22121_ (_13801_, _13394_, _08758_);
  or _22122_ (_13803_, _13801_, _13800_);
  and _22123_ (_13804_, _13803_, _08917_);
  and _22124_ (_13805_, _13408_, _08759_);
  and _22125_ (_13806_, _13404_, _08758_);
  or _22126_ (_13807_, _13806_, _13805_);
  and _22127_ (_13808_, _13807_, _08925_);
  or _22128_ (_13810_, _13808_, _13804_);
  or _22129_ (_13811_, _13810_, _13799_);
  nor _22130_ (_13813_, _13811_, _13794_);
  nor _22131_ (_13814_, _13813_, _08908_);
  or _22132_ (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _13814_, _13790_);
  and _22133_ (_13816_, _08908_, word_in[27]);
  and _22134_ (_13818_, _13435_, _08759_);
  and _22135_ (_13819_, _13431_, _08758_);
  or _22136_ (_13820_, _13819_, _13818_);
  and _22137_ (_13821_, _13820_, _08880_);
  and _22138_ (_13823_, _13425_, _08759_);
  and _22139_ (_13824_, _13420_, _08758_);
  or _22140_ (_13825_, _13824_, _13823_);
  and _22141_ (_13826_, _13825_, _08885_);
  and _22142_ (_13827_, _13445_, _08759_);
  and _22143_ (_13828_, _13441_, _08758_);
  or _22144_ (_13829_, _13828_, _13827_);
  and _22145_ (_13830_, _13829_, _08917_);
  and _22146_ (_13831_, _13456_, _08759_);
  and _22147_ (_13832_, _13452_, _08758_);
  or _22148_ (_13833_, _13832_, _13831_);
  and _22149_ (_13834_, _13833_, _08925_);
  or _22150_ (_13835_, _13834_, _13830_);
  or _22151_ (_13836_, _13835_, _13826_);
  nor _22152_ (_13837_, _13836_, _13821_);
  nor _22153_ (_13838_, _13837_, _08908_);
  or _22154_ (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _13838_, _13816_);
  and _22155_ (_13839_, _08908_, word_in[28]);
  and _22156_ (_13840_, _13472_, _08759_);
  and _22157_ (_13841_, _13468_, _08758_);
  or _22158_ (_13842_, _13841_, _13840_);
  and _22159_ (_13843_, _13842_, _08885_);
  and _22160_ (_13844_, _13482_, _08759_);
  and _22161_ (_13845_, _13478_, _08758_);
  or _22162_ (_13846_, _13845_, _13844_);
  and _22163_ (_13847_, _13846_, _08880_);
  and _22164_ (_13848_, _13492_, _08759_);
  and _22165_ (_13849_, _13488_, _08758_);
  or _22166_ (_13850_, _13849_, _13848_);
  and _22167_ (_13851_, _13850_, _08917_);
  and _22168_ (_13852_, _13502_, _08759_);
  and _22169_ (_13853_, _13498_, _08758_);
  or _22170_ (_13854_, _13853_, _13852_);
  and _22171_ (_13855_, _13854_, _08925_);
  or _22172_ (_13856_, _13855_, _13851_);
  or _22173_ (_13857_, _13856_, _13847_);
  nor _22174_ (_13858_, _13857_, _13843_);
  nor _22175_ (_13859_, _13858_, _08908_);
  or _22176_ (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _13859_, _13839_);
  and _22177_ (_13860_, _08908_, word_in[29]);
  and _22178_ (_13861_, _13517_, _08759_);
  and _22179_ (_13862_, _13513_, _08758_);
  or _22180_ (_13863_, _13862_, _13861_);
  and _22181_ (_13864_, _13863_, _08885_);
  and _22182_ (_13865_, _13527_, _08759_);
  and _22183_ (_13866_, _13523_, _08758_);
  or _22184_ (_13867_, _13866_, _13865_);
  and _22185_ (_13868_, _13867_, _08880_);
  and _22186_ (_13869_, _13537_, _08759_);
  and _22187_ (_13870_, _13533_, _08758_);
  or _22188_ (_13871_, _13870_, _13869_);
  and _22189_ (_13873_, _13871_, _08917_);
  and _22190_ (_13874_, _13547_, _08759_);
  and _22191_ (_13875_, _13543_, _08758_);
  or _22192_ (_13876_, _13875_, _13874_);
  and _22193_ (_13877_, _13876_, _08925_);
  or _22194_ (_13878_, _13877_, _13873_);
  or _22195_ (_13879_, _13878_, _13868_);
  nor _22196_ (_13880_, _13879_, _13864_);
  nor _22197_ (_13881_, _13880_, _08908_);
  or _22198_ (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _13881_, _13860_);
  and _22199_ (_13882_, _08908_, word_in[30]);
  and _22200_ (_13883_, _13572_, _08759_);
  and _22201_ (_13885_, _13568_, _08758_);
  or _22202_ (_13886_, _13885_, _13883_);
  and _22203_ (_13887_, _13886_, _08880_);
  and _22204_ (_13888_, _13562_, _08759_);
  and _22205_ (_13889_, _13558_, _08758_);
  or _22206_ (_13890_, _13889_, _13888_);
  and _22207_ (_13891_, _13890_, _08885_);
  and _22208_ (_13892_, _13584_, _08759_);
  and _22209_ (_13893_, _13579_, _08758_);
  or _22210_ (_13894_, _13893_, _13892_);
  and _22211_ (_13895_, _13894_, _08917_);
  and _22212_ (_13896_, _13595_, _08759_);
  and _22213_ (_13897_, _13590_, _08758_);
  or _22214_ (_13898_, _13897_, _13896_);
  and _22215_ (_13899_, _13898_, _08925_);
  or _22216_ (_13900_, _13899_, _13895_);
  or _22217_ (_13901_, _13900_, _13891_);
  nor _22218_ (_13902_, _13901_, _13887_);
  nor _22219_ (_13903_, _13902_, _08908_);
  or _22220_ (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _13903_, _13882_);
  and _22221_ (_11200_, _08085_, _06989_);
  and _22222_ (_11222_, _09182_, _06989_);
  and _22223_ (_11228_, _07978_, _06989_);
  and _22224_ (_11259_, _08231_, _06989_);
  and _22225_ (_11268_, _08317_, _06989_);
  nor _22226_ (_13904_, _07027_, _07662_);
  and _22227_ (_13905_, _07027_, _07662_);
  or _22228_ (_13906_, _13905_, _13904_);
  and _22229_ (_11307_, _13906_, _06989_);
  and _22230_ (_11318_, _07691_, _06989_);
  and _22231_ (_11323_, _07684_, _06989_);
  and _22232_ (_11357_, _08197_, _06989_);
  and _22233_ (_11362_, _08302_, _06989_);
  and _22234_ (_11384_, _08380_, _06989_);
  and _22235_ (_11434_, _09280_, _06989_);
  or _22236_ (_13909_, _09389_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or _22237_ (_13911_, _09516_, _09418_);
  and _22238_ (_11465_, _13911_, _13909_);
  and _22239_ (_11487_, _09349_, _06989_);
  or _22240_ (_13912_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  or _22241_ (_13913_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and _22242_ (_13915_, _13913_, _06989_);
  and _22243_ (_11544_, _13915_, _13912_);
  and _22244_ (_13916_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and _22245_ (_13917_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or _22246_ (_13918_, _13917_, _13916_);
  and _22247_ (_11592_, _13918_, _06989_);
  and _22248_ (_11633_, _08402_, _06989_);
  and _22249_ (_13920_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _22250_ (_13921_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _22251_ (_13922_, _08139_, _13921_);
  or _22252_ (_13923_, _13922_, _13920_);
  and _22253_ (_11677_, _13923_, _06989_);
  and _22254_ (_13924_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor _22255_ (_13925_, _07493_, _11081_);
  or _22256_ (_13926_, _13925_, _13924_);
  and _22257_ (_11826_, _13926_, _06989_);
  or _22258_ (_13927_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  or _22259_ (_13928_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  and _22260_ (_13929_, _13928_, _06989_);
  and _22261_ (_11831_, _13929_, _13927_);
  and _22262_ (_13930_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and _22263_ (_13931_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  or _22264_ (_13932_, _13931_, _13930_);
  and _22265_ (_11847_, _13932_, _06989_);
  or _22266_ (_13933_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  or _22267_ (_13934_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and _22268_ (_13935_, _13934_, _06989_);
  and _22269_ (_11854_, _13935_, _13933_);
  nand _22270_ (_13936_, _11529_, _10146_);
  or _22271_ (_13937_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and _22272_ (_13938_, _13937_, _06989_);
  and _22273_ (_11893_, _13938_, _13936_);
  and _22274_ (_11967_, _07816_, _06989_);
  and _22275_ (_11997_, _08396_, _06989_);
  and _22276_ (_12000_, _09179_, _06989_);
  nor _22277_ (_13939_, _07262_, _07118_);
  and _22278_ (_13940_, _07262_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or _22279_ (_13941_, _13940_, _13939_);
  and _22280_ (_12039_, _13941_, _06989_);
  and _22281_ (_13942_, _09393_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and _22282_ (_13943_, _13942_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and _22283_ (_13944_, _13943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and _22284_ (_13945_, _13944_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and _22285_ (_13946_, _13945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or _22286_ (_13947_, _13946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand _22287_ (_13948_, _13946_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and _22288_ (_13949_, _13948_, _13947_);
  and _22289_ (_13950_, _07453_, _07085_);
  and _22290_ (_13951_, _06985_, _07089_);
  and _22291_ (_13952_, _13951_, _13950_);
  nor _22292_ (_13953_, _13952_, rst);
  and _22293_ (_12052_, _13953_, _13949_);
  and _22294_ (_13955_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor _22295_ (_13956_, _07493_, _12556_);
  or _22296_ (_13957_, _13956_, _13955_);
  and _22297_ (_12057_, _13957_, _06989_);
  and _22298_ (_13958_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.pres_ow );
  and _22299_ (_13959_, _13958_, _09392_);
  nor _22300_ (_13960_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _22301_ (_13961_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _22302_ (_13962_, _13961_, _13960_);
  nor _22303_ (_13963_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor _22304_ (_13964_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor _22305_ (_13965_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _22306_ (_13966_, _13965_, _13964_);
  and _22307_ (_13967_, _13966_, _13963_);
  and _22308_ (_13968_, _13967_, _13962_);
  not _22309_ (_13969_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor _22310_ (_13970_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _22311_ (_13971_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and _22312_ (_13972_, _13971_, _13970_);
  and _22313_ (_13973_, _13972_, _13969_);
  and _22314_ (_13974_, _13973_, _13968_);
  not _22315_ (_13975_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor _22316_ (_13976_, _13972_, _13975_);
  or _22317_ (_13977_, _13976_, _13974_);
  and _22318_ (_13978_, _13977_, _13943_);
  nand _22319_ (_13979_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _22320_ (_13980_, _13979_, _13942_);
  nor _22321_ (_13981_, _13980_, _13978_);
  nor _22322_ (_13982_, _13981_, _13959_);
  and _22323_ (_13983_, _13968_, _13959_);
  or _22324_ (_13984_, _13983_, _13982_);
  and _22325_ (_12060_, _13984_, _13953_);
  and _22326_ (_13985_, _07090_, _06983_);
  and _22327_ (_13986_, _13985_, _13950_);
  nand _22328_ (_13987_, _13974_, _13942_);
  nand _22329_ (_13988_, _13987_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor _22330_ (_13989_, _13988_, _13983_);
  or _22331_ (_13990_, _13989_, _13986_);
  and _22332_ (_12075_, _13990_, _06989_);
  not _22333_ (_13991_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and _22334_ (_13992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not _22335_ (_13993_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _22336_ (_13994_, _07462_, _13993_);
  not _22337_ (_13995_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor _22338_ (_13996_, _13995_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _22339_ (_13997_, _13996_, _13994_);
  nor _22340_ (_13998_, _13997_, _13992_);
  nand _22341_ (_13999_, _13998_, _13991_);
  nor _22342_ (_14000_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor _22343_ (_14001_, _14000_, _13998_);
  nand _22344_ (_14002_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand _22345_ (_14003_, _14002_, _14001_);
  and _22346_ (_14004_, _14003_, _06989_);
  and _22347_ (_12082_, _14004_, _13999_);
  and _22348_ (_12085_, _14001_, _06989_);
  and _22349_ (_14005_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  not _22350_ (_14007_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor _22351_ (_14008_, _07493_, _14007_);
  or _22352_ (_14010_, _14008_, _14005_);
  and _22353_ (_12104_, _14010_, _06989_);
  and _22354_ (_14011_, _09072_, _06539_);
  and _22355_ (_14012_, _14011_, _07454_);
  or _22356_ (_14013_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _22357_ (_14015_, _14013_, _06989_);
  and _22358_ (_14016_, _09239_, _06539_);
  nand _22359_ (_14017_, _14016_, _07040_);
  and _22360_ (_12115_, _14017_, _14015_);
  and _22361_ (_14018_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  not _22362_ (_14020_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor _22363_ (_14021_, _07493_, _14020_);
  or _22364_ (_14023_, _14021_, _14018_);
  and _22365_ (_12121_, _14023_, _06989_);
  nor _22366_ (_14025_, _06447_, _06434_);
  and _22367_ (_14026_, _06477_, _06463_);
  and _22368_ (_14027_, _14026_, _06500_);
  and _22369_ (_14028_, _14027_, _14025_);
  and _22370_ (_14029_, _14028_, _06539_);
  nand _22371_ (_14030_, _14029_, _06968_);
  and _22372_ (_14031_, _13950_, _06986_);
  not _22373_ (_14032_, _14031_);
  or _22374_ (_14033_, _14029_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and _22375_ (_14034_, _14033_, _14032_);
  and _22376_ (_14035_, _14034_, _14030_);
  nor _22377_ (_14036_, _14032_, _07040_);
  or _22378_ (_14037_, _14036_, _14035_);
  and _22379_ (_12128_, _14037_, _06989_);
  and _22380_ (_12133_, _08212_, _06989_);
  and _22381_ (_14038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not _22382_ (_14039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _22383_ (_14040_, _07462_, _14039_);
  or _22384_ (_14041_, _14040_, _13996_);
  nor _22385_ (_14042_, _14041_, _14038_);
  or _22386_ (_14043_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand _22387_ (_14044_, _14043_, _06989_);
  nor _22388_ (_12160_, _14044_, _14042_);
  nor _22389_ (_12170_, _07461_, rst);
  or _22390_ (_14045_, _09403_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  not _22391_ (_14046_, rxd_i);
  nand _22392_ (_14047_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _14046_);
  nand _22393_ (_14048_, _14047_, _09403_);
  and _22394_ (_14049_, _14048_, _09393_);
  and _22395_ (_14050_, _14049_, _14045_);
  or _22396_ (_14051_, _09414_, _09411_);
  or _22397_ (_14052_, _14051_, _14050_);
  and _22398_ (_12208_, _14052_, _09418_);
  and _22399_ (_14053_, _09763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _22400_ (_14054_, _14053_, _09396_);
  and _22401_ (_14055_, _09762_, _14054_);
  not _22402_ (_14056_, _09395_);
  nor _22403_ (_14057_, _14053_, _14056_);
  or _22404_ (_14058_, _14057_, _09760_);
  and _22405_ (_14060_, _14058_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or _22406_ (_14061_, _14060_, _14055_);
  and _22407_ (_12211_, _14061_, _06989_);
  and _22408_ (_14062_, _09764_, _09397_);
  and _22409_ (_14063_, _09762_, _14062_);
  nand _22410_ (_14065_, _14063_, _14046_);
  or _22411_ (_14066_, _14063_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and _22412_ (_14067_, _14066_, _06989_);
  and _22413_ (_12214_, _14067_, _14065_);
  not _22414_ (_14068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor _22415_ (_14069_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _09405_);
  not _22416_ (_14070_, _14069_);
  nor _22417_ (_14071_, _09392_, _09389_);
  and _22418_ (_14073_, _14071_, _14070_);
  and _22419_ (_14074_, _14073_, _14056_);
  nor _22420_ (_14076_, _14074_, _14068_);
  and _22421_ (_14077_, _14074_, rxd_i);
  or _22422_ (_14078_, _14077_, rst);
  or _22423_ (_12220_, _14078_, _14076_);
  or _22424_ (_14079_, _09420_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or _22425_ (_14080_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _22426_ (_14081_, _14080_, _09392_);
  or _22427_ (_14083_, _14081_, _09395_);
  nand _22428_ (_14084_, _14083_, _14079_);
  nand _22429_ (_12229_, _14084_, _09418_);
  nand _22430_ (_14086_, _07669_, _07027_);
  or _22431_ (_14088_, _07027_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and _22432_ (_14089_, _14088_, _06989_);
  and _22433_ (_12373_, _14089_, _14086_);
  and _22434_ (_12387_, _09086_, _06989_);
  and _22435_ (_14091_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  not _22436_ (_14092_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor _22437_ (_14093_, _07493_, _14092_);
  or _22438_ (_14094_, _14093_, _14091_);
  and _22439_ (_12405_, _14094_, _06989_);
  or _22440_ (_14095_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  or _22441_ (_14096_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and _22442_ (_14097_, _14096_, _06989_);
  and _22443_ (_12414_, _14097_, _14095_);
  and _22444_ (_14098_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not _22445_ (_14099_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor _22446_ (_14100_, _07493_, _14099_);
  or _22447_ (_14101_, _14100_, _14098_);
  and _22448_ (_12423_, _14101_, _06989_);
  and _22449_ (_14102_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or _22450_ (_12440_, _14102_, _09477_);
  and _22451_ (_14103_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  not _22452_ (_14104_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor _22453_ (_14106_, _07493_, _14104_);
  or _22454_ (_14107_, _14106_, _14103_);
  and _22455_ (_12441_, _14107_, _06989_);
  and _22456_ (_14109_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  not _22457_ (_14110_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor _22458_ (_14112_, _07493_, _14110_);
  or _22459_ (_14113_, _14112_, _14109_);
  and _22460_ (_12445_, _14113_, _06989_);
  and _22461_ (_14114_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and _22462_ (_14116_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or _22463_ (_14117_, _14116_, _14114_);
  and _22464_ (_12475_, _14117_, _06989_);
  or _22465_ (_14119_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or _22466_ (_14120_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and _22467_ (_14122_, _14120_, _06989_);
  and _22468_ (_12478_, _14122_, _14119_);
  nor _22469_ (_14124_, _07486_, _07260_);
  and _22470_ (_14125_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or _22471_ (_14126_, _14125_, _14124_);
  and _22472_ (_12548_, _14126_, _06989_);
  nor _22473_ (_14128_, _07486_, _07118_);
  and _22474_ (_14129_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or _22475_ (_14130_, _14129_, _14128_);
  and _22476_ (_12655_, _14130_, _06989_);
  nor _22477_ (_14131_, _12938_, _10970_);
  and _22478_ (_14132_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or _22479_ (_14133_, _14132_, _14131_);
  and _22480_ (_12672_, _14133_, _06989_);
  nor _22481_ (_14134_, _12938_, _07118_);
  and _22482_ (_14135_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or _22483_ (_14136_, _14135_, _14134_);
  and _22484_ (_12693_, _14136_, _06989_);
  and _22485_ (_14137_, _07262_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor _22486_ (_14138_, _07262_, _07040_);
  or _22487_ (_14140_, _14138_, _14137_);
  and _22488_ (_12810_, _14140_, _06989_);
  and _22489_ (_14141_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or _22490_ (_12863_, _14141_, _09391_);
  and _22491_ (_14143_, _07135_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and _22492_ (_14144_, _09488_, _09009_);
  or _22493_ (_14145_, _14144_, _14143_);
  and _22494_ (_12941_, _14145_, _06989_);
  and _22495_ (_12965_, _06989_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  not _22496_ (_14146_, _09010_);
  and _22497_ (_14147_, _14146_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor _22498_ (_14148_, _14146_, _07317_);
  or _22499_ (_14149_, _14148_, _14147_);
  and _22500_ (_12976_, _14149_, _06989_);
  or _22501_ (_14150_, _14056_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or _22502_ (_14151_, _14150_, _09401_);
  and _22503_ (_14152_, _14151_, _09481_);
  or _22504_ (_14153_, _14152_, rxd_i);
  and _22505_ (_14154_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], rxd_i);
  nor _22506_ (_14155_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  and _22507_ (_14156_, _14155_, _09395_);
  and _22508_ (_14157_, _14156_, _09400_);
  nor _22509_ (_14158_, _14157_, _09426_);
  and _22510_ (_14159_, _14158_, _14153_);
  or _22511_ (_14160_, _14159_, _09389_);
  nor _22512_ (_14161_, _09420_, _09389_);
  or _22513_ (_14162_, _14161_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and _22514_ (_14163_, _14162_, _06989_);
  and _22515_ (_13093_, _14163_, _14160_);
  and _22516_ (_14164_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor _22517_ (_14165_, _07493_, _12549_);
  or _22518_ (_14166_, _14165_, _14164_);
  and _22519_ (_13103_, _14166_, _06989_);
  and _22520_ (_13114_, _06989_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  and _22521_ (_13118_, _07643_, _06989_);
  and _22522_ (_14167_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  not _22523_ (_14168_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor _22524_ (_14169_, _07493_, _14168_);
  or _22525_ (_14170_, _14169_, _14167_);
  and _22526_ (_13137_, _14170_, _06989_);
  nand _22527_ (_14171_, _10146_, _07260_);
  or _22528_ (_14172_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and _22529_ (_14173_, _14172_, _06989_);
  and _22530_ (_13146_, _14173_, _14171_);
  and _22531_ (_14174_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and _22532_ (_14175_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or _22533_ (_14176_, _14175_, _14174_);
  and _22534_ (_13154_, _14176_, _06989_);
  nor _22535_ (_14177_, _11529_, _09614_);
  and _22536_ (_14178_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or _22537_ (_14179_, _14178_, _06982_);
  or _22538_ (_14180_, _14179_, _14177_);
  or _22539_ (_14181_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and _22540_ (_14182_, _14181_, _06989_);
  and _22541_ (_13157_, _14182_, _14180_);
  and _22542_ (_14183_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not _22543_ (_14184_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor _22544_ (_14185_, _07493_, _14184_);
  or _22545_ (_14186_, _14185_, _14183_);
  and _22546_ (_13207_, _14186_, _06989_);
  or _22547_ (_14187_, _09607_, _06982_);
  or _22548_ (_14188_, _14187_, _12943_);
  and _22549_ (_14189_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and _22550_ (_14190_, _08994_, _06981_);
  and _22551_ (_14191_, _14190_, _11821_);
  or _22552_ (_14192_, _14191_, _14189_);
  and _22553_ (_13272_, _14192_, _06989_);
  and _22554_ (_14193_, _07135_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  nor _22555_ (_14194_, _09489_, _07040_);
  or _22556_ (_14195_, _14194_, _14193_);
  and _22557_ (_13343_, _14195_, _06989_);
  and _22558_ (_14196_, _06538_, _06513_);
  and _22559_ (_14197_, _14028_, _14196_);
  nand _22560_ (_14198_, _14197_, _06968_);
  or _22561_ (_14199_, _14197_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _22562_ (_14200_, _14199_, _14032_);
  and _22563_ (_14201_, _14200_, _14198_);
  nor _22564_ (_14202_, _14032_, _10970_);
  or _22565_ (_14203_, _14202_, _14201_);
  and _22566_ (_13365_, _14203_, _06989_);
  not _22567_ (_14204_, _11799_);
  nor _22568_ (_14205_, _14204_, _11748_);
  and _22569_ (_14206_, _11724_, _11688_);
  not _22570_ (_14207_, _11613_);
  and _22571_ (_14208_, _11652_, _14207_);
  and _22572_ (_14209_, _14208_, _14206_);
  and _22573_ (_14210_, _11857_, _11556_);
  and _22574_ (_14211_, _14210_, _14209_);
  and _22575_ (_14212_, _14211_, _14205_);
  and _22576_ (_14213_, _14212_, _09071_);
  nor _22577_ (_14214_, _11652_, _11613_);
  and _22578_ (_14215_, _14206_, _14214_);
  and _22579_ (_14217_, _11799_, _11748_);
  nor _22580_ (_14218_, _11857_, _11556_);
  and _22581_ (_14219_, _14218_, _14217_);
  and _22582_ (_14220_, _14219_, _14215_);
  and _22583_ (_14221_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  not _22584_ (_14222_, _11556_);
  and _22585_ (_14223_, _11857_, _14222_);
  and _22586_ (_14224_, _14217_, _14223_);
  and _22587_ (_14226_, _14224_, _14215_);
  and _22588_ (_14228_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _22589_ (_14229_, _14228_, _14221_);
  and _22590_ (_14230_, _14223_, _14205_);
  and _22591_ (_14231_, _14230_, _14215_);
  and _22592_ (_14232_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and _22593_ (_14233_, _14204_, _11748_);
  and _22594_ (_14234_, _14233_, _14218_);
  and _22595_ (_14235_, _14234_, _14215_);
  and _22596_ (_14236_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _22597_ (_14237_, _14236_, _14232_);
  or _22598_ (_14238_, _14237_, _14229_);
  and _22599_ (_14239_, _14224_, _14209_);
  and _22600_ (_14240_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _22601_ (_14241_, _11799_, _11748_);
  and _22602_ (_14242_, _14241_, _14223_);
  and _22603_ (_14243_, _14242_, _14215_);
  and _22604_ (_14244_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or _22605_ (_14245_, _14244_, _14240_);
  not _22606_ (_14246_, _11688_);
  and _22607_ (_14247_, _14208_, _14246_);
  and _22608_ (_14248_, _14247_, _11724_);
  and _22609_ (_14249_, _14248_, _14224_);
  and _22610_ (_14250_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  not _22611_ (_14251_, _11724_);
  and _22612_ (_14252_, _14247_, _14251_);
  not _22613_ (_14253_, _11857_);
  and _22614_ (_14254_, _14241_, _14253_);
  and _22615_ (_14256_, _14254_, _11556_);
  and _22616_ (_14257_, _14256_, _14252_);
  and _22617_ (_14258_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _22618_ (_14259_, _14258_, _14250_);
  or _22619_ (_14260_, _14259_, _14245_);
  or _22620_ (_14261_, _14260_, _14238_);
  and _22621_ (_14262_, _14233_, _14223_);
  and _22622_ (_14263_, _14262_, _14209_);
  and _22623_ (_14265_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _22624_ (_14266_, _14242_, _14209_);
  and _22625_ (_14267_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _22626_ (_14268_, _14267_, _14265_);
  and _22627_ (_14269_, _14234_, _14209_);
  and _22628_ (_14270_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _22629_ (_14271_, _14209_, _14230_);
  and _22630_ (_14272_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or _22631_ (_14273_, _14272_, _14270_);
  or _22632_ (_14274_, _14273_, _14268_);
  and _22633_ (_14275_, _14208_, _11688_);
  and _22634_ (_14276_, _14275_, _14251_);
  and _22635_ (_14277_, _14276_, _14224_);
  and _22636_ (_14278_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and _22637_ (_14279_, _14276_, _14262_);
  and _22638_ (_14280_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or _22639_ (_14281_, _14280_, _14278_);
  and _22640_ (_14282_, _14219_, _14209_);
  and _22641_ (_14283_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _22642_ (_14284_, _14256_, _14209_);
  and _22643_ (_14285_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or _22644_ (_14286_, _14285_, _14283_);
  or _22645_ (_14287_, _14286_, _14281_);
  or _22646_ (_14288_, _14287_, _14274_);
  or _22647_ (_14289_, _14288_, _14261_);
  and _22648_ (_14290_, _14217_, _14210_);
  and _22649_ (_14291_, _14290_, _14251_);
  and _22650_ (_14292_, _14214_, _14246_);
  and _22651_ (_14293_, _14292_, _14291_);
  and _22652_ (_14294_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _22653_ (_14295_, _14233_, _14210_);
  and _22654_ (_14296_, _14295_, _14209_);
  and _22655_ (_14297_, _14296_, _11627_);
  or _22656_ (_14298_, _14297_, _14294_);
  and _22657_ (_14299_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and _22658_ (_14300_, _14241_, _14210_);
  and _22659_ (_14301_, _14300_, _14209_);
  and _22660_ (_14302_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or _22661_ (_14303_, _14302_, _14299_);
  or _22662_ (_14304_, _14303_, _14298_);
  and _22663_ (_14305_, _14252_, _14290_);
  nor _22664_ (_14306_, _11460_, _11401_);
  nor _22665_ (_14307_, _11330_, _11299_);
  and _22666_ (_14308_, _14307_, _11295_);
  nor _22667_ (_14309_, _14308_, _11473_);
  nor _22668_ (_14310_, _11912_, _11452_);
  and _22669_ (_14311_, _14310_, _14309_);
  and _22670_ (_14312_, _14311_, _14306_);
  and _22671_ (_14313_, _11908_, _11403_);
  not _22672_ (_14314_, _14313_);
  and _22673_ (_14315_, _14314_, _11457_);
  and _22674_ (_14316_, _11396_, _11364_);
  and _22675_ (_14317_, _11478_, _11322_);
  nor _22676_ (_14318_, _14317_, _14316_);
  and _22677_ (_14319_, _11382_, _11375_);
  and _22678_ (_14320_, _11462_, _11321_);
  nor _22679_ (_14321_, _14320_, _14319_);
  and _22680_ (_14322_, _14321_, _14318_);
  and _22681_ (_14323_, _14322_, _14315_);
  and _22682_ (_14324_, _14323_, _14312_);
  and _22683_ (_14325_, _14324_, _11443_);
  nor _22684_ (_14326_, _14325_, _11283_);
  or _22685_ (_14327_, _14326_, p3_in[6]);
  not _22686_ (_14328_, _14326_);
  or _22687_ (_14329_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _22688_ (_14330_, _14329_, _14327_);
  and _22689_ (_14331_, _14330_, _14305_);
  and _22690_ (_14332_, _14290_, _11724_);
  and _22691_ (_14333_, _14332_, _14247_);
  or _22692_ (_14334_, _14326_, p2_in[6]);
  or _22693_ (_14335_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _22694_ (_14336_, _14335_, _14334_);
  and _22695_ (_14337_, _14336_, _14333_);
  or _22696_ (_14338_, _14337_, _14331_);
  and _22697_ (_14339_, _14290_, _14209_);
  or _22698_ (_14340_, _14326_, p0_in[6]);
  or _22699_ (_14341_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _22700_ (_14342_, _14341_, _14340_);
  and _22701_ (_14343_, _14342_, _14339_);
  and _22702_ (_14344_, _14291_, _14275_);
  or _22703_ (_14345_, _14326_, p1_in[6]);
  or _22704_ (_14346_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _22705_ (_14347_, _14346_, _14345_);
  and _22706_ (_14348_, _14347_, _14344_);
  or _22707_ (_14349_, _14348_, _14343_);
  or _22708_ (_14350_, _14349_, _14338_);
  or _22709_ (_14351_, _14350_, _14304_);
  and _22710_ (_14352_, _14332_, _14292_);
  and _22711_ (_14353_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and _22712_ (_14354_, _14214_, _11688_);
  and _22713_ (_14355_, _14291_, _14354_);
  and _22714_ (_14356_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or _22715_ (_14357_, _14356_, _14353_);
  or _22716_ (_14358_, _14357_, _14351_);
  or _22717_ (_14359_, _14358_, _14289_);
  and _22718_ (_14360_, _14355_, _11951_);
  and _22719_ (_14361_, _14352_, _07699_);
  and _22720_ (_14362_, _14241_, _14211_);
  and _22721_ (_14363_, _14362_, _09071_);
  or _22722_ (_14364_, _14363_, _14361_);
  nor _22723_ (_14365_, _14364_, _14360_);
  nor _22724_ (_14366_, _14365_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not _22725_ (_14367_, _14366_);
  and _22726_ (_14368_, _14352_, _07705_);
  not _22727_ (_14369_, _06500_);
  nor _22728_ (_14370_, _14254_, _14369_);
  and _22729_ (_14371_, _14370_, _11730_);
  nor _22730_ (_14372_, _14371_, _14368_);
  and _22731_ (_14373_, _14372_, _11866_);
  and _22732_ (_14374_, _14373_, _14367_);
  and _22733_ (_14375_, _14374_, _14359_);
  not _22734_ (_14376_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  not _22735_ (_14377_, _14374_);
  nor _22736_ (_14378_, _14226_, _14220_);
  nor _22737_ (_14379_, _14235_, _14231_);
  and _22738_ (_14380_, _14379_, _14378_);
  nor _22739_ (_14381_, _14243_, _14239_);
  nor _22740_ (_14382_, _14257_, _14249_);
  and _22741_ (_14383_, _14382_, _14381_);
  and _22742_ (_14384_, _14383_, _14380_);
  nor _22743_ (_14385_, _14266_, _14263_);
  nor _22744_ (_14386_, _14271_, _14269_);
  and _22745_ (_14387_, _14386_, _14385_);
  nor _22746_ (_14388_, _14279_, _14277_);
  nor _22747_ (_14389_, _14284_, _14282_);
  and _22748_ (_14390_, _14389_, _14388_);
  and _22749_ (_14391_, _14390_, _14387_);
  and _22750_ (_14392_, _14391_, _14384_);
  nor _22751_ (_14394_, _14355_, _14352_);
  and _22752_ (_14395_, _14290_, _14208_);
  not _22753_ (_14396_, _14395_);
  nor _22754_ (_14397_, _14301_, _14212_);
  nor _22755_ (_14398_, _14296_, _14293_);
  and _22756_ (_14399_, _14398_, _14397_);
  and _22757_ (_14400_, _14399_, _14396_);
  and _22758_ (_14401_, _14400_, _14394_);
  and _22759_ (_14402_, _14401_, _14392_);
  nor _22760_ (_14404_, _14402_, _14377_);
  nor _22761_ (_14405_, _14404_, _14376_);
  or _22762_ (_14406_, _14405_, _14375_);
  or _22763_ (_14407_, _14406_, _14213_);
  nand _22764_ (_14408_, _14213_, _09145_);
  and _22765_ (_14409_, _14408_, _06989_);
  and _22766_ (_13423_, _14409_, _14407_);
  and _22767_ (_14410_, _07262_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and _22768_ (_14411_, _09009_, _07261_);
  or _22769_ (_14412_, _14411_, _14410_);
  and _22770_ (_13446_, _14412_, _06989_);
  and _22771_ (_13463_, _07814_, _06989_);
  and _22772_ (_14413_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _22773_ (_14414_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _22774_ (_14415_, _14414_, _14413_);
  and _22775_ (_14416_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _22776_ (_14417_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _22777_ (_14418_, _14417_, _14416_);
  or _22778_ (_14419_, _14418_, _14415_);
  and _22779_ (_14420_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and _22780_ (_14421_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or _22781_ (_14422_, _14421_, _14420_);
  and _22782_ (_14423_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _22783_ (_14424_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _22784_ (_14425_, _14424_, _14423_);
  or _22785_ (_14426_, _14425_, _14422_);
  or _22786_ (_14427_, _14426_, _14419_);
  and _22787_ (_14428_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _22788_ (_14429_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _22789_ (_14430_, _14429_, _14428_);
  and _22790_ (_14431_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _22791_ (_14432_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or _22792_ (_14433_, _14432_, _14431_);
  or _22793_ (_14434_, _14433_, _14430_);
  and _22794_ (_14435_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and _22795_ (_14436_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or _22796_ (_14437_, _14436_, _14435_);
  and _22797_ (_14438_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _22798_ (_14439_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or _22799_ (_14440_, _14439_, _14438_);
  or _22800_ (_14441_, _14440_, _14437_);
  or _22801_ (_14442_, _14441_, _14434_);
  or _22802_ (_14443_, _14442_, _14427_);
  and _22803_ (_14444_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and _22804_ (_14445_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or _22805_ (_14446_, _14445_, _14444_);
  and _22806_ (_14447_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and _22807_ (_14448_, _14296_, _11549_);
  or _22808_ (_14449_, _14448_, _14447_);
  or _22809_ (_14450_, _14449_, _14446_);
  or _22810_ (_14451_, _14326_, p2_in[3]);
  or _22811_ (_14452_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _22812_ (_14453_, _14452_, _14451_);
  and _22813_ (_14454_, _14453_, _14333_);
  or _22814_ (_14455_, _14326_, p3_in[3]);
  or _22815_ (_14457_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _22816_ (_14458_, _14457_, _14455_);
  and _22817_ (_14459_, _14458_, _14305_);
  or _22818_ (_14460_, _14459_, _14454_);
  or _22819_ (_14461_, _14326_, p0_in[3]);
  or _22820_ (_14462_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _22821_ (_14463_, _14462_, _14461_);
  and _22822_ (_14464_, _14463_, _14339_);
  or _22823_ (_14465_, _14326_, p1_in[3]);
  or _22824_ (_14466_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _22825_ (_14467_, _14466_, _14465_);
  and _22826_ (_14468_, _14467_, _14344_);
  or _22827_ (_14469_, _14468_, _14464_);
  or _22828_ (_14470_, _14469_, _14460_);
  or _22829_ (_14471_, _14470_, _14450_);
  and _22830_ (_14472_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and _22831_ (_14473_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or _22832_ (_14474_, _14473_, _14472_);
  or _22833_ (_14475_, _14474_, _14471_);
  or _22834_ (_14476_, _14475_, _14443_);
  not _22835_ (_14477_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nor _22836_ (_14478_, _14404_, _14477_);
  or _22837_ (_14479_, _14478_, _14476_);
  or _22838_ (_14480_, _14374_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and _22839_ (_14481_, _14480_, _14479_);
  or _22840_ (_14482_, _14481_, _14213_);
  not _22841_ (_14483_, _14213_);
  or _22842_ (_14484_, _14483_, _08433_);
  and _22843_ (_14485_, _14484_, _06989_);
  and _22844_ (_13573_, _14485_, _14482_);
  not _22845_ (_14486_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nor _22846_ (_14487_, _14404_, _14486_);
  nand _22847_ (_14488_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  nand _22848_ (_14489_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and _22849_ (_14490_, _14489_, _14488_);
  nand _22850_ (_14491_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nand _22851_ (_14492_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _22852_ (_14493_, _14492_, _14491_);
  and _22853_ (_14494_, _14493_, _14490_);
  nand _22854_ (_14495_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand _22855_ (_14496_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _22856_ (_14497_, _14496_, _14495_);
  nand _22857_ (_14498_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nand _22858_ (_14499_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _22859_ (_14500_, _14499_, _14498_);
  and _22860_ (_14501_, _14500_, _14497_);
  and _22861_ (_14502_, _14501_, _14494_);
  nand _22862_ (_14503_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nand _22863_ (_14504_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _22864_ (_14505_, _14504_, _14503_);
  nand _22865_ (_14506_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nand _22866_ (_14507_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _22867_ (_14508_, _14507_, _14506_);
  and _22868_ (_14509_, _14508_, _14505_);
  nand _22869_ (_14510_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nand _22870_ (_14511_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  and _22871_ (_14512_, _14511_, _14510_);
  nand _22872_ (_14513_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _22873_ (_14514_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _22874_ (_14515_, _14514_, _14513_);
  and _22875_ (_14516_, _14515_, _14512_);
  and _22876_ (_14517_, _14516_, _14509_);
  and _22877_ (_14518_, _14517_, _14502_);
  nand _22878_ (_14519_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _22879_ (_14520_, _14296_, _11852_);
  and _22880_ (_14521_, _14520_, _14519_);
  nand _22881_ (_14522_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  nand _22882_ (_14523_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and _22883_ (_14524_, _14523_, _14522_);
  and _22884_ (_14525_, _14524_, _14521_);
  nor _22885_ (_14526_, _14326_, p0_in[2]);
  not _22886_ (_14527_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _22887_ (_14528_, _14326_, _14527_);
  nor _22888_ (_14529_, _14528_, _14526_);
  nand _22889_ (_14530_, _14529_, _14339_);
  nor _22890_ (_14531_, _14326_, p1_in[2]);
  not _22891_ (_14532_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _22892_ (_14533_, _14326_, _14532_);
  nor _22893_ (_14534_, _14533_, _14531_);
  nand _22894_ (_14535_, _14534_, _14344_);
  and _22895_ (_14536_, _14535_, _14530_);
  nor _22896_ (_14537_, _14326_, p3_in[2]);
  not _22897_ (_14538_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _22898_ (_14539_, _14326_, _14538_);
  nor _22899_ (_14540_, _14539_, _14537_);
  nand _22900_ (_14541_, _14540_, _14305_);
  or _22901_ (_14542_, _14326_, p2_in[2]);
  or _22902_ (_14543_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _22903_ (_14544_, _14543_, _14542_);
  nand _22904_ (_14545_, _14544_, _14333_);
  and _22905_ (_14546_, _14545_, _14541_);
  and _22906_ (_14547_, _14546_, _14536_);
  and _22907_ (_14548_, _14547_, _14525_);
  nand _22908_ (_14549_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand _22909_ (_14550_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and _22910_ (_14551_, _14550_, _14549_);
  and _22911_ (_14552_, _14551_, _14548_);
  nand _22912_ (_14553_, _14552_, _14518_);
  nand _22913_ (_14554_, _14553_, _14374_);
  nand _22914_ (_14555_, _14554_, _14483_);
  or _22915_ (_14556_, _14555_, _14487_);
  nand _22916_ (_14557_, _14213_, _09227_);
  and _22917_ (_14558_, _14557_, _06989_);
  and _22918_ (_13580_, _14558_, _14556_);
  and _22919_ (_14559_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _22920_ (_14560_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _22921_ (_14561_, _14560_, _14559_);
  and _22922_ (_14562_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _22923_ (_14563_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _22924_ (_14564_, _14563_, _14562_);
  or _22925_ (_14565_, _14564_, _14561_);
  and _22926_ (_14566_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _22927_ (_14567_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _22928_ (_14568_, _14567_, _14566_);
  and _22929_ (_14569_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _22930_ (_14570_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or _22931_ (_14571_, _14570_, _14569_);
  or _22932_ (_14573_, _14571_, _14568_);
  or _22933_ (_14574_, _14573_, _14565_);
  and _22934_ (_14575_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _22935_ (_14576_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _22936_ (_14577_, _14576_, _14575_);
  and _22937_ (_14578_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _22938_ (_14579_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _22939_ (_14580_, _14579_, _14578_);
  or _22940_ (_14581_, _14580_, _14577_);
  and _22941_ (_14582_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and _22942_ (_14584_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _22943_ (_14586_, _14584_, _14582_);
  and _22944_ (_14587_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _22945_ (_14588_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or _22946_ (_14589_, _14588_, _14587_);
  or _22947_ (_14590_, _14589_, _14586_);
  or _22948_ (_14591_, _14590_, _14581_);
  or _22949_ (_14592_, _14591_, _14574_);
  and _22950_ (_14593_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _22951_ (_14594_, _14296_, _11740_);
  or _22952_ (_14595_, _14594_, _14593_);
  and _22953_ (_14596_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and _22954_ (_14597_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or _22955_ (_14598_, _14597_, _14596_);
  or _22956_ (_14599_, _14598_, _14595_);
  or _22957_ (_14600_, _14326_, p0_in[1]);
  or _22958_ (_14601_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _22959_ (_14602_, _14601_, _14600_);
  and _22960_ (_14603_, _14602_, _14339_);
  or _22961_ (_14604_, _14326_, p1_in[1]);
  or _22962_ (_14605_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _22963_ (_14606_, _14605_, _14604_);
  and _22964_ (_14608_, _14606_, _14344_);
  or _22965_ (_14609_, _14608_, _14603_);
  or _22966_ (_14610_, _14326_, p3_in[1]);
  or _22967_ (_14611_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _22968_ (_14612_, _14611_, _14610_);
  and _22969_ (_14613_, _14612_, _14305_);
  or _22970_ (_14614_, _14326_, p2_in[1]);
  or _22971_ (_14615_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _22972_ (_14616_, _14615_, _14614_);
  and _22973_ (_14617_, _14616_, _14333_);
  or _22974_ (_14618_, _14617_, _14613_);
  or _22975_ (_14619_, _14618_, _14609_);
  or _22976_ (_14620_, _14619_, _14599_);
  and _22977_ (_14621_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _22978_ (_14622_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _22979_ (_14623_, _14622_, _14621_);
  or _22980_ (_14624_, _14623_, _14620_);
  or _22981_ (_14625_, _14624_, _14592_);
  not _22982_ (_14626_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nor _22983_ (_14627_, _14404_, _14626_);
  or _22984_ (_14628_, _14627_, _14625_);
  or _22985_ (_14629_, _14374_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and _22986_ (_14630_, _14629_, _14628_);
  or _22987_ (_14631_, _14630_, _14213_);
  or _22988_ (_14632_, _14483_, _08030_);
  and _22989_ (_14633_, _14632_, _06989_);
  and _22990_ (_13592_, _14633_, _14631_);
  and _22991_ (_14634_, _07135_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor _22992_ (_14635_, _09489_, _07317_);
  or _22993_ (_14636_, _14635_, _14634_);
  and _22994_ (_13597_, _14636_, _06989_);
  or _22995_ (_14637_, _12278_, _09077_);
  or _22996_ (_14638_, _09079_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and _22997_ (_14639_, _14638_, _06989_);
  and _22998_ (_13649_, _14639_, _14637_);
  and _22999_ (_14640_, _09240_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _23000_ (_14641_, _12278_, _09292_);
  or _23001_ (_00001_, _14641_, _14640_);
  or _23002_ (_00002_, _00001_, _09071_);
  or _23003_ (_00003_, _12314_, _09369_);
  and _23004_ (_00004_, _00003_, _06989_);
  and _23005_ (_13651_, _00004_, _00002_);
  and _23006_ (_00005_, _13951_, _07454_);
  or _23007_ (_00006_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _23008_ (_00007_, _00006_, _06989_);
  nand _23009_ (_00008_, _00005_, _11529_);
  and _23010_ (_13707_, _00008_, _00007_);
  and _23011_ (_00010_, _13985_, _07454_);
  nand _23012_ (_00011_, _00010_, _09008_);
  or _23013_ (_00012_, _00010_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _23014_ (_00013_, _00012_, _06989_);
  and _23015_ (_13710_, _00013_, _00011_);
  or _23016_ (_00014_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and _23017_ (_00015_, _00014_, _06989_);
  nand _23018_ (_00016_, _00005_, _07317_);
  and _23019_ (_13729_, _00016_, _00015_);
  or _23020_ (_00017_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _23021_ (_00019_, _00017_, _06989_);
  nand _23022_ (_00020_, _00005_, _07260_);
  and _23023_ (_13735_, _00020_, _00019_);
  nand _23024_ (_00021_, _00010_, _09598_);
  or _23025_ (_00022_, _00010_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _23026_ (_00023_, _00022_, _06989_);
  and _23027_ (_13745_, _00023_, _00021_);
  and _23028_ (_00025_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or _23029_ (_13758_, _00025_, _09434_);
  and _23030_ (_00027_, _07454_, _07045_);
  nand _23031_ (_00029_, _00027_, _07118_);
  and _23032_ (_00030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _23033_ (_00032_, _00030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23034_ (_00033_, _00032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _23035_ (_00034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _23036_ (_00035_, _00034_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _23037_ (_00036_, t0_i);
  and _23038_ (_00037_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and _23039_ (_00038_, _00037_, _00036_);
  or _23040_ (_00039_, _00038_, _00035_);
  and _23041_ (_00040_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _23042_ (_00041_, _00040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and _23043_ (_00042_, _00041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _23044_ (_00043_, _00042_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _23045_ (_00044_, _00043_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _23046_ (_00045_, _00044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _23047_ (_00046_, _00045_, _00033_);
  and _23048_ (_00047_, _00046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _23049_ (_00049_, _00047_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _23050_ (_00051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not _23051_ (_00052_, _00051_);
  and _23052_ (_00053_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _23053_ (_00054_, _00053_, _00033_);
  and _23054_ (_00056_, _00054_, _00045_);
  nor _23055_ (_00057_, _00056_, _00052_);
  and _23056_ (_00058_, _00057_, _00049_);
  not _23057_ (_00059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nor _23058_ (_00060_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _00059_);
  and _23059_ (_00061_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _00059_);
  or _23060_ (_00062_, _00061_, _00060_);
  not _23061_ (_00063_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _23062_ (_00064_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and _23063_ (_00065_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and _23064_ (_00066_, _00065_, _00064_);
  and _23065_ (_00067_, _00066_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _23066_ (_00068_, _00067_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _23067_ (_00069_, _00068_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _23068_ (_00070_, _00069_, _00040_);
  and _23069_ (_00071_, _00070_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _23070_ (_00072_, _00071_, _00033_);
  and _23071_ (_00073_, _00072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _23072_ (_00074_, _00073_, _00059_);
  nor _23073_ (_00075_, _00074_, _00063_);
  and _23074_ (_00076_, _00074_, _00063_);
  or _23075_ (_00077_, _00076_, _00075_);
  and _23076_ (_00078_, _00077_, _00062_);
  and _23077_ (_00079_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and _23078_ (_00080_, _00079_, _00033_);
  and _23079_ (_00081_, _00080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _23080_ (_00082_, _00081_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _23081_ (_00083_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _23082_ (_00084_, _00080_, _00053_);
  not _23083_ (_00085_, _00084_);
  and _23084_ (_00086_, _00085_, _00083_);
  and _23085_ (_00087_, _00086_, _00082_);
  or _23086_ (_00088_, _00087_, _00078_);
  or _23087_ (_00089_, _00088_, _00058_);
  or _23088_ (_00090_, _00089_, _00027_);
  and _23089_ (_00091_, _09075_, _06985_);
  not _23090_ (_00092_, _00091_);
  and _23091_ (_00093_, _00092_, _00090_);
  and _23092_ (_00094_, _00093_, _00029_);
  and _23093_ (_00095_, _00091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or _23094_ (_00096_, _00095_, _00094_);
  and _23095_ (_13766_, _00096_, _06989_);
  not _23096_ (_00097_, _00027_);
  nor _23097_ (_00098_, _00097_, _10970_);
  and _23098_ (_00099_, _00056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _23099_ (_00100_, _00056_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _23100_ (_00101_, _00100_, _00051_);
  nor _23101_ (_00102_, _00101_, _00099_);
  and _23102_ (_00103_, _00054_, _00071_);
  or _23103_ (_00104_, _00103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _23104_ (_00105_, _00103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not _23105_ (_00106_, _00105_);
  and _23106_ (_00107_, _00106_, _00061_);
  and _23107_ (_00108_, _00107_, _00104_);
  and _23108_ (_00109_, _00080_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _23109_ (_00110_, _00109_, _00053_);
  or _23110_ (_00112_, _00110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand _23111_ (_00114_, _00110_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _23112_ (_00115_, _00114_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and _23113_ (_00116_, _00115_, _00112_);
  or _23114_ (_00118_, _00116_, _00108_);
  nor _23115_ (_00120_, _00118_, _00102_);
  nor _23116_ (_00122_, _00120_, _00027_);
  or _23117_ (_00124_, _00122_, _00091_);
  or _23118_ (_00125_, _00124_, _00098_);
  or _23119_ (_00126_, _00092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _23120_ (_00127_, _00126_, _06989_);
  and _23121_ (_13768_, _00127_, _00125_);
  and _23122_ (_00129_, _00071_, _00059_);
  nor _23123_ (_00131_, _00129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _23124_ (_00132_, _00129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _23125_ (_00133_, _00132_, _00131_);
  and _23126_ (_00134_, _00133_, _00062_);
  and _23127_ (_00135_, _00079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _23128_ (_00137_, _00079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _23129_ (_00139_, _00137_, _00083_);
  nor _23130_ (_00141_, _00139_, _00135_);
  and _23131_ (_00142_, _00045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _23132_ (_00143_, _00045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor _23133_ (_00144_, _00143_, _00142_);
  and _23134_ (_00145_, _00144_, _00051_);
  or _23135_ (_00146_, _00145_, _00141_);
  or _23136_ (_00147_, _00146_, _00134_);
  or _23137_ (_00149_, _00147_, _00027_);
  and _23138_ (_00150_, _00027_, _09598_);
  nor _23139_ (_00151_, _00150_, _00091_);
  and _23140_ (_00152_, _00151_, _00149_);
  and _23141_ (_00153_, _00091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _23142_ (_00154_, _00153_, _00152_);
  and _23143_ (_13788_, _00154_, _06989_);
  nand _23144_ (_00155_, _00091_, _10970_);
  or _23145_ (_00156_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _23146_ (_00157_, _00045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or _23147_ (_00158_, _00157_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor _23148_ (_00159_, _00051_, _00070_);
  or _23149_ (_00161_, _00159_, _00027_);
  and _23150_ (_00163_, _00161_, _00158_);
  and _23151_ (_00164_, _00051_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _23152_ (_00165_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and _23153_ (_00166_, _00165_, _00040_);
  and _23154_ (_00167_, _00166_, _00067_);
  and _23155_ (_00168_, _00167_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _23156_ (_00169_, _00168_, _00060_);
  and _23157_ (_00170_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or _23158_ (_00171_, _00170_, _00164_);
  or _23159_ (_00172_, _00171_, _00163_);
  and _23160_ (_00173_, _00172_, _00156_);
  or _23161_ (_00174_, _00173_, _00091_);
  and _23162_ (_00175_, _00174_, _06989_);
  and _23163_ (_13798_, _00175_, _00155_);
  and _23164_ (_00176_, _00052_, _00045_);
  nand _23165_ (_00177_, _00176_, _00097_);
  and _23166_ (_00178_, _00177_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  not _23167_ (_00180_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _23168_ (_00182_, _00176_, _00180_);
  and _23169_ (_00183_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor _23170_ (_00184_, _00183_, _00182_);
  nor _23171_ (_00185_, _00184_, _00027_);
  or _23172_ (_00186_, _00185_, _00178_);
  and _23173_ (_00187_, _00186_, _00092_);
  nor _23174_ (_00189_, _00092_, _07118_);
  or _23175_ (_00190_, _00189_, _00187_);
  and _23176_ (_13802_, _00190_, _06989_);
  nand _23177_ (_00191_, _00027_, _11529_);
  and _23178_ (_00192_, _00071_, _00030_);
  or _23179_ (_00193_, _00192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _23180_ (_00194_, _00168_, _00032_);
  and _23181_ (_00195_, _00194_, _00061_);
  and _23182_ (_00196_, _00195_, _00193_);
  not _23183_ (_00197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and _23184_ (_00198_, _00067_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and _23185_ (_00199_, _00040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _23186_ (_00200_, _00199_, _00198_);
  and _23187_ (_00201_, _00200_, _00197_);
  nor _23188_ (_00202_, _00200_, _00197_);
  or _23189_ (_00203_, _00202_, _00201_);
  and _23190_ (_00204_, _00203_, _00051_);
  and _23191_ (_00205_, _00079_, _00030_);
  and _23192_ (_00206_, _00205_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nor _23193_ (_00207_, _00206_, _00197_);
  and _23194_ (_00208_, _00206_, _00197_);
  or _23195_ (_00209_, _00208_, _00207_);
  and _23196_ (_00210_, _00209_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _23197_ (_00211_, _00210_, _00204_);
  or _23198_ (_00212_, _00211_, _00196_);
  nor _23199_ (_00214_, _00212_, _00027_);
  nor _23200_ (_00215_, _00214_, _00091_);
  and _23201_ (_00216_, _00215_, _00191_);
  and _23202_ (_00217_, _00091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or _23203_ (_00218_, _00217_, _00216_);
  and _23204_ (_13809_, _00218_, _06989_);
  nand _23205_ (_00220_, _00027_, _07260_);
  or _23206_ (_00221_, _00046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _23207_ (_00223_, _00221_, _00051_);
  nor _23208_ (_00224_, _00223_, _00047_);
  or _23209_ (_00225_, _00072_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not _23210_ (_00226_, _00073_);
  and _23211_ (_00227_, _00226_, _00061_);
  and _23212_ (_00229_, _00227_, _00225_);
  or _23213_ (_00231_, _00109_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and _23214_ (_00232_, _00231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand _23215_ (_00233_, _00081_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _23216_ (_00234_, _00233_, _00232_);
  or _23217_ (_00235_, _00234_, _00229_);
  or _23218_ (_00236_, _00235_, _00224_);
  nor _23219_ (_00237_, _00236_, _00027_);
  nor _23220_ (_00238_, _00237_, _00091_);
  and _23221_ (_00239_, _00238_, _00220_);
  and _23222_ (_00240_, _00091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _23223_ (_00241_, _00240_, _00239_);
  and _23224_ (_13812_, _00241_, _06989_);
  nand _23225_ (_00242_, _00027_, _07317_);
  nand _23226_ (_00243_, _00045_, _00030_);
  nor _23227_ (_00244_, _00243_, _00197_);
  or _23228_ (_00245_, _00244_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand _23229_ (_00246_, _00244_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _23230_ (_00247_, _00051_, _00246_);
  and _23231_ (_00248_, _00247_, _00245_);
  and _23232_ (_00249_, _00079_, _00032_);
  or _23233_ (_00251_, _00249_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _23234_ (_00253_, _00080_);
  and _23235_ (_00255_, _00083_, _00253_);
  and _23236_ (_00257_, _00255_, _00251_);
  and _23237_ (_00259_, _00129_, _00032_);
  or _23238_ (_00260_, _00259_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _23239_ (_00262_, _00072_);
  or _23240_ (_00263_, _00262_, _00060_);
  and _23241_ (_00264_, _00263_, _00062_);
  and _23242_ (_00265_, _00264_, _00260_);
  or _23243_ (_00266_, _00265_, _00257_);
  or _23244_ (_00267_, _00266_, _00248_);
  or _23245_ (_00268_, _00267_, _00027_);
  and _23246_ (_00269_, _00268_, _00242_);
  or _23247_ (_00270_, _00269_, _00091_);
  or _23248_ (_00271_, _00092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and _23249_ (_00273_, _00271_, _06989_);
  and _23250_ (_13815_, _00273_, _00270_);
  or _23251_ (_00274_, _00132_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not _23252_ (_00276_, _00192_);
  or _23253_ (_00277_, _00276_, _00060_);
  and _23254_ (_00278_, _00277_, _00062_);
  and _23255_ (_00279_, _00278_, _00274_);
  or _23256_ (_00280_, _00135_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not _23257_ (_00281_, _00205_);
  and _23258_ (_00282_, _00083_, _00281_);
  and _23259_ (_00283_, _00282_, _00280_);
  or _23260_ (_00284_, _00142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _23261_ (_00285_, _00051_, _00243_);
  and _23262_ (_00286_, _00285_, _00284_);
  or _23263_ (_00287_, _00286_, _00283_);
  or _23264_ (_00288_, _00287_, _00279_);
  or _23265_ (_00290_, _00288_, _00027_);
  nand _23266_ (_00291_, _00027_, _09008_);
  and _23267_ (_00292_, _00291_, _00290_);
  or _23268_ (_00293_, _00292_, _00091_);
  or _23269_ (_00294_, _00092_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and _23270_ (_00295_, _00294_, _06989_);
  and _23271_ (_13817_, _00295_, _00293_);
  and _23272_ (_00296_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and _23273_ (_00297_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or _23274_ (_00298_, _00297_, _00296_);
  and _23275_ (_13822_, _00298_, _06989_);
  and _23276_ (_00299_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and _23277_ (_00300_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or _23278_ (_00301_, _00300_, _00299_);
  and _23279_ (_13872_, _00301_, _06989_);
  nand _23280_ (_00302_, _00044_, _00097_);
  and _23281_ (_00303_, _00302_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nand _23282_ (_00304_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not _23283_ (_00305_, _00043_);
  or _23284_ (_00306_, _00305_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and _23285_ (_00307_, _00306_, _00304_);
  nor _23286_ (_00308_, _00307_, _00027_);
  or _23287_ (_00309_, _00308_, _00303_);
  and _23288_ (_00311_, _00309_, _00092_);
  nor _23289_ (_00312_, _00092_, _07317_);
  or _23290_ (_00313_, _00312_, _00311_);
  and _23291_ (_13907_, _00313_, _06989_);
  or _23292_ (_00314_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _23293_ (_00315_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or _23294_ (_00316_, _00044_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nand _23295_ (_00317_, _00045_, _00097_);
  and _23296_ (_00319_, _00317_, _00316_);
  or _23297_ (_00320_, _00319_, _00315_);
  and _23298_ (_00322_, _00320_, _00314_);
  or _23299_ (_00323_, _00322_, _00091_);
  nand _23300_ (_00324_, _00091_, _07260_);
  and _23301_ (_00326_, _00324_, _06989_);
  and _23302_ (_13908_, _00326_, _00323_);
  or _23303_ (_00328_, _00305_, _00027_);
  and _23304_ (_00329_, _00328_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nand _23305_ (_00330_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand _23306_ (_00331_, _00305_, _00042_);
  and _23307_ (_00332_, _00331_, _00330_);
  nor _23308_ (_00333_, _00332_, _00027_);
  or _23309_ (_00335_, _00333_, _00329_);
  and _23310_ (_00336_, _00335_, _00092_);
  nor _23311_ (_00337_, _00092_, _11529_);
  or _23312_ (_00338_, _00337_, _00336_);
  and _23313_ (_13910_, _00338_, _06989_);
  or _23314_ (_00339_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _23315_ (_00340_, _00339_, _06989_);
  nand _23316_ (_00341_, _00005_, _10970_);
  and _23317_ (_13914_, _00341_, _00340_);
  or _23318_ (_00342_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23319_ (_00343_, _00342_, _06989_);
  nand _23320_ (_00344_, _00005_, _07118_);
  and _23321_ (_13919_, _00344_, _00343_);
  and _23322_ (_00346_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and _23323_ (_00347_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  or _23324_ (_00349_, _00347_, _00346_);
  and _23325_ (_13954_, _00349_, _06989_);
  or _23326_ (_00350_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _23327_ (_00351_, _00040_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor _23328_ (_00352_, _00351_, _00041_);
  and _23329_ (_00353_, _00071_, _00060_);
  and _23330_ (_00354_, _00353_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or _23331_ (_00355_, _00354_, _00352_);
  or _23332_ (_00356_, _00355_, _00027_);
  and _23333_ (_00357_, _00356_, _00350_);
  or _23334_ (_00358_, _00357_, _00091_);
  nand _23335_ (_00359_, _00091_, _09598_);
  and _23336_ (_00360_, _00359_, _06989_);
  and _23337_ (_14006_, _00360_, _00358_);
  nor _23338_ (_00361_, _00041_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor _23339_ (_00362_, _00361_, _00042_);
  and _23340_ (_00363_, _00169_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor _23341_ (_00364_, _00363_, _00362_);
  nor _23342_ (_00365_, _00364_, _00027_);
  and _23343_ (_00366_, _00027_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or _23344_ (_00367_, _00366_, _00365_);
  and _23345_ (_00368_, _00367_, _00092_);
  and _23346_ (_00369_, _00091_, _09009_);
  or _23347_ (_00370_, _00369_, _00368_);
  and _23348_ (_14009_, _00370_, _06989_);
  nand _23349_ (_00371_, _10146_, _07040_);
  or _23350_ (_00372_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and _23351_ (_00373_, _00372_, _06989_);
  and _23352_ (_14014_, _00373_, _00371_);
  and _23353_ (_00374_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and _23354_ (_00375_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or _23355_ (_00376_, _00375_, _00374_);
  and _23356_ (_14019_, _00376_, _06989_);
  nor _23357_ (_00377_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and _23358_ (_14022_, _00377_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and _23359_ (_00378_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and _23360_ (_00379_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or _23361_ (_00380_, _00379_, _00378_);
  and _23362_ (_14024_, _00380_, _06989_);
  and _23363_ (_00381_, _07454_, _07049_);
  not _23364_ (_00382_, _00381_);
  nor _23365_ (_00383_, _00382_, _10970_);
  nor _23366_ (_00384_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not _23367_ (_00385_, _00384_);
  and _23368_ (_00386_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _23369_ (_00388_, _00386_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not _23370_ (_00389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _23371_ (_00390_, _00389_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  not _23372_ (_00391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _23373_ (_00392_, _00391_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not _23374_ (_00393_, t1_i);
  and _23375_ (_00394_, _00393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and _23376_ (_00395_, _00394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or _23377_ (_00396_, _00395_, _00392_);
  and _23378_ (_00397_, _00396_, _00390_);
  and _23379_ (_00398_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23380_ (_00399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _23381_ (_00400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and _23382_ (_00401_, _00400_, _00399_);
  and _23383_ (_00402_, _00401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _23384_ (_00403_, _00402_, _00398_);
  and _23385_ (_00404_, _00403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23386_ (_00405_, _00404_, _00397_);
  and _23387_ (_00406_, _00405_, _00388_);
  and _23388_ (_00407_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _23389_ (_00408_, _00407_, _00385_);
  not _23390_ (_00409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23391_ (_00410_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _00409_);
  not _23392_ (_00411_, _00410_);
  and _23393_ (_00412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _23394_ (_00413_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _23395_ (_00414_, _00413_, _00412_);
  and _23396_ (_00415_, _00414_, _00401_);
  and _23397_ (_00416_, _00415_, _00398_);
  and _23398_ (_00417_, _00416_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23399_ (_00418_, _00417_, _00397_);
  and _23400_ (_00419_, _00418_, _00388_);
  and _23401_ (_00420_, _00419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor _23402_ (_00421_, _00420_, _00411_);
  or _23403_ (_00422_, _00421_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _23404_ (_00423_, _00412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and _23405_ (_00424_, _00421_, _00423_);
  or _23406_ (_00425_, _00424_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _23407_ (_00426_, _00425_, _00422_);
  or _23408_ (_00427_, _00426_, _00408_);
  or _23409_ (_00428_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _23410_ (_00429_, _09560_, _07454_);
  nor _23411_ (_00430_, _00429_, _00381_);
  and _23412_ (_00431_, _00430_, _00428_);
  and _23413_ (_00432_, _00431_, _00427_);
  and _23414_ (_00433_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _23415_ (_00434_, _00433_, _00432_);
  or _23416_ (_00435_, _00434_, _00383_);
  and _23417_ (_14059_, _00435_, _06989_);
  nor _23418_ (_00436_, _00382_, _07118_);
  not _23419_ (_00437_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _23420_ (_00438_, _00402_, _00397_);
  and _23421_ (_00439_, _00423_, _00438_);
  and _23422_ (_00440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _23423_ (_00441_, _00440_, _00398_);
  and _23424_ (_00443_, _00441_, _00410_);
  and _23425_ (_00444_, _00443_, _00439_);
  and _23426_ (_00446_, _00403_, _00397_);
  and _23427_ (_00447_, _00440_, _00446_);
  and _23428_ (_00448_, _00447_, _00384_);
  nor _23429_ (_00449_, _00448_, _00444_);
  or _23430_ (_00450_, _00449_, _00437_);
  nor _23431_ (_00451_, _00450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and _23432_ (_00452_, _00450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _23433_ (_00454_, _00452_, _00451_);
  and _23434_ (_00455_, _00454_, _00430_);
  and _23435_ (_00456_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or _23436_ (_00458_, _00456_, _00455_);
  or _23437_ (_00459_, _00458_, _00436_);
  and _23438_ (_14064_, _00459_, _06989_);
  nor _23439_ (_00460_, _00382_, _07317_);
  and _23440_ (_00461_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _23441_ (_00462_, _00418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _23442_ (_00463_, _00418_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and _23443_ (_00464_, _00463_, _00462_);
  and _23444_ (_00466_, _00464_, _00410_);
  not _23445_ (_00467_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23446_ (_00468_, _00384_, _00467_);
  nor _23447_ (_00469_, _00446_, _00385_);
  or _23448_ (_00470_, _00469_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or _23449_ (_00471_, _00470_, _00468_);
  and _23450_ (_00472_, _00471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nand _23451_ (_00473_, _00405_, _00384_);
  nor _23452_ (_00474_, _00473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or _23453_ (_00475_, _00474_, _00472_);
  or _23454_ (_00476_, _00475_, _00466_);
  and _23455_ (_00477_, _00476_, _00430_);
  or _23456_ (_00478_, _00477_, _00461_);
  or _23457_ (_00479_, _00478_, _00460_);
  and _23458_ (_14072_, _00479_, _06989_);
  nor _23459_ (_00480_, _00382_, _07260_);
  nand _23460_ (_00481_, _00449_, _00437_);
  and _23461_ (_00482_, _00481_, _00450_);
  and _23462_ (_00483_, _00482_, _00430_);
  and _23463_ (_00484_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or _23464_ (_00485_, _00484_, _00483_);
  or _23465_ (_00486_, _00485_, _00480_);
  and _23466_ (_14075_, _00486_, _06989_);
  not _23467_ (_00487_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and _23468_ (_00488_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and _23469_ (_00489_, _00488_, _00487_);
  and _23470_ (_00490_, _00489_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor _23471_ (_00491_, _00488_, _00487_);
  or _23472_ (_00492_, _00491_, _00489_);
  nand _23473_ (_00493_, _00492_, _06989_);
  nor _23474_ (_14082_, _00493_, _00490_);
  and _23475_ (_00495_, _09529_, _07454_);
  and _23476_ (_00496_, _00495_, _06983_);
  and _23477_ (_00497_, _00438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _23478_ (_00498_, _00497_, _00423_);
  nand _23479_ (_00499_, _00498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _23480_ (_00500_, _00498_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23481_ (_00501_, _00500_, _00410_);
  and _23482_ (_00503_, _00501_, _00499_);
  and _23483_ (_00504_, _00497_, _00469_);
  or _23484_ (_00505_, _00504_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and _23485_ (_00506_, _00505_, _00470_);
  nor _23486_ (_00507_, _00506_, _00503_);
  or _23487_ (_00508_, _00507_, _00381_);
  or _23488_ (_00509_, _00382_, _09008_);
  and _23489_ (_00510_, _00509_, _00508_);
  nor _23490_ (_00511_, _00510_, _00496_);
  and _23491_ (_00512_, _00496_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or _23492_ (_00513_, _00512_, _00511_);
  and _23493_ (_14085_, _00513_, _06989_);
  or _23494_ (_00514_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor _23495_ (_00515_, _00488_, rst);
  and _23496_ (_14087_, _00515_, _00514_);
  nor _23497_ (_00516_, _00382_, _11529_);
  nor _23498_ (_00517_, _00418_, _00411_);
  or _23499_ (_00518_, _00517_, _00471_);
  and _23500_ (_00519_, _00518_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and _23501_ (_00520_, _00410_, _00467_);
  and _23502_ (_00521_, _00520_, _00423_);
  or _23503_ (_00522_, _00521_, _00468_);
  and _23504_ (_00523_, _00522_, _00446_);
  or _23505_ (_00524_, _00523_, _00519_);
  and _23506_ (_00525_, _00524_, _00430_);
  and _23507_ (_00526_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or _23508_ (_00527_, _00526_, _00525_);
  or _23509_ (_00528_, _00527_, _00516_);
  and _23510_ (_14090_, _00528_, _06989_);
  and _23511_ (_00530_, _09530_, _07454_);
  nand _23512_ (_00531_, _00530_, _07118_);
  and _23513_ (_00532_, _00438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  not _23514_ (_00533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and _23515_ (_00534_, _00533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _23516_ (_00535_, _00534_, _00410_);
  nor _23517_ (_00536_, _00438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _23518_ (_00537_, _00536_, _00535_);
  nor _23519_ (_00538_, _00537_, _00532_);
  and _23520_ (_00539_, _00534_, _00439_);
  and _23521_ (_00540_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor _23522_ (_00541_, _00540_, _00538_);
  nor _23523_ (_00542_, _00541_, _00381_);
  nor _23524_ (_00543_, _00535_, _00381_);
  not _23525_ (_00544_, _00543_);
  and _23526_ (_00545_, _00544_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  or _23527_ (_00546_, _00545_, _00542_);
  or _23528_ (_00547_, _00546_, _00530_);
  and _23529_ (_00548_, _00547_, _06989_);
  and _23530_ (_14105_, _00548_, _00531_);
  and _23531_ (_00549_, _00532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor _23532_ (_00550_, _00532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or _23533_ (_00551_, _00550_, _00549_);
  nand _23534_ (_00552_, _00551_, _00543_);
  or _23535_ (_00553_, _00543_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and _23536_ (_00554_, _00553_, _00552_);
  and _23537_ (_00555_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or _23538_ (_00556_, _00555_, _00429_);
  and _23539_ (_00557_, _00556_, _00382_);
  or _23540_ (_00558_, _00557_, _00554_);
  and _23541_ (_00559_, _00558_, _06989_);
  nand _23542_ (_00560_, _00530_, _10970_);
  and _23543_ (_14108_, _00560_, _00559_);
  nand _23544_ (_00561_, _00530_, _07260_);
  and _23545_ (_00562_, _00397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _23546_ (_00563_, _00562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and _23547_ (_00564_, _00563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and _23548_ (_00565_, _00564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _23549_ (_00566_, _00565_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _23550_ (_00567_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor _23551_ (_00568_, _00567_, _00438_);
  and _23552_ (_00569_, _00568_, _00566_);
  and _23553_ (_00571_, _00534_, _00397_);
  and _23554_ (_00572_, _00571_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and _23555_ (_00573_, _00572_, _00415_);
  nor _23556_ (_00574_, _00573_, _00569_);
  nor _23557_ (_00576_, _00574_, _00381_);
  or _23558_ (_00577_, _00567_, _00381_);
  and _23559_ (_00578_, _00577_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  or _23560_ (_00579_, _00578_, _00576_);
  or _23561_ (_00580_, _00579_, _00530_);
  and _23562_ (_00581_, _00580_, _06989_);
  and _23563_ (_14111_, _00581_, _00561_);
  and _23564_ (_00582_, _00577_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or _23565_ (_00583_, _00563_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  nor _23566_ (_00584_, _00564_, _00567_);
  and _23567_ (_00585_, _00584_, _00583_);
  and _23568_ (_00586_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor _23569_ (_00587_, _00586_, _00585_);
  nor _23570_ (_00589_, _00587_, _00381_);
  or _23571_ (_00590_, _00589_, _00582_);
  or _23572_ (_00591_, _00590_, _00530_);
  nand _23573_ (_00592_, _00530_, _11529_);
  and _23574_ (_00593_, _00592_, _06989_);
  and _23575_ (_14115_, _00593_, _00591_);
  not _23576_ (_00594_, _00496_);
  and _23577_ (_00595_, _00577_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or _23578_ (_00597_, _00564_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor _23579_ (_00598_, _00565_, _00567_);
  and _23580_ (_00599_, _00598_, _00597_);
  and _23581_ (_00600_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor _23582_ (_00601_, _00600_, _00599_);
  nor _23583_ (_00602_, _00601_, _00381_);
  or _23584_ (_00603_, _00602_, _00595_);
  and _23585_ (_00604_, _00603_, _00594_);
  nor _23586_ (_00605_, _00594_, _07317_);
  or _23587_ (_00606_, _00605_, _00604_);
  and _23588_ (_14118_, _00606_, _06989_);
  and _23589_ (_00607_, _00577_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or _23590_ (_00608_, _00562_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  nor _23591_ (_00609_, _00563_, _00567_);
  and _23592_ (_00610_, _00609_, _00608_);
  and _23593_ (_00611_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor _23594_ (_00612_, _00611_, _00610_);
  nor _23595_ (_00613_, _00612_, _00381_);
  or _23596_ (_00614_, _00613_, _00530_);
  or _23597_ (_00615_, _00614_, _00607_);
  nand _23598_ (_00616_, _00530_, _09008_);
  and _23599_ (_00617_, _00616_, _06989_);
  and _23600_ (_14121_, _00617_, _00615_);
  and _23601_ (_00618_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not _23602_ (_00619_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _23603_ (_00620_, _08139_, _00619_);
  or _23604_ (_00621_, _00620_, _00618_);
  and _23605_ (_14123_, _00621_, _06989_);
  or _23606_ (_00622_, _00439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _23607_ (_00623_, _00498_, _00411_);
  and _23608_ (_00624_, _00623_, _00622_);
  or _23609_ (_00625_, _00438_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _23610_ (_00626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor _23611_ (_00627_, _00497_, _00385_);
  or _23612_ (_00628_, _00627_, _00626_);
  and _23613_ (_00629_, _00628_, _00625_);
  nor _23614_ (_00630_, _00629_, _00624_);
  and _23615_ (_00631_, _00630_, _00430_);
  nand _23616_ (_00632_, _00381_, _09598_);
  not _23617_ (_00633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nand _23618_ (_00634_, _00530_, _00633_);
  and _23619_ (_00635_, _00634_, _06989_);
  nand _23620_ (_00636_, _00635_, _00632_);
  nor _23621_ (_14127_, _00636_, _00631_);
  and _23622_ (_00637_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or _23623_ (_14139_, _00637_, _09441_);
  nor _23624_ (_14216_, _11613_, rst);
  and _23625_ (_00640_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _23626_ (_00641_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _23627_ (_00642_, _00641_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _23628_ (_00643_, _00641_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor _23629_ (_00644_, _00643_, _00642_);
  or _23630_ (_00645_, _00644_, _00640_);
  and _23631_ (_14225_, _00645_, _06989_);
  not _23632_ (_00646_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  nor _23633_ (_00648_, _00640_, _00646_);
  nor _23634_ (_00649_, _00648_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and _23635_ (_00650_, _00648_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or _23636_ (_00651_, _00650_, _00649_);
  nor _23637_ (_14227_, _00651_, rst);
  and _23638_ (_00652_, _00640_, _00646_);
  nor _23639_ (_00653_, _00652_, _00648_);
  and _23640_ (_14255_, _00653_, _06989_);
  and _23641_ (_00654_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not _23642_ (_00655_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _23643_ (_00656_, _08139_, _00655_);
  or _23644_ (_00657_, _00656_, _00654_);
  and _23645_ (_14264_, _00657_, _06989_);
  or _23646_ (_00658_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not _23647_ (_00659_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _23648_ (_00660_, _08139_, _00659_);
  and _23649_ (_00661_, _00660_, _06989_);
  and _23650_ (_14403_, _00661_, _00658_);
  not _23651_ (_00662_, _00567_);
  and _23652_ (_00664_, _00662_, _00397_);
  nand _23653_ (_00665_, _00664_, _00382_);
  and _23654_ (_00666_, _00665_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  not _23655_ (_00668_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and _23656_ (_00669_, _00664_, _00668_);
  and _23657_ (_00670_, _00534_, _00498_);
  nor _23658_ (_00671_, _00670_, _00669_);
  nor _23659_ (_00672_, _00671_, _00381_);
  or _23660_ (_00673_, _00672_, _00666_);
  or _23661_ (_00674_, _00673_, _00530_);
  nand _23662_ (_00675_, _00530_, _09598_);
  and _23663_ (_00676_, _00675_, _06989_);
  and _23664_ (_14456_, _00676_, _00674_);
  nand _23665_ (_00677_, _10146_, _09008_);
  or _23666_ (_00678_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and _23667_ (_00680_, _00678_, _06989_);
  and _23668_ (_14572_, _00680_, _00677_);
  and _23669_ (_00682_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not _23670_ (_00683_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _23671_ (_00684_, _08139_, _00683_);
  or _23672_ (_00685_, _00684_, _00682_);
  and _23673_ (_14583_, _00685_, _06989_);
  or _23674_ (_00686_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not _23675_ (_00687_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _23676_ (_00688_, _08139_, _00687_);
  and _23677_ (_00689_, _00688_, _06989_);
  and _23678_ (_14585_, _00689_, _00686_);
  and _23679_ (_00690_, _08036_, _07084_);
  and _23680_ (_00691_, _00690_, _14026_);
  and _23681_ (_00692_, _00691_, _06539_);
  nand _23682_ (_00693_, _00692_, _06968_);
  or _23683_ (_00694_, _00692_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _23684_ (_00695_, _00694_, _06485_);
  and _23685_ (_00696_, _00695_, _00693_);
  and _23686_ (_00697_, _13950_, _07125_);
  nand _23687_ (_00698_, _00697_, _07040_);
  or _23688_ (_00699_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and _23689_ (_00700_, _00699_, _06983_);
  and _23690_ (_00701_, _00700_, _00698_);
  not _23691_ (_00702_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  nor _23692_ (_00703_, _06484_, _00702_);
  or _23693_ (_00704_, _00703_, rst);
  or _23694_ (_00706_, _00704_, _00701_);
  or _23695_ (_14607_, _00706_, _00696_);
  and _23696_ (_00707_, _09022_, _06500_);
  and _23697_ (_00708_, _00707_, _14025_);
  and _23698_ (_00709_, _00708_, _14196_);
  nand _23699_ (_00710_, _00709_, _06968_);
  or _23700_ (_00711_, _00709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nor _23701_ (_00712_, _06477_, _06434_);
  and _23702_ (_00713_, _00712_, _07453_);
  and _23703_ (_00714_, _00713_, _14011_);
  not _23704_ (_00715_, _00714_);
  and _23705_ (_00716_, _00715_, _00711_);
  and _23706_ (_00717_, _00716_, _00710_);
  nor _23707_ (_00718_, _00715_, _10970_);
  or _23708_ (_00719_, _00718_, _00717_);
  and _23709_ (_00009_, _00719_, _06989_);
  and _23710_ (_00720_, _08037_, _14026_);
  and _23711_ (_00721_, _00720_, _06539_);
  nand _23712_ (_00722_, _00721_, _06968_);
  or _23713_ (_00723_, _00721_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _23714_ (_00724_, _00723_, _06485_);
  and _23715_ (_00725_, _00724_, _00722_);
  and _23716_ (_00726_, _07454_, _07125_);
  nand _23717_ (_00727_, _00726_, _07040_);
  or _23718_ (_00728_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and _23719_ (_00729_, _00728_, _06983_);
  and _23720_ (_00730_, _00729_, _00727_);
  not _23721_ (_00731_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  nor _23722_ (_00732_, _06484_, _00731_);
  or _23723_ (_00733_, _00732_, rst);
  or _23724_ (_00734_, _00733_, _00730_);
  or _23725_ (_00018_, _00734_, _00725_);
  and _23726_ (_00735_, _00708_, _07048_);
  nand _23727_ (_00736_, _00735_, _06968_);
  or _23728_ (_00737_, _00735_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _23729_ (_00738_, _00737_, _00715_);
  and _23730_ (_00739_, _00738_, _00736_);
  nor _23731_ (_00740_, _00715_, _07118_);
  or _23732_ (_00741_, _00740_, _00739_);
  and _23733_ (_00024_, _00741_, _06989_);
  and _23734_ (_00742_, _00708_, _07044_);
  nand _23735_ (_00743_, _00742_, _06968_);
  or _23736_ (_00744_, _00742_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _23737_ (_00745_, _00744_, _00715_);
  and _23738_ (_00746_, _00745_, _00743_);
  nor _23739_ (_00747_, _00715_, _07260_);
  or _23740_ (_00748_, _00747_, _00746_);
  and _23741_ (_00026_, _00748_, _06989_);
  or _23742_ (_00749_, _08435_, _07043_);
  nor _23743_ (_00750_, _00749_, _07217_);
  or _23744_ (_00751_, _00750_, _08437_);
  and _23745_ (_00752_, _00751_, _00708_);
  nand _23746_ (_00753_, _00708_, _06525_);
  and _23747_ (_00754_, _00753_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _23748_ (_00755_, _00754_, _00714_);
  or _23749_ (_00756_, _00755_, _00752_);
  nand _23750_ (_00757_, _00714_, _07317_);
  and _23751_ (_00758_, _00757_, _06989_);
  and _23752_ (_00028_, _00758_, _00756_);
  not _23753_ (_00759_, _09074_);
  nor _23754_ (_00760_, _06968_, _00759_);
  and _23755_ (_00761_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _23756_ (_00762_, _00761_, _00760_);
  and _23757_ (_00763_, _00762_, _00708_);
  not _23758_ (_00764_, _00749_);
  nand _23759_ (_00765_, _00708_, _00764_);
  and _23760_ (_00766_, _00765_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or _23761_ (_00767_, _00766_, _00714_);
  or _23762_ (_00768_, _00767_, _00763_);
  nand _23763_ (_00769_, _00714_, _11529_);
  and _23764_ (_00770_, _00769_, _06989_);
  and _23765_ (_00031_, _00770_, _00768_);
  and _23766_ (_00771_, _00708_, _07089_);
  or _23767_ (_00772_, _00771_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and _23768_ (_00773_, _00772_, _00715_);
  nand _23769_ (_00774_, _00771_, _06968_);
  and _23770_ (_00775_, _00774_, _00773_);
  nor _23771_ (_00776_, _00715_, _09008_);
  or _23772_ (_00777_, _00776_, _00775_);
  and _23773_ (_00048_, _00777_, _06989_);
  and _23774_ (_00778_, _00708_, _06979_);
  or _23775_ (_00779_, _00778_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _23776_ (_00780_, _00779_, _00715_);
  nand _23777_ (_00781_, _00778_, _06968_);
  and _23778_ (_00782_, _00781_, _00780_);
  and _23779_ (_00783_, _00714_, _09599_);
  or _23780_ (_00784_, _00783_, _00782_);
  and _23781_ (_00050_, _00784_, _06989_);
  or _23782_ (_00785_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  nand _23783_ (_00786_, _07493_, _07495_);
  and _23784_ (_00787_, _00786_, _06989_);
  and _23785_ (_00055_, _00787_, _00785_);
  not _23786_ (_00788_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nor _23787_ (_00789_, _00749_, _00788_);
  or _23788_ (_00790_, _00789_, _08437_);
  and _23789_ (_00791_, _00707_, _06449_);
  and _23790_ (_00792_, _00791_, _00790_);
  and _23791_ (_00793_, _09029_, _06986_);
  and _23792_ (_00795_, _00791_, _06525_);
  nor _23793_ (_00796_, _00795_, _00788_);
  or _23794_ (_00797_, _00796_, _00793_);
  or _23795_ (_00798_, _00797_, _00792_);
  nand _23796_ (_00799_, _00793_, _07317_);
  and _23797_ (_00800_, _00799_, _06989_);
  and _23798_ (_00111_, _00800_, _00798_);
  and _23799_ (_00801_, _00791_, _14196_);
  nand _23800_ (_00802_, _00801_, _06968_);
  not _23801_ (_00803_, _00793_);
  or _23802_ (_00804_, _00801_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and _23803_ (_00805_, _00804_, _00803_);
  and _23804_ (_00806_, _00805_, _00802_);
  nor _23805_ (_00807_, _00803_, _10970_);
  or _23806_ (_00808_, _00807_, _00806_);
  and _23807_ (_00113_, _00808_, _06989_);
  and _23808_ (_00809_, _00791_, _07048_);
  nand _23809_ (_00810_, _00809_, _06968_);
  or _23810_ (_00811_, _00809_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and _23811_ (_00812_, _00811_, _00803_);
  and _23812_ (_00813_, _00812_, _00810_);
  nor _23813_ (_00814_, _00803_, _07118_);
  or _23814_ (_00815_, _00814_, _00813_);
  and _23815_ (_00117_, _00815_, _06989_);
  and _23816_ (_00816_, _00791_, _08349_);
  nor _23817_ (_00817_, _06978_, _06525_);
  not _23818_ (_00818_, _00791_);
  or _23819_ (_00819_, _00818_, _00817_);
  or _23820_ (_00820_, _00819_, _00795_);
  and _23821_ (_00821_, _00820_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or _23822_ (_00822_, _00821_, _00793_);
  or _23823_ (_00823_, _00822_, _00816_);
  nand _23824_ (_00824_, _00793_, _07260_);
  and _23825_ (_00825_, _00824_, _06989_);
  and _23826_ (_00119_, _00825_, _00823_);
  and _23827_ (_00826_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _08578_);
  and _23828_ (_00827_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [2]);
  or _23829_ (_00828_, _00827_, _00826_);
  and _23830_ (_00121_, _00828_, _06989_);
  and _23831_ (_00829_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _23832_ (_00830_, _00829_, _00760_);
  and _23833_ (_00831_, _00830_, _00791_);
  nand _23834_ (_00832_, _00791_, _00764_);
  and _23835_ (_00833_, _00832_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or _23836_ (_00834_, _00833_, _00793_);
  or _23837_ (_00835_, _00834_, _00831_);
  nand _23838_ (_00836_, _00793_, _11529_);
  and _23839_ (_00837_, _00836_, _06989_);
  and _23840_ (_00123_, _00837_, _00835_);
  and _23841_ (_00838_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _08578_);
  and _23842_ (_00839_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _23843_ (_00840_, _00839_, _00838_);
  and _23844_ (_00128_, _00840_, _06989_);
  and _23845_ (_00841_, _08578_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and _23846_ (_00842_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [5]);
  or _23847_ (_00843_, _00842_, _00841_);
  and _23848_ (_00130_, _00843_, _06989_);
  and _23849_ (_00844_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _08578_);
  and _23850_ (_00845_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _23851_ (_00846_, _00845_, _00844_);
  and _23852_ (_00136_, _00846_, _06989_);
  and _23853_ (_00847_, _00791_, _07089_);
  or _23854_ (_00848_, _00847_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and _23855_ (_00849_, _00848_, _00803_);
  nand _23856_ (_00850_, _00847_, _06968_);
  and _23857_ (_00851_, _00850_, _00849_);
  nor _23858_ (_00852_, _00803_, _09008_);
  or _23859_ (_00853_, _00852_, _00851_);
  and _23860_ (_00138_, _00853_, _06989_);
  and _23861_ (_00854_, _00791_, _06979_);
  or _23862_ (_00855_, _00854_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and _23863_ (_00856_, _00855_, _00803_);
  nand _23864_ (_00857_, _00854_, _06968_);
  and _23865_ (_00858_, _00857_, _00856_);
  and _23866_ (_00859_, _00793_, _09599_);
  or _23867_ (_00860_, _00859_, _00858_);
  and _23868_ (_00140_, _00860_, _06989_);
  and _23869_ (_00861_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _08578_);
  and _23870_ (_00862_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _23871_ (_00863_, _00862_, _00861_);
  and _23872_ (_00148_, _00863_, _06989_);
  and _23873_ (_00864_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _08578_);
  and _23874_ (_00865_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _23875_ (_00866_, _00865_, _00864_);
  and _23876_ (_00160_, _00866_, _06989_);
  and _23877_ (_00867_, _14027_, _06449_);
  and _23878_ (_00868_, _00867_, _07044_);
  nand _23879_ (_00869_, _00868_, _06968_);
  or _23880_ (_00870_, _00868_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _23881_ (_00871_, _00870_, _07460_);
  and _23882_ (_00872_, _00871_, _00869_);
  nor _23883_ (_00873_, _07460_, _07260_);
  or _23884_ (_00874_, _00873_, _00872_);
  and _23885_ (_00162_, _00874_, _06989_);
  and _23886_ (_00875_, _00867_, _09074_);
  nand _23887_ (_00876_, _00875_, _06968_);
  or _23888_ (_00877_, _00875_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _23889_ (_00878_, _00877_, _07460_);
  and _23890_ (_00879_, _00878_, _00876_);
  nor _23891_ (_00880_, _11529_, _07460_);
  or _23892_ (_00881_, _00880_, _00879_);
  and _23893_ (_00179_, _00881_, _06989_);
  and _23894_ (_00882_, _00867_, _06979_);
  or _23895_ (_00883_, _00882_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _23896_ (_00884_, _00883_, _07460_);
  nand _23897_ (_00885_, _00882_, _06968_);
  and _23898_ (_00886_, _00885_, _00884_);
  and _23899_ (_00887_, _09599_, _07459_);
  or _23900_ (_00888_, _00887_, _00886_);
  and _23901_ (_00181_, _00888_, _06989_);
  and _23902_ (_00889_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or _23903_ (_00890_, _00889_, _09510_);
  and _23904_ (_00188_, _00890_, _06989_);
  nor _23905_ (_00891_, _14042_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or _23906_ (_00892_, _00891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand _23907_ (_00893_, _00891_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and _23908_ (_00894_, _00893_, _06989_);
  and _23909_ (_00213_, _00894_, _00892_);
  nor _23910_ (_00895_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _23911_ (_00896_, _00895_, _09393_);
  and _23912_ (_00897_, _00896_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not _23913_ (_00898_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor _23914_ (_00899_, _00896_, _00898_);
  or _23915_ (_00900_, _00899_, _00897_);
  or _23916_ (_00901_, _00900_, _14028_);
  or _23917_ (_00902_, _09074_, _00898_);
  nand _23918_ (_00903_, _00902_, _14028_);
  or _23919_ (_00904_, _00903_, _00760_);
  and _23920_ (_00905_, _00904_, _00901_);
  or _23921_ (_00906_, _00905_, _14031_);
  nand _23922_ (_00907_, _14031_, _11529_);
  and _23923_ (_00908_, _00907_, _06989_);
  and _23924_ (_00219_, _00908_, _00906_);
  nor _23925_ (_00909_, _07161_, _07166_);
  nand _23926_ (_00910_, _00909_, _07274_);
  and _23927_ (_00911_, _00909_, _07196_);
  or _23928_ (_00912_, _00911_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and _23929_ (_00913_, _00912_, _06989_);
  and _23930_ (_00222_, _00913_, _00910_);
  nand _23931_ (_00914_, _07277_, _07274_);
  and _23932_ (_00915_, _07277_, _07196_);
  or _23933_ (_00916_, _00915_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and _23934_ (_00917_, _00916_, _06989_);
  and _23935_ (_00228_, _00917_, _00914_);
  and _23936_ (_00918_, _13972_, _13943_);
  nor _23937_ (_00919_, _00918_, _13959_);
  and _23938_ (_00920_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _23939_ (_00921_, _00920_, _13953_);
  and _23940_ (_00922_, _13952_, _06989_);
  and _23941_ (_00923_, _00922_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or _23942_ (_00230_, _00923_, _00921_);
  nor _23943_ (_00924_, _11413_, rst);
  and _23944_ (_00250_, _00924_, _11964_);
  or _23945_ (_00925_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23946_ (_00926_, _00925_, _07202_);
  or _23947_ (_00927_, _00926_, _07208_);
  and _23948_ (_00928_, _07212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23949_ (_00929_, _00928_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23950_ (_00930_, _07215_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23951_ (_00931_, _00930_, _07218_);
  and _23952_ (_00932_, _00931_, _00929_);
  nand _23953_ (_00933_, _07474_, _07218_);
  nand _23954_ (_00934_, _00933_, _07207_);
  or _23955_ (_00935_, _00934_, _00932_);
  and _23956_ (_00936_, _00935_, _00927_);
  and _23957_ (_00937_, _07474_, _07201_);
  or _23958_ (_00938_, _00937_, _07222_);
  or _23959_ (_00939_, _00938_, _00936_);
  not _23960_ (_00940_, _07222_);
  or _23961_ (_00941_, _00940_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23962_ (_00942_, _00941_, _00939_);
  and _23963_ (_00943_, _00942_, _07197_);
  and _23964_ (_00944_, _00925_, _07187_);
  or _23965_ (_00945_, _00944_, _07194_);
  and _23966_ (_00946_, _07175_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _23967_ (_00947_, _00946_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23968_ (_00948_, _07179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor _23969_ (_00949_, _00948_, _07182_);
  and _23970_ (_00950_, _00949_, _00947_);
  nand _23971_ (_00951_, _07474_, _07182_);
  nand _23972_ (_00952_, _00951_, _07193_);
  or _23973_ (_00953_, _00952_, _00950_);
  and _23974_ (_00954_, _00953_, _00945_);
  and _23975_ (_00955_, _07474_, _07186_);
  or _23976_ (_00956_, _00955_, _00954_);
  and _23977_ (_00957_, _00956_, _07196_);
  or _23978_ (_00958_, _00957_, _07161_);
  or _23979_ (_00959_, _00958_, _00943_);
  or _23980_ (_00960_, _07164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and _23981_ (_00961_, _00960_, _06989_);
  and _23982_ (_00252_, _00961_, _00959_);
  not _23983_ (_00962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _23984_ (_00963_, _00928_, _00962_);
  nand _23985_ (_00964_, _00963_, _00931_);
  or _23986_ (_00965_, _07465_, _07219_);
  and _23987_ (_00966_, _00965_, _00964_);
  or _23988_ (_00967_, _00966_, _07206_);
  not _23989_ (_00968_, _07204_);
  not _23990_ (_00969_, _07206_);
  or _23991_ (_00970_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or _23992_ (_00971_, _00970_, _00969_);
  and _23993_ (_00972_, _00971_, _00968_);
  and _23994_ (_00973_, _00972_, _00967_);
  and _23995_ (_00974_, _07465_, _07204_);
  or _23996_ (_00975_, _00974_, _07201_);
  or _23997_ (_00976_, _00975_, _00973_);
  or _23998_ (_00977_, _00970_, _07202_);
  nand _23999_ (_00978_, _00977_, _00976_);
  nand _24000_ (_00979_, _00978_, _07274_);
  not _24001_ (_00980_, _07189_);
  or _24002_ (_00981_, _07465_, _00980_);
  or _24003_ (_00982_, _00946_, _00962_);
  nand _24004_ (_00983_, _00982_, _00949_);
  not _24005_ (_00984_, _07191_);
  or _24006_ (_00985_, _07465_, _07183_);
  and _24007_ (_00986_, _00985_, _00984_);
  and _24008_ (_00987_, _00986_, _00983_);
  and _24009_ (_00988_, _00970_, _07191_);
  or _24010_ (_00989_, _00988_, _07189_);
  or _24011_ (_00990_, _00989_, _00987_);
  and _24012_ (_00991_, _00990_, _00981_);
  or _24013_ (_00992_, _00991_, _07186_);
  or _24014_ (_00993_, _00970_, _07187_);
  and _24015_ (_00994_, _00993_, _00992_);
  or _24016_ (_00995_, _00994_, _07197_);
  and _24017_ (_00996_, _00995_, _00979_);
  or _24018_ (_00997_, _00996_, _07161_);
  nor _24019_ (_00998_, _07223_, _07161_);
  or _24020_ (_00999_, _00998_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and _24021_ (_01001_, _00999_, _06989_);
  and _24022_ (_00254_, _01001_, _00997_);
  or _24023_ (_01002_, _00642_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and _24024_ (_00256_, _01002_, _06989_);
  nor _24025_ (_00258_, _12740_, rst);
  nand _24026_ (_01003_, _11351_, _06989_);
  nor _24027_ (_00261_, _01003_, _11417_);
  or _24028_ (_01004_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _24029_ (_01005_, _01004_, _07202_);
  or _24030_ (_01006_, _01005_, _07208_);
  and _24031_ (_01007_, _07212_, _07166_);
  or _24032_ (_01008_, _01007_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _24033_ (_01009_, _07215_, _07166_);
  nor _24034_ (_01010_, _01009_, _07218_);
  and _24035_ (_01011_, _01010_, _01008_);
  nand _24036_ (_01012_, _07473_, _07218_);
  nand _24037_ (_01013_, _01012_, _07207_);
  or _24038_ (_01014_, _01013_, _01011_);
  and _24039_ (_01015_, _01014_, _01006_);
  and _24040_ (_01016_, _07473_, _07201_);
  or _24041_ (_01017_, _01016_, _07222_);
  or _24042_ (_01018_, _01017_, _01015_);
  or _24043_ (_01019_, _00940_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _24044_ (_01020_, _01019_, _01018_);
  and _24045_ (_01021_, _01020_, _07197_);
  and _24046_ (_01022_, _01004_, _07187_);
  or _24047_ (_01024_, _01022_, _07194_);
  and _24048_ (_01025_, _07175_, _07166_);
  or _24049_ (_01026_, _01025_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _24050_ (_01027_, _07179_, _07166_);
  nor _24051_ (_01028_, _01027_, _07182_);
  and _24052_ (_01029_, _01028_, _01026_);
  nand _24053_ (_01030_, _07473_, _07182_);
  nand _24054_ (_01031_, _01030_, _07193_);
  or _24055_ (_01032_, _01031_, _01029_);
  and _24056_ (_01033_, _01032_, _01024_);
  and _24057_ (_01034_, _07473_, _07186_);
  or _24058_ (_01035_, _01034_, _01033_);
  and _24059_ (_01036_, _01035_, _07196_);
  or _24060_ (_01037_, _01036_, _07161_);
  or _24061_ (_01038_, _01037_, _01021_);
  or _24062_ (_01039_, _07164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and _24063_ (_01040_, _01039_, _06989_);
  and _24064_ (_00272_, _01040_, _01038_);
  nor _24065_ (_01041_, _07196_, _07161_);
  and _24066_ (_01042_, _07222_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  not _24067_ (_01043_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _24068_ (_01044_, _01007_, _01043_);
  nand _24069_ (_01045_, _01044_, _01010_);
  or _24070_ (_01046_, _07464_, _07219_);
  and _24071_ (_01047_, _01046_, _01045_);
  or _24072_ (_01048_, _01047_, _07206_);
  or _24073_ (_01049_, _07166_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _24074_ (_01050_, _01049_, _00969_);
  and _24075_ (_01051_, _01050_, _00968_);
  and _24076_ (_01052_, _01051_, _01048_);
  and _24077_ (_01053_, _07464_, _07204_);
  or _24078_ (_01054_, _01053_, _07201_);
  or _24079_ (_01055_, _01054_, _01052_);
  nor _24080_ (_01056_, _01049_, _07202_);
  nor _24081_ (_01057_, _01056_, _07222_);
  and _24082_ (_01058_, _01057_, _01055_);
  or _24083_ (_01059_, _01058_, _01042_);
  and _24084_ (_01060_, _01059_, _01041_);
  or _24085_ (_01061_, _07189_, _07182_);
  or _24086_ (_01062_, _01061_, _07175_);
  and _24087_ (_01063_, _01062_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or _24088_ (_01064_, _01063_, _07179_);
  nand _24089_ (_01065_, _07182_, _07166_);
  and _24090_ (_01066_, _01065_, _01064_);
  or _24091_ (_01067_, _01066_, _07191_);
  nand _24092_ (_01068_, _07189_, _07166_);
  and _24093_ (_01069_, _01068_, _01067_);
  or _24094_ (_01070_, _07186_, _07161_);
  or _24095_ (_01071_, _01070_, _01069_);
  or _24096_ (_01072_, _07277_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or _24097_ (_01073_, \oc8051_top_1.oc8051_memory_interface1.reti , _07165_);
  or _24098_ (_01074_, _01073_, _07170_);
  and _24099_ (_01075_, _01074_, _01072_);
  and _24100_ (_01076_, _01075_, _01071_);
  or _24101_ (_01077_, _01076_, _01060_);
  and _24102_ (_00275_, _01077_, _06989_);
  nand _24103_ (_01078_, _07277_, _07223_);
  or _24104_ (_01079_, _01041_, _07166_);
  and _24105_ (_01080_, _01079_, _06989_);
  and _24106_ (_00289_, _01080_, _01078_);
  and _24107_ (_01081_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _06989_);
  and _24108_ (_00310_, _01081_, _07161_);
  nor _24109_ (_01082_, _07216_, _07199_);
  and _24110_ (_01083_, _07219_, _07208_);
  nand _24111_ (_01084_, _01083_, _01082_);
  nor _24112_ (_01085_, _01084_, _07196_);
  and _24113_ (_01086_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  or _24114_ (_01087_, _07182_, _07161_);
  nor _24115_ (_01088_, _01087_, _07171_);
  not _24116_ (_01089_, _07194_);
  nor _24117_ (_01090_, _01089_, _07180_);
  and _24118_ (_01091_, _01090_, _01088_);
  or _24119_ (_01092_, _01091_, _01086_);
  or _24120_ (_01093_, _01092_, _01085_);
  and _24121_ (_00318_, _01093_, _06989_);
  or _24122_ (_01094_, _07218_, _07206_);
  and _24123_ (_01095_, _07216_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _24124_ (_01096_, _01095_, _01094_);
  and _24125_ (_01097_, _01096_, _00968_);
  and _24126_ (_01098_, _07274_, _07202_);
  and _24127_ (_01099_, _01098_, _01097_);
  or _24128_ (_01100_, _07191_, _07182_);
  and _24129_ (_01101_, _07180_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or _24130_ (_01102_, _01101_, _01100_);
  and _24131_ (_01103_, _01102_, _00980_);
  and _24132_ (_01104_, _07196_, _07187_);
  and _24133_ (_01105_, _01104_, _01103_);
  or _24134_ (_01106_, _01105_, _07161_);
  or _24135_ (_01107_, _01106_, _01099_);
  or _24136_ (_01108_, _07164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _24137_ (_01109_, _01108_, _06989_);
  and _24138_ (_00321_, _01109_, _01107_);
  nor _24139_ (_01110_, _07212_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _24140_ (_01111_, _01110_, _07215_);
  or _24141_ (_01112_, _01111_, _07218_);
  and _24142_ (_01113_, _01112_, _00969_);
  or _24143_ (_01114_, _01113_, _07204_);
  and _24144_ (_01115_, _01114_, _01098_);
  nor _24145_ (_01116_, _07175_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor _24146_ (_01117_, _01116_, _07179_);
  or _24147_ (_01118_, _01117_, _07182_);
  and _24148_ (_01119_, _01118_, _00984_);
  or _24149_ (_01120_, _01119_, _07189_);
  and _24150_ (_01121_, _01120_, _01104_);
  or _24151_ (_01122_, _01121_, _07161_);
  or _24152_ (_01123_, _01122_, _01115_);
  or _24153_ (_01124_, _07164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _24154_ (_01125_, _01124_, _06989_);
  and _24155_ (_00325_, _01125_, _01123_);
  and _24156_ (_00327_, _12822_, _07161_);
  and _24157_ (_01126_, _14028_, _07048_);
  nand _24158_ (_01127_, _01126_, _06968_);
  or _24159_ (_01128_, _01126_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _24160_ (_01129_, _01128_, _14032_);
  and _24161_ (_01130_, _01129_, _01127_);
  nor _24162_ (_01131_, _14032_, _07118_);
  or _24163_ (_01132_, _01131_, _01130_);
  and _24164_ (_00334_, _01132_, _06989_);
  and _24165_ (_01133_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or _24166_ (_01134_, _01133_, _00998_);
  and _24167_ (_00345_, _01134_, _06989_);
  and _24168_ (_01135_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or _24169_ (_01136_, _01135_, _00998_);
  and _24170_ (_00348_, _01136_, _06989_);
  or _24171_ (_01137_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  nand _24172_ (_01138_, _07493_, _09525_);
  and _24173_ (_01139_, _01138_, _06989_);
  and _24174_ (_00387_, _01139_, _01137_);
  and _24175_ (_01140_, _12937_, _09009_);
  and _24176_ (_01141_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  or _24177_ (_01142_, _01141_, _01140_);
  and _24178_ (_00442_, _01142_, _06989_);
  or _24179_ (_01143_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  not _24180_ (_01144_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _24181_ (_01145_, _08139_, _01144_);
  and _24182_ (_01146_, _01145_, _06989_);
  and _24183_ (_00445_, _01146_, _01143_);
  and _24184_ (_01147_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or _24185_ (_00453_, _01147_, _09459_);
  or _24186_ (_01148_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  not _24187_ (_01149_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand _24188_ (_01150_, _08139_, _01149_);
  and _24189_ (_01151_, _01150_, _06989_);
  and _24190_ (_00457_, _01151_, _01148_);
  and _24191_ (_01152_, _09418_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or _24192_ (_00465_, _01152_, _09466_);
  nor _24193_ (_01153_, _12938_, _07317_);
  and _24194_ (_01154_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or _24195_ (_01155_, _01154_, _01153_);
  and _24196_ (_00494_, _01155_, _06989_);
  and _24197_ (_01156_, _00690_, _09022_);
  and _24198_ (_01157_, _01156_, _06539_);
  nand _24199_ (_01158_, _01157_, _06968_);
  or _24200_ (_01159_, _01157_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and _24201_ (_01160_, _01159_, _06485_);
  and _24202_ (_01161_, _01160_, _01158_);
  and _24203_ (_01162_, _00713_, _07125_);
  not _24204_ (_01163_, _01162_);
  nor _24205_ (_01164_, _01163_, _07040_);
  not _24206_ (_01165_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  nor _24207_ (_01166_, _01162_, _01165_);
  or _24208_ (_01167_, _01166_, _01164_);
  and _24209_ (_01168_, _01167_, _06983_);
  nor _24210_ (_01169_, _06484_, _01165_);
  or _24211_ (_01170_, _01169_, rst);
  or _24212_ (_01171_, _01170_, _01168_);
  or _24213_ (_00502_, _01171_, _01161_);
  and _24214_ (_01172_, _14190_, _07429_);
  and _24215_ (_01173_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  or _24216_ (_01174_, _01173_, _01172_);
  and _24217_ (_00529_, _01174_, _06989_);
  and _24218_ (_01175_, _14028_, _08349_);
  not _24219_ (_01176_, _14028_);
  or _24220_ (_01177_, _00817_, _01176_);
  and _24221_ (_01179_, _14028_, _06525_);
  or _24222_ (_01180_, _01179_, _01177_);
  and _24223_ (_01181_, _01180_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or _24224_ (_01182_, _01181_, _14031_);
  or _24225_ (_01183_, _01182_, _01175_);
  nand _24226_ (_01184_, _14031_, _07260_);
  and _24227_ (_01185_, _01184_, _06989_);
  and _24228_ (_00570_, _01185_, _01183_);
  or _24229_ (_01186_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not _24230_ (_01188_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand _24231_ (_01189_, _08139_, _01188_);
  and _24232_ (_01190_, _01189_, _06989_);
  and _24233_ (_00575_, _01190_, _01186_);
  or _24234_ (_01191_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  not _24235_ (_01192_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _24236_ (_01193_, _08139_, _01192_);
  and _24237_ (_01194_, _01193_, _06989_);
  and _24238_ (_00588_, _01194_, _01191_);
  nor _24239_ (_00596_, _11513_, rst);
  and _24240_ (_01195_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor _24241_ (_01196_, _08139_, _01192_);
  or _24242_ (_01197_, _01196_, _01195_);
  and _24243_ (_00638_, _01197_, _06989_);
  not _24244_ (_01198_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor _24245_ (_01199_, _00749_, _01198_);
  or _24246_ (_01200_, _01199_, _08437_);
  and _24247_ (_01202_, _01200_, _14028_);
  nor _24248_ (_01203_, _01179_, _01198_);
  or _24249_ (_01204_, _01203_, _14031_);
  or _24250_ (_01205_, _01204_, _01202_);
  nand _24251_ (_01206_, _14031_, _07317_);
  and _24252_ (_01207_, _01206_, _06989_);
  and _24253_ (_00639_, _01207_, _01205_);
  nor _24254_ (_01209_, _10961_, _07335_);
  nor _24255_ (_01210_, _10950_, _07349_);
  and _24256_ (_01211_, _10950_, _07349_);
  nor _24257_ (_01212_, _01211_, _01210_);
  and _24258_ (_01213_, _01212_, _01209_);
  nor _24259_ (_01214_, _01212_, _01209_);
  nor _24260_ (_01215_, _01214_, _01213_);
  or _24261_ (_01216_, _01215_, _07490_);
  or _24262_ (_01217_, _07325_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and _24263_ (_01218_, _01217_, _10964_);
  and _24264_ (_00647_, _01218_, _01216_);
  or _24265_ (_01219_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  not _24266_ (_01220_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _24267_ (_01221_, _08139_, _01220_);
  and _24268_ (_01222_, _01221_, _06989_);
  and _24269_ (_00663_, _01222_, _01219_);
  and _24270_ (_01223_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor _24271_ (_01224_, _08139_, _01220_);
  or _24272_ (_01225_, _01224_, _01223_);
  and _24273_ (_00667_, _01225_, _06989_);
  or _24274_ (_01226_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  not _24275_ (_01227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _24276_ (_01228_, _08139_, _01227_);
  and _24277_ (_01229_, _01228_, _06989_);
  and _24278_ (_00679_, _01229_, _01226_);
  and _24279_ (_01230_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not _24280_ (_01231_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _24281_ (_01232_, _08139_, _01231_);
  or _24282_ (_01233_, _01232_, _01230_);
  and _24283_ (_00681_, _01233_, _06989_);
  or _24284_ (_01234_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand _24285_ (_01235_, _07493_, _14104_);
  and _24286_ (_01236_, _01235_, _06989_);
  and _24287_ (_00705_, _01236_, _01234_);
  nor _24288_ (_01237_, _13945_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor _24289_ (_01238_, _01237_, _13946_);
  and _24290_ (_00794_, _01238_, _13953_);
  and _24291_ (_01239_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or _24292_ (_01241_, _01239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and _24293_ (_01000_, _01241_, _06989_);
  and _24294_ (_01242_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or _24295_ (_01243_, _01242_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and _24296_ (_01023_, _01243_, _06989_);
  not _24297_ (_01244_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nor _24298_ (_01245_, _14404_, _01244_);
  nand _24299_ (_01246_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand _24300_ (_01247_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _24301_ (_01248_, _01247_, _01246_);
  nand _24302_ (_01249_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nand _24303_ (_01251_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and _24304_ (_01252_, _01251_, _01249_);
  and _24305_ (_01253_, _01252_, _01248_);
  nand _24306_ (_01254_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  nand _24307_ (_01255_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _24308_ (_01256_, _01255_, _01254_);
  nand _24309_ (_01257_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nand _24310_ (_01258_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and _24311_ (_01259_, _01258_, _01257_);
  and _24312_ (_01260_, _01259_, _01256_);
  and _24313_ (_01261_, _01260_, _01253_);
  nand _24314_ (_01262_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nand _24315_ (_01263_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _24316_ (_01264_, _01263_, _01262_);
  nand _24317_ (_01265_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nand _24318_ (_01266_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and _24319_ (_01267_, _01266_, _01265_);
  and _24320_ (_01268_, _01267_, _01264_);
  nand _24321_ (_01269_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  nand _24322_ (_01270_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and _24323_ (_01271_, _01270_, _01269_);
  nand _24324_ (_01272_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  nand _24325_ (_01273_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and _24326_ (_01274_, _01273_, _01272_);
  and _24327_ (_01275_, _01274_, _01271_);
  and _24328_ (_01276_, _01275_, _01268_);
  and _24329_ (_01277_, _01276_, _01261_);
  nand _24330_ (_01278_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand _24331_ (_01279_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  and _24332_ (_01280_, _01279_, _01278_);
  nand _24333_ (_01281_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _24334_ (_01282_, _14296_, _11683_);
  and _24335_ (_01283_, _01282_, _01281_);
  and _24336_ (_01284_, _01283_, _01280_);
  nor _24337_ (_01285_, _14326_, p0_in[5]);
  not _24338_ (_01286_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _24339_ (_01287_, _14326_, _01286_);
  nor _24340_ (_01288_, _01287_, _01285_);
  nand _24341_ (_01289_, _01288_, _14339_);
  nor _24342_ (_01290_, _14326_, p1_in[5]);
  not _24343_ (_01291_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _24344_ (_01292_, _14326_, _01291_);
  nor _24345_ (_01293_, _01292_, _01290_);
  nand _24346_ (_01294_, _01293_, _14344_);
  and _24347_ (_01295_, _01294_, _01289_);
  or _24348_ (_01296_, _14326_, p2_in[5]);
  or _24349_ (_01297_, _14328_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _24350_ (_01298_, _01297_, _01296_);
  nand _24351_ (_01299_, _01298_, _14333_);
  nor _24352_ (_01300_, _14326_, p3_in[5]);
  not _24353_ (_01301_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _24354_ (_01302_, _14326_, _01301_);
  nor _24355_ (_01303_, _01302_, _01300_);
  nand _24356_ (_01304_, _01303_, _14305_);
  and _24357_ (_01305_, _01304_, _01299_);
  and _24358_ (_01306_, _01305_, _01295_);
  and _24359_ (_01307_, _01306_, _01284_);
  nand _24360_ (_01308_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  nand _24361_ (_01309_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and _24362_ (_01310_, _01309_, _01308_);
  and _24363_ (_01311_, _01310_, _01307_);
  nand _24364_ (_01312_, _01311_, _01277_);
  and _24365_ (_01313_, _01312_, _14374_);
  or _24366_ (_01314_, _01313_, _14213_);
  or _24367_ (_01315_, _01314_, _01245_);
  or _24368_ (_01316_, _14483_, _08268_);
  and _24369_ (_01317_, _01316_, _06989_);
  and _24370_ (_01187_, _01317_, _01315_);
  and _24371_ (_01318_, _00690_, _08038_);
  nand _24372_ (_01319_, _01318_, _06979_);
  or _24373_ (_01320_, _01319_, _08268_);
  not _24374_ (_01321_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand _24375_ (_01322_, _01319_, _01321_);
  and _24376_ (_01323_, _01322_, _06983_);
  and _24377_ (_01324_, _01323_, _01320_);
  nor _24378_ (_01325_, _06484_, _01321_);
  and _24379_ (_01326_, _01318_, _07048_);
  nand _24380_ (_01327_, _01326_, _06968_);
  or _24381_ (_01328_, _01326_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and _24382_ (_01329_, _01328_, _06485_);
  and _24383_ (_01330_, _01329_, _01327_);
  or _24384_ (_01331_, _01330_, _01325_);
  or _24385_ (_01332_, _01331_, _01324_);
  and _24386_ (_01201_, _01332_, _06989_);
  nor _24387_ (_01333_, _11529_, _07262_);
  and _24388_ (_01334_, _10974_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or _24389_ (_01335_, _01334_, _01333_);
  and _24390_ (_01208_, _01335_, _06989_);
  and _24391_ (_01336_, _09599_, _09488_);
  and _24392_ (_01337_, _09489_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or _24393_ (_01338_, _01337_, _01336_);
  and _24394_ (_01240_, _01338_, _06989_);
  and _24395_ (_01339_, _09599_, _09605_);
  and _24396_ (_01340_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or _24397_ (_01341_, _01340_, _06982_);
  or _24398_ (_01342_, _01341_, _01339_);
  or _24399_ (_01343_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and _24400_ (_01344_, _01343_, _06989_);
  and _24401_ (_01250_, _01344_, _01342_);
  and _24402_ (_01345_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  not _24403_ (_01346_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _24404_ (_01347_, _08139_, _01346_);
  or _24405_ (_01348_, _01347_, _01345_);
  and _24406_ (_01627_, _01348_, _06989_);
  and _24407_ (_01349_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not _24408_ (_01350_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _24409_ (_01351_, _08139_, _01350_);
  or _24410_ (_01352_, _01351_, _01349_);
  and _24411_ (_01629_, _01352_, _06989_);
  or _24412_ (_01353_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _24413_ (_01354_, _01353_, _14028_);
  nand _24414_ (_01355_, _08032_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand _24415_ (_01356_, _01355_, _14028_);
  or _24416_ (_01357_, _01356_, _08033_);
  and _24417_ (_01358_, _01357_, _01354_);
  or _24418_ (_01359_, _01358_, _14031_);
  nand _24419_ (_01360_, _14031_, _09008_);
  and _24420_ (_01361_, _01360_, _06989_);
  and _24421_ (_01649_, _01361_, _01359_);
  and _24422_ (_01363_, _14190_, _07410_);
  and _24423_ (_01364_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or _24424_ (_01365_, _01364_, _01363_);
  and _24425_ (_01662_, _01365_, _06989_);
  nor _24426_ (_01366_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and _24427_ (_01367_, _01366_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  not _24428_ (_01368_, _01367_);
  or _24429_ (_01369_, _01368_, _08433_);
  or _24430_ (_01370_, _01367_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and _24431_ (_01371_, _01370_, _06989_);
  and _24432_ (_01669_, _01371_, _01369_);
  not _24433_ (_01372_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or _24434_ (_01373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01372_);
  or _24435_ (_01374_, _01373_, _09392_);
  and _24436_ (_01375_, _01374_, _00895_);
  or _24437_ (_01376_, _01375_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _24438_ (_01377_, _01376_, _14028_);
  or _24439_ (_01378_, _06979_, _09407_);
  nand _24440_ (_01379_, _01378_, _14028_);
  or _24441_ (_01380_, _01379_, _08127_);
  and _24442_ (_01381_, _01380_, _01377_);
  or _24443_ (_01382_, _01381_, _14031_);
  nand _24444_ (_01383_, _14031_, _09598_);
  and _24445_ (_01384_, _01383_, _06989_);
  and _24446_ (_01673_, _01384_, _01382_);
  and _24447_ (_01385_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or _24448_ (_01386_, _01385_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and _24449_ (_01695_, _01386_, _06989_);
  and _24450_ (_01387_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or _24451_ (_01388_, _01387_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and _24452_ (_01697_, _01388_, _06989_);
  nand _24453_ (_01389_, _01367_, _09227_);
  or _24454_ (_01390_, _01367_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and _24455_ (_01391_, _01390_, _06989_);
  and _24456_ (_01711_, _01391_, _01389_);
  and _24457_ (_01392_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and _24458_ (_01393_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or _24459_ (_01394_, _01393_, _01392_);
  and _24460_ (_01721_, _01394_, _06989_);
  and _24461_ (_01395_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or _24462_ (_01396_, _01395_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and _24463_ (_01732_, _01396_, _06989_);
  and _24464_ (_01397_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or _24465_ (_01398_, _01397_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and _24466_ (_01734_, _01398_, _06989_);
  or _24467_ (_01399_, _01368_, _08030_);
  or _24468_ (_01400_, _01367_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and _24469_ (_01401_, _01400_, _06989_);
  and _24470_ (_01762_, _01401_, _01399_);
  and _24471_ (_01402_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and _24472_ (_01403_, _14190_, _11646_);
  or _24473_ (_01404_, _01403_, _01402_);
  and _24474_ (_01770_, _01404_, _06989_);
  and _24475_ (_01405_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor _24476_ (_01406_, _07486_, _07040_);
  or _24477_ (_01407_, _01406_, _01405_);
  and _24478_ (_01800_, _01407_, _06989_);
  or _24479_ (_01408_, _01368_, _08123_);
  or _24480_ (_01409_, _01367_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and _24481_ (_01410_, _01409_, _06989_);
  and _24482_ (_01803_, _01410_, _01408_);
  and _24483_ (_01411_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and _24484_ (_01412_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or _24485_ (_01413_, _01412_, _01411_);
  and _24486_ (_01817_, _01413_, _06989_);
  nor _24487_ (_01821_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  not _24488_ (_01414_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nor _24489_ (_01415_, _14404_, _01414_);
  nand _24490_ (_01416_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand _24491_ (_01417_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _24492_ (_01418_, _01417_, _01416_);
  nand _24493_ (_01419_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nand _24494_ (_01420_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _24495_ (_01421_, _01420_, _01419_);
  and _24496_ (_01422_, _01421_, _01418_);
  nand _24497_ (_01423_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  nand _24498_ (_01424_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _24499_ (_01425_, _01424_, _01423_);
  nand _24500_ (_01426_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nand _24501_ (_01427_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and _24502_ (_01428_, _01427_, _01426_);
  and _24503_ (_01429_, _01428_, _01425_);
  and _24504_ (_01430_, _01429_, _01422_);
  nand _24505_ (_01431_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nand _24506_ (_01432_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and _24507_ (_01433_, _01432_, _01431_);
  nand _24508_ (_01434_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand _24509_ (_01435_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and _24510_ (_01436_, _01435_, _01434_);
  and _24511_ (_01437_, _01436_, _01433_);
  nand _24512_ (_01438_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nand _24513_ (_01439_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  and _24514_ (_01440_, _01439_, _01438_);
  nand _24515_ (_01441_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nand _24516_ (_01442_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _24517_ (_01443_, _01442_, _01441_);
  and _24518_ (_01444_, _01443_, _01440_);
  and _24519_ (_01445_, _01444_, _01437_);
  and _24520_ (_01446_, _01445_, _01430_);
  nand _24521_ (_01447_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _24522_ (_01448_, _14296_, _11698_);
  and _24523_ (_01449_, _01448_, _01447_);
  nand _24524_ (_01450_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  nand _24525_ (_01451_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and _24526_ (_01452_, _01451_, _01450_);
  and _24527_ (_01453_, _01452_, _01449_);
  nor _24528_ (_01454_, _14326_, p1_in[4]);
  not _24529_ (_01455_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _24530_ (_01456_, _14326_, _01455_);
  nor _24531_ (_01457_, _01456_, _01454_);
  nand _24532_ (_01458_, _01457_, _14344_);
  nor _24533_ (_01459_, _14326_, p0_in[4]);
  not _24534_ (_01460_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _24535_ (_01461_, _14326_, _01460_);
  nor _24536_ (_01462_, _01461_, _01459_);
  nand _24537_ (_01463_, _01462_, _14339_);
  and _24538_ (_01464_, _01463_, _01458_);
  nor _24539_ (_01465_, _14326_, p3_in[4]);
  not _24540_ (_01466_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _24541_ (_01467_, _14326_, _01466_);
  nor _24542_ (_01468_, _01467_, _01465_);
  nand _24543_ (_01469_, _01468_, _14305_);
  nor _24544_ (_01470_, _14326_, p2_in[4]);
  not _24545_ (_01471_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _24546_ (_01472_, _14326_, _01471_);
  nor _24547_ (_01473_, _01472_, _01470_);
  nand _24548_ (_01474_, _01473_, _14333_);
  and _24549_ (_01475_, _01474_, _01469_);
  and _24550_ (_01476_, _01475_, _01464_);
  and _24551_ (_01477_, _01476_, _01453_);
  nand _24552_ (_01478_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nand _24553_ (_01479_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _24554_ (_01480_, _01479_, _01478_);
  and _24555_ (_01481_, _01480_, _01477_);
  nand _24556_ (_01482_, _01481_, _01446_);
  nand _24557_ (_01483_, _01482_, _14374_);
  nand _24558_ (_01484_, _01483_, _14483_);
  or _24559_ (_01485_, _01484_, _01415_);
  or _24560_ (_01486_, _14483_, _08346_);
  and _24561_ (_01487_, _01486_, _06989_);
  and _24562_ (_01823_, _01487_, _01485_);
  nand _24563_ (_01488_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand _24564_ (_01489_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _24565_ (_01490_, _01489_, _01488_);
  nand _24566_ (_01491_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _24567_ (_01492_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _24568_ (_01493_, _01492_, _01491_);
  and _24569_ (_01494_, _01493_, _01490_);
  nand _24570_ (_01495_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  nand _24571_ (_01496_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _24572_ (_01497_, _01496_, _01495_);
  nand _24573_ (_01498_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  nand _24574_ (_01499_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and _24575_ (_01500_, _01499_, _01498_);
  and _24576_ (_01501_, _01500_, _01497_);
  and _24577_ (_01502_, _01501_, _01494_);
  nand _24578_ (_01503_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nand _24579_ (_01504_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and _24580_ (_01505_, _01504_, _01503_);
  nand _24581_ (_01506_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nand _24582_ (_01507_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and _24583_ (_01508_, _01507_, _01506_);
  and _24584_ (_01509_, _01508_, _01505_);
  nand _24585_ (_01510_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand _24586_ (_01511_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  and _24587_ (_01512_, _01511_, _01510_);
  nand _24588_ (_01513_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand _24589_ (_01514_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _24590_ (_01515_, _01514_, _01513_);
  and _24591_ (_01516_, _01515_, _01512_);
  and _24592_ (_01517_, _01516_, _01509_);
  and _24593_ (_01518_, _01517_, _01502_);
  nand _24594_ (_01519_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  nand _24595_ (_01520_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  and _24596_ (_01521_, _01520_, _01519_);
  nand _24597_ (_01522_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _24598_ (_01523_, _14296_, _11795_);
  and _24599_ (_01524_, _01523_, _01522_);
  and _24600_ (_01525_, _01524_, _01521_);
  nor _24601_ (_01527_, _14326_, p2_in[0]);
  not _24602_ (_01528_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _24603_ (_01529_, _14326_, _01528_);
  nor _24604_ (_01530_, _01529_, _01527_);
  nand _24605_ (_01531_, _01530_, _14333_);
  nor _24606_ (_01532_, _14326_, p3_in[0]);
  not _24607_ (_01533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _24608_ (_01534_, _14326_, _01533_);
  nor _24609_ (_01535_, _01534_, _01532_);
  nand _24610_ (_01536_, _01535_, _14305_);
  and _24611_ (_01537_, _01536_, _01531_);
  nor _24612_ (_01538_, _14326_, p0_in[0]);
  not _24613_ (_01539_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _24614_ (_01540_, _14326_, _01539_);
  nor _24615_ (_01541_, _01540_, _01538_);
  nand _24616_ (_01542_, _01541_, _14339_);
  nor _24617_ (_01543_, _14326_, p1_in[0]);
  not _24618_ (_01544_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _24619_ (_01545_, _14326_, _01544_);
  nor _24620_ (_01546_, _01545_, _01543_);
  nand _24621_ (_01547_, _01546_, _14344_);
  and _24622_ (_01548_, _01547_, _01542_);
  and _24623_ (_01549_, _01548_, _01537_);
  and _24624_ (_01550_, _01549_, _01525_);
  nand _24625_ (_01551_, _08359_, _08279_);
  or _24626_ (_01552_, _08359_, _08279_);
  nand _24627_ (_01553_, _01552_, _01551_);
  or _24628_ (_01554_, _09145_, _07710_);
  not _24629_ (_01555_, _14196_);
  nor _24630_ (_01556_, _06968_, _01555_);
  nor _24631_ (_01557_, _14196_, _06813_);
  nor _24632_ (_01558_, _01557_, _01556_);
  nor _24633_ (_01559_, _01558_, _08043_);
  nor _24634_ (_01560_, _11948_, _06813_);
  or _24635_ (_01561_, _01560_, _07699_);
  nor _24636_ (_01562_, _01561_, _01559_);
  nand _24637_ (_01563_, _01562_, _01554_);
  and _24638_ (_01564_, _09285_, _07699_);
  not _24639_ (_01565_, _01564_);
  and _24640_ (_01566_, _01565_, _01563_);
  or _24641_ (_01567_, _01566_, _12316_);
  nand _24642_ (_01568_, _01566_, _12316_);
  and _24643_ (_01569_, _01568_, _01567_);
  nand _24644_ (_01570_, _01569_, _01553_);
  or _24645_ (_01571_, _01569_, _01553_);
  nand _24646_ (_01572_, _01571_, _01570_);
  nand _24647_ (_01573_, _08138_, _08052_);
  or _24648_ (_01574_, _08138_, _08052_);
  nand _24649_ (_01575_, _01574_, _01573_);
  or _24650_ (_01576_, _09227_, _07710_);
  nor _24651_ (_01577_, _09074_, _06703_);
  nor _24652_ (_01578_, _01577_, _00760_);
  nor _24653_ (_01579_, _01578_, _08043_);
  nor _24654_ (_01580_, _11948_, _06703_);
  or _24655_ (_01581_, _01580_, _07699_);
  nor _24656_ (_01582_, _01581_, _01579_);
  nand _24657_ (_01583_, _01582_, _01576_);
  and _24658_ (_01584_, _09356_, _07699_);
  not _24659_ (_01585_, _01584_);
  and _24660_ (_01586_, _01585_, _01583_);
  or _24661_ (_01587_, _01586_, _08447_);
  nand _24662_ (_01588_, _01586_, _08447_);
  and _24663_ (_01589_, _01588_, _01587_);
  nand _24664_ (_01590_, _01589_, _01575_);
  or _24665_ (_01591_, _01589_, _01575_);
  nand _24666_ (_01592_, _01591_, _01590_);
  nand _24667_ (_01593_, _01592_, _01572_);
  or _24668_ (_01594_, _01592_, _01572_);
  and _24669_ (_01595_, _01594_, _01593_);
  nand _24670_ (_01596_, _01595_, _14355_);
  nand _24671_ (_01597_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and _24672_ (_01598_, _01597_, _01596_);
  and _24673_ (_01599_, _01598_, _01550_);
  and _24674_ (_01600_, _01599_, _01518_);
  nor _24675_ (_01601_, _01600_, _14377_);
  not _24676_ (_01602_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nor _24677_ (_01603_, _14404_, _01602_);
  or _24678_ (_01604_, _01603_, _14213_);
  or _24679_ (_01605_, _01604_, _01601_);
  or _24680_ (_01606_, _14483_, _08123_);
  and _24681_ (_01607_, _01606_, _06989_);
  and _24682_ (_01825_, _01607_, _01605_);
  and _24683_ (_01608_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor _24684_ (_01609_, _08139_, _00687_);
  or _24685_ (_01610_, _01609_, _01608_);
  and _24686_ (_01835_, _01610_, _06989_);
  not _24687_ (_01611_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not _24688_ (_01612_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _24689_ (_01613_, _11004_, _01612_);
  and _24690_ (_01614_, _01613_, _01611_);
  nor _24691_ (_01615_, _01613_, _01611_);
  nor _24692_ (_01616_, _01615_, _01614_);
  not _24693_ (_01617_, _01616_);
  nor _24694_ (_01618_, _11004_, _01612_);
  or _24695_ (_01619_, _01618_, _01613_);
  and _24696_ (_01620_, _01619_, _11055_);
  and _24697_ (_01621_, _01620_, _01617_);
  nor _24698_ (_01622_, _01620_, _01617_);
  nor _24699_ (_01623_, _01622_, _01621_);
  or _24700_ (_01624_, _01623_, _08477_);
  or _24701_ (_01625_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _24702_ (_01626_, _01625_, _10964_);
  and _24703_ (_01628_, _01626_, _01624_);
  and _24704_ (_01630_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _24705_ (_01860_, _01630_, _01628_);
  not _24706_ (_01631_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not _24707_ (_01632_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not _24708_ (_01633_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and _24709_ (_01634_, _01614_, _01633_);
  and _24710_ (_01635_, _01634_, _01632_);
  nor _24711_ (_01636_, _01635_, _01631_);
  and _24712_ (_01637_, _01635_, _01631_);
  nor _24713_ (_01638_, _01637_, _01636_);
  not _24714_ (_01639_, _01638_);
  nor _24715_ (_01640_, _01634_, _01632_);
  or _24716_ (_01641_, _01640_, _01635_);
  nor _24717_ (_01642_, _01614_, _01633_);
  nor _24718_ (_01643_, _01642_, _01634_);
  not _24719_ (_01644_, _01643_);
  and _24720_ (_01645_, _01644_, _01621_);
  and _24721_ (_01646_, _01645_, _01641_);
  and _24722_ (_01647_, _01646_, _01639_);
  nor _24723_ (_01648_, _01646_, _01639_);
  nor _24724_ (_01650_, _01648_, _01647_);
  or _24725_ (_01651_, _01650_, _08477_);
  or _24726_ (_01652_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and _24727_ (_01653_, _01652_, _10964_);
  and _24728_ (_01654_, _01653_, _01651_);
  and _24729_ (_01655_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _24730_ (_01865_, _01655_, _01654_);
  nor _24731_ (_01656_, _01645_, _01641_);
  nor _24732_ (_01657_, _01656_, _01646_);
  or _24733_ (_01658_, _01657_, _08477_);
  or _24734_ (_01659_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _24735_ (_01660_, _01659_, _10964_);
  and _24736_ (_01661_, _01660_, _01658_);
  and _24737_ (_01663_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or _24738_ (_01870_, _01663_, _01661_);
  nor _24739_ (_01664_, _13943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor _24740_ (_01665_, _01664_, _13944_);
  and _24741_ (_01896_, _01665_, _13953_);
  and _24742_ (_01666_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _24743_ (_01667_, _08139_, _00659_);
  or _24744_ (_01668_, _01667_, _01666_);
  and _24745_ (_02001_, _01668_, _06989_);
  nor _24746_ (_01670_, _01644_, _01621_);
  nor _24747_ (_01671_, _01670_, _01645_);
  or _24748_ (_01672_, _01671_, _08477_);
  or _24749_ (_01674_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and _24750_ (_01675_, _01674_, _10964_);
  and _24751_ (_01676_, _01675_, _01672_);
  and _24752_ (_01677_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or _24753_ (_02024_, _01677_, _01676_);
  nor _24754_ (_01678_, _01619_, _11055_);
  nor _24755_ (_01679_, _01678_, _01620_);
  or _24756_ (_01680_, _01679_, _08477_);
  or _24757_ (_01681_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and _24758_ (_01682_, _01681_, _10964_);
  and _24759_ (_01683_, _01682_, _01680_);
  and _24760_ (_01684_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _24761_ (_02056_, _01684_, _01683_);
  and _24762_ (_01685_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _24763_ (_01686_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor _24764_ (_01687_, _08139_, _01686_);
  or _24765_ (_01688_, _01687_, _01685_);
  and _24766_ (_02058_, _01688_, _06989_);
  or _24767_ (_01689_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _24768_ (_01690_, _08139_, _08171_);
  and _24769_ (_01691_, _01690_, _06989_);
  and _24770_ (_02100_, _01691_, _01689_);
  or _24771_ (_01692_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and _24772_ (_01693_, _01692_, _06989_);
  nand _24773_ (_01694_, _14016_, _07118_);
  and _24774_ (_02185_, _01694_, _01693_);
  or _24775_ (_01696_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and _24776_ (_01698_, _01696_, _06989_);
  nand _24777_ (_01699_, _14016_, _10970_);
  and _24778_ (_02212_, _01699_, _01698_);
  or _24779_ (_01700_, _09760_, _09398_);
  or _24780_ (_01701_, _09762_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and _24781_ (_01702_, _01701_, _06989_);
  and _24782_ (_02225_, _01702_, _01700_);
  or _24783_ (_01703_, _14055_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand _24784_ (_01704_, _14055_, _14046_);
  and _24785_ (_01705_, _01704_, _06989_);
  and _24786_ (_02284_, _01705_, _01703_);
  or _24787_ (_01706_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and _24788_ (_01707_, _01706_, _06989_);
  nand _24789_ (_01708_, _14016_, _07260_);
  and _24790_ (_02286_, _01708_, _01707_);
  nor _24791_ (_01709_, _10970_, _09489_);
  nor _24792_ (_01710_, _07131_, _06982_);
  or _24793_ (_01712_, _01710_, _07134_);
  and _24794_ (_01713_, _01712_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  or _24795_ (_01714_, _01713_, _01709_);
  and _24796_ (_02294_, _01714_, _06989_);
  nor _24797_ (_01715_, _07260_, _09614_);
  and _24798_ (_01716_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or _24799_ (_01717_, _01716_, _06982_);
  or _24800_ (_01718_, _01717_, _01715_);
  or _24801_ (_01719_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and _24802_ (_01720_, _01719_, _06989_);
  and _24803_ (_02297_, _01720_, _01718_);
  or _24804_ (_01722_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and _24805_ (_01723_, _01722_, _06989_);
  nand _24806_ (_01724_, _14016_, _07317_);
  and _24807_ (_02300_, _01724_, _01723_);
  and _24808_ (_02542_, _01566_, _06989_);
  or _24809_ (_01725_, _01319_, _08433_);
  not _24810_ (_01726_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand _24811_ (_01727_, _01319_, _01726_);
  and _24812_ (_01728_, _01727_, _06983_);
  and _24813_ (_01729_, _01728_, _01725_);
  nor _24814_ (_01730_, _06484_, _01726_);
  nand _24815_ (_01731_, _01318_, _06525_);
  and _24816_ (_01733_, _01731_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor _24817_ (_01735_, _00749_, _01726_);
  or _24818_ (_01736_, _01735_, _08437_);
  and _24819_ (_01737_, _01736_, _01318_);
  or _24820_ (_01738_, _01737_, _01733_);
  and _24821_ (_01739_, _01738_, _06485_);
  or _24822_ (_01740_, _01739_, _01730_);
  or _24823_ (_01741_, _01740_, _01729_);
  and _24824_ (_02563_, _01741_, _06989_);
  and _24825_ (_02576_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _06989_);
  or _24826_ (_01742_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand _24827_ (_01743_, _07493_, _14099_);
  and _24828_ (_01744_, _01743_, _06989_);
  and _24829_ (_02578_, _01744_, _01742_);
  or _24830_ (_01745_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  or _24831_ (_01746_, _11273_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  and _24832_ (_01747_, _01746_, _06989_);
  and _24833_ (_02597_, _01747_, _01745_);
  or _24834_ (_01748_, _01319_, _08346_);
  not _24835_ (_01749_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand _24836_ (_01750_, _01319_, _01749_);
  and _24837_ (_01751_, _01750_, _06983_);
  and _24838_ (_01752_, _01751_, _01748_);
  nor _24839_ (_01753_, _06484_, _01749_);
  and _24840_ (_01754_, _01318_, _07044_);
  nand _24841_ (_01755_, _01754_, _06968_);
  or _24842_ (_01756_, _01754_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and _24843_ (_01757_, _01756_, _06485_);
  and _24844_ (_01758_, _01757_, _01755_);
  or _24845_ (_01759_, _01758_, _01753_);
  or _24846_ (_01760_, _01759_, _01752_);
  and _24847_ (_02622_, _01760_, _06989_);
  and _24848_ (_01761_, _09599_, _07261_);
  and _24849_ (_01763_, _10974_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  or _24850_ (_01764_, _01763_, _01761_);
  and _24851_ (_02650_, _01764_, _06989_);
  or _24852_ (_01765_, _00005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and _24853_ (_01766_, _01765_, _06989_);
  nand _24854_ (_01767_, _00005_, _07040_);
  and _24855_ (_02668_, _01767_, _01766_);
  nand _24856_ (_01768_, _00027_, _07040_);
  and _24857_ (_01769_, _00105_, _00059_);
  or _24858_ (_01771_, _01769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _24859_ (_01772_, _01769_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _24860_ (_01773_, _01772_, _01771_);
  and _24861_ (_01774_, _01773_, _00062_);
  and _24862_ (_01775_, _00084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and _24863_ (_01776_, _01775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _24864_ (_01777_, _01775_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _24865_ (_01778_, _01777_, _00083_);
  nor _24866_ (_01779_, _01778_, _01776_);
  or _24867_ (_01780_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _24868_ (_01781_, _01780_, _00051_);
  and _24869_ (_01782_, _00099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor _24870_ (_01783_, _01782_, _01781_);
  or _24871_ (_01784_, _01783_, _01779_);
  or _24872_ (_01785_, _01784_, _01774_);
  or _24873_ (_01786_, _01785_, _00027_);
  and _24874_ (_01787_, _01786_, _00092_);
  and _24875_ (_01788_, _01787_, _01768_);
  and _24876_ (_01789_, _00091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _24877_ (_01790_, _01789_, _01788_);
  and _24878_ (_02671_, _01790_, _06989_);
  not _24879_ (_01791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor _24880_ (_01792_, _00079_, _01791_);
  or _24881_ (_01793_, _01792_, _01776_);
  and _24882_ (_01794_, _01793_, _00083_);
  or _24883_ (_01795_, _00027_, rst);
  nor _24884_ (_01796_, _01795_, _00091_);
  and _24885_ (_02677_, _01796_, _01794_);
  nand _24886_ (_01797_, _00091_, _07040_);
  and _24887_ (_01798_, _00353_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and _24888_ (_01799_, _00052_, _00070_);
  nand _24889_ (_01801_, _01799_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or _24890_ (_01802_, _01799_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _24891_ (_01804_, _01802_, _01801_);
  or _24892_ (_01805_, _01804_, _01798_);
  or _24893_ (_01806_, _01805_, _00027_);
  or _24894_ (_01807_, _00097_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _24895_ (_01808_, _01807_, _01806_);
  or _24896_ (_01809_, _01808_, _00091_);
  and _24897_ (_01810_, _01809_, _06989_);
  and _24898_ (_02680_, _01810_, _01797_);
  not _24899_ (_01811_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor _24900_ (_01812_, _00040_, _01811_);
  or _24901_ (_01813_, _01812_, _01782_);
  and _24902_ (_01814_, _01813_, _00051_);
  and _24903_ (_01815_, _00105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or _24904_ (_01816_, _01815_, _01812_);
  and _24905_ (_01818_, _01816_, _00061_);
  or _24906_ (_01819_, _01812_, _00071_);
  and _24907_ (_01820_, _01819_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or _24908_ (_01822_, _01820_, _01818_);
  or _24909_ (_01824_, _01822_, _01814_);
  and _24910_ (_02683_, _01824_, _01796_);
  not _24911_ (_01826_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor _24912_ (_01827_, _00397_, _01826_);
  and _24913_ (_01828_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and _24914_ (_01829_, _01828_, _00419_);
  or _24915_ (_01830_, _01829_, _01827_);
  and _24916_ (_01831_, _01830_, _00410_);
  nand _24917_ (_01832_, _00397_, _00533_);
  and _24918_ (_01833_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and _24919_ (_01834_, _01833_, _01832_);
  or _24920_ (_01836_, _01834_, _00539_);
  and _24921_ (_01837_, _01828_, _00406_);
  or _24922_ (_01838_, _01837_, _01827_);
  and _24923_ (_01839_, _01838_, _00384_);
  or _24924_ (_01840_, _01839_, _01836_);
  or _24925_ (_01841_, _01840_, _01831_);
  and _24926_ (_01842_, _00430_, _06989_);
  and _24927_ (_02684_, _01842_, _01841_);
  and _24928_ (_02689_, t0_i, _06989_);
  nor _24929_ (_01843_, _00382_, _07040_);
  and _24930_ (_01844_, _00429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _24931_ (_01845_, _00407_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _24932_ (_01846_, _00407_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and _24933_ (_01847_, _01846_, _01845_);
  and _24934_ (_01848_, _01847_, _00384_);
  and _24935_ (_01849_, _00422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _24936_ (_01850_, _00420_, _00410_);
  nor _24937_ (_01851_, _01850_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _24938_ (_01852_, _01851_, _01849_);
  or _24939_ (_01853_, _01852_, _01848_);
  and _24940_ (_01854_, _01853_, _00430_);
  or _24941_ (_01855_, _01854_, _01844_);
  or _24942_ (_01856_, _01855_, _01843_);
  and _24943_ (_02692_, _01856_, _06989_);
  or _24944_ (_01857_, _00549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor _24945_ (_01858_, _00535_, _00439_);
  and _24946_ (_01859_, _01858_, _01857_);
  and _24947_ (_01861_, _00539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or _24948_ (_01862_, _01861_, _01859_);
  and _24949_ (_01863_, _01862_, _00430_);
  not _24950_ (_01864_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  or _24951_ (_01866_, _00429_, _01864_);
  nor _24952_ (_01867_, _01866_, _00543_);
  or _24953_ (_01868_, _01867_, _01863_);
  nor _24954_ (_01869_, _00594_, _07040_);
  or _24955_ (_01871_, _01869_, _01868_);
  and _24956_ (_02695_, _01871_, _06989_);
  and _24957_ (_02698_, t1_i, _06989_);
  nand _24958_ (_01872_, _14012_, _11529_);
  or _24959_ (_01873_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and _24960_ (_01874_, _01873_, _06989_);
  and _24961_ (_02703_, _01874_, _01872_);
  nand _24962_ (_01875_, _14012_, _09008_);
  or _24963_ (_01876_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and _24964_ (_01877_, _01876_, _06989_);
  and _24965_ (_02705_, _01877_, _01875_);
  nand _24966_ (_01878_, _14012_, _09598_);
  or _24967_ (_01879_, _14012_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and _24968_ (_01880_, _01879_, _06989_);
  and _24969_ (_02723_, _01880_, _01878_);
  nand _24970_ (_01881_, _12937_, _07040_);
  or _24971_ (_01882_, _12937_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and _24972_ (_01883_, _01882_, _06989_);
  and _24973_ (_02737_, _01883_, _01881_);
  or _24974_ (_01884_, _01319_, _11966_);
  not _24975_ (_01885_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand _24976_ (_01886_, _01319_, _01885_);
  and _24977_ (_01887_, _01886_, _06983_);
  and _24978_ (_01888_, _01887_, _01884_);
  nor _24979_ (_01889_, _06484_, _01885_);
  and _24980_ (_01890_, _01318_, _14196_);
  nand _24981_ (_01891_, _01890_, _06968_);
  or _24982_ (_01892_, _01890_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and _24983_ (_01893_, _01892_, _06485_);
  and _24984_ (_01894_, _01893_, _01891_);
  or _24985_ (_01895_, _01894_, _01889_);
  or _24986_ (_01897_, _01895_, _01888_);
  and _24987_ (_02756_, _01897_, _06989_);
  not _24988_ (_01898_, _09227_);
  or _24989_ (_01899_, _01319_, _01898_);
  not _24990_ (_01900_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand _24991_ (_01901_, _01319_, _01900_);
  and _24992_ (_01902_, _01901_, _06983_);
  and _24993_ (_01903_, _01902_, _01899_);
  nor _24994_ (_01904_, _06484_, _01900_);
  nand _24995_ (_01905_, _01318_, _00764_);
  and _24996_ (_01906_, _01905_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and _24997_ (_01907_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _24998_ (_01908_, _01907_, _00760_);
  and _24999_ (_01909_, _01908_, _01318_);
  or _25000_ (_01910_, _01909_, _01906_);
  and _25001_ (_01911_, _01910_, _06485_);
  or _25002_ (_01912_, _01911_, _01904_);
  or _25003_ (_01913_, _01912_, _01903_);
  and _25004_ (_02759_, _01913_, _06989_);
  or _25005_ (_01914_, _01319_, _08030_);
  not _25006_ (_01915_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand _25007_ (_01916_, _01319_, _01915_);
  and _25008_ (_01917_, _01916_, _06983_);
  and _25009_ (_01918_, _01917_, _01914_);
  nor _25010_ (_01919_, _06484_, _01915_);
  and _25011_ (_01920_, _01318_, _07089_);
  nand _25012_ (_01921_, _01920_, _06968_);
  or _25013_ (_01922_, _01920_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and _25014_ (_01923_, _01922_, _06485_);
  and _25015_ (_01924_, _01923_, _01921_);
  or _25016_ (_01925_, _01924_, _01919_);
  or _25017_ (_01926_, _01925_, _01918_);
  and _25018_ (_02805_, _01926_, _06989_);
  and _25019_ (_01927_, _01156_, _07089_);
  nand _25020_ (_01928_, _01927_, _06968_);
  or _25021_ (_01929_, _01927_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and _25022_ (_01930_, _01929_, _06485_);
  and _25023_ (_01931_, _01930_, _01928_);
  nor _25024_ (_01932_, _01163_, _09008_);
  and _25025_ (_01933_, _01163_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _25026_ (_01934_, _01933_, _01932_);
  and _25027_ (_01935_, _01934_, _06983_);
  and _25028_ (_01936_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or _25029_ (_01937_, _01936_, rst);
  or _25030_ (_01938_, _01937_, _01935_);
  or _25031_ (_02899_, _01938_, _01931_);
  and _25032_ (_01939_, _01156_, _07048_);
  nand _25033_ (_01940_, _01939_, _06968_);
  or _25034_ (_01941_, _01939_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and _25035_ (_01942_, _01941_, _06485_);
  and _25036_ (_01943_, _01942_, _01940_);
  nor _25037_ (_01944_, _01163_, _07118_);
  nor _25038_ (_01945_, _01162_, _01301_);
  or _25039_ (_01946_, _01945_, _01944_);
  and _25040_ (_01947_, _01946_, _06983_);
  nor _25041_ (_01948_, _06484_, _01301_);
  or _25042_ (_01949_, _01948_, rst);
  or _25043_ (_01950_, _01949_, _01947_);
  or _25044_ (_02900_, _01950_, _01943_);
  and _25045_ (_01951_, _09023_, _07089_);
  nand _25046_ (_01952_, _01951_, _06968_);
  or _25047_ (_01953_, _01951_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and _25048_ (_01954_, _01953_, _06485_);
  and _25049_ (_01955_, _01954_, _01952_);
  nor _25050_ (_01956_, _09031_, _09008_);
  and _25051_ (_01957_, _09031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _25052_ (_01958_, _01957_, _01956_);
  and _25053_ (_01959_, _01958_, _06983_);
  and _25054_ (_01960_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or _25055_ (_01961_, _01960_, rst);
  or _25056_ (_01962_, _01961_, _01959_);
  or _25057_ (_02903_, _01962_, _01955_);
  and _25058_ (_01963_, _09023_, _07048_);
  nand _25059_ (_01964_, _01963_, _06968_);
  or _25060_ (_01965_, _01963_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and _25061_ (_01966_, _01965_, _06485_);
  and _25062_ (_01967_, _01966_, _01964_);
  nor _25063_ (_01968_, _09031_, _07118_);
  and _25064_ (_01969_, _09031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _25065_ (_01970_, _01969_, _01968_);
  and _25066_ (_01971_, _01970_, _06983_);
  and _25067_ (_01972_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or _25068_ (_01973_, _01972_, rst);
  or _25069_ (_01974_, _01973_, _01971_);
  or _25070_ (_02905_, _01974_, _01967_);
  and _25071_ (_01975_, _00691_, _09074_);
  nand _25072_ (_01976_, _01975_, _06968_);
  or _25073_ (_01977_, _01975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _25074_ (_01978_, _01977_, _06485_);
  and _25075_ (_01979_, _01978_, _01976_);
  nand _25076_ (_01980_, _11529_, _00697_);
  or _25077_ (_01981_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and _25078_ (_01982_, _01981_, _06983_);
  and _25079_ (_01983_, _01982_, _01980_);
  nor _25080_ (_01984_, _06484_, _14532_);
  or _25081_ (_01985_, _01984_, rst);
  or _25082_ (_01986_, _01985_, _01983_);
  or _25083_ (_02907_, _01986_, _01979_);
  and _25084_ (_01987_, _00720_, _07048_);
  nand _25085_ (_01988_, _01987_, _06968_);
  or _25086_ (_01989_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _25087_ (_01990_, _01989_, _06485_);
  and _25088_ (_01991_, _01990_, _01988_);
  nand _25089_ (_01992_, _00726_, _07118_);
  or _25090_ (_01993_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and _25091_ (_01994_, _01993_, _06983_);
  and _25092_ (_01995_, _01994_, _01992_);
  nor _25093_ (_01996_, _06484_, _01286_);
  or _25094_ (_01997_, _01996_, rst);
  or _25095_ (_01998_, _01997_, _01995_);
  or _25096_ (_02909_, _01998_, _01991_);
  and _25097_ (_01999_, _00720_, _07089_);
  nand _25098_ (_02000_, _01999_, _06968_);
  or _25099_ (_02002_, _01999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _25100_ (_02003_, _02002_, _06485_);
  and _25101_ (_02004_, _02003_, _02000_);
  nand _25102_ (_02005_, _00726_, _09008_);
  or _25103_ (_02006_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and _25104_ (_02007_, _02006_, _06983_);
  and _25105_ (_02008_, _02007_, _02005_);
  and _25106_ (_02009_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or _25107_ (_02010_, _02009_, rst);
  or _25108_ (_02011_, _02010_, _02008_);
  or _25109_ (_02911_, _02011_, _02004_);
  and _25110_ (_02012_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor _25111_ (_02013_, _08139_, _01227_);
  or _25112_ (_02014_, _02013_, _02012_);
  and _25113_ (_02922_, _02014_, _06989_);
  nand _25114_ (_02015_, _01162_, _06968_);
  or _25115_ (_02016_, _01162_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and _25116_ (_02017_, _02016_, _06485_);
  and _25117_ (_02018_, _02017_, _02015_);
  and _25118_ (_02019_, _01162_, _09599_);
  nor _25119_ (_02020_, _01162_, _01533_);
  or _25120_ (_02021_, _02020_, _02019_);
  and _25121_ (_02022_, _02021_, _06983_);
  nor _25122_ (_02023_, _06484_, _01533_);
  or _25123_ (_02025_, _02023_, rst);
  or _25124_ (_02026_, _02025_, _02022_);
  or _25125_ (_02928_, _02026_, _02018_);
  and _25126_ (_02027_, _01156_, _08436_);
  nand _25127_ (_02028_, _02027_, _06968_);
  or _25128_ (_02029_, _02027_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and _25129_ (_02030_, _02029_, _06485_);
  and _25130_ (_02031_, _02030_, _02028_);
  nor _25131_ (_02032_, _01163_, _07317_);
  and _25132_ (_02033_, _01163_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _25133_ (_02034_, _02033_, _02032_);
  and _25134_ (_02035_, _02034_, _06983_);
  and _25135_ (_02036_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or _25136_ (_02037_, _02036_, rst);
  or _25137_ (_02038_, _02037_, _02035_);
  or _25138_ (_02930_, _02038_, _02031_);
  and _25139_ (_02039_, _00691_, _14196_);
  nand _25140_ (_02040_, _02039_, _06968_);
  or _25141_ (_02041_, _02039_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _25142_ (_02042_, _02041_, _06485_);
  and _25143_ (_02043_, _02042_, _02040_);
  nand _25144_ (_02044_, _10970_, _00697_);
  or _25145_ (_02045_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and _25146_ (_02046_, _02045_, _06983_);
  and _25147_ (_02047_, _02046_, _02044_);
  and _25148_ (_02048_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or _25149_ (_02049_, _02048_, rst);
  or _25150_ (_02050_, _02049_, _02047_);
  or _25151_ (_02933_, _02050_, _02043_);
  and _25152_ (_02051_, _00691_, _06979_);
  nand _25153_ (_02052_, _02051_, _06968_);
  or _25154_ (_02053_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and _25155_ (_02054_, _02053_, _06485_);
  and _25156_ (_02055_, _02054_, _02052_);
  nand _25157_ (_02057_, _09598_, _00697_);
  and _25158_ (_02059_, _02053_, _06983_);
  and _25159_ (_02060_, _02059_, _02057_);
  nor _25160_ (_02061_, _06484_, _01544_);
  or _25161_ (_02062_, _02061_, rst);
  or _25162_ (_02063_, _02062_, _02060_);
  or _25163_ (_02935_, _02063_, _02055_);
  or _25164_ (_02064_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and _25165_ (_02065_, _02064_, _06485_);
  and _25166_ (_02066_, _00720_, _06979_);
  nand _25167_ (_02067_, _02066_, _06968_);
  and _25168_ (_02068_, _02067_, _02065_);
  nand _25169_ (_02069_, _09598_, _00726_);
  and _25170_ (_02070_, _02064_, _06983_);
  and _25171_ (_02071_, _02070_, _02069_);
  nor _25172_ (_02072_, _06484_, _01539_);
  or _25173_ (_02073_, _02072_, rst);
  or _25174_ (_02074_, _02073_, _02071_);
  or _25175_ (_02937_, _02074_, _02068_);
  nand _25176_ (_02075_, _00720_, _06525_);
  and _25177_ (_02076_, _02075_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _25178_ (_02077_, _00764_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _25179_ (_02078_, _02077_, _08437_);
  and _25180_ (_02079_, _02078_, _00720_);
  or _25181_ (_02080_, _02079_, _02076_);
  and _25182_ (_02081_, _02080_, _06485_);
  nand _25183_ (_02082_, _00726_, _07317_);
  or _25184_ (_02083_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and _25185_ (_02084_, _02083_, _06983_);
  and _25186_ (_02085_, _02084_, _02082_);
  and _25187_ (_02086_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or _25188_ (_02087_, _02086_, rst);
  or _25189_ (_02088_, _02087_, _02085_);
  or _25190_ (_02939_, _02088_, _02081_);
  and _25191_ (_02089_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor _25192_ (_02090_, _08139_, _01144_);
  or _25193_ (_02091_, _02090_, _02089_);
  and _25194_ (_02962_, _02091_, _06989_);
  and _25195_ (_02092_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor _25196_ (_02093_, _08139_, _01149_);
  or _25197_ (_02094_, _02093_, _02092_);
  and _25198_ (_02965_, _02094_, _06989_);
  and _25199_ (_03047_, _01586_, _06989_);
  and _25200_ (_02095_, _00691_, _07048_);
  nand _25201_ (_02096_, _02095_, _06968_);
  or _25202_ (_02097_, _02095_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _25203_ (_02098_, _02097_, _06485_);
  and _25204_ (_02099_, _02098_, _02096_);
  nand _25205_ (_02101_, _00697_, _07118_);
  or _25206_ (_02102_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and _25207_ (_02103_, _02102_, _06983_);
  and _25208_ (_02104_, _02103_, _02101_);
  nor _25209_ (_02105_, _06484_, _01291_);
  or _25210_ (_02106_, _02105_, rst);
  or _25211_ (_02107_, _02106_, _02104_);
  or _25212_ (_03053_, _02107_, _02099_);
  and _25213_ (_02108_, _00691_, _07044_);
  nand _25214_ (_02109_, _02108_, _06968_);
  or _25215_ (_02110_, _02108_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _25216_ (_02111_, _02110_, _06485_);
  and _25217_ (_02112_, _02111_, _02109_);
  nand _25218_ (_02113_, _00697_, _07260_);
  or _25219_ (_02114_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and _25220_ (_02115_, _02114_, _06983_);
  and _25221_ (_02116_, _02115_, _02113_);
  nor _25222_ (_02117_, _06484_, _01455_);
  or _25223_ (_02118_, _02117_, rst);
  or _25224_ (_02119_, _02118_, _02116_);
  or _25225_ (_03055_, _02119_, _02112_);
  and _25226_ (_02120_, _09023_, _07044_);
  nand _25227_ (_02121_, _02120_, _06968_);
  or _25228_ (_02122_, _02120_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and _25229_ (_02123_, _02122_, _06485_);
  and _25230_ (_02124_, _02123_, _02121_);
  nor _25231_ (_02125_, _09031_, _07260_);
  nor _25232_ (_02126_, _09030_, _01471_);
  or _25233_ (_02127_, _02126_, _02125_);
  and _25234_ (_02128_, _02127_, _06983_);
  nor _25235_ (_02129_, _06484_, _01471_);
  or _25236_ (_02130_, _02129_, rst);
  or _25237_ (_02131_, _02130_, _02128_);
  or _25238_ (_03057_, _02131_, _02124_);
  and _25239_ (_02132_, _09023_, _08436_);
  nand _25240_ (_02133_, _02132_, _06968_);
  or _25241_ (_02134_, _02132_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and _25242_ (_02135_, _02134_, _06485_);
  and _25243_ (_02136_, _02135_, _02133_);
  nor _25244_ (_02137_, _09031_, _07317_);
  and _25245_ (_02138_, _09031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _25246_ (_02139_, _02138_, _02137_);
  and _25247_ (_02140_, _02139_, _06983_);
  and _25248_ (_02141_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or _25249_ (_02142_, _02141_, rst);
  or _25250_ (_02143_, _02142_, _02140_);
  or _25251_ (_03058_, _02143_, _02136_);
  nand _25252_ (_02144_, _12937_, _09598_);
  or _25253_ (_02145_, _12937_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and _25254_ (_02146_, _02145_, _02144_);
  and _25255_ (_03072_, _02146_, _06989_);
  and _25256_ (_02147_, _00720_, _14196_);
  nand _25257_ (_02148_, _02147_, _06968_);
  or _25258_ (_02149_, _02147_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _25259_ (_02150_, _02149_, _06485_);
  and _25260_ (_02151_, _02150_, _02148_);
  nand _25261_ (_02152_, _10970_, _00726_);
  or _25262_ (_02153_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and _25263_ (_02154_, _02153_, _06983_);
  and _25264_ (_02155_, _02154_, _02152_);
  and _25265_ (_02156_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or _25266_ (_02157_, _02156_, rst);
  or _25267_ (_02158_, _02157_, _02155_);
  or _25268_ (_03077_, _02158_, _02151_);
  and _25269_ (_02159_, _00720_, _07044_);
  nand _25270_ (_02160_, _02159_, _06968_);
  or _25271_ (_02161_, _02159_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _25272_ (_02162_, _02161_, _06485_);
  and _25273_ (_02163_, _02162_, _02160_);
  nand _25274_ (_02164_, _00726_, _07260_);
  or _25275_ (_02165_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and _25276_ (_02166_, _02165_, _06983_);
  and _25277_ (_02167_, _02166_, _02164_);
  nor _25278_ (_02168_, _06484_, _01460_);
  or _25279_ (_02169_, _02168_, rst);
  or _25280_ (_02170_, _02169_, _02167_);
  or _25281_ (_03079_, _02170_, _02163_);
  nand _25282_ (_02171_, _00720_, _00764_);
  and _25283_ (_02172_, _02171_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _25284_ (_02173_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or _25285_ (_02174_, _02173_, _00760_);
  and _25286_ (_02175_, _02174_, _00720_);
  or _25287_ (_02176_, _02175_, _02172_);
  and _25288_ (_02177_, _02176_, _06485_);
  nand _25289_ (_02178_, _11529_, _00726_);
  or _25290_ (_02179_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and _25291_ (_02180_, _02179_, _06983_);
  and _25292_ (_02181_, _02180_, _02178_);
  nor _25293_ (_02182_, _06484_, _14527_);
  or _25294_ (_02183_, _02182_, rst);
  or _25295_ (_02184_, _02183_, _02181_);
  or _25296_ (_03081_, _02184_, _02177_);
  and _25297_ (_02186_, _00691_, _08436_);
  nand _25298_ (_02187_, _02186_, _06968_);
  or _25299_ (_02188_, _02186_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _25300_ (_02189_, _02188_, _06485_);
  and _25301_ (_02190_, _02189_, _02187_);
  nand _25302_ (_02191_, _00697_, _07317_);
  or _25303_ (_02192_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and _25304_ (_02193_, _02192_, _06983_);
  and _25305_ (_02194_, _02193_, _02191_);
  and _25306_ (_02195_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or _25307_ (_02196_, _02195_, rst);
  or _25308_ (_02197_, _02196_, _02194_);
  or _25309_ (_03083_, _02197_, _02190_);
  and _25310_ (_02198_, _09023_, _14196_);
  nand _25311_ (_02199_, _02198_, _06968_);
  or _25312_ (_02200_, _02198_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and _25313_ (_02201_, _02200_, _06485_);
  and _25314_ (_02202_, _02201_, _02199_);
  nor _25315_ (_02203_, _10970_, _09031_);
  and _25316_ (_02204_, _09031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _25317_ (_02205_, _02204_, _02203_);
  and _25318_ (_02206_, _02205_, _06983_);
  and _25319_ (_02207_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or _25320_ (_02208_, _02207_, rst);
  or _25321_ (_02209_, _02208_, _02206_);
  or _25322_ (_03085_, _02209_, _02202_);
  and _25323_ (_02210_, _00691_, _07089_);
  nand _25324_ (_02211_, _02210_, _06968_);
  or _25325_ (_02213_, _02210_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _25326_ (_02214_, _02213_, _06485_);
  and _25327_ (_02215_, _02214_, _02211_);
  nand _25328_ (_02216_, _00697_, _09008_);
  or _25329_ (_02217_, _00697_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and _25330_ (_02218_, _02217_, _06983_);
  and _25331_ (_02219_, _02218_, _02216_);
  and _25332_ (_02220_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or _25333_ (_02221_, _02220_, rst);
  or _25334_ (_02222_, _02221_, _02219_);
  or _25335_ (_03087_, _02222_, _02215_);
  and _25336_ (_02223_, _09023_, _09074_);
  nand _25337_ (_02224_, _02223_, _06968_);
  or _25338_ (_02226_, _02223_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and _25339_ (_02227_, _02226_, _06485_);
  and _25340_ (_02228_, _02227_, _02224_);
  nor _25341_ (_02229_, _11529_, _09031_);
  and _25342_ (_02230_, _09031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _25343_ (_02231_, _02230_, _02229_);
  and _25344_ (_02232_, _02231_, _06983_);
  and _25345_ (_02233_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or _25346_ (_02234_, _02233_, rst);
  or _25347_ (_02235_, _02234_, _02232_);
  or _25348_ (_03089_, _02235_, _02228_);
  nand _25349_ (_02236_, _09030_, _06968_);
  or _25350_ (_02237_, _09030_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and _25351_ (_02238_, _02237_, _06485_);
  and _25352_ (_02239_, _02238_, _02236_);
  and _25353_ (_02240_, _09599_, _09030_);
  nor _25354_ (_02241_, _09030_, _01528_);
  or _25355_ (_02242_, _02241_, _02240_);
  and _25356_ (_02243_, _02242_, _06983_);
  nor _25357_ (_02244_, _06484_, _01528_);
  or _25358_ (_02245_, _02244_, rst);
  or _25359_ (_02246_, _02245_, _02243_);
  or _25360_ (_03091_, _02246_, _02239_);
  and _25361_ (_02247_, _01156_, _14196_);
  nand _25362_ (_02248_, _02247_, _06968_);
  or _25363_ (_02249_, _02247_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and _25364_ (_02250_, _02249_, _06485_);
  and _25365_ (_02251_, _02250_, _02248_);
  nor _25366_ (_02252_, _01163_, _10970_);
  and _25367_ (_02253_, _01163_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _25368_ (_02254_, _02253_, _02252_);
  and _25369_ (_02255_, _02254_, _06983_);
  and _25370_ (_02256_, _11804_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or _25371_ (_02257_, _02256_, rst);
  or _25372_ (_02258_, _02257_, _02255_);
  or _25373_ (_03093_, _02258_, _02251_);
  and _25374_ (_02259_, _01156_, _07044_);
  nand _25375_ (_02260_, _02259_, _06968_);
  or _25376_ (_02261_, _02259_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and _25377_ (_02262_, _02261_, _06485_);
  and _25378_ (_02263_, _02262_, _02260_);
  nor _25379_ (_02264_, _01163_, _07260_);
  nor _25380_ (_02265_, _01162_, _01466_);
  or _25381_ (_02266_, _02265_, _02264_);
  and _25382_ (_02267_, _02266_, _06983_);
  nor _25383_ (_02268_, _06484_, _01466_);
  or _25384_ (_02269_, _02268_, rst);
  or _25385_ (_02270_, _02269_, _02267_);
  or _25386_ (_03095_, _02270_, _02263_);
  and _25387_ (_02271_, _01156_, _09074_);
  nand _25388_ (_02272_, _02271_, _06968_);
  or _25389_ (_02273_, _02271_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and _25390_ (_02274_, _02273_, _06485_);
  and _25391_ (_02275_, _02274_, _02272_);
  nor _25392_ (_02276_, _01163_, _11529_);
  nor _25393_ (_02277_, _01162_, _14538_);
  or _25394_ (_02278_, _02277_, _02276_);
  and _25395_ (_02279_, _02278_, _06983_);
  nor _25396_ (_02280_, _06484_, _14538_);
  or _25397_ (_02281_, _02280_, rst);
  or _25398_ (_02282_, _02281_, _02279_);
  or _25399_ (_03098_, _02282_, _02275_);
  and _25400_ (_02283_, _11954_, _07048_);
  or _25401_ (_02285_, _02283_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _25402_ (_02287_, _02285_, _07292_);
  nand _25403_ (_02288_, _02283_, _06968_);
  and _25404_ (_02289_, _02288_, _02287_);
  nor _25405_ (_02290_, _07292_, _07118_);
  or _25406_ (_02291_, _02290_, _02289_);
  and _25407_ (_03127_, _02291_, _06989_);
  and _25408_ (_03135_, _01367_, _06989_);
  and _25409_ (_03420_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _06989_);
  and _25410_ (_02292_, _03420_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or _25411_ (_03146_, _02292_, _03135_);
  or _25412_ (_02293_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand _25413_ (_02295_, _07493_, _14110_);
  and _25414_ (_02296_, _02295_, _06989_);
  and _25415_ (_03150_, _02296_, _02293_);
  nand _25416_ (_02298_, _07321_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and _25417_ (_03156_, _02298_, _06989_);
  nand _25418_ (_02299_, _11951_, _06968_);
  nor _25419_ (_02301_, _11951_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor _25420_ (_02302_, _02301_, _11954_);
  and _25421_ (_02303_, _02302_, _02299_);
  or _25422_ (_02304_, _02303_, _07291_);
  and _25423_ (_02305_, _06540_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _25424_ (_02306_, _02305_, _06969_);
  and _25425_ (_02307_, _02306_, _11954_);
  or _25426_ (_02308_, _02307_, _02304_);
  nand _25427_ (_02309_, _07291_, _07040_);
  and _25428_ (_02310_, _02309_, _06989_);
  and _25429_ (_03209_, _02310_, _02308_);
  and _25430_ (_03313_, _08080_, _06989_);
  nor _25431_ (_02311_, _07493_, _07490_);
  nor _25432_ (_02312_, _01213_, _01210_);
  nor _25433_ (_02313_, _02312_, _07490_);
  and _25434_ (_02314_, _02313_, _07331_);
  nor _25435_ (_02315_, _02313_, _07331_);
  nor _25436_ (_02316_, _02315_, _02314_);
  nor _25437_ (_02317_, _02316_, _02311_);
  and _25438_ (_02318_, _07350_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand _25439_ (_02319_, _02318_, _02311_);
  nor _25440_ (_02320_, _02319_, _10959_);
  or _25441_ (_02321_, _02320_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _25442_ (_02322_, _02321_, _02317_);
  and _25443_ (_03315_, _02322_, _06989_);
  nor _25444_ (_02323_, _12938_, _07260_);
  and _25445_ (_02324_, _12945_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or _25446_ (_02325_, _02324_, _02323_);
  and _25447_ (_03327_, _02325_, _06989_);
  and _25448_ (_02326_, _12829_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or _25449_ (_02327_, _02326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and _25450_ (_03329_, _02327_, _06989_);
  nor _25451_ (_02328_, _12829_, rst);
  not _25452_ (_02329_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nand _25453_ (_02330_, _07325_, _02329_);
  and _25454_ (_03350_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _06989_);
  and _25455_ (_02331_, _03350_, _02330_);
  or _25456_ (_03331_, _02331_, _02328_);
  and _25457_ (_02332_, _14190_, _09599_);
  and _25458_ (_02333_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  or _25459_ (_02334_, _02333_, _02332_);
  and _25460_ (_03345_, _02334_, _06989_);
  and _25461_ (_02335_, _14146_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor _25462_ (_02336_, _14146_, _07260_);
  or _25463_ (_02337_, _02336_, _02335_);
  and _25464_ (_03354_, _02337_, _06989_);
  and _25465_ (_02338_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and _25466_ (_02339_, _14190_, _09009_);
  or _25467_ (_02340_, _02339_, _02338_);
  and _25468_ (_03364_, _02340_, _06989_);
  nor _25469_ (_02341_, _11042_, _11040_);
  nor _25470_ (_02342_, _02341_, _11043_);
  or _25471_ (_02343_, _02342_, _08477_);
  or _25472_ (_02344_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and _25473_ (_02345_, _02344_, _10964_);
  and _25474_ (_02346_, _02345_, _02343_);
  and _25475_ (_02347_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or _25476_ (_03372_, _02347_, _02346_);
  nor _25477_ (_02348_, _11037_, _11035_);
  nor _25478_ (_02349_, _02348_, _11038_);
  or _25479_ (_02350_, _02349_, _08477_);
  or _25480_ (_02351_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and _25481_ (_02352_, _02351_, _10964_);
  and _25482_ (_02353_, _02352_, _02350_);
  and _25483_ (_02354_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or _25484_ (_03374_, _02354_, _02353_);
  nor _25485_ (_02355_, _11034_, _11032_);
  nor _25486_ (_02356_, _02355_, _11035_);
  or _25487_ (_02357_, _02356_, _08477_);
  or _25488_ (_02358_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and _25489_ (_02359_, _02358_, _10964_);
  and _25490_ (_02360_, _02359_, _02357_);
  and _25491_ (_02361_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or _25492_ (_03399_, _02361_, _02360_);
  not _25493_ (_02362_, _00653_);
  and _25494_ (_02363_, _02362_, _00651_);
  and _25495_ (_02364_, _00256_, _00645_);
  and _25496_ (_03413_, _02364_, _02363_);
  nor _25497_ (_02365_, _13944_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor _25498_ (_02366_, _02365_, _13945_);
  and _25499_ (_03422_, _02366_, _13953_);
  and _25500_ (_02367_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _08578_);
  and _25501_ (_02368_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or _25502_ (_02369_, _02368_, _02367_);
  and _25503_ (_03428_, _02369_, _06989_);
  and _25504_ (_02370_, _14188_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and _25505_ (_02371_, _14190_, _07119_);
  or _25506_ (_02372_, _02371_, _02370_);
  and _25507_ (_03439_, _02372_, _06989_);
  and _25508_ (_02373_, _08525_, _08459_);
  and _25509_ (_02374_, _02373_, _08557_);
  not _25510_ (_02375_, _08542_);
  and _25511_ (_02376_, _02375_, _08509_);
  and _25512_ (_02377_, _02376_, _08572_);
  and _25513_ (_02378_, _07326_, _06989_);
  and _25514_ (_02379_, _02378_, _08492_);
  and _25515_ (_02380_, _02379_, _07356_);
  and _25516_ (_02381_, _02380_, _02377_);
  and _25517_ (_03444_, _02381_, _02374_);
  and _25518_ (_02382_, _07486_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nor _25519_ (_02383_, _10970_, _07486_);
  or _25520_ (_02384_, _02383_, _02382_);
  and _25521_ (_03447_, _02384_, _06989_);
  and _25522_ (_03456_, _11518_, _06989_);
  and _25523_ (_03475_, _11605_, _06989_);
  and _25524_ (_02385_, _14058_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and _25525_ (_02386_, _09763_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and _25526_ (_02387_, _02386_, _14057_);
  or _25527_ (_02388_, _02387_, _02385_);
  and _25528_ (_03479_, _02388_, _06989_);
  and _25529_ (_02389_, _07161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  or _25530_ (_02390_, _00909_, _07278_);
  nand _25531_ (_02391_, _07209_, _07166_);
  or _25532_ (_02392_, _02391_, _07196_);
  and _25533_ (_02393_, _02392_, _02390_);
  or _25534_ (_02394_, _02393_, _02389_);
  and _25535_ (_02395_, _07271_, _07269_);
  or _25536_ (_02396_, _02395_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor _25537_ (_02397_, _07470_, rst);
  and _25538_ (_02398_, _02397_, _02396_);
  and _25539_ (_03486_, _02398_, _02394_);
  or _25540_ (_02399_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  nand _25541_ (_02400_, _07493_, _11224_);
  and _25542_ (_02401_, _02400_, _06989_);
  and _25543_ (_03489_, _02401_, _02399_);
  and _25544_ (_02402_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and _25545_ (_02403_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or _25546_ (_02404_, _02403_, _02402_);
  and _25547_ (_03512_, _02404_, _06989_);
  and _25548_ (_02405_, _11908_, _11359_);
  and _25549_ (_02406_, _11911_, _11364_);
  and _25550_ (_02407_, _11359_, _11287_);
  or _25551_ (_02408_, _02407_, _02406_);
  and _25552_ (_02409_, _11911_, _11306_);
  or _25553_ (_02410_, _02409_, _11405_);
  or _25554_ (_02411_, _02410_, _02408_);
  or _25555_ (_02412_, _02411_, _02405_);
  and _25556_ (_02413_, _11339_, _11313_);
  and _25557_ (_02414_, _11332_, _11430_);
  or _25558_ (_02415_, _02414_, _11435_);
  or _25559_ (_02416_, _02415_, _02413_);
  or _25560_ (_02417_, _11332_, _11478_);
  and _25561_ (_02418_, _02417_, _11389_);
  and _25562_ (_02419_, _11354_, _11290_);
  or _25563_ (_02420_, _02419_, _02418_);
  or _25564_ (_02421_, _02420_, _02416_);
  and _25565_ (_02422_, _11908_, _11451_);
  and _25566_ (_02423_, _11908_, _11313_);
  or _25567_ (_02424_, _02423_, _02422_);
  or _25568_ (_02425_, _02424_, _11385_);
  and _25569_ (_02426_, _11430_, _11287_);
  or _25570_ (_02427_, _02426_, _11468_);
  or _25571_ (_02428_, _02427_, _11404_);
  or _25572_ (_02429_, _02428_, _02425_);
  or _25573_ (_02430_, _02429_, _02421_);
  and _25574_ (_02431_, _11332_, _11472_);
  and _25575_ (_02432_, _11332_, _11356_);
  and _25576_ (_02433_, _11332_, _11375_);
  or _25577_ (_02434_, _02433_, _02432_);
  or _25578_ (_02435_, _02434_, _02431_);
  or _25579_ (_02436_, _14313_, _11320_);
  and _25580_ (_02437_, _11332_, _11324_);
  or _25581_ (_02438_, _02437_, _14317_);
  not _25582_ (_02439_, _11397_);
  nand _25583_ (_02440_, _02439_, _11391_);
  or _25584_ (_02441_, _02440_, _02438_);
  or _25585_ (_02442_, _02441_, _02436_);
  or _25586_ (_02443_, _02442_, _02435_);
  or _25587_ (_02444_, _02443_, _02430_);
  or _25588_ (_02445_, _02444_, _02412_);
  and _25589_ (_02446_, _02445_, _07325_);
  and _25590_ (_02447_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not _25591_ (_02448_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and _25592_ (_02449_, _11353_, _02448_);
  and _25593_ (_02450_, _11290_, _11306_);
  not _25594_ (_02451_, _11467_);
  nor _25595_ (_02452_, _11339_, _11289_);
  nor _25596_ (_02453_, _02452_, _02451_);
  nor _25597_ (_02454_, _02453_, _02450_);
  not _25598_ (_02455_, _02454_);
  and _25599_ (_02456_, _02455_, _02449_);
  or _25600_ (_02457_, _02456_, _02447_);
  or _25601_ (_02458_, _02457_, _02446_);
  and _25602_ (_03518_, _02458_, _06989_);
  and _25603_ (_02459_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and _25604_ (_02460_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  or _25605_ (_02461_, _02460_, _02459_);
  and _25606_ (_03521_, _02461_, _06989_);
  nor _25607_ (_03539_, _11579_, rst);
  and _25608_ (_02462_, \oc8051_top_1.oc8051_sfr1.wait_data , _06989_);
  and _25609_ (_02463_, _02462_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and _25610_ (_02464_, _02422_, _07383_);
  and _25611_ (_02465_, _11925_, _11382_);
  or _25612_ (_02466_, _02465_, _02464_);
  and _25613_ (_02467_, _11478_, _11373_);
  or _25614_ (_02468_, _02467_, _14317_);
  or _25615_ (_02469_, _11467_, _11359_);
  and _25616_ (_02470_, _02469_, _11332_);
  or _25617_ (_02471_, _02470_, _02468_);
  or _25618_ (_02472_, _02471_, _02466_);
  or _25619_ (_02473_, _14320_, _11395_);
  and _25620_ (_02474_, _02450_, _11316_);
  or _25621_ (_02475_, _02474_, _02473_);
  and _25622_ (_02476_, _14313_, _07383_);
  and _25623_ (_02477_, _02423_, _07383_);
  or _25624_ (_02478_, _02477_, _02476_);
  or _25625_ (_02479_, _02478_, _02475_);
  and _25626_ (_02480_, _11332_, _11399_);
  or _25627_ (_02481_, _11919_, _02480_);
  nor _25628_ (_02482_, _02481_, _11400_);
  nand _25629_ (_02483_, _02482_, _11454_);
  or _25630_ (_02484_, _02483_, _02416_);
  or _25631_ (_02485_, _02484_, _02479_);
  or _25632_ (_02486_, _02485_, _02472_);
  and _25633_ (_02487_, _07325_, _06989_);
  and _25634_ (_02488_, _02487_, _02486_);
  or _25635_ (_03541_, _02488_, _02463_);
  nor _25636_ (_03549_, _07294_, rst);
  and _25637_ (_02489_, _11358_, _11342_);
  not _25638_ (_02490_, _11335_);
  and _25639_ (_02491_, _02490_, _02449_);
  and _25640_ (_02492_, _11941_, _11312_);
  and _25641_ (_02493_, _11940_, _11312_);
  or _25642_ (_02494_, _02493_, _02492_);
  and _25643_ (_02495_, _02494_, _11342_);
  or _25644_ (_02496_, _02495_, _02491_);
  or _25645_ (_02497_, _02496_, _02489_);
  and _25646_ (_02498_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _25647_ (_02499_, _11478_, _11306_);
  or _25648_ (_02500_, _02499_, _11456_);
  and _25649_ (_02501_, _11925_, _11289_);
  or _25650_ (_02502_, _02501_, _11449_);
  or _25651_ (_02503_, _11473_, _11425_);
  or _25652_ (_02504_, _02503_, _02492_);
  or _25653_ (_02505_, _02504_, _02502_);
  and _25654_ (_02506_, _11469_, _11388_);
  or _25655_ (_02507_, _11461_, _11453_);
  or _25656_ (_02508_, _02507_, _02506_);
  nor _25657_ (_02509_, _11477_, _11423_);
  nand _25658_ (_02510_, _02509_, _11440_);
  or _25659_ (_02511_, _02510_, _02508_);
  or _25660_ (_02512_, _02511_, _02505_);
  or _25661_ (_02513_, _02493_, _11380_);
  or _25662_ (_02514_, _02513_, _02512_);
  or _25663_ (_02515_, _02514_, _02500_);
  and _25664_ (_02516_, _02515_, _07325_);
  or _25665_ (_02517_, _02516_, _02498_);
  or _25666_ (_02518_, _02517_, _02497_);
  and _25667_ (_03557_, _02518_, _06989_);
  and _25668_ (_02519_, _06894_, _06845_);
  and _25669_ (_02520_, _06790_, _06548_);
  and _25670_ (_02521_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  nand _25671_ (_02522_, _06951_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand _25672_ (_02523_, _02522_, _02521_);
  or _25673_ (_02524_, _02523_, _02520_);
  or _25674_ (_02525_, _02524_, _02519_);
  nor _25675_ (_02526_, _02521_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor _25676_ (_02527_, _02526_, _11954_);
  and _25677_ (_02528_, _02527_, _02525_);
  or _25678_ (_02529_, _02528_, _07291_);
  nor _25679_ (_02530_, _14196_, _08412_);
  or _25680_ (_02531_, _02530_, _01556_);
  and _25681_ (_02532_, _02531_, _11954_);
  or _25682_ (_02533_, _02532_, _02529_);
  nand _25683_ (_02534_, _10970_, _07291_);
  and _25684_ (_02535_, _02534_, _06989_);
  and _25685_ (_03561_, _02535_, _02533_);
  and _25686_ (_02536_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25687_ (_02537_, _02536_, _02496_);
  nor _25688_ (_02538_, _11942_, _11316_);
  and _25689_ (_02539_, _11477_, _11316_);
  and _25690_ (_02540_, _11394_, _11319_);
  and _25691_ (_02541_, _11396_, _11388_);
  or _25692_ (_02543_, _02541_, _11401_);
  or _25693_ (_02544_, _02543_, _02540_);
  or _25694_ (_02545_, _02544_, _02539_);
  or _25695_ (_02546_, _02545_, _11395_);
  or _25696_ (_02547_, _02546_, _02538_);
  and _25697_ (_02548_, _02547_, _07325_);
  or _25698_ (_02549_, _02548_, _02537_);
  and _25699_ (_03566_, _02549_, _06989_);
  and _25700_ (_02550_, _11332_, _11451_);
  or _25701_ (_02551_, _02550_, _02414_);
  or _25702_ (_02552_, _02408_, _02419_);
  and _25703_ (_02553_, _11389_, _11312_);
  and _25704_ (_02554_, _02553_, _11422_);
  or _25705_ (_02555_, _02541_, _02493_);
  or _25706_ (_02556_, _02555_, _02554_);
  and _25707_ (_02557_, _11403_, _11382_);
  or _25708_ (_02558_, _02437_, _02557_);
  or _25709_ (_02559_, _02558_, _02556_);
  or _25710_ (_02560_, _02559_, _02552_);
  or _25711_ (_02561_, _02560_, _02551_);
  or _25712_ (_02562_, _02410_, _11404_);
  and _25713_ (_02564_, _11911_, _11388_);
  or _25714_ (_02565_, _11397_, _11325_);
  or _25715_ (_02566_, _02565_, _02564_);
  and _25716_ (_02567_, _11356_, _11382_);
  and _25717_ (_02568_, _11908_, _11927_);
  or _25718_ (_02569_, _02568_, _02567_);
  or _25719_ (_02570_, _02569_, _02566_);
  or _25720_ (_02571_, _02570_, _02562_);
  or _25721_ (_02572_, _02571_, _02561_);
  and _25722_ (_02573_, _11332_, _11438_);
  or _25723_ (_02574_, _02573_, _02423_);
  and _25724_ (_02575_, _11359_, _11312_);
  and _25725_ (_02577_, _02575_, _11908_);
  or _25726_ (_02579_, _02577_, _14313_);
  or _25727_ (_02580_, _02579_, _02574_);
  and _25728_ (_02581_, _11332_, _11467_);
  or _25729_ (_02582_, _02581_, _11909_);
  and _25730_ (_02583_, _02553_, _11332_);
  or _25731_ (_02584_, _02583_, _11333_);
  or _25732_ (_02585_, _02584_, _02582_);
  or _25733_ (_02586_, _02585_, _02435_);
  or _25734_ (_02587_, _02450_, _11334_);
  or _25735_ (_02588_, _02587_, _02586_);
  or _25736_ (_02589_, _02588_, _02580_);
  or _25737_ (_02590_, _02589_, _02572_);
  and _25738_ (_02591_, _02590_, _07325_);
  and _25739_ (_02592_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or _25740_ (_02593_, _02456_, _11347_);
  or _25741_ (_02594_, _02593_, _02592_);
  or _25742_ (_02595_, _02594_, _02591_);
  and _25743_ (_03579_, _02595_, _06989_);
  or _25744_ (_02596_, _02553_, _11324_);
  and _25745_ (_02598_, _02596_, _11422_);
  or _25746_ (_02599_, _02565_, _02598_);
  and _25747_ (_02600_, _11451_, _11290_);
  and _25748_ (_02601_, _11430_, _11290_);
  or _25749_ (_02602_, _02601_, _02600_);
  or _25750_ (_02603_, _02602_, _11456_);
  or _25751_ (_02604_, _02603_, _02599_);
  and _25752_ (_02605_, _02541_, _11299_);
  or _25753_ (_02606_, _02605_, _02413_);
  and _25754_ (_02607_, _02553_, _11287_);
  or _25755_ (_02608_, _02607_, _02606_);
  or _25756_ (_02609_, _11334_, _11314_);
  or _25757_ (_02610_, _02609_, _02562_);
  or _25758_ (_02611_, _02610_, _02608_);
  or _25759_ (_02612_, _02611_, _02604_);
  or _25760_ (_02613_, _02574_, _11447_);
  or _25761_ (_02614_, _02613_, _02586_);
  or _25762_ (_02615_, _02614_, _02612_);
  or _25763_ (_02616_, _02615_, _02552_);
  and _25764_ (_02617_, _02616_, _07325_);
  and _25765_ (_02618_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or _25766_ (_02619_, _02618_, _02593_);
  or _25767_ (_02620_, _02619_, _02617_);
  and _25768_ (_03598_, _02620_, _06989_);
  nand _25769_ (_02621_, _01555_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand _25770_ (_02623_, _02621_, _06501_);
  or _25771_ (_02624_, _02623_, _01556_);
  not _25772_ (_02625_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and _25773_ (_02626_, _07075_, _02625_);
  or _25774_ (_02627_, _02626_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _25775_ (_02628_, _02627_, _06501_);
  and _25776_ (_02629_, _02628_, _02624_);
  or _25777_ (_02630_, _02629_, _06987_);
  nand _25778_ (_02631_, _10970_, _06987_);
  and _25779_ (_02632_, _02631_, _06989_);
  and _25780_ (_03617_, _02632_, _02630_);
  and _25781_ (_02633_, _07048_, _06501_);
  nand _25782_ (_02634_, _02633_, _06968_);
  not _25783_ (_02635_, _06987_);
  or _25784_ (_02636_, _02633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and _25785_ (_02637_, _02636_, _02635_);
  and _25786_ (_02638_, _02637_, _02634_);
  nor _25787_ (_02639_, _07118_, _02635_);
  or _25788_ (_02640_, _02639_, _02638_);
  and _25789_ (_03619_, _02640_, _06989_);
  and _25790_ (_02641_, _07044_, _06501_);
  nand _25791_ (_02642_, _02641_, _06968_);
  or _25792_ (_02643_, _02641_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and _25793_ (_02644_, _02643_, _02635_);
  and _25794_ (_02645_, _02644_, _02642_);
  nor _25795_ (_02646_, _07260_, _02635_);
  or _25796_ (_02647_, _02646_, _02645_);
  and _25797_ (_03622_, _02647_, _06989_);
  nor _25798_ (_03634_, _11349_, rst);
  nand _25799_ (_02648_, _02487_, _11389_);
  or _25800_ (_03636_, _02648_, _02452_);
  and _25801_ (_02649_, _10851_, _10812_);
  and _25802_ (_02651_, _10841_, _10834_);
  and _25803_ (_02652_, _10824_, _10854_);
  and _25804_ (_02653_, _10917_, _02652_);
  or _25805_ (_02654_, _02653_, _02651_);
  or _25806_ (_02655_, _02654_, _02649_);
  or _25807_ (_02656_, _10904_, _10860_);
  and _25808_ (_02657_, _10917_, _10818_);
  and _25809_ (_02658_, _10870_, _10851_);
  or _25810_ (_02659_, _02658_, _02657_);
  or _25811_ (_02660_, _02659_, _02656_);
  nor _25812_ (_02661_, _02660_, _02655_);
  nand _25813_ (_02662_, _02661_, _10941_);
  and _25814_ (_02663_, _10871_, _10837_);
  not _25815_ (_02664_, _10906_);
  nand _25816_ (_02665_, _10951_, _02664_);
  or _25817_ (_02666_, _02665_, _02663_);
  or _25818_ (_02667_, _10912_, _10831_);
  or _25819_ (_02669_, _10828_, _10816_);
  or _25820_ (_02670_, _02669_, _02667_);
  or _25821_ (_02672_, _10911_, _10878_);
  or _25822_ (_02673_, _02672_, _02670_);
  or _25823_ (_02674_, _02673_, _02666_);
  or _25824_ (_02675_, _02674_, _02662_);
  and _25825_ (_02676_, _02675_, _07326_);
  and _25826_ (_02678_, _07323_, _06406_);
  and _25827_ (_02679_, _02678_, _11340_);
  nor _25828_ (_02681_, _02679_, _02448_);
  or _25829_ (_02682_, _02681_, rst);
  or _25830_ (_03638_, _02682_, _02676_);
  or _25831_ (_02685_, _08463_, _11345_);
  or _25832_ (_02686_, _07324_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and _25833_ (_02687_, _02686_, _06989_);
  and _25834_ (_03641_, _02687_, _02685_);
  and _25835_ (_02688_, _02462_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and _25836_ (_02690_, _11375_, _11289_);
  and _25837_ (_02691_, _11438_, _11290_);
  or _25838_ (_02693_, _02691_, _02581_);
  or _25839_ (_02694_, _02693_, _02690_);
  or _25840_ (_02696_, _11439_, _11369_);
  and _25841_ (_02697_, _11360_, _11316_);
  or _25842_ (_02699_, _11936_, _02697_);
  or _25843_ (_02700_, _02699_, _02696_);
  or _25844_ (_02701_, _11913_, _11358_);
  or _25845_ (_02702_, _02701_, _02474_);
  or _25846_ (_02704_, _02702_, _02700_);
  or _25847_ (_02706_, _02704_, _02694_);
  and _25848_ (_02707_, _02706_, _02487_);
  or _25849_ (_03643_, _02707_, _02688_);
  or _25850_ (_02708_, _02413_, _11320_);
  and _25851_ (_02709_, _11908_, _11438_);
  and _25852_ (_02710_, _11478_, _11374_);
  or _25853_ (_02711_, _02710_, _11395_);
  or _25854_ (_02712_, _02711_, _02709_);
  or _25855_ (_02713_, _02712_, _02708_);
  and _25856_ (_02714_, _02713_, _07325_);
  and _25857_ (_02715_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25858_ (_02716_, _02715_, _02491_);
  or _25859_ (_02717_, _02716_, _02714_);
  and _25860_ (_03645_, _02717_, _06989_);
  and _25861_ (_02718_, _02462_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and _25862_ (_02719_, _11908_, _11356_);
  or _25863_ (_02720_, _02503_, _02431_);
  or _25864_ (_02721_, _02720_, _02719_);
  not _25865_ (_02722_, _11402_);
  and _25866_ (_02724_, _11355_, _11287_);
  or _25867_ (_02725_, _02724_, _11912_);
  or _25868_ (_02726_, _02725_, _02722_);
  or _25869_ (_02727_, _02481_, _02477_);
  or _25870_ (_02728_, _02727_, _02708_);
  or _25871_ (_02729_, _02728_, _02726_);
  or _25872_ (_02730_, _02729_, _02721_);
  and _25873_ (_02731_, _02730_, _02487_);
  or _25874_ (_03648_, _02731_, _02718_);
  or _25875_ (_02732_, _11052_, _11014_);
  and _25876_ (_02733_, _02732_, _11053_);
  or _25877_ (_02734_, _02733_, _08477_);
  or _25878_ (_02735_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and _25879_ (_02736_, _02735_, _10964_);
  and _25880_ (_02738_, _02736_, _02734_);
  and _25881_ (_02739_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or _25882_ (_03651_, _02739_, _02738_);
  and _25883_ (_02740_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _25884_ (_02741_, _11461_, _07325_);
  or _25885_ (_02742_, _02741_, _02740_);
  or _25886_ (_02743_, _02742_, _02491_);
  and _25887_ (_03655_, _02743_, _06989_);
  or _25888_ (_02744_, _02494_, _02474_);
  and _25889_ (_02745_, _02744_, _11282_);
  or _25890_ (_02746_, _02456_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25891_ (_02747_, _02746_, _02495_);
  or _25892_ (_02748_, _02747_, _02745_);
  or _25893_ (_02749_, _06406_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and _25894_ (_02750_, _02749_, _06989_);
  and _25895_ (_03657_, _02750_, _02748_);
  and _25896_ (_02751_, _02462_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or _25897_ (_02752_, _11355_, _11374_);
  and _25898_ (_02753_, _02752_, _11911_);
  or _25899_ (_02754_, _11425_, _11320_);
  or _25900_ (_02755_, _02754_, _02753_);
  or _25901_ (_02757_, _02690_, _02719_);
  and _25902_ (_02758_, _11438_, _11394_);
  and _25903_ (_02760_, _11356_, _11394_);
  or _25904_ (_02761_, _02760_, _02758_);
  or _25905_ (_02762_, _02761_, _02757_);
  or _25906_ (_02763_, _02710_, _11437_);
  or _25907_ (_02764_, _11474_, _11453_);
  or _25908_ (_02765_, _02764_, _02763_);
  or _25909_ (_02766_, _02765_, _02762_);
  or _25910_ (_02767_, _02766_, _02755_);
  and _25911_ (_02768_, _02767_, _02487_);
  or _25912_ (_03659_, _02768_, _02751_);
  and _25913_ (_02769_, _02462_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  not _25914_ (_02770_, _11432_);
  or _25915_ (_02771_, _02414_, _02770_);
  or _25916_ (_02772_, _02709_, _02422_);
  or _25917_ (_02773_, _02419_, _11426_);
  or _25918_ (_02774_, _02773_, _02772_);
  nand _25919_ (_02775_, _14306_, _11436_);
  or _25920_ (_02776_, _02775_, _02774_);
  or _25921_ (_02777_, _02776_, _02771_);
  or _25922_ (_02778_, _02473_, _02468_);
  or _25923_ (_02779_, _02778_, _02725_);
  or _25924_ (_02780_, _02779_, _02721_);
  or _25925_ (_02781_, _02780_, _02777_);
  and _25926_ (_02782_, _02781_, _02487_);
  or _25927_ (_03662_, _02782_, _02769_);
  or _25928_ (_02783_, _02405_, _02407_);
  or _25929_ (_02784_, _02410_, _11397_);
  or _25930_ (_02785_, _02784_, _02783_);
  or _25931_ (_02786_, _02785_, _02423_);
  and _25932_ (_02787_, _02786_, _07325_);
  and _25933_ (_02788_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25934_ (_02789_, _02788_, _11346_);
  or _25935_ (_02790_, _02789_, _02787_);
  and _25936_ (_03664_, _02790_, _06989_);
  or _25937_ (_02791_, _11456_, _11380_);
  or _25938_ (_02792_, _02725_, _02711_);
  or _25939_ (_02793_, _02493_, _11479_);
  or _25940_ (_02794_, _02793_, _02564_);
  or _25941_ (_02795_, _02794_, _02792_);
  or _25942_ (_02796_, _02795_, _02791_);
  or _25943_ (_02797_, _02796_, _02512_);
  or _25944_ (_02798_, _02797_, _02544_);
  and _25945_ (_02799_, _02798_, _07325_);
  and _25946_ (_02800_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or _25947_ (_02801_, _02800_, _02497_);
  or _25948_ (_02802_, _02801_, _02799_);
  and _25949_ (_03666_, _02802_, _06989_);
  and _25950_ (_02803_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _25951_ (_02804_, _02803_, _09580_);
  and _25952_ (_02806_, _07071_, _07054_);
  or _25953_ (_02807_, _02806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand _25954_ (_02808_, _07071_, _07055_);
  and _25955_ (_02809_, _02808_, _02807_);
  or _25956_ (_02810_, _02809_, _02804_);
  and _25957_ (_02811_, _02810_, _09574_);
  and _25958_ (_02812_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _25959_ (_02813_, _02812_, _07046_);
  or _25960_ (_02814_, _02813_, _02811_);
  nand _25961_ (_02815_, _07260_, _07046_);
  and _25962_ (_02816_, _02815_, _09590_);
  and _25963_ (_02817_, _02816_, _02814_);
  and _25964_ (_02818_, _07050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _25965_ (_02819_, _02818_, _02817_);
  and _25966_ (_03669_, _02819_, _06989_);
  and _25967_ (_02820_, _07071_, _07053_);
  nor _25968_ (_02821_, _02820_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor _25969_ (_02822_, _02821_, _02806_);
  and _25970_ (_02823_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _25971_ (_02824_, _02823_, _09580_);
  or _25972_ (_02825_, _02824_, _02822_);
  and _25973_ (_02826_, _02825_, _09574_);
  and _25974_ (_02827_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _25975_ (_02828_, _02827_, _07046_);
  or _25976_ (_02829_, _02828_, _02826_);
  nand _25977_ (_02830_, _07317_, _07046_);
  and _25978_ (_02831_, _02830_, _09590_);
  and _25979_ (_02832_, _02831_, _02829_);
  and _25980_ (_02833_, _07050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _25981_ (_02834_, _02833_, _02832_);
  and _25982_ (_03672_, _02834_, _06989_);
  and _25983_ (_02835_, _07071_, _07052_);
  nor _25984_ (_02836_, _02835_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor _25985_ (_02837_, _02836_, _02820_);
  and _25986_ (_02838_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _25987_ (_02839_, _02838_, _09580_);
  or _25988_ (_02840_, _02839_, _02837_);
  and _25989_ (_02841_, _02840_, _09574_);
  and _25990_ (_02842_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _25991_ (_02843_, _02842_, _07046_);
  or _25992_ (_02844_, _02843_, _02841_);
  nand _25993_ (_02845_, _11529_, _07046_);
  and _25994_ (_02846_, _02845_, _09590_);
  and _25995_ (_02847_, _02846_, _02844_);
  and _25996_ (_02848_, _07050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _25997_ (_02849_, _02848_, _02847_);
  and _25998_ (_03675_, _02849_, _06989_);
  and _25999_ (_02850_, _07071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor _26000_ (_02851_, _02850_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor _26001_ (_02852_, _02851_, _02835_);
  and _26002_ (_02853_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and _26003_ (_02854_, _02853_, _09580_);
  or _26004_ (_02855_, _02854_, _02852_);
  and _26005_ (_02856_, _02855_, _09574_);
  and _26006_ (_02857_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _26007_ (_02858_, _02857_, _07046_);
  or _26008_ (_02859_, _02858_, _02856_);
  nand _26009_ (_02860_, _09008_, _07046_);
  and _26010_ (_02861_, _02860_, _09590_);
  and _26011_ (_02862_, _02861_, _02859_);
  and _26012_ (_02863_, _07050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or _26013_ (_02864_, _02863_, _02862_);
  and _26014_ (_03679_, _02864_, _06989_);
  or _26015_ (_02865_, _11051_, _11018_);
  nor _26016_ (_02866_, _11052_, _08477_);
  and _26017_ (_02867_, _02866_, _02865_);
  nor _26018_ (_02868_, _08476_, _06798_);
  or _26019_ (_02869_, _02868_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or _26020_ (_02870_, _02869_, _02867_);
  or _26021_ (_02871_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _02329_);
  and _26022_ (_02872_, _02871_, _06989_);
  and _26023_ (_03682_, _02872_, _02870_);
  or _26024_ (_02873_, _01319_, _08123_);
  not _26025_ (_02874_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand _26026_ (_02875_, _01319_, _02874_);
  and _26027_ (_02876_, _02875_, _06983_);
  and _26028_ (_02877_, _02876_, _02873_);
  nor _26029_ (_02878_, _06484_, _02874_);
  or _26030_ (_02879_, _01319_, _08126_);
  and _26031_ (_02880_, _02875_, _06485_);
  and _26032_ (_02881_, _02880_, _02879_);
  or _26033_ (_02882_, _02881_, _02878_);
  or _26034_ (_02883_, _02882_, _02877_);
  and _26035_ (_03687_, _02883_, _06989_);
  not _26036_ (_02884_, _02487_);
  or _26037_ (_03693_, _02884_, _02454_);
  and _26038_ (_02885_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand _26039_ (_02886_, _02885_, _07066_);
  nand _26040_ (_02887_, _02886_, _02850_);
  or _26041_ (_02888_, _07071_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _26042_ (_02889_, _02888_, _09574_);
  and _26043_ (_02890_, _02889_, _02887_);
  and _26044_ (_02891_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _26045_ (_02892_, _02891_, _07046_);
  or _26046_ (_02893_, _02892_, _02890_);
  nand _26047_ (_02894_, _09598_, _07046_);
  and _26048_ (_02895_, _02894_, _02893_);
  or _26049_ (_02896_, _02895_, _07050_);
  or _26050_ (_02897_, _09590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _26051_ (_02898_, _02897_, _06989_);
  and _26052_ (_03698_, _02898_, _02896_);
  or _26053_ (_02901_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand _26054_ (_02902_, _07493_, _14007_);
  and _26055_ (_02904_, _02902_, _06989_);
  and _26056_ (_03706_, _02904_, _02901_);
  or _26057_ (_02906_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand _26058_ (_02908_, _07493_, _14020_);
  and _26059_ (_02910_, _02908_, _06989_);
  and _26060_ (_03712_, _02910_, _02906_);
  and _26061_ (_02912_, _11389_, _11339_);
  nor _26062_ (_02913_, _02912_, _02450_);
  or _26063_ (_03715_, _02913_, _02884_);
  and _26064_ (_02914_, _02462_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or _26065_ (_02915_, _11433_, _11429_);
  or _26066_ (_02916_, _11455_, _11426_);
  or _26067_ (_02917_, _02916_, _02915_);
  and _26068_ (_02918_, _02407_, _11312_);
  and _26069_ (_02919_, _11399_, _11290_);
  and _26070_ (_02920_, _11405_, _11312_);
  or _26071_ (_02921_, _02920_, _02919_);
  or _26072_ (_02923_, _02921_, _02918_);
  or _26073_ (_02924_, _02923_, _02755_);
  or _26074_ (_02925_, _02924_, _02917_);
  or _26075_ (_02926_, _02434_, _11423_);
  and _26076_ (_02927_, _02752_, _11934_);
  or _26077_ (_02929_, _02710_, _02409_);
  and _26078_ (_02931_, _11359_, _11934_);
  or _26079_ (_02932_, _02931_, _02929_);
  or _26080_ (_02934_, _02932_, _02927_);
  and _26081_ (_02936_, _02405_, _11312_);
  or _26082_ (_02938_, _02936_, _02423_);
  or _26083_ (_02940_, _02938_, _02761_);
  and _26084_ (_02941_, _11394_, _11313_);
  or _26085_ (_02942_, _11453_, _02941_);
  or _26086_ (_02943_, _02942_, _11449_);
  or _26087_ (_02944_, _02943_, _02940_);
  or _26088_ (_02945_, _02944_, _02934_);
  or _26089_ (_02946_, _02945_, _02926_);
  or _26090_ (_02947_, _02946_, _02925_);
  and _26091_ (_02948_, _02947_, _02487_);
  or _26092_ (_03719_, _02948_, _02914_);
  or _26093_ (_02949_, _02663_, _02651_);
  or _26094_ (_02950_, _02653_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or _26095_ (_02951_, _02950_, _02949_);
  and _26096_ (_02952_, _02951_, _02679_);
  nor _26097_ (_02953_, _02678_, _11340_);
  or _26098_ (_02954_, _02953_, rst);
  or _26099_ (_03721_, _02954_, _02952_);
  nor _26100_ (_02955_, _11050_, _11022_);
  nor _26101_ (_02956_, _02955_, _11051_);
  or _26102_ (_02957_, _02956_, _08477_);
  or _26103_ (_02958_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and _26104_ (_02959_, _02958_, _10964_);
  and _26105_ (_02960_, _02959_, _02957_);
  and _26106_ (_02961_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or _26107_ (_03723_, _02961_, _02960_);
  and _26108_ (_02963_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  not _26109_ (_02964_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor _26110_ (_02966_, _01637_, _02964_);
  and _26111_ (_02967_, _01637_, _02964_);
  nor _26112_ (_02968_, _02967_, _02966_);
  and _26113_ (_02969_, _02968_, _01647_);
  nor _26114_ (_02970_, _02968_, _01647_);
  or _26115_ (_02971_, _02970_, _02969_);
  or _26116_ (_02972_, _02971_, _08477_);
  or _26117_ (_02973_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _26118_ (_02974_, _02973_, _10964_);
  and _26119_ (_02975_, _02974_, _02972_);
  or _26120_ (_03726_, _02975_, _02963_);
  and _26121_ (_02976_, _12716_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _26122_ (_02977_, _02976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand _26123_ (_02978_, _02977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or _26124_ (_02979_, _02977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _26125_ (_02980_, _02979_, _02978_);
  or _26126_ (_02981_, _02980_, _11964_);
  and _26127_ (_02982_, _02981_, _06989_);
  and _26128_ (_02983_, _12278_, _11413_);
  and _26129_ (_02984_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and _26130_ (_02985_, _11974_, _11608_);
  or _26131_ (_02986_, _02985_, _02984_);
  and _26132_ (_02987_, _12314_, _11968_);
  or _26133_ (_02988_, _02987_, _02986_);
  or _26134_ (_02989_, _02988_, _02983_);
  or _26135_ (_02990_, _12751_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or _26136_ (_02991_, _02990_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or _26137_ (_02992_, _02991_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _26138_ (_02993_, _02992_, _12742_);
  or _26139_ (_02994_, _12757_, _08182_);
  nor _26140_ (_02995_, _02994_, _08187_);
  nand _26141_ (_02996_, _02995_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _26142_ (_02997_, _02996_, _12753_);
  nand _26143_ (_02998_, _02997_, _02993_);
  nand _26144_ (_02999_, _02998_, _12303_);
  or _26145_ (_03000_, _02998_, _12303_);
  and _26146_ (_03001_, _03000_, _02999_);
  and _26147_ (_03002_, _03001_, _12722_);
  or _26148_ (_03003_, _03002_, _02989_);
  and _26149_ (_03004_, _12793_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and _26150_ (_03005_, _03004_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or _26151_ (_03006_, _03005_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand _26152_ (_03007_, _03005_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and _26153_ (_03008_, _03007_, _03006_);
  and _26154_ (_03009_, _03008_, _12783_);
  or _26155_ (_03010_, _03009_, _12781_);
  or _26156_ (_03011_, _03010_, _03003_);
  and _26157_ (_03742_, _03011_, _02982_);
  and _26158_ (_03755_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _06989_);
  nor _26159_ (_03758_, _12156_, rst);
  nand _26160_ (_03012_, _10970_, _09531_);
  not _26161_ (_03013_, _09537_);
  and _26162_ (_03014_, _03013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _26163_ (_03015_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or _26164_ (_03016_, _03015_, _03014_);
  or _26165_ (_03017_, _03016_, _09531_);
  and _26166_ (_03018_, _03017_, _06989_);
  and _26167_ (_03761_, _03018_, _03012_);
  nand _26168_ (_03019_, _10146_, _09598_);
  or _26169_ (_03020_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and _26170_ (_03021_, _03020_, _06989_);
  and _26171_ (_03764_, _03021_, _03019_);
  nor _26172_ (_03766_, _11492_, rst);
  or _26173_ (_03022_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or _26174_ (_03023_, _03013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and _26175_ (_03024_, _03023_, _03022_);
  or _26176_ (_03025_, _03024_, _09561_);
  nand _26177_ (_03026_, _09561_, _09008_);
  and _26178_ (_03027_, _03026_, _06989_);
  and _26179_ (_03791_, _03027_, _03025_);
  and _26180_ (_03028_, _11954_, _07044_);
  or _26181_ (_03029_, _03028_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _26182_ (_03030_, _03029_, _07292_);
  nand _26183_ (_03031_, _03028_, _06968_);
  and _26184_ (_03032_, _03031_, _03030_);
  or _26185_ (_03033_, _03032_, _07293_);
  and _26186_ (_03793_, _03033_, _06989_);
  nor _26187_ (_03795_, _11415_, rst);
  nand _26188_ (_03034_, _09531_, _07118_);
  and _26189_ (_03035_, _03013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _26190_ (_03036_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _26191_ (_03037_, _03036_, _03035_);
  or _26192_ (_03038_, _03037_, _09531_);
  and _26193_ (_03039_, _03038_, _06989_);
  and _26194_ (_03799_, _03039_, _03034_);
  nand _26195_ (_03040_, _09531_, _07260_);
  and _26196_ (_03041_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and _26197_ (_03042_, _03013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or _26198_ (_03043_, _03042_, _03041_);
  or _26199_ (_03044_, _03043_, _09531_);
  and _26200_ (_03045_, _03044_, _06989_);
  and _26201_ (_03802_, _03045_, _03040_);
  not _26202_ (_03046_, _09561_);
  or _26203_ (_03048_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  not _26204_ (_03049_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand _26205_ (_03050_, _09537_, _03049_);
  and _26206_ (_03051_, _03050_, _03048_);
  and _26207_ (_03052_, _03051_, _03046_);
  nor _26208_ (_03054_, _03046_, _07317_);
  or _26209_ (_03056_, _03054_, _03052_);
  and _26210_ (_03805_, _03056_, _06989_);
  nor _26211_ (_03808_, _12013_, rst);
  nor _26212_ (_03810_, _12036_, rst);
  and _26213_ (_03059_, _02462_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or _26214_ (_03060_, _02568_, _02709_);
  or _26215_ (_03061_, _03060_, _11395_);
  nand _26216_ (_03062_, _02575_, _11290_);
  nand _26217_ (_03063_, _03062_, _11326_);
  or _26218_ (_03064_, _03063_, _03061_);
  or _26219_ (_03065_, _02587_, _02408_);
  or _26220_ (_03066_, _03065_, _02579_);
  nand _26221_ (_03067_, _11457_, _11406_);
  or _26222_ (_03068_, _02467_, _11387_);
  or _26223_ (_03069_, _03068_, _02433_);
  and _26224_ (_03070_, _11356_, _11290_);
  or _26225_ (_03071_, _03070_, _11435_);
  or _26226_ (_03073_, _03071_, _03069_);
  or _26227_ (_03074_, _03073_, _03067_);
  or _26228_ (_03075_, _03074_, _03066_);
  or _26229_ (_03076_, _03075_, _03064_);
  not _26230_ (_03078_, _11429_);
  and _26231_ (_03080_, _11430_, _11382_);
  nor _26232_ (_03082_, _03080_, _02601_);
  and _26233_ (_03084_, _03082_, _03078_);
  not _26234_ (_03086_, _03084_);
  or _26235_ (_03088_, _02414_, _03086_);
  or _26236_ (_03090_, _03088_, _11283_);
  or _26237_ (_03092_, _03090_, _03076_);
  or _26238_ (_03094_, _11334_, _11282_);
  nor _26239_ (_03096_, \oc8051_top_1.oc8051_sfr1.wait_data , rst);
  and _26240_ (_03097_, _03096_, _03094_);
  and _26241_ (_03099_, _03097_, _03092_);
  or _26242_ (_03815_, _03099_, _03059_);
  or _26243_ (_03100_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or _26244_ (_03101_, _03013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _26245_ (_03102_, _03101_, _03100_);
  or _26246_ (_03103_, _03102_, _09531_);
  nand _26247_ (_03104_, _11529_, _09531_);
  and _26248_ (_03105_, _03104_, _06989_);
  and _26249_ (_03821_, _03105_, _03103_);
  and _26250_ (_03106_, _11954_, _08436_);
  or _26251_ (_03107_, _03106_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _26252_ (_03108_, _03107_, _07292_);
  nand _26253_ (_03109_, _03106_, _06968_);
  and _26254_ (_03110_, _03109_, _03108_);
  or _26255_ (_03111_, _03110_, _07318_);
  and _26256_ (_03825_, _03111_, _06989_);
  or _26257_ (_03112_, _07360_, _11345_);
  or _26258_ (_03113_, _07324_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and _26259_ (_03114_, _03113_, _06989_);
  and _26260_ (_03829_, _03114_, _03112_);
  nor _26261_ (_03115_, _11049_, _11044_);
  nor _26262_ (_03116_, _03115_, _11050_);
  or _26263_ (_03117_, _03116_, _08477_);
  or _26264_ (_03118_, _08476_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and _26265_ (_03119_, _03118_, _10964_);
  and _26266_ (_03120_, _03119_, _03117_);
  and _26267_ (_03121_, _10977_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or _26268_ (_03831_, _03121_, _03120_);
  or _26269_ (_03122_, _08496_, _11345_);
  or _26270_ (_03123_, _07324_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and _26271_ (_03124_, _03123_, _06989_);
  and _26272_ (_03833_, _03124_, _03122_);
  nand _26273_ (_03125_, _08512_, _07324_);
  or _26274_ (_03126_, _07324_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and _26275_ (_03128_, _03126_, _06989_);
  and _26276_ (_03835_, _03128_, _03125_);
  or _26277_ (_03129_, _08529_, _11345_);
  or _26278_ (_03130_, _07324_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and _26279_ (_03131_, _03130_, _06989_);
  and _26280_ (_03837_, _03131_, _03129_);
  or _26281_ (_03132_, _08545_, _11345_);
  or _26282_ (_03133_, _07324_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and _26283_ (_03134_, _03133_, _06989_);
  and _26284_ (_03839_, _03134_, _03132_);
  or _26285_ (_03136_, _08561_, _11345_);
  or _26286_ (_03137_, _07324_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and _26287_ (_03138_, _03137_, _06989_);
  and _26288_ (_03841_, _03138_, _03136_);
  nand _26289_ (_03139_, _08576_, _07324_);
  or _26290_ (_03140_, _07324_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and _26291_ (_03141_, _03140_, _06989_);
  and _26292_ (_03854_, _03141_, _03139_);
  or _26293_ (_03142_, _09537_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not _26294_ (_03143_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand _26295_ (_03144_, _09537_, _03143_);
  and _26296_ (_03145_, _03144_, _03142_);
  or _26297_ (_03147_, _03145_, _09561_);
  nand _26298_ (_03148_, _09598_, _09561_);
  and _26299_ (_03149_, _03148_, _06989_);
  and _26300_ (_03862_, _03149_, _03147_);
  or _26301_ (_03151_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _26302_ (_03152_, _08085_, _07978_);
  or _26303_ (_03153_, _03152_, _09182_);
  or _26304_ (_03154_, _03153_, _08402_);
  or _26305_ (_03155_, _03154_, _08231_);
  or _26306_ (_03157_, _03155_, _09092_);
  and _26307_ (_03158_, _03157_, _07027_);
  and _26308_ (_03159_, _06898_, _06848_);
  not _26309_ (_03160_, _06898_);
  and _26310_ (_03161_, _06900_, _03160_);
  or _26311_ (_03162_, _03161_, _03159_);
  and _26312_ (_03163_, _03162_, _06845_);
  nand _26313_ (_03164_, _06834_, _06599_);
  and _26314_ (_03165_, _06837_, _06548_);
  and _26315_ (_03166_, _03165_, _03164_);
  and _26316_ (_03167_, _07024_, _06652_);
  and _26317_ (_03168_, _03167_, _06622_);
  and _26318_ (_03169_, _03168_, _07634_);
  nand _26319_ (_03170_, _03169_, _08152_);
  nand _26320_ (_03171_, _03170_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or _26321_ (_03172_, _03171_, _03166_);
  nor _26322_ (_03173_, _03172_, _03163_);
  and _26323_ (_03174_, _03173_, _08318_);
  nand _26324_ (_03175_, _03174_, _12250_);
  or _26325_ (_03176_, _03175_, _03158_);
  and _26326_ (_03177_, _03176_, _03151_);
  or _26327_ (_03178_, _03177_, _11954_);
  not _26328_ (_03179_, _11954_);
  and _26329_ (_03180_, _00759_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _26330_ (_03181_, _03180_, _03179_);
  or _26331_ (_03182_, _03181_, _00760_);
  and _26332_ (_03183_, _03182_, _03178_);
  or _26333_ (_03184_, _03183_, _07291_);
  nand _26334_ (_03185_, _11529_, _07291_);
  and _26335_ (_03186_, _03185_, _06989_);
  and _26336_ (_03864_, _03186_, _03184_);
  or _26337_ (_03187_, _02583_, _11437_);
  or _26338_ (_03188_, _03187_, _02919_);
  or _26339_ (_03189_, _03188_, _02726_);
  not _26340_ (_03190_, _14315_);
  or _26341_ (_03191_, _02720_, _03190_);
  or _26342_ (_03192_, _03191_, _03189_);
  or _26343_ (_03193_, _02941_, _11395_);
  or _26344_ (_03194_, _02709_, _02423_);
  or _26345_ (_03195_, _03194_, _03193_);
  or _26346_ (_03196_, _02929_, _02582_);
  or _26347_ (_03197_, _03196_, _03195_);
  and _26348_ (_03198_, _11359_, _11290_);
  or _26349_ (_03199_, _02719_, _02406_);
  or _26350_ (_03200_, _03199_, _03198_);
  or _26351_ (_03201_, _11334_, _11433_);
  or _26352_ (_03202_, _11919_, _14316_);
  or _26353_ (_03203_, _03202_, _03201_);
  or _26354_ (_03204_, _03203_, _03200_);
  or _26355_ (_03205_, _03204_, _03197_);
  or _26356_ (_03206_, _03205_, _03192_);
  and _26357_ (_03207_, _03206_, _03097_);
  and _26358_ (_03208_, _02462_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  or _26359_ (_03869_, _03208_, _03207_);
  and _26360_ (_03210_, _11954_, _07089_);
  or _26361_ (_03211_, _03210_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and _26362_ (_03212_, _03211_, _07292_);
  nand _26363_ (_03213_, _03210_, _06968_);
  and _26364_ (_03214_, _03213_, _03212_);
  nor _26365_ (_03215_, _09008_, _07292_);
  or _26366_ (_03216_, _03215_, _03214_);
  and _26367_ (_03873_, _03216_, _06989_);
  and _26368_ (_03217_, _11355_, _11290_);
  or _26369_ (_03218_, _02406_, _14313_);
  or _26370_ (_03219_, _03218_, _03217_);
  or _26371_ (_03220_, _03219_, _02720_);
  or _26372_ (_03221_, _03188_, _02792_);
  or _26373_ (_03222_, _03221_, _03220_);
  or _26374_ (_03223_, _11456_, _11401_);
  or _26375_ (_03224_, _11453_, _14316_);
  or _26376_ (_03225_, _03224_, _03223_);
  or _26377_ (_03226_, _03225_, _02916_);
  or _26378_ (_03227_, _03226_, _02926_);
  or _26379_ (_03228_, _03227_, _03222_);
  and _26380_ (_03229_, _03228_, _07325_);
  and _26381_ (_03230_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and _26382_ (_03231_, _11333_, _06406_);
  or _26383_ (_03232_, _03231_, _03230_);
  or _26384_ (_03233_, _03232_, _03229_);
  and _26385_ (_03879_, _03233_, _06989_);
  nand _26386_ (_03234_, _09536_, _07317_);
  and _26387_ (_03235_, _09534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and _26388_ (_03236_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or _26389_ (_03237_, _03236_, _03235_);
  or _26390_ (_03238_, _03237_, _09536_);
  and _26391_ (_03239_, _03238_, _09552_);
  and _26392_ (_03240_, _03239_, _03234_);
  and _26393_ (_03241_, _09531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or _26394_ (_03242_, _03241_, _03240_);
  and _26395_ (_03917_, _03242_, _06989_);
  not _26396_ (_03243_, _09536_);
  or _26397_ (_03244_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  not _26398_ (_03245_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nand _26399_ (_03246_, _09533_, _03245_);
  nand _26400_ (_03247_, _03246_, _03244_);
  nand _26401_ (_03248_, _03247_, _03243_);
  nand _26402_ (_03249_, _10970_, _09536_);
  and _26403_ (_03250_, _03249_, _03248_);
  or _26404_ (_03251_, _03250_, _09561_);
  not _26405_ (_03252_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nand _26406_ (_03253_, _09561_, _03252_);
  and _26407_ (_03254_, _03253_, _06989_);
  and _26408_ (_03920_, _03254_, _03251_);
  nand _26409_ (_03255_, _09536_, _07118_);
  not _26410_ (_03256_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor _26411_ (_03257_, _09533_, _03256_);
  and _26412_ (_03258_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or _26413_ (_03259_, _03258_, _03257_);
  or _26414_ (_03260_, _03259_, _09536_);
  and _26415_ (_03261_, _03260_, _09552_);
  and _26416_ (_03262_, _03261_, _03255_);
  and _26417_ (_03263_, _09531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or _26418_ (_03264_, _03263_, _03262_);
  and _26419_ (_03926_, _03264_, _06989_);
  nand _26420_ (_03265_, _09536_, _07260_);
  and _26421_ (_03266_, _09534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and _26422_ (_03267_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or _26423_ (_03268_, _03267_, _03266_);
  or _26424_ (_03269_, _03268_, _09536_);
  and _26425_ (_03270_, _03269_, _09552_);
  and _26426_ (_03271_, _03270_, _03265_);
  and _26427_ (_03272_, _09531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or _26428_ (_03273_, _03272_, _03271_);
  and _26429_ (_03929_, _03273_, _06989_);
  nand _26430_ (_03274_, _11529_, _09536_);
  and _26431_ (_03275_, _09534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and _26432_ (_03276_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or _26433_ (_03277_, _03276_, _03275_);
  or _26434_ (_03278_, _03277_, _09536_);
  and _26435_ (_03279_, _03278_, _09552_);
  and _26436_ (_03280_, _03279_, _03274_);
  and _26437_ (_03281_, _09531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or _26438_ (_03282_, _03281_, _03280_);
  and _26439_ (_03942_, _03282_, _06989_);
  and _26440_ (_03283_, _08999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _26441_ (_03284_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and _26442_ (_03285_, _03284_, _09002_);
  and _26443_ (_03286_, _11821_, _09010_);
  or _26444_ (_03287_, _03286_, _03285_);
  or _26445_ (_03288_, _03287_, _03283_);
  and _26446_ (_03957_, _03288_, _06989_);
  nand _26447_ (_03289_, _09536_, _09008_);
  or _26448_ (_03290_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _26449_ (_03291_, _09534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and _26450_ (_03292_, _03291_, _03290_);
  or _26451_ (_03293_, _03292_, _09536_);
  and _26452_ (_03294_, _03293_, _09552_);
  and _26453_ (_03295_, _03294_, _03289_);
  and _26454_ (_03296_, _09531_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or _26455_ (_03297_, _03296_, _03295_);
  and _26456_ (_03966_, _03297_, _06989_);
  nand _26457_ (_03298_, _09598_, _09536_);
  or _26458_ (_03299_, _09533_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or _26459_ (_03300_, _09534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and _26460_ (_03301_, _03300_, _03299_);
  or _26461_ (_03302_, _03301_, _09536_);
  and _26462_ (_03303_, _03302_, _03298_);
  or _26463_ (_03304_, _03303_, _09561_);
  or _26464_ (_03305_, _03046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and _26465_ (_03306_, _03305_, _06989_);
  and _26466_ (_03971_, _03306_, _03304_);
  or _26467_ (_03307_, _08994_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand _26468_ (_03308_, _08994_, _07040_);
  and _26469_ (_03309_, _03308_, _03307_);
  or _26470_ (_03310_, _03309_, _06982_);
  or _26471_ (_03311_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  and _26472_ (_03312_, _03311_, _06989_);
  and _26473_ (_03992_, _03312_, _03310_);
  and _26474_ (_03314_, _02462_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  nor _26475_ (_03316_, _11909_, _11474_);
  nand _26476_ (_03317_, _03316_, _11920_);
  or _26477_ (_03318_, _02931_, _02927_);
  or _26478_ (_03319_, _03318_, _03317_);
  or _26479_ (_03320_, _02433_, _02423_);
  or _26480_ (_03321_, _02919_, _02691_);
  or _26481_ (_03322_, _03321_, _03320_);
  or _26482_ (_03323_, _03322_, _02785_);
  or _26483_ (_03324_, _03323_, _02917_);
  or _26484_ (_03325_, _03324_, _03319_);
  and _26485_ (_03326_, _03325_, _02487_);
  or _26486_ (_03995_, _03326_, _03314_);
  nor _26487_ (_03328_, _14146_, _07118_);
  and _26488_ (_03330_, _08999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _26489_ (_03332_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  and _26490_ (_03333_, _03332_, _09002_);
  or _26491_ (_03334_, _03333_, _03330_);
  or _26492_ (_03335_, _03334_, _03328_);
  and _26493_ (_04003_, _03335_, _06989_);
  nor _26494_ (_04007_, _12061_, rst);
  nor _26495_ (_03336_, _09614_, _07040_);
  and _26496_ (_03337_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or _26497_ (_03338_, _03337_, _06982_);
  or _26498_ (_03339_, _03338_, _03336_);
  or _26499_ (_03340_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and _26500_ (_03341_, _03340_, _06989_);
  and _26501_ (_04034_, _03341_, _03339_);
  or _26502_ (_03342_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand _26503_ (_03343_, _07493_, _14092_);
  and _26504_ (_03344_, _03343_, _06989_);
  and _26505_ (_04059_, _03344_, _03342_);
  and _26506_ (_03346_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and _26507_ (_03347_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  or _26508_ (_03348_, _03347_, _03346_);
  and _26509_ (_04061_, _03348_, _06989_);
  and _26510_ (_03349_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and _26511_ (_03351_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  or _26512_ (_03352_, _03351_, _03349_);
  and _26513_ (_04068_, _03352_, _06989_);
  and _26514_ (_04086_, _06989_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  and _26515_ (_03353_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or _26516_ (_03355_, _07024_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand _26517_ (_03356_, _03355_, _06989_);
  nor _26518_ (_04099_, _03356_, _03353_);
  and _26519_ (_04104_, _08314_, _06989_);
  and _26520_ (_03357_, _09610_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor _26521_ (_03358_, _11529_, _07486_);
  and _26522_ (_03359_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and _26523_ (_03360_, _03359_, _09615_);
  or _26524_ (_03361_, _03360_, _03358_);
  or _26525_ (_03362_, _03361_, _03357_);
  and _26526_ (_04112_, _03362_, _06989_);
  and _26527_ (_03363_, _11277_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and _26528_ (_03365_, _03363_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _26529_ (_03366_, _03365_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _26530_ (_03367_, _03366_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or _26531_ (_03368_, _03367_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nand _26532_ (_03369_, _03367_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and _26533_ (_03370_, _03369_, _03368_);
  or _26534_ (_03371_, _03370_, _11964_);
  and _26535_ (_03373_, _03371_, _06989_);
  and _26536_ (_03375_, _12750_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or _26537_ (_03376_, _03375_, _12752_);
  or _26538_ (_03377_, _12756_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and _26539_ (_03378_, _03377_, _12757_);
  or _26540_ (_03379_, _03378_, _12742_);
  and _26541_ (_03380_, _03379_, _12722_);
  and _26542_ (_03381_, _03380_, _03376_);
  nor _26543_ (_03382_, _12790_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor _26544_ (_03383_, _03382_, _12791_);
  and _26545_ (_03384_, _03383_, _12783_);
  and _26546_ (_03385_, _11413_, _08433_);
  nor _26547_ (_03386_, _12797_, _08385_);
  and _26548_ (_03387_, _11974_, _11514_);
  and _26549_ (_03388_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or _26550_ (_03389_, _03388_, _03387_);
  or _26551_ (_03390_, _03389_, _03386_);
  or _26552_ (_03391_, _03390_, _03385_);
  or _26553_ (_03392_, _03391_, _03384_);
  or _26554_ (_03393_, _03392_, _12781_);
  or _26555_ (_03394_, _03393_, _03381_);
  and _26556_ (_04114_, _03394_, _03373_);
  nand _26557_ (_03395_, _10970_, _10146_);
  or _26558_ (_03396_, _10146_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and _26559_ (_03397_, _03396_, _06989_);
  and _26560_ (_04117_, _03397_, _03395_);
  nor _26561_ (_03398_, _03366_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor _26562_ (_03400_, _03398_, _03367_);
  or _26563_ (_03401_, _03400_, _11964_);
  and _26564_ (_03402_, _03401_, _06989_);
  nor _26565_ (_03403_, _12797_, _09356_);
  nor _26566_ (_03404_, _11989_, _09227_);
  and _26567_ (_03405_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and _26568_ (_03406_, _11974_, _11842_);
  and _26569_ (_03407_, _12176_, _08463_);
  or _26570_ (_03408_, _03407_, _03406_);
  or _26571_ (_03409_, _03408_, _03405_);
  or _26572_ (_03410_, _03409_, _03404_);
  or _26573_ (_03411_, _03410_, _03403_);
  and _26574_ (_03412_, _12749_, _12742_);
  and _26575_ (_03414_, _12754_, _12747_);
  nor _26576_ (_03415_, _03414_, _12742_);
  or _26577_ (_03416_, _03415_, _03412_);
  nand _26578_ (_03417_, _03416_, _08175_);
  or _26579_ (_03418_, _03416_, _08175_);
  and _26580_ (_03419_, _03418_, _03417_);
  and _26581_ (_03421_, _03419_, _12722_);
  or _26582_ (_03423_, _03421_, _03411_);
  or _26583_ (_03424_, _03423_, _12781_);
  and _26584_ (_04122_, _03424_, _03402_);
  nor _26585_ (_03425_, _03365_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor _26586_ (_03426_, _03425_, _03366_);
  or _26587_ (_03427_, _03426_, _11964_);
  and _26588_ (_03429_, _03427_, _06989_);
  and _26589_ (_03430_, _12747_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or _26590_ (_03431_, _03430_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and _26591_ (_03432_, _03431_, _03415_);
  nand _26592_ (_03433_, _12748_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand _26593_ (_03434_, _03433_, _12749_);
  and _26594_ (_03435_, _03434_, _12742_);
  or _26595_ (_03436_, _03435_, _03432_);
  and _26596_ (_03437_, _03436_, _12722_);
  and _26597_ (_03438_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and _26598_ (_03440_, _11974_, _11744_);
  or _26599_ (_03441_, _03440_, _03438_);
  nor _26600_ (_03442_, _12797_, _07696_);
  or _26601_ (_03443_, _03442_, _03441_);
  and _26602_ (_03445_, _11413_, _08030_);
  and _26603_ (_03446_, _12783_, _10835_);
  or _26604_ (_03448_, _03446_, _03445_);
  or _26605_ (_03449_, _03448_, _03443_);
  or _26606_ (_03450_, _03449_, _03437_);
  or _26607_ (_03451_, _03450_, _12781_);
  and _26608_ (_04130_, _03451_, _03429_);
  nor _26609_ (_03452_, _03363_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor _26610_ (_03453_, _03452_, _03365_);
  or _26611_ (_03454_, _03453_, _11964_);
  and _26612_ (_03455_, _03454_, _06989_);
  and _26613_ (_03457_, _11413_, _08123_);
  nand _26614_ (_03458_, _12747_, _07646_);
  or _26615_ (_03459_, _12747_, _07646_);
  and _26616_ (_03460_, _03459_, _03458_);
  and _26617_ (_03461_, _03460_, _12742_);
  nor _26618_ (_03462_, _03460_, _12742_);
  or _26619_ (_03463_, _03462_, _03461_);
  and _26620_ (_03464_, _03463_, _12171_);
  and _26621_ (_03465_, _12167_, _08075_);
  and _26622_ (_03466_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and _26623_ (_03467_, _11974_, _11786_);
  or _26624_ (_03468_, _03467_, _03466_);
  and _26625_ (_03469_, _12176_, _08561_);
  nor _26626_ (_03470_, _03469_, _03468_);
  nand _26627_ (_03471_, _03470_, _11964_);
  or _26628_ (_03472_, _03471_, _03465_);
  or _26629_ (_03473_, _03472_, _03464_);
  or _26630_ (_03474_, _03473_, _03457_);
  and _26631_ (_04134_, _03474_, _03455_);
  nor _26632_ (_03476_, _11277_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _26633_ (_03477_, _03476_, _03363_);
  or _26634_ (_03478_, _03477_, _11964_);
  and _26635_ (_03480_, _03478_, _06989_);
  and _26636_ (_03481_, _12278_, _11986_);
  and _26637_ (_03482_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor _26638_ (_03483_, _12740_, _11988_);
  and _26639_ (_03484_, _12783_, _11608_);
  or _26640_ (_03485_, _03484_, _03483_);
  or _26641_ (_03487_, _03485_, _03482_);
  or _26642_ (_03488_, _12744_, _12743_);
  not _26643_ (_03490_, _03488_);
  nand _26644_ (_03491_, _03490_, _12745_);
  or _26645_ (_03492_, _03490_, _12745_);
  and _26646_ (_03493_, _03492_, _12722_);
  and _26647_ (_03494_, _03493_, _03491_);
  or _26648_ (_03495_, _03494_, _03487_);
  or _26649_ (_03496_, _03495_, _03481_);
  or _26650_ (_03497_, _03496_, _12781_);
  and _26651_ (_04137_, _03497_, _03480_);
  not _26652_ (_03498_, _00919_);
  and _26653_ (_03499_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and _26654_ (_03500_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _26655_ (_03501_, _03500_, _03499_);
  and _26656_ (_03502_, _03501_, _13953_);
  and _26657_ (_03503_, _13952_, _09393_);
  or _26658_ (_03504_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _13995_);
  and _26659_ (_03505_, _03504_, _06989_);
  and _26660_ (_03506_, _03505_, _03503_);
  or _26661_ (_04187_, _03506_, _03502_);
  nor _26662_ (_03507_, _03353_, _07526_);
  and _26663_ (_03508_, _03353_, _07526_);
  or _26664_ (_03509_, _03508_, _03507_);
  and _26665_ (_04196_, _03509_, _06989_);
  and _26666_ (_04199_, _12244_, _06989_);
  and _26667_ (_04206_, _06989_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nor _26668_ (_03510_, _14146_, _07040_);
  and _26669_ (_03511_, _08999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _26670_ (_03513_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  and _26671_ (_03514_, _03513_, _09002_);
  or _26672_ (_03515_, _03514_, _03511_);
  or _26673_ (_03516_, _03515_, _03510_);
  and _26674_ (_04207_, _03516_, _06989_);
  or _26675_ (_03517_, _09605_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nand _26676_ (_03519_, _09008_, _09605_);
  and _26677_ (_03520_, _03519_, _03517_);
  or _26678_ (_03522_, _03520_, _06982_);
  or _26679_ (_03523_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and _26680_ (_03524_, _03523_, _06989_);
  and _26681_ (_04211_, _03524_, _03522_);
  nor _26682_ (_03525_, _07317_, _09614_);
  and _26683_ (_03526_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or _26684_ (_03527_, _03526_, _06982_);
  or _26685_ (_03528_, _03527_, _03525_);
  or _26686_ (_03529_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and _26687_ (_03530_, _03529_, _06989_);
  and _26688_ (_04214_, _03530_, _03528_);
  nor _26689_ (_03531_, _10970_, _09614_);
  and _26690_ (_03532_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or _26691_ (_03533_, _03532_, _06982_);
  or _26692_ (_03534_, _03533_, _03531_);
  or _26693_ (_03535_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and _26694_ (_03536_, _03535_, _06989_);
  and _26695_ (_04216_, _03536_, _03534_);
  nor _26696_ (_03537_, _11724_, _14222_);
  and _26697_ (_03538_, _03537_, _14354_);
  or _26698_ (_03540_, _01595_, _14253_);
  or _26699_ (_03542_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and _26700_ (_03543_, _03542_, _14217_);
  and _26701_ (_03544_, _03543_, _03540_);
  and _26702_ (_03545_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and _26703_ (_03546_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or _26704_ (_03547_, _03546_, _03545_);
  and _26705_ (_03548_, _03547_, _14241_);
  nor _26706_ (_03550_, _11857_, _08412_);
  and _26707_ (_03551_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or _26708_ (_03552_, _03551_, _03550_);
  and _26709_ (_03553_, _03552_, _14205_);
  and _26710_ (_03554_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and _26711_ (_03555_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or _26712_ (_03556_, _03555_, _03554_);
  and _26713_ (_03558_, _03556_, _14233_);
  or _26714_ (_03559_, _03558_, _03553_);
  or _26715_ (_03560_, _03559_, _03548_);
  or _26716_ (_03562_, _03560_, _03544_);
  and _26717_ (_03563_, _03562_, _03538_);
  and _26718_ (_03564_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and _26719_ (_03565_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _26720_ (_03567_, _03565_, _03564_);
  and _26721_ (_03568_, _03567_, _14233_);
  and _26722_ (_03569_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and _26723_ (_03570_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _26724_ (_03571_, _03570_, _03569_);
  and _26725_ (_03572_, _03571_, _14205_);
  and _26726_ (_03573_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and _26727_ (_03574_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or _26728_ (_03575_, _03574_, _03573_);
  and _26729_ (_03576_, _03575_, _14217_);
  or _26730_ (_03577_, _03576_, _03572_);
  and _26731_ (_03578_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and _26732_ (_03580_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or _26733_ (_03581_, _03580_, _03578_);
  and _26734_ (_03582_, _03581_, _14241_);
  or _26735_ (_03583_, _03582_, _03577_);
  or _26736_ (_03584_, _03583_, _03568_);
  and _26737_ (_03585_, _03584_, _14209_);
  and _26738_ (_03586_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and _26739_ (_03587_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or _26740_ (_03588_, _03587_, _03586_);
  and _26741_ (_03589_, _03588_, _14241_);
  and _26742_ (_03590_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and _26743_ (_03591_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or _26744_ (_03592_, _03591_, _03590_);
  and _26745_ (_03593_, _03592_, _14205_);
  nor _26746_ (_03594_, _11857_, _07176_);
  and _26747_ (_03595_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or _26748_ (_03596_, _03595_, _03594_);
  and _26749_ (_03597_, _03596_, _14217_);
  or _26750_ (_03599_, _03597_, _03593_);
  nor _26751_ (_03600_, _11857_, _07172_);
  and _26752_ (_03601_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or _26753_ (_03602_, _03601_, _03600_);
  and _26754_ (_03603_, _03602_, _14233_);
  or _26755_ (_03604_, _03603_, _03599_);
  or _26756_ (_03605_, _03604_, _03589_);
  and _26757_ (_03606_, _03605_, _14248_);
  nor _26758_ (_03607_, _11857_, _07213_);
  and _26759_ (_03608_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or _26760_ (_03609_, _03608_, _03607_);
  and _26761_ (_03610_, _03609_, _14217_);
  and _26762_ (_03611_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _26763_ (_03612_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or _26764_ (_03613_, _03612_, _03611_);
  and _26765_ (_03614_, _03613_, _14241_);
  or _26766_ (_03615_, _03614_, _03610_);
  and _26767_ (_03616_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and _26768_ (_03618_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or _26769_ (_03620_, _03618_, _03616_);
  and _26770_ (_03621_, _03620_, _14205_);
  and _26771_ (_03623_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  nor _26772_ (_03624_, _11857_, _07211_);
  or _26773_ (_03625_, _03624_, _03623_);
  and _26774_ (_03626_, _03625_, _14233_);
  or _26775_ (_03627_, _03626_, _03621_);
  or _26776_ (_03628_, _03627_, _03615_);
  and _26777_ (_03629_, _03628_, _14252_);
  or _26778_ (_03630_, _03629_, _03606_);
  or _26779_ (_03631_, _03630_, _03585_);
  and _26780_ (_03632_, _03631_, _14222_);
  and _26781_ (_03633_, _14209_, _11556_);
  nor _26782_ (_03635_, _14326_, p0_in[7]);
  and _26783_ (_03637_, _14326_, _00731_);
  nor _26784_ (_03639_, _03637_, _03635_);
  and _26785_ (_03640_, _03639_, _14253_);
  and _26786_ (_03642_, _14463_, _11857_);
  or _26787_ (_03644_, _03642_, _03640_);
  and _26788_ (_03646_, _03644_, _14241_);
  and _26789_ (_03647_, _14602_, _11857_);
  and _26790_ (_03649_, _01288_, _14253_);
  or _26791_ (_03650_, _03649_, _03647_);
  and _26792_ (_03652_, _03650_, _14233_);
  and _26793_ (_03653_, _14529_, _11857_);
  and _26794_ (_03654_, _14342_, _14253_);
  or _26795_ (_03656_, _03654_, _03653_);
  and _26796_ (_03658_, _03656_, _14205_);
  and _26797_ (_03660_, _01462_, _14253_);
  and _26798_ (_03661_, _01541_, _11857_);
  or _26799_ (_03663_, _03661_, _03660_);
  and _26800_ (_03665_, _03663_, _14217_);
  or _26801_ (_03667_, _03665_, _03658_);
  or _26802_ (_03668_, _03667_, _03652_);
  or _26803_ (_03670_, _03668_, _03646_);
  and _26804_ (_03671_, _03670_, _03633_);
  and _26805_ (_03673_, _11724_, _11556_);
  and _26806_ (_03674_, _03673_, _14292_);
  nor _26807_ (_03676_, _11857_, _06649_);
  and _26808_ (_03677_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or _26809_ (_03678_, _03677_, _03676_);
  and _26810_ (_03680_, _03678_, _14217_);
  nor _26811_ (_03681_, _11857_, _06813_);
  and _26812_ (_03683_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or _26813_ (_03684_, _03683_, _03681_);
  and _26814_ (_03685_, _03684_, _14205_);
  or _26815_ (_03686_, _03685_, _03680_);
  nor _26816_ (_03688_, _11857_, _06619_);
  and _26817_ (_03689_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or _26818_ (_03690_, _03689_, _03688_);
  and _26819_ (_03691_, _03690_, _14233_);
  nor _26820_ (_03692_, _11857_, _06592_);
  and _26821_ (_03694_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or _26822_ (_03695_, _03694_, _03692_);
  and _26823_ (_03696_, _03695_, _14241_);
  or _26824_ (_03697_, _03696_, _03691_);
  or _26825_ (_03699_, _03697_, _03686_);
  and _26826_ (_03700_, _03699_, _03674_);
  or _26827_ (_03701_, _03700_, _03671_);
  and _26828_ (_03702_, _11863_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and _26829_ (_03703_, _14214_, _14222_);
  and _26830_ (_03704_, _03703_, _14206_);
  and _26831_ (_03705_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and _26832_ (_03707_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or _26833_ (_03708_, _03707_, _03705_);
  and _26834_ (_03709_, _03708_, _14205_);
  nor _26835_ (_03710_, _11857_, _13993_);
  and _26836_ (_03711_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or _26837_ (_03713_, _03711_, _03710_);
  and _26838_ (_03714_, _03713_, _14217_);
  or _26839_ (_03716_, _03714_, _03709_);
  and _26840_ (_03717_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  nor _26841_ (_03718_, _11857_, _06970_);
  or _26842_ (_03720_, _03718_, _03717_);
  and _26843_ (_03722_, _03720_, _14241_);
  nor _26844_ (_03724_, _11857_, _14039_);
  and _26845_ (_03725_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or _26846_ (_03727_, _03725_, _03724_);
  and _26847_ (_03728_, _03727_, _14233_);
  or _26848_ (_03729_, _03728_, _03722_);
  or _26849_ (_03730_, _03729_, _03716_);
  and _26850_ (_03731_, _03730_, _03704_);
  or _26851_ (_03732_, _03731_, _03702_);
  or _26852_ (_03733_, _03732_, _03701_);
  and _26853_ (_03734_, _01535_, _11857_);
  and _26854_ (_03735_, _01468_, _14253_);
  or _26855_ (_03736_, _03735_, _03734_);
  and _26856_ (_03737_, _03736_, _14217_);
  and _26857_ (_03738_, _14612_, _11857_);
  and _26858_ (_03739_, _01303_, _14253_);
  or _26859_ (_03740_, _03739_, _03738_);
  and _26860_ (_03741_, _03740_, _14233_);
  or _26861_ (_03743_, _03741_, _11724_);
  or _26862_ (_03744_, _03743_, _03737_);
  and _26863_ (_03745_, _14540_, _14205_);
  and _26864_ (_03746_, _14458_, _14241_);
  or _26865_ (_03747_, _03746_, _03745_);
  and _26866_ (_03748_, _03747_, _11857_);
  and _26867_ (_03749_, _14330_, _14205_);
  nor _26868_ (_03750_, _14326_, p3_in[7]);
  and _26869_ (_03751_, _14326_, _01165_);
  nor _26870_ (_03752_, _03751_, _03750_);
  and _26871_ (_03753_, _03752_, _14241_);
  or _26872_ (_03754_, _03753_, _03749_);
  and _26873_ (_03756_, _03754_, _14253_);
  or _26874_ (_03757_, _03756_, _03748_);
  or _26875_ (_03759_, _03757_, _03744_);
  and _26876_ (_03760_, _14247_, _11556_);
  and _26877_ (_03762_, _14544_, _11857_);
  and _26878_ (_03763_, _14336_, _14253_);
  or _26879_ (_03765_, _03763_, _03762_);
  and _26880_ (_03767_, _03765_, _14205_);
  and _26881_ (_03768_, _14616_, _11857_);
  and _26882_ (_03769_, _01298_, _14253_);
  or _26883_ (_03770_, _03769_, _03768_);
  and _26884_ (_03771_, _03770_, _14233_);
  or _26885_ (_03772_, _03771_, _14251_);
  or _26886_ (_03773_, _03772_, _03767_);
  and _26887_ (_03774_, _14453_, _14241_);
  and _26888_ (_03775_, _01530_, _14217_);
  or _26889_ (_03776_, _03775_, _03774_);
  and _26890_ (_03777_, _03776_, _11857_);
  nor _26891_ (_03778_, _14326_, p2_in[7]);
  and _26892_ (_03779_, _14326_, _09033_);
  nor _26893_ (_03780_, _03779_, _03778_);
  and _26894_ (_03781_, _03780_, _14241_);
  and _26895_ (_03782_, _01473_, _14217_);
  or _26896_ (_03783_, _03782_, _03781_);
  and _26897_ (_03784_, _03783_, _14253_);
  or _26898_ (_03785_, _03784_, _03777_);
  or _26899_ (_03786_, _03785_, _03773_);
  and _26900_ (_03787_, _03786_, _03760_);
  and _26901_ (_03788_, _03787_, _03759_);
  nor _26902_ (_03789_, _11857_, _01372_);
  and _26903_ (_03790_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or _26904_ (_03792_, _03790_, _03789_);
  and _26905_ (_03794_, _03792_, _14233_);
  or _26906_ (_03796_, _03794_, _11556_);
  and _26907_ (_03797_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and _26908_ (_03798_, _14253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or _26909_ (_03800_, _03798_, _03797_);
  and _26910_ (_03801_, _03800_, _14205_);
  nor _26911_ (_03803_, _11857_, _09405_);
  and _26912_ (_03804_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or _26913_ (_03806_, _03804_, _03803_);
  and _26914_ (_03807_, _03806_, _14217_);
  and _26915_ (_03809_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  nor _26916_ (_03811_, _11857_, _13995_);
  or _26917_ (_03812_, _03811_, _03809_);
  and _26918_ (_03813_, _03812_, _14241_);
  or _26919_ (_03814_, _03813_, _03807_);
  or _26920_ (_03816_, _03814_, _03801_);
  or _26921_ (_03817_, _03816_, _03796_);
  and _26922_ (_03818_, _14534_, _11857_);
  and _26923_ (_03819_, _14347_, _14253_);
  or _26924_ (_03820_, _03819_, _03818_);
  and _26925_ (_03822_, _03820_, _14205_);
  and _26926_ (_03823_, _14606_, _11857_);
  and _26927_ (_03824_, _01293_, _14253_);
  or _26928_ (_03826_, _03824_, _03823_);
  and _26929_ (_03827_, _03826_, _14233_);
  or _26930_ (_03828_, _03827_, _14222_);
  or _26931_ (_03830_, _03828_, _03822_);
  nor _26932_ (_03832_, _14326_, p1_in[7]);
  and _26933_ (_03834_, _14326_, _00702_);
  nor _26934_ (_03836_, _03834_, _03832_);
  and _26935_ (_03838_, _03836_, _14241_);
  and _26936_ (_03840_, _01457_, _14217_);
  or _26937_ (_03842_, _03840_, _03838_);
  and _26938_ (_03843_, _03842_, _14253_);
  and _26939_ (_03844_, _14467_, _14241_);
  and _26940_ (_03845_, _01546_, _14217_);
  or _26941_ (_03846_, _03845_, _03844_);
  and _26942_ (_03847_, _03846_, _11857_);
  or _26943_ (_03848_, _03847_, _03843_);
  or _26944_ (_03849_, _03848_, _03830_);
  and _26945_ (_03850_, _03849_, _14276_);
  and _26946_ (_03851_, _03850_, _03817_);
  and _26947_ (_03852_, _03537_, _14292_);
  nor _26948_ (_03853_, _03852_, _03538_);
  nor _26949_ (_03855_, _03704_, _03674_);
  and _26950_ (_03856_, _03855_, _03853_);
  nor _26951_ (_03857_, _14275_, _14222_);
  nor _26952_ (_03858_, _14208_, _11556_);
  or _26953_ (_03859_, _03858_, _03857_);
  not _26954_ (_03860_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor _26955_ (_03861_, _03760_, _03860_);
  and _26956_ (_03863_, _03861_, _03859_);
  and _26957_ (_03865_, _03863_, _03856_);
  nor _26958_ (_03866_, _11857_, _01749_);
  and _26959_ (_03867_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or _26960_ (_03868_, _03867_, _03866_);
  and _26961_ (_03870_, _03868_, _14217_);
  nor _26962_ (_03871_, _11857_, _01885_);
  and _26963_ (_03872_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or _26964_ (_03874_, _03872_, _03871_);
  and _26965_ (_03875_, _03874_, _14205_);
  or _26966_ (_03876_, _03875_, _03870_);
  nor _26967_ (_03877_, _11857_, _01321_);
  and _26968_ (_03878_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or _26969_ (_03880_, _03878_, _03877_);
  and _26970_ (_03881_, _03880_, _14233_);
  not _26971_ (_03882_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor _26972_ (_03883_, _11857_, _03882_);
  and _26973_ (_03884_, _11857_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or _26974_ (_03885_, _03884_, _03883_);
  and _26975_ (_03886_, _03885_, _14241_);
  or _26976_ (_03887_, _03886_, _03881_);
  or _26977_ (_03888_, _03887_, _03876_);
  and _26978_ (_03889_, _03888_, _03852_);
  or _26979_ (_03890_, _03889_, _03865_);
  or _26980_ (_03891_, _03890_, _03851_);
  or _26981_ (_03892_, _03891_, _03788_);
  or _26982_ (_03893_, _03892_, _03733_);
  or _26983_ (_03894_, _03893_, _03632_);
  or _26984_ (_03895_, _03894_, _03563_);
  and _26985_ (_03896_, _03674_, _07705_);
  nor _26986_ (_03897_, _03896_, _11873_);
  nand _26987_ (_03898_, _03702_, _06968_);
  and _26988_ (_03899_, _03898_, _03897_);
  and _26989_ (_03900_, _03899_, _03895_);
  and _26990_ (_03901_, _11857_, _09009_);
  nor _26991_ (_03902_, _11857_, _07118_);
  or _26992_ (_03903_, _03902_, _03901_);
  and _26993_ (_03904_, _03903_, _14233_);
  and _26994_ (_03905_, _11857_, _11821_);
  nor _26995_ (_03906_, _11857_, _10970_);
  or _26996_ (_03907_, _03906_, _03905_);
  and _26997_ (_03908_, _03907_, _14205_);
  nor _26998_ (_03909_, _11857_, _07260_);
  and _26999_ (_03910_, _11857_, _09599_);
  or _27000_ (_03911_, _03910_, _03909_);
  and _27001_ (_03912_, _03911_, _14217_);
  or _27002_ (_03913_, _03912_, _03908_);
  nor _27003_ (_03914_, _11857_, _07040_);
  and _27004_ (_03915_, _11857_, _07410_);
  or _27005_ (_03916_, _03915_, _03914_);
  and _27006_ (_03918_, _03916_, _14241_);
  or _27007_ (_03919_, _03918_, _03913_);
  nor _27008_ (_03921_, _03919_, _03904_);
  nor _27009_ (_03922_, _03921_, _03897_);
  or _27010_ (_03923_, _03922_, _03900_);
  and _27011_ (_04219_, _03923_, _06989_);
  nor _27012_ (_03924_, _00489_, rst);
  or _27013_ (_03925_, _00488_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand _27014_ (_03927_, _00488_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and _27015_ (_03928_, _03927_, _03925_);
  and _27016_ (_04224_, _03928_, _03924_);
  and _27017_ (_04227_, _00490_, _06989_);
  nor _27018_ (_03930_, _02976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor _27019_ (_03931_, _03930_, _02977_);
  or _27020_ (_03932_, _03931_, _11964_);
  and _27021_ (_03933_, _03932_, _06989_);
  and _27022_ (_03934_, _02995_, _09270_);
  nor _27023_ (_03935_, _02995_, _09270_);
  or _27024_ (_03936_, _03935_, _03934_);
  and _27025_ (_03937_, _03936_, _12753_);
  nand _27026_ (_03938_, _02991_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand _27027_ (_03939_, _03938_, _02992_);
  and _27028_ (_03940_, _03939_, _12742_);
  or _27029_ (_03941_, _03940_, _03937_);
  and _27030_ (_03943_, _03941_, _12722_);
  nor _27031_ (_03944_, _03004_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor _27032_ (_03945_, _03944_, _03005_);
  and _27033_ (_03946_, _03945_, _12783_);
  nor _27034_ (_03947_, _11989_, _09145_);
  nor _27035_ (_03948_, _12797_, _09285_);
  and _27036_ (_03949_, _11974_, _11618_);
  and _27037_ (_03950_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or _27038_ (_03951_, _03950_, _03949_);
  or _27039_ (_03952_, _03951_, _03948_);
  or _27040_ (_03953_, _03952_, _03947_);
  or _27041_ (_03954_, _03953_, _03946_);
  or _27042_ (_03955_, _03954_, _12781_);
  or _27043_ (_03956_, _03955_, _03943_);
  and _27044_ (_04233_, _03956_, _03933_);
  nor _27045_ (_03958_, _12716_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor _27046_ (_03959_, _03958_, _02976_);
  or _27047_ (_03960_, _03959_, _11964_);
  and _27048_ (_03961_, _03960_, _06989_);
  or _27049_ (_03962_, _12793_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not _27050_ (_03963_, _03004_);
  and _27051_ (_03964_, _03963_, _12783_);
  and _27052_ (_03965_, _03964_, _03962_);
  and _27053_ (_03967_, _11413_, _08268_);
  nor _27054_ (_03968_, _12797_, _08202_);
  and _27055_ (_03969_, _11985_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and _27056_ (_03970_, _11974_, _11671_);
  or _27057_ (_03972_, _03970_, _03969_);
  or _27058_ (_03973_, _03972_, _03968_);
  or _27059_ (_03974_, _03973_, _03967_);
  or _27060_ (_03975_, _02990_, _12753_);
  or _27061_ (_03976_, _02994_, _12742_);
  and _27062_ (_03977_, _03976_, _03975_);
  nand _27063_ (_03978_, _03977_, _08187_);
  or _27064_ (_03979_, _03977_, _08187_);
  and _27065_ (_03980_, _03979_, _03978_);
  and _27066_ (_03981_, _03980_, _12722_);
  or _27067_ (_03982_, _03981_, _03974_);
  or _27068_ (_03983_, _03982_, _03965_);
  or _27069_ (_03984_, _03983_, _12781_);
  and _27070_ (_04236_, _03984_, _03961_);
  and _27071_ (_03986_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _27072_ (_03987_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or _27073_ (_03988_, _03987_, _03986_);
  or _27074_ (_03989_, _03988_, _13986_);
  and _27075_ (_03990_, _03989_, _06989_);
  nand _27076_ (_03991_, _03503_, _07040_);
  and _27077_ (_04282_, _03991_, _03990_);
  or _27078_ (_03993_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand _27079_ (_03994_, _07493_, _14184_);
  and _27080_ (_03996_, _03994_, _06989_);
  and _27081_ (_04306_, _03996_, _03993_);
  and _27082_ (_03997_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and _27083_ (_03998_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or _27084_ (_03999_, _03998_, _03997_);
  and _27085_ (_04000_, _03999_, _13953_);
  nand _27086_ (_04001_, _09392_, _07040_);
  nand _27087_ (_04002_, _10970_, _09393_);
  and _27088_ (_04004_, _04002_, _00922_);
  and _27089_ (_04005_, _04004_, _04001_);
  or _27090_ (_04334_, _04005_, _04000_);
  and _27091_ (_04006_, _13952_, _09392_);
  and _27092_ (_04008_, _04006_, _11646_);
  and _27093_ (_04009_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and _27094_ (_04010_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor _27095_ (_04011_, _04010_, _04009_);
  nor _27096_ (_04012_, _04011_, _13986_);
  and _27097_ (_04013_, _03503_, _07119_);
  or _27098_ (_04014_, _04013_, _04012_);
  or _27099_ (_04015_, _04014_, _04008_);
  and _27100_ (_04339_, _04015_, _06989_);
  not _27101_ (_04016_, _11353_);
  and _27102_ (_04017_, _02701_, _04016_);
  nor _27103_ (_04018_, _02697_, _11474_);
  nand _27104_ (_04019_, _04018_, _11440_);
  or _27105_ (_04020_, _04019_, _11449_);
  or _27106_ (_04021_, _04020_, _02917_);
  and _27107_ (_04022_, _04021_, _11282_);
  or _27108_ (_04023_, _04022_, _04017_);
  and _27109_ (_04353_, _04023_, _06989_);
  nor _27110_ (_04024_, _14213_, rst);
  and _27111_ (_04025_, _12278_, _06989_);
  or _27112_ (_04026_, _04025_, _04024_);
  not _27113_ (_04027_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nor _27114_ (_04028_, _14404_, _04027_);
  nand _27115_ (_04029_, _14226_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand _27116_ (_04030_, _14220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and _27117_ (_04031_, _04030_, _04029_);
  nand _27118_ (_04032_, _14231_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nand _27119_ (_04033_, _14235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and _27120_ (_04035_, _04033_, _04032_);
  and _27121_ (_04036_, _04035_, _04031_);
  nand _27122_ (_04037_, _14239_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  nand _27123_ (_04038_, _14243_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and _27124_ (_04039_, _04038_, _04037_);
  nand _27125_ (_04040_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nand _27126_ (_04041_, _14257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _27127_ (_04042_, _04041_, _04040_);
  and _27128_ (_04043_, _04042_, _04039_);
  and _27129_ (_04044_, _04043_, _04036_);
  nand _27130_ (_04045_, _14263_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  nand _27131_ (_04046_, _14266_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and _27132_ (_04047_, _04046_, _04045_);
  nand _27133_ (_04048_, _14269_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand _27134_ (_04049_, _14271_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and _27135_ (_04050_, _04049_, _04048_);
  and _27136_ (_04051_, _04050_, _04047_);
  nand _27137_ (_04052_, _14277_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nand _27138_ (_04053_, _14279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and _27139_ (_04054_, _04053_, _04052_);
  nand _27140_ (_04055_, _14282_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand _27141_ (_04056_, _14284_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and _27142_ (_04057_, _04056_, _04055_);
  and _27143_ (_04058_, _04057_, _04054_);
  and _27144_ (_04060_, _04058_, _04051_);
  and _27145_ (_04062_, _04060_, _04044_);
  nand _27146_ (_04063_, _14293_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nand _27147_ (_04064_, _14296_, _11605_);
  and _27148_ (_04065_, _04064_, _04063_);
  nand _27149_ (_04066_, _14212_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  nand _27150_ (_04067_, _14301_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  and _27151_ (_04069_, _04067_, _04066_);
  and _27152_ (_04070_, _04069_, _04065_);
  nand _27153_ (_04071_, _03780_, _14333_);
  nand _27154_ (_04072_, _03752_, _14305_);
  and _27155_ (_04073_, _04072_, _04071_);
  nand _27156_ (_04074_, _03639_, _14339_);
  nand _27157_ (_04075_, _03836_, _14344_);
  and _27158_ (_04076_, _04075_, _04074_);
  and _27159_ (_04077_, _04076_, _04073_);
  and _27160_ (_04078_, _04077_, _04070_);
  nand _27161_ (_04079_, _14355_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nand _27162_ (_04080_, _14352_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and _27163_ (_04081_, _04080_, _04079_);
  and _27164_ (_04082_, _04081_, _04078_);
  nand _27165_ (_04083_, _04082_, _04062_);
  nand _27166_ (_04084_, _04083_, _14374_);
  nand _27167_ (_04085_, _04084_, _14483_);
  or _27168_ (_04087_, _04085_, _04028_);
  and _27169_ (_04355_, _04087_, _04026_);
  or _27170_ (_04088_, _07493_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand _27171_ (_04089_, _07493_, _14168_);
  and _27172_ (_04090_, _04089_, _06989_);
  and _27173_ (_04360_, _04090_, _04088_);
  or _27174_ (_04091_, _01319_, _12278_);
  nand _27175_ (_04092_, _01319_, _03882_);
  and _27176_ (_04093_, _04092_, _06983_);
  and _27177_ (_04094_, _04093_, _04091_);
  nor _27178_ (_04095_, _06484_, _03882_);
  and _27179_ (_04096_, _01318_, _06539_);
  nand _27180_ (_04097_, _04096_, _06968_);
  or _27181_ (_04098_, _04096_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and _27182_ (_04100_, _04098_, _06485_);
  and _27183_ (_04101_, _04100_, _04097_);
  or _27184_ (_04102_, _04101_, _04095_);
  or _27185_ (_04103_, _04102_, _04094_);
  and _27186_ (_04485_, _04103_, _06989_);
  nor _27187_ (_04487_, _11841_, rst);
  nor _27188_ (_04105_, _09614_, _07118_);
  and _27189_ (_04106_, _09614_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or _27190_ (_04107_, _04106_, _06982_);
  or _27191_ (_04108_, _04107_, _04105_);
  or _27192_ (_04109_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and _27193_ (_04110_, _04109_, _06989_);
  and _27194_ (_04524_, _04110_, _04108_);
  nand _27195_ (_04111_, _06513_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor _27196_ (_04113_, _04111_, _06538_);
  or _27197_ (_04115_, _04113_, _01556_);
  and _27198_ (_04116_, _04115_, _00867_);
  nand _27199_ (_04118_, _00867_, _06513_);
  and _27200_ (_04119_, _04118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or _27201_ (_04120_, _04119_, _07459_);
  or _27202_ (_04121_, _04120_, _04116_);
  nand _27203_ (_04123_, _10970_, _07459_);
  and _27204_ (_04124_, _04123_, _06989_);
  and _27205_ (_04527_, _04124_, _04121_);
  and _27206_ (_04125_, _00791_, _06539_);
  nand _27207_ (_04126_, _04125_, _06968_);
  or _27208_ (_04127_, _04125_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and _27209_ (_04128_, _04127_, _00803_);
  and _27210_ (_04129_, _04128_, _04126_);
  nor _27211_ (_04131_, _00803_, _07040_);
  or _27212_ (_04132_, _04131_, _04129_);
  and _27213_ (_04529_, _04132_, _06989_);
  and _27214_ (_04133_, _07493_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and _27215_ (_04135_, _11273_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  or _27216_ (_04136_, _04135_, _04133_);
  and _27217_ (_04532_, _04136_, _06989_);
  and _27218_ (_04138_, _00708_, _06539_);
  nand _27219_ (_04139_, _04138_, _06968_);
  or _27220_ (_04140_, _04138_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and _27221_ (_04141_, _04140_, _00715_);
  and _27222_ (_04142_, _04141_, _04139_);
  nor _27223_ (_04143_, _00715_, _07040_);
  or _27224_ (_04144_, _04143_, _04142_);
  and _27225_ (_04539_, _04144_, _06989_);
  and _27226_ (_04145_, _08436_, _06501_);
  nand _27227_ (_04146_, _04145_, _06968_);
  or _27228_ (_04147_, _04145_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and _27229_ (_04148_, _04147_, _02635_);
  and _27230_ (_04149_, _04148_, _04146_);
  nor _27231_ (_04150_, _07317_, _02635_);
  or _27232_ (_04151_, _04150_, _04149_);
  and _27233_ (_04544_, _04151_, _06989_);
  and _27234_ (_04152_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _27235_ (_04153_, _04152_, _00760_);
  and _27236_ (_04154_, _04153_, _06501_);
  nand _27237_ (_04155_, _00764_, _06501_);
  and _27238_ (_04156_, _04155_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or _27239_ (_04157_, _04156_, _06987_);
  or _27240_ (_04158_, _04157_, _04154_);
  nand _27241_ (_04159_, _11529_, _06987_);
  and _27242_ (_04160_, _04159_, _06989_);
  and _27243_ (_04547_, _04160_, _04158_);
  and _27244_ (_04161_, _07089_, _06501_);
  nand _27245_ (_04162_, _04161_, _06968_);
  or _27246_ (_04163_, _04161_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and _27247_ (_04164_, _04163_, _02635_);
  and _27248_ (_04165_, _04164_, _04162_);
  nor _27249_ (_04166_, _09008_, _02635_);
  or _27250_ (_04167_, _04166_, _04165_);
  and _27251_ (_04550_, _04167_, _06989_);
  and _27252_ (_04168_, _06979_, _06501_);
  nand _27253_ (_04169_, _04168_, _06968_);
  or _27254_ (_04170_, _04168_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and _27255_ (_04171_, _04170_, _02635_);
  and _27256_ (_04172_, _04171_, _04169_);
  and _27257_ (_04173_, _09599_, _06987_);
  or _27258_ (_04174_, _04173_, _04172_);
  and _27259_ (_04555_, _04174_, _06989_);
  and _27260_ (_04175_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and _27261_ (_04176_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor _27262_ (_04177_, _04176_, _04175_);
  nor _27263_ (_04178_, _04177_, _13986_);
  and _27264_ (_04179_, _03503_, _07429_);
  or _27265_ (_04180_, _04179_, _04178_);
  and _27266_ (_04181_, _13986_, _09392_);
  and _27267_ (_04182_, _04181_, _07119_);
  or _27268_ (_04183_, _04182_, _04180_);
  and _27269_ (_04557_, _04183_, _06989_);
  and _27270_ (_04184_, _04006_, _07429_);
  and _27271_ (_04185_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and _27272_ (_04186_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor _27273_ (_04188_, _04186_, _04185_);
  nor _27274_ (_04189_, _04188_, _13986_);
  and _27275_ (_04190_, _03503_, _07410_);
  or _27276_ (_04191_, _04190_, _04189_);
  or _27277_ (_04192_, _04191_, _04184_);
  and _27278_ (_04560_, _04192_, _06989_);
  and _27279_ (_04193_, _04006_, _07410_);
  and _27280_ (_04194_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and _27281_ (_04195_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor _27282_ (_04197_, _04195_, _04194_);
  nor _27283_ (_04198_, _04197_, _13986_);
  and _27284_ (_04200_, _03503_, _11821_);
  or _27285_ (_04201_, _04200_, _04198_);
  or _27286_ (_04202_, _04201_, _04193_);
  and _27287_ (_04563_, _04202_, _06989_);
  and _27288_ (_04203_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor _27289_ (_04204_, _08139_, _01188_);
  or _27290_ (_04205_, _04204_, _04203_);
  and _27291_ (_04566_, _04205_, _06989_);
  and _27292_ (_04208_, _11986_, _08346_);
  or _27293_ (_04209_, _12134_, _12131_);
  and _27294_ (_04210_, _12171_, _12135_);
  and _27295_ (_04212_, _04210_, _04209_);
  nor _27296_ (_04213_, _12036_, _11988_);
  and _27297_ (_04215_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and _27298_ (_04217_, _12176_, _11718_);
  or _27299_ (_04218_, _04217_, _04215_);
  or _27300_ (_04220_, _04218_, _04213_);
  nor _27301_ (_04221_, _04220_, _04212_);
  nand _27302_ (_04222_, _04221_, _11964_);
  or _27303_ (_04223_, _04222_, _04208_);
  nor _27304_ (_04225_, _08595_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor _27305_ (_04226_, _04225_, _12673_);
  or _27306_ (_04228_, _04226_, _11964_);
  and _27307_ (_04229_, _04228_, _06989_);
  and _27308_ (_04568_, _04229_, _04223_);
  and _27309_ (_04570_, _04024_, _14377_);
  or _27310_ (_04230_, _11964_, _08596_);
  and _27311_ (_04231_, _11986_, _08433_);
  and _27312_ (_04232_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor _27313_ (_04234_, _12061_, _11988_);
  and _27314_ (_04235_, _12783_, _11514_);
  or _27315_ (_04237_, _04235_, _04234_);
  or _27316_ (_04238_, _04237_, _04232_);
  or _27317_ (_04239_, _12064_, _12065_);
  nor _27318_ (_04240_, _04239_, _12129_);
  and _27319_ (_04241_, _04239_, _12129_);
  or _27320_ (_04242_, _04241_, _04240_);
  and _27321_ (_04243_, _04242_, _12722_);
  or _27322_ (_04244_, _04243_, _04238_);
  or _27323_ (_04245_, _04244_, _04231_);
  or _27324_ (_04246_, _04245_, _12781_);
  and _27325_ (_04247_, _04246_, _06989_);
  and _27326_ (_04572_, _04247_, _04230_);
  and _27327_ (_04248_, _12691_, _08588_);
  and _27328_ (_04249_, _11986_, _01898_);
  and _27329_ (_04250_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor _27330_ (_04251_, _11988_, _11207_);
  and _27331_ (_04252_, _12783_, _11842_);
  or _27332_ (_04253_, _04252_, _04251_);
  or _27333_ (_04254_, _04253_, _04250_);
  nor _27334_ (_04255_, _12126_, _12124_);
  nor _27335_ (_04256_, _04255_, _12127_);
  and _27336_ (_04257_, _04256_, _12722_);
  or _27337_ (_04258_, _04257_, _04254_);
  or _27338_ (_04259_, _04258_, _04249_);
  and _27339_ (_04260_, _04259_, _11964_);
  or _27340_ (_04261_, _04260_, _04248_);
  and _27341_ (_04582_, _04261_, _06989_);
  and _27342_ (_04262_, _12691_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _27343_ (_04263_, _11986_, _08030_);
  or _27344_ (_04264_, _12120_, _12118_);
  and _27345_ (_04265_, _12171_, _12123_);
  and _27346_ (_04266_, _04265_, _04264_);
  and _27347_ (_04267_, _12091_, _11974_);
  and _27348_ (_04268_, _11413_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and _27349_ (_04269_, _12176_, _11744_);
  or _27350_ (_04270_, _04269_, _04268_);
  or _27351_ (_04271_, _04270_, _04267_);
  or _27352_ (_04272_, _04271_, _04266_);
  or _27353_ (_04273_, _04272_, _04263_);
  and _27354_ (_04274_, _04273_, _11964_);
  or _27355_ (_04275_, _04274_, _04262_);
  and _27356_ (_04585_, _04275_, _06989_);
  and _27357_ (_04276_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and _27358_ (_04277_, _04276_, _09580_);
  nor _27359_ (_04278_, _07140_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  nor _27360_ (_04279_, _04278_, _07141_);
  or _27361_ (_04280_, _04279_, _04277_);
  and _27362_ (_04281_, _04280_, _09574_);
  and _27363_ (_04283_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or _27364_ (_04284_, _04283_, _07046_);
  or _27365_ (_04285_, _04284_, _04281_);
  not _27366_ (_04286_, _07046_);
  or _27367_ (_04287_, _04286_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and _27368_ (_04288_, _04287_, _09590_);
  and _27369_ (_04289_, _04288_, _04285_);
  nor _27370_ (_04290_, _10970_, _09590_);
  or _27371_ (_04291_, _04290_, _04289_);
  and _27372_ (_04592_, _04291_, _06989_);
  nor _27373_ (_04292_, _07118_, _09590_);
  and _27374_ (_04293_, _07071_, _07063_);
  nor _27375_ (_04294_, _04293_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nor _27376_ (_04295_, _04294_, _07140_);
  or _27377_ (_04296_, _04295_, _07077_);
  and _27378_ (_04297_, _07147_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _27379_ (_04298_, _04297_, _07066_);
  or _27380_ (_04299_, _04298_, _04296_);
  or _27381_ (_04300_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and _27382_ (_04301_, _04300_, _07051_);
  and _27383_ (_04302_, _04301_, _04299_);
  and _27384_ (_04303_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or _27385_ (_04304_, _04303_, _04302_);
  or _27386_ (_04305_, _04304_, _04292_);
  and _27387_ (_04594_, _04305_, _06989_);
  nand _27388_ (_04799_, _11794_, _06989_);
  nand _27389_ (_04801_, _11739_, _06989_);
  nand _27390_ (_04805_, _11851_, _06989_);
  nor _27391_ (_04813_, _11548_, rst);
  nor _27392_ (_04815_, _11697_, rst);
  nor _27393_ (_04817_, _11682_, rst);
  nor _27394_ (_04819_, _11626_, rst);
  nor _27395_ (_04307_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not _27396_ (_04308_, _04307_);
  and _27397_ (_04309_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _27398_ (_04310_, _04309_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _27399_ (_04311_, _04309_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _27400_ (_04312_, _04311_, _04310_);
  not _27401_ (_04313_, _04312_);
  and _27402_ (_04314_, _04310_, _01350_);
  nor _27403_ (_04315_, _04310_, _01350_);
  nor _27404_ (_04316_, _04315_, _04314_);
  nor _27405_ (_04317_, _04316_, _08593_);
  and _27406_ (_04318_, _04316_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor _27407_ (_04319_, _04318_, _04317_);
  nor _27408_ (_04320_, _04319_, _04313_);
  and _27409_ (_04321_, _04316_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor _27410_ (_04322_, _04316_, _08621_);
  nor _27411_ (_04323_, _04322_, _04321_);
  nor _27412_ (_04324_, _04323_, _04312_);
  nor _27413_ (_04325_, _04324_, _04320_);
  nor _27414_ (_04326_, _04325_, _04308_);
  and _27415_ (_04327_, _13921_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not _27416_ (_04328_, _04327_);
  not _27417_ (_04329_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nor _27418_ (_04330_, _04316_, _04329_);
  and _27419_ (_04331_, _04316_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _27420_ (_04332_, _04331_, _04330_);
  nor _27421_ (_04333_, _04332_, _04313_);
  and _27422_ (_04335_, _04316_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not _27423_ (_04336_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _27424_ (_04337_, _04316_, _04336_);
  nor _27425_ (_04338_, _04337_, _04335_);
  nor _27426_ (_04340_, _04338_, _04312_);
  nor _27427_ (_04341_, _04340_, _04333_);
  nor _27428_ (_04342_, _04341_, _04328_);
  nor _27429_ (_04343_, _04342_, _04326_);
  not _27430_ (_04344_, _04309_);
  nor _27431_ (_04345_, _04316_, _08647_);
  and _27432_ (_04346_, _04316_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _27433_ (_04347_, _04346_, _04345_);
  nor _27434_ (_04348_, _04347_, _04313_);
  and _27435_ (_04349_, _04316_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor _27436_ (_04350_, _04316_, _09234_);
  nor _27437_ (_04351_, _04350_, _04349_);
  nor _27438_ (_04352_, _04351_, _04312_);
  nor _27439_ (_04354_, _04352_, _04348_);
  nor _27440_ (_04356_, _04354_, _04344_);
  and _27441_ (_04357_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _12949_);
  not _27442_ (_04358_, _04357_);
  not _27443_ (_04359_, \oc8051_symbolic_cxrom1.regvalid [14]);
  nor _27444_ (_04361_, _04316_, _04359_);
  and _27445_ (_04362_, _04316_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _27446_ (_04363_, _04362_, _04361_);
  nor _27447_ (_04364_, _04363_, _04313_);
  and _27448_ (_04365_, _04316_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not _27449_ (_04366_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor _27450_ (_04367_, _04316_, _04366_);
  nor _27451_ (_04368_, _04367_, _04365_);
  nor _27452_ (_04369_, _04368_, _04312_);
  nor _27453_ (_04370_, _04369_, _04364_);
  nor _27454_ (_04371_, _04370_, _04358_);
  nor _27455_ (_04372_, _04371_, _04356_);
  and _27456_ (_04373_, _04372_, _04343_);
  and _27457_ (_04374_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and _27458_ (_04375_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor _27459_ (_04376_, _04375_, _04374_);
  and _27460_ (_04377_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and _27461_ (_04378_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor _27462_ (_04379_, _04378_, _04377_);
  and _27463_ (_04380_, _04379_, _04376_);
  and _27464_ (_04381_, _04380_, _04313_);
  not _27465_ (_04382_, _04316_);
  and _27466_ (_04383_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and _27467_ (_04384_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor _27468_ (_04385_, _04384_, _04383_);
  and _27469_ (_04386_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and _27470_ (_04387_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor _27471_ (_04388_, _04387_, _04386_);
  and _27472_ (_04389_, _04388_, _04385_);
  and _27473_ (_04390_, _04389_, _04312_);
  or _27474_ (_04391_, _04390_, _04382_);
  nor _27475_ (_04392_, _04391_, _04381_);
  and _27476_ (_04393_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and _27477_ (_04394_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor _27478_ (_04395_, _04394_, _04393_);
  and _27479_ (_04396_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and _27480_ (_04397_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor _27481_ (_04398_, _04397_, _04396_);
  and _27482_ (_04399_, _04398_, _04395_);
  nor _27483_ (_04400_, _04399_, _04312_);
  and _27484_ (_04401_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and _27485_ (_04402_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor _27486_ (_04403_, _04402_, _04401_);
  and _27487_ (_04404_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and _27488_ (_04405_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor _27489_ (_04406_, _04405_, _04404_);
  and _27490_ (_04407_, _04406_, _04403_);
  nor _27491_ (_04408_, _04407_, _04313_);
  or _27492_ (_04409_, _04408_, _04400_);
  and _27493_ (_04410_, _04409_, _04382_);
  nor _27494_ (_04411_, _04410_, _04392_);
  nor _27495_ (_04412_, _04411_, _04373_);
  or _27496_ (_04413_, _04412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand _27497_ (_04414_, _04412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _27498_ (_04415_, _04414_, _04413_);
  not _27499_ (_04416_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not _27500_ (_04417_, _04373_);
  and _27501_ (_04418_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and _27502_ (_04419_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor _27503_ (_04420_, _04419_, _04418_);
  and _27504_ (_04421_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and _27505_ (_04422_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor _27506_ (_04423_, _04422_, _04421_);
  and _27507_ (_04424_, _04423_, _04420_);
  and _27508_ (_04425_, _04424_, _04313_);
  and _27509_ (_04426_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and _27510_ (_04427_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor _27511_ (_04428_, _04427_, _04426_);
  and _27512_ (_04429_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and _27513_ (_04430_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor _27514_ (_04431_, _04430_, _04429_);
  and _27515_ (_04432_, _04431_, _04428_);
  and _27516_ (_04433_, _04432_, _04312_);
  nor _27517_ (_04434_, _04433_, _04425_);
  nor _27518_ (_04435_, _04434_, _04382_);
  and _27519_ (_04436_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and _27520_ (_04437_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor _27521_ (_04438_, _04437_, _04436_);
  and _27522_ (_04439_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and _27523_ (_04440_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor _27524_ (_04441_, _04440_, _04439_);
  and _27525_ (_04442_, _04441_, _04438_);
  and _27526_ (_04443_, _04442_, _04313_);
  and _27527_ (_04444_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and _27528_ (_04445_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor _27529_ (_04446_, _04445_, _04444_);
  and _27530_ (_04447_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and _27531_ (_04448_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor _27532_ (_04449_, _04448_, _04447_);
  and _27533_ (_04450_, _04449_, _04446_);
  and _27534_ (_04451_, _04450_, _04312_);
  nor _27535_ (_04452_, _04451_, _04443_);
  nor _27536_ (_04453_, _04452_, _04316_);
  nor _27537_ (_04454_, _04453_, _04435_);
  and _27538_ (_04455_, _04454_, _04417_);
  and _27539_ (_04456_, _04455_, _04416_);
  nor _27540_ (_04457_, _04455_, _04416_);
  or _27541_ (_04458_, _04457_, _04456_);
  or _27542_ (_04459_, _04458_, _04415_);
  and _27543_ (_04460_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and _27544_ (_04461_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor _27545_ (_04462_, _04461_, _04460_);
  and _27546_ (_04463_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and _27547_ (_04464_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor _27548_ (_04465_, _04464_, _04463_);
  and _27549_ (_04466_, _04465_, _04462_);
  and _27550_ (_04467_, _04466_, _04313_);
  and _27551_ (_04468_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and _27552_ (_04469_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor _27553_ (_04470_, _04469_, _04468_);
  and _27554_ (_04471_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and _27555_ (_04472_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor _27556_ (_04473_, _04472_, _04471_);
  and _27557_ (_04474_, _04473_, _04470_);
  and _27558_ (_04475_, _04474_, _04312_);
  nor _27559_ (_04476_, _04475_, _04467_);
  nor _27560_ (_04477_, _04476_, _04382_);
  and _27561_ (_04478_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and _27562_ (_04479_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor _27563_ (_04480_, _04479_, _04478_);
  and _27564_ (_04481_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and _27565_ (_04482_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor _27566_ (_04483_, _04482_, _04481_);
  and _27567_ (_04484_, _04483_, _04480_);
  and _27568_ (_04486_, _04484_, _04313_);
  and _27569_ (_04488_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and _27570_ (_04489_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor _27571_ (_04490_, _04489_, _04488_);
  and _27572_ (_04491_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and _27573_ (_04492_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor _27574_ (_04493_, _04492_, _04491_);
  and _27575_ (_04494_, _04493_, _04490_);
  and _27576_ (_04495_, _04494_, _04312_);
  nor _27577_ (_04496_, _04495_, _04486_);
  nor _27578_ (_04497_, _04496_, _04316_);
  nor _27579_ (_04498_, _04497_, _04477_);
  and _27580_ (_04499_, _04498_, _04417_);
  or _27581_ (_04500_, _04499_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand _27582_ (_04501_, _04499_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _27583_ (_04502_, _04501_, _04500_);
  not _27584_ (_04503_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _27585_ (_04504_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and _27586_ (_04505_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor _27587_ (_04506_, _04505_, _04504_);
  and _27588_ (_04507_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and _27589_ (_04508_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor _27590_ (_04509_, _04508_, _04507_);
  and _27591_ (_04510_, _04509_, _04506_);
  and _27592_ (_04511_, _04510_, _04313_);
  and _27593_ (_04512_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and _27594_ (_04513_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor _27595_ (_04514_, _04513_, _04512_);
  and _27596_ (_04515_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and _27597_ (_04516_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor _27598_ (_04517_, _04516_, _04515_);
  and _27599_ (_04518_, _04517_, _04514_);
  and _27600_ (_04519_, _04518_, _04312_);
  or _27601_ (_04520_, _04519_, _04382_);
  nor _27602_ (_04521_, _04520_, _04511_);
  and _27603_ (_04522_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and _27604_ (_04523_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor _27605_ (_04525_, _04523_, _04522_);
  and _27606_ (_04526_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and _27607_ (_04528_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor _27608_ (_04530_, _04528_, _04526_);
  and _27609_ (_04531_, _04530_, _04525_);
  nor _27610_ (_04533_, _04531_, _04312_);
  and _27611_ (_04534_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and _27612_ (_04535_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor _27613_ (_04536_, _04535_, _04534_);
  and _27614_ (_04537_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and _27615_ (_04538_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor _27616_ (_04540_, _04538_, _04537_);
  and _27617_ (_04541_, _04540_, _04536_);
  nor _27618_ (_04542_, _04541_, _04313_);
  or _27619_ (_04543_, _04542_, _04533_);
  and _27620_ (_04545_, _04543_, _04382_);
  nor _27621_ (_04546_, _04545_, _04521_);
  nor _27622_ (_04548_, _04546_, _04373_);
  nor _27623_ (_04549_, _04548_, _04503_);
  and _27624_ (_04551_, _04548_, _04503_);
  or _27625_ (_04552_, _04551_, _04549_);
  or _27626_ (_04553_, _04552_, _04502_);
  or _27627_ (_04554_, _04553_, _04459_);
  and _27628_ (_04556_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and _27629_ (_04558_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor _27630_ (_04559_, _04558_, _04556_);
  and _27631_ (_04561_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and _27632_ (_04562_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor _27633_ (_04564_, _04562_, _04561_);
  and _27634_ (_04565_, _04564_, _04559_);
  and _27635_ (_04567_, _04565_, _04313_);
  and _27636_ (_04569_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and _27637_ (_04571_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor _27638_ (_04573_, _04571_, _04569_);
  and _27639_ (_04574_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and _27640_ (_04575_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor _27641_ (_04576_, _04575_, _04574_);
  and _27642_ (_04577_, _04576_, _04573_);
  and _27643_ (_04578_, _04577_, _04312_);
  or _27644_ (_04579_, _04578_, _04316_);
  nor _27645_ (_04580_, _04579_, _04567_);
  and _27646_ (_04581_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and _27647_ (_04583_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor _27648_ (_04584_, _04583_, _04581_);
  and _27649_ (_04586_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and _27650_ (_04587_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor _27651_ (_04588_, _04587_, _04586_);
  and _27652_ (_04589_, _04588_, _04584_);
  nor _27653_ (_04590_, _04589_, _04312_);
  and _27654_ (_04591_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and _27655_ (_04593_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor _27656_ (_04595_, _04593_, _04591_);
  and _27657_ (_04596_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and _27658_ (_04597_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor _27659_ (_04598_, _04597_, _04596_);
  and _27660_ (_04599_, _04598_, _04595_);
  nor _27661_ (_04600_, _04599_, _04313_);
  or _27662_ (_04601_, _04600_, _04590_);
  and _27663_ (_04602_, _04601_, _04316_);
  nor _27664_ (_04603_, _04602_, _04580_);
  nor _27665_ (_04604_, _04603_, _04373_);
  or _27666_ (_04605_, _04604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand _27667_ (_04606_, _04604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _27668_ (_04607_, _04606_, _04605_);
  not _27669_ (_04608_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _27670_ (_04609_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and _27671_ (_04610_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor _27672_ (_04611_, _04610_, _04609_);
  and _27673_ (_04612_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and _27674_ (_04613_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor _27675_ (_04614_, _04613_, _04612_);
  and _27676_ (_04615_, _04614_, _04611_);
  and _27677_ (_04616_, _04615_, _04313_);
  and _27678_ (_04617_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and _27679_ (_04618_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor _27680_ (_04619_, _04618_, _04617_);
  and _27681_ (_04620_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and _27682_ (_04621_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor _27683_ (_04622_, _04621_, _04620_);
  and _27684_ (_04623_, _04622_, _04619_);
  and _27685_ (_04624_, _04623_, _04312_);
  or _27686_ (_04625_, _04624_, _04382_);
  nor _27687_ (_04626_, _04625_, _04616_);
  and _27688_ (_04627_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and _27689_ (_04628_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor _27690_ (_04629_, _04628_, _04627_);
  and _27691_ (_04630_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and _27692_ (_04631_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor _27693_ (_04632_, _04631_, _04630_);
  and _27694_ (_04633_, _04632_, _04629_);
  and _27695_ (_04634_, _04633_, _04313_);
  and _27696_ (_04635_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and _27697_ (_04636_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor _27698_ (_04637_, _04636_, _04635_);
  and _27699_ (_04638_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and _27700_ (_04639_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor _27701_ (_04640_, _04639_, _04638_);
  and _27702_ (_04641_, _04640_, _04637_);
  and _27703_ (_04642_, _04641_, _04312_);
  or _27704_ (_04643_, _04642_, _04316_);
  nor _27705_ (_04644_, _04643_, _04634_);
  nor _27706_ (_04645_, _04644_, _04626_);
  nor _27707_ (_04646_, _04645_, _04373_);
  and _27708_ (_04647_, _04646_, _04608_);
  nor _27709_ (_04648_, _04646_, _04608_);
  or _27710_ (_04649_, _04648_, _04647_);
  or _27711_ (_04650_, _04649_, _04607_);
  and _27712_ (_04651_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _27713_ (_04652_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor _27714_ (_04653_, _04652_, _04651_);
  and _27715_ (_04654_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and _27716_ (_04655_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor _27717_ (_04656_, _04655_, _04654_);
  and _27718_ (_04657_, _04656_, _04653_);
  and _27719_ (_04658_, _04657_, _04313_);
  and _27720_ (_04659_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and _27721_ (_04660_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor _27722_ (_04661_, _04660_, _04659_);
  and _27723_ (_04662_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _27724_ (_04663_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor _27725_ (_04664_, _04663_, _04662_);
  and _27726_ (_04665_, _04664_, _04661_);
  and _27727_ (_04666_, _04665_, _04312_);
  or _27728_ (_04667_, _04666_, _04382_);
  nor _27729_ (_04668_, _04667_, _04658_);
  and _27730_ (_04669_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _27731_ (_04670_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor _27732_ (_04671_, _04670_, _04669_);
  and _27733_ (_04672_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and _27734_ (_04673_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor _27735_ (_04674_, _04673_, _04672_);
  and _27736_ (_04675_, _04674_, _04671_);
  and _27737_ (_04676_, _04675_, _04313_);
  and _27738_ (_04677_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _27739_ (_04678_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor _27740_ (_04679_, _04678_, _04677_);
  and _27741_ (_04680_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and _27742_ (_04681_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor _27743_ (_04682_, _04681_, _04680_);
  and _27744_ (_04683_, _04682_, _04679_);
  and _27745_ (_04684_, _04683_, _04312_);
  or _27746_ (_04685_, _04684_, _04316_);
  nor _27747_ (_04686_, _04685_, _04676_);
  nor _27748_ (_04687_, _04686_, _04668_);
  nor _27749_ (_04688_, _04687_, _04373_);
  nor _27750_ (_04689_, _04688_, _01149_);
  and _27751_ (_04690_, _04688_, _01149_);
  or _27752_ (_04691_, _04690_, _04689_);
  and _27753_ (_04692_, _04357_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and _27754_ (_04693_, _04309_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor _27755_ (_04694_, _04693_, _04692_);
  and _27756_ (_04695_, _04327_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and _27757_ (_04696_, _04307_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor _27758_ (_04697_, _04696_, _04695_);
  and _27759_ (_04698_, _04697_, _04694_);
  and _27760_ (_04699_, _04698_, _04313_);
  and _27761_ (_04700_, _04327_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and _27762_ (_04701_, _04307_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor _27763_ (_04702_, _04701_, _04700_);
  and _27764_ (_04703_, _04357_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and _27765_ (_04704_, _04309_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor _27766_ (_04705_, _04704_, _04703_);
  and _27767_ (_04706_, _04705_, _04702_);
  and _27768_ (_04707_, _04706_, _04312_);
  or _27769_ (_04708_, _04707_, _04316_);
  nor _27770_ (_04709_, _04708_, _04699_);
  and _27771_ (_04710_, _04327_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and _27772_ (_04711_, _04357_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor _27773_ (_04712_, _04711_, _04710_);
  and _27774_ (_04713_, _04307_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and _27775_ (_04714_, _04309_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor _27776_ (_04715_, _04714_, _04713_);
  and _27777_ (_04716_, _04715_, _04712_);
  nor _27778_ (_04717_, _04716_, _04312_);
  and _27779_ (_04718_, _04357_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and _27780_ (_04719_, _04309_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor _27781_ (_04720_, _04719_, _04718_);
  and _27782_ (_04721_, _04327_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and _27783_ (_04722_, _04307_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor _27784_ (_04723_, _04722_, _04721_);
  and _27785_ (_04724_, _04723_, _04720_);
  nor _27786_ (_04725_, _04724_, _04313_);
  or _27787_ (_04726_, _04725_, _04717_);
  and _27788_ (_04727_, _04726_, _04316_);
  nor _27789_ (_04728_, _04727_, _04709_);
  nor _27790_ (_04729_, _04728_, _04373_);
  nor _27791_ (_04730_, _04729_, _01188_);
  and _27792_ (_04731_, _04729_, _01188_);
  or _27793_ (_04732_, _04731_, _04730_);
  or _27794_ (_04733_, _04732_, _04691_);
  or _27795_ (_04734_, _04733_, _04650_);
  or _27796_ (_04735_, _04734_, _04554_);
  and _27797_ (_04736_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27798_ (_04737_, _04736_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _27799_ (_04738_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and _27800_ (_04739_, _04738_, _04737_);
  and _27801_ (_04740_, _04739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  and _27802_ (_04741_, _04740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _27803_ (_04742_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and _27804_ (_04743_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _27805_ (_04744_, _04743_, _04742_);
  and _27806_ (_04745_, _04744_, _04741_);
  and _27807_ (_04746_, _04745_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _27808_ (_04747_, _04746_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _27809_ (_04748_, _04747_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  and _27810_ (_04749_, _04748_, _00655_);
  nor _27811_ (_04750_, _04748_, _00655_);
  or _27812_ (_04751_, _04750_, _04749_);
  nor _27813_ (_04752_, _04751_, _00619_);
  and _27814_ (_04753_, _04751_, _00619_);
  or _27815_ (_04754_, _04753_, _04752_);
  and _27816_ (_04755_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _27817_ (_04756_, _04755_, _04738_);
  and _27818_ (_04757_, _04756_, _04737_);
  and _27819_ (_04758_, _04757_, _04744_);
  and _27820_ (_04759_, _04758_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _27821_ (_04760_, _04759_, _00683_);
  and _27822_ (_04761_, _04759_, _00683_);
  or _27823_ (_04762_, _04761_, _04760_);
  nor _27824_ (_04763_, _04762_, _01686_);
  and _27825_ (_04764_, _04762_, _01686_);
  or _27826_ (_04765_, _04764_, _04763_);
  nor _27827_ (_04766_, _04745_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _27828_ (_04767_, _04766_, _04746_);
  or _27829_ (_04768_, _04767_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand _27830_ (_04769_, _04767_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  and _27831_ (_04770_, _04769_, _04768_);
  or _27832_ (_04771_, _04770_, _04765_);
  nor _27833_ (_04772_, _04747_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _27834_ (_04773_, _04772_, _04748_);
  or _27835_ (_04774_, _04773_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand _27836_ (_04775_, _04773_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _27837_ (_04776_, _04775_, _04774_);
  or _27838_ (_04777_, _04776_, _04771_);
  or _27839_ (_04778_, _04777_, _04754_);
  and _27840_ (_04779_, _12949_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _27841_ (_04780_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08593_);
  nor _27842_ (_04781_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  nor _27843_ (_04782_, _04781_, _04780_);
  and _27844_ (_04783_, _04782_, _04779_);
  nor _27845_ (_04784_, _04783_, _13921_);
  nor _27846_ (_04785_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and _27847_ (_04786_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04329_);
  or _27848_ (_04787_, _04786_, _01231_);
  nor _27849_ (_04788_, _04787_, _04785_);
  and _27850_ (_04789_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04336_);
  nor _27851_ (_04790_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  nor _27852_ (_04791_, _04790_, _04789_);
  and _27853_ (_04792_, _04791_, _01231_);
  nor _27854_ (_04793_, _04792_, _04788_);
  nor _27855_ (_04794_, _04793_, _12949_);
  nor _27856_ (_04795_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor _27857_ (_04796_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  and _27858_ (_04797_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08621_);
  nor _27859_ (_04798_, _04797_, _04796_);
  and _27860_ (_04800_, _04798_, _04795_);
  nor _27861_ (_04802_, _04800_, _04794_);
  and _27862_ (_04803_, _04802_, _04784_);
  nor _27863_ (_04804_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and _27864_ (_04806_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04359_);
  or _27865_ (_04807_, _04806_, _01231_);
  nor _27866_ (_04808_, _04807_, _04804_);
  and _27867_ (_04809_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04366_);
  nor _27868_ (_04810_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _27869_ (_04811_, _04810_, _04809_);
  and _27870_ (_04812_, _04811_, _01231_);
  nor _27871_ (_04814_, _04812_, _04808_);
  nor _27872_ (_04816_, _04814_, _12949_);
  nor _27873_ (_04818_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [0]);
  and _27874_ (_04820_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _09234_);
  nor _27875_ (_04821_, _04820_, _04818_);
  and _27876_ (_04822_, _04821_, _04795_);
  and _27877_ (_04823_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08647_);
  nor _27878_ (_04824_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _27879_ (_04825_, _04824_, _04823_);
  and _27880_ (_04826_, _04825_, _04779_);
  or _27881_ (_04827_, _04826_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _27882_ (_04828_, _04827_, _04822_);
  nor _27883_ (_04829_, _04828_, _04816_);
  nor _27884_ (_04830_, _04829_, _04803_);
  nor _27885_ (_04831_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27886_ (_04832_, _09847_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27887_ (_04833_, _04832_, _04831_);
  and _27888_ (_04834_, _04833_, _04795_);
  nor _27889_ (_04836_, _04834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _27890_ (_04837_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27891_ (_04838_, _10325_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27892_ (_04839_, _04838_, _04837_);
  and _27893_ (_04840_, _04839_, _04779_);
  not _27894_ (_04841_, _04840_);
  nor _27895_ (_04842_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27896_ (_04844_, _10100_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27897_ (_04845_, _04844_, _04842_);
  and _27898_ (_04846_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _01231_);
  and _27899_ (_04847_, _04846_, _04845_);
  nor _27900_ (_04849_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27901_ (_04850_, _10537_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27902_ (_04851_, _04850_, _04849_);
  and _27903_ (_04852_, _04851_, _04736_);
  nor _27904_ (_04853_, _04852_, _04847_);
  and _27905_ (_04854_, _04853_, _04841_);
  and _27906_ (_04855_, _04854_, _04836_);
  nor _27907_ (_04856_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27908_ (_04857_, _10759_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27909_ (_04858_, _04857_, _04856_);
  and _27910_ (_04859_, _04858_, _04795_);
  nor _27911_ (_04860_, _04859_, _01350_);
  nor _27912_ (_04861_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27913_ (_04862_, _12513_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27914_ (_04863_, _04862_, _04861_);
  and _27915_ (_04864_, _04863_, _04779_);
  not _27916_ (_04865_, _04864_);
  nor _27917_ (_04866_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27918_ (_04867_, _12209_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27919_ (_04868_, _04867_, _04866_);
  and _27920_ (_04869_, _04868_, _04846_);
  nor _27921_ (_04870_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27922_ (_04871_, _12899_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27923_ (_04873_, _04871_, _04870_);
  and _27924_ (_04874_, _04873_, _04736_);
  nor _27925_ (_04875_, _04874_, _04869_);
  and _27926_ (_04876_, _04875_, _04865_);
  and _27927_ (_04877_, _04876_, _04860_);
  nor _27928_ (_04878_, _04877_, _04855_);
  and _27929_ (_04879_, _04878_, _04830_);
  nor _27930_ (_04880_, _04879_, _01144_);
  and _27931_ (_04881_, _04879_, _01144_);
  or _27932_ (_04882_, _04881_, _04880_);
  nor _27933_ (_04883_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27934_ (_04884_, _10113_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27935_ (_04885_, _04884_, _04883_);
  and _27936_ (_04886_, _04885_, _04846_);
  nor _27937_ (_04887_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27938_ (_04888_, _10338_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27939_ (_04890_, _04888_, _04887_);
  and _27940_ (_04891_, _04890_, _04779_);
  nor _27941_ (_04892_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27942_ (_04893_, _09860_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27943_ (_04894_, _04893_, _04892_);
  and _27944_ (_04895_, _04894_, _04795_);
  nor _27945_ (_04897_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27946_ (_04898_, _10548_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27947_ (_04899_, _04898_, _04897_);
  and _27948_ (_04900_, _04899_, _04736_);
  or _27949_ (_04901_, _04900_, _04895_);
  or _27950_ (_04902_, _04901_, _04891_);
  or _27951_ (_04903_, _04902_, _04886_);
  and _27952_ (_04904_, _04903_, _01350_);
  nor _27953_ (_04905_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27954_ (_04906_, _12225_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27955_ (_04907_, _04906_, _04905_);
  and _27956_ (_04908_, _04907_, _04846_);
  nor _27957_ (_04910_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27958_ (_04911_, _12524_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27959_ (_04912_, _04911_, _04910_);
  and _27960_ (_04913_, _04912_, _04779_);
  nor _27961_ (_04914_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27962_ (_04915_, _10771_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27963_ (_04917_, _04915_, _04914_);
  and _27964_ (_04918_, _04917_, _04795_);
  nor _27965_ (_04919_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _27966_ (_04921_, _12914_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _27967_ (_04923_, _04921_, _04919_);
  and _27968_ (_04925_, _04923_, _04736_);
  or _27969_ (_04926_, _04925_, _04918_);
  or _27970_ (_04927_, _04926_, _04913_);
  or _27971_ (_04928_, _04927_, _04908_);
  and _27972_ (_04929_, _04928_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _27973_ (_04930_, _04929_, _04904_);
  and _27974_ (_04931_, _04930_, _04830_);
  nor _27975_ (_04932_, _04931_, _01227_);
  and _27976_ (_04933_, _04931_, _01227_);
  or _27977_ (_04934_, _04933_, _04932_);
  or _27978_ (_04935_, _04934_, _04882_);
  and _27979_ (_04936_, _04741_, _04742_);
  and _27980_ (_04937_, _04936_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _27981_ (_04938_, _04937_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _27982_ (_04939_, _04937_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _27983_ (_04940_, _04939_, _04938_);
  nor _27984_ (_04942_, _04940_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _27985_ (_04944_, _04940_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor _27986_ (_04946_, _04944_, _04942_);
  nor _27987_ (_04947_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and _27988_ (_04948_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08682_);
  nor _27989_ (_04949_, _04948_, _04947_);
  and _27990_ (_04950_, _04949_, _04846_);
  nor _27991_ (_04951_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and _27992_ (_04952_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08687_);
  nor _27993_ (_04953_, _04952_, _04951_);
  and _27994_ (_04954_, _04953_, _04736_);
  nor _27995_ (_04955_, _04954_, _04950_);
  nor _27996_ (_04956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and _27997_ (_04957_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08693_);
  nor _27998_ (_04958_, _04957_, _04956_);
  and _27999_ (_04959_, _04958_, _04779_);
  nor _28000_ (_04960_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and _28001_ (_04961_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08698_);
  nor _28002_ (_04962_, _04961_, _04960_);
  and _28003_ (_04963_, _04962_, _04795_);
  nor _28004_ (_04964_, _04963_, _04959_);
  and _28005_ (_04965_, _04964_, _04955_);
  nor _28006_ (_04966_, _04965_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not _28007_ (_04967_, _04966_);
  nor _28008_ (_04968_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and _28009_ (_04969_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08663_);
  nor _28010_ (_04970_, _04969_, _04968_);
  and _28011_ (_04971_, _04970_, _04846_);
  nor _28012_ (_04972_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and _28013_ (_04973_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08669_);
  nor _28014_ (_04974_, _04973_, _04972_);
  and _28015_ (_04975_, _04974_, _04779_);
  nor _28016_ (_04976_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and _28017_ (_04977_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08674_);
  nor _28018_ (_04979_, _04977_, _04976_);
  and _28019_ (_04980_, _04979_, _04795_);
  nor _28020_ (_04981_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and _28021_ (_04982_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08657_);
  nor _28022_ (_04983_, _04982_, _04981_);
  and _28023_ (_04984_, _04983_, _04736_);
  or _28024_ (_04985_, _04984_, _04980_);
  or _28025_ (_04986_, _04985_, _04975_);
  nor _28026_ (_04987_, _04986_, _04971_);
  or _28027_ (_04988_, _04987_, _01350_);
  and _28028_ (_04989_, _04988_, _04967_);
  not _28029_ (_04991_, _04989_);
  and _28030_ (_04992_, _04991_, _04830_);
  nor _28031_ (_04993_, _04992_, _01220_);
  and _28032_ (_04994_, _04992_, _01220_);
  or _28033_ (_04995_, _04994_, _04993_);
  or _28034_ (_04996_, _04995_, _04946_);
  or _28035_ (_04997_, _04996_, _04935_);
  or _28036_ (_04998_, _04997_, _04778_);
  or _28037_ (_04999_, _04998_, _04735_);
  or _28038_ (_05000_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  not _28039_ (_05001_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _28040_ (_05003_, _05001_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and _28041_ (_05004_, _05003_, _05000_);
  and _28042_ (_05005_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _04503_);
  and _28043_ (_05006_, _05005_, _05004_);
  or _28044_ (_05007_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and _28045_ (_05008_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _28046_ (_05009_, _05001_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _28047_ (_05010_, _05009_, _05008_);
  and _28048_ (_05011_, _05010_, _05007_);
  or _28049_ (_05012_, _05011_, _05006_);
  not _28050_ (_05013_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor _28051_ (_05014_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _28052_ (_05015_, _05014_, _04503_);
  nor _28053_ (_05016_, _05015_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _28054_ (_05017_, _05015_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _28055_ (_05019_, _05017_, _05016_);
  and _28056_ (_05020_, _05019_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _28057_ (_05021_, _05014_, _04503_);
  nor _28058_ (_05022_, _05021_, _05015_);
  or _28059_ (_05023_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _08615_);
  nand _28060_ (_05024_, _05023_, _05022_);
  or _28061_ (_05025_, _05024_, _05020_);
  and _28062_ (_05026_, _05025_, _05013_);
  nand _28063_ (_05027_, _05019_, _04336_);
  or _28064_ (_05028_, _05019_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _28065_ (_05029_, _05028_, _05027_);
  or _28066_ (_05030_, _05022_, _05029_);
  and _28067_ (_05031_, _05030_, _05026_);
  or _28068_ (_05032_, _05031_, _05012_);
  and _28069_ (_05034_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _28070_ (_05035_, _05001_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _28071_ (_05036_, _05035_, _05034_);
  and _28072_ (_05037_, _05036_, _04503_);
  and _28073_ (_05038_, _05001_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and _28074_ (_05039_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or _28075_ (_05040_, _05039_, _05038_);
  and _28076_ (_05041_, _05040_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _28077_ (_05042_, _05041_, _05037_);
  and _28078_ (_05043_, _05042_, _05013_);
  and _28079_ (_05044_, _05008_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _28080_ (_05045_, _05044_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _28081_ (_05046_, _05044_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _28082_ (_05047_, _05046_, _05045_);
  nand _28083_ (_05048_, _05047_, _08593_);
  and _28084_ (_05049_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor _28085_ (_05050_, _05049_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor _28086_ (_05051_, _05050_, _05044_);
  and _28087_ (_05052_, _05051_, _05000_);
  and _28088_ (_05053_, _05052_, _05048_);
  nand _28089_ (_05054_, _05047_, _08621_);
  not _28090_ (_05055_, _05051_);
  or _28091_ (_05056_, _05047_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and _28092_ (_05057_, _05056_, _05055_);
  and _28093_ (_05058_, _05057_, _05054_);
  or _28094_ (_05059_, _05058_, _05053_);
  and _28095_ (_05060_, _05059_, _05043_);
  nand _28096_ (_05061_, _05047_, _04329_);
  or _28097_ (_05062_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and _28098_ (_05063_, _05062_, _05051_);
  and _28099_ (_05064_, _05063_, _05061_);
  nand _28100_ (_05065_, _05047_, _04336_);
  or _28101_ (_05066_, _05047_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and _28102_ (_05067_, _05066_, _05055_);
  and _28103_ (_05068_, _05067_, _05065_);
  or _28104_ (_05069_, _05068_, _05064_);
  and _28105_ (_05070_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  and _28106_ (_05071_, _05001_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or _28107_ (_05072_, _05071_, _04503_);
  or _28108_ (_05073_, _05072_, _05070_);
  or _28109_ (_05074_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or _28110_ (_05075_, _05001_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and _28111_ (_05076_, _05075_, _05074_);
  or _28112_ (_05077_, _05076_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _28113_ (_05078_, _05077_, _05073_);
  and _28114_ (_05079_, _05078_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _28115_ (_05080_, _05040_, _05005_);
  or _28116_ (_05081_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or _28117_ (_05082_, _05001_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and _28118_ (_05083_, _05082_, _05008_);
  and _28119_ (_05084_, _05083_, _05081_);
  or _28120_ (_05085_, _05084_, _05080_);
  and _28121_ (_05086_, _05085_, _05079_);
  and _28122_ (_05087_, _05086_, _05069_);
  or _28123_ (_05088_, _05087_, _05060_);
  or _28124_ (_05089_, _05085_, _05078_);
  and _28125_ (_05090_, _05089_, _04416_);
  and _28126_ (_05091_, _05090_, _05088_);
  and _28127_ (_05092_, _05091_, _05032_);
  or _28128_ (_05093_, _05013_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or _28129_ (_05094_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and _28130_ (_05095_, _05094_, _05093_);
  or _28131_ (_05096_, _05095_, _05019_);
  or _28132_ (_05097_, _05013_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or _28133_ (_05098_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand _28134_ (_05099_, _05098_, _05097_);
  and _28135_ (_05100_, _05099_, _05019_);
  nor _28136_ (_05101_, _05100_, _05022_);
  and _28137_ (_05102_, _05101_, _05096_);
  and _28138_ (_05103_, _05019_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or _28139_ (_05104_, _05038_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or _28140_ (_05105_, _05104_, _05103_);
  and _28141_ (_05106_, _05019_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or _28142_ (_05107_, _05071_, _05013_);
  or _28143_ (_05108_, _05107_, _05106_);
  and _28144_ (_05109_, _05108_, _05022_);
  and _28145_ (_05110_, _05109_, _05105_);
  or _28146_ (_05111_, _05110_, _05102_);
  nand _28147_ (_05112_, _05047_, _04359_);
  or _28148_ (_05113_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  and _28149_ (_05114_, _05113_, _05112_);
  or _28150_ (_05115_, _05114_, _05055_);
  or _28151_ (_05116_, _05047_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand _28152_ (_05117_, _05047_, _04366_);
  and _28153_ (_05118_, _05117_, _05116_);
  or _28154_ (_05119_, _05118_, _05051_);
  and _28155_ (_05120_, _05119_, _05115_);
  or _28156_ (_05121_, _05120_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and _28157_ (_05122_, _05047_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _28158_ (_05123_, _05047_, _08639_);
  or _28159_ (_05124_, _05123_, _05122_);
  and _28160_ (_05125_, _05124_, _05055_);
  nand _28161_ (_05126_, _05047_, _08647_);
  or _28162_ (_05127_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  and _28163_ (_05128_, _05127_, _05051_);
  and _28164_ (_05129_, _05128_, _05126_);
  or _28165_ (_05130_, _05129_, _05013_);
  or _28166_ (_05131_, _05130_, _05125_);
  or _28167_ (_05132_, _05001_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and _28168_ (_05133_, _05062_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _28169_ (_05134_, _05133_, _05132_);
  or _28170_ (_05135_, _05001_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or _28171_ (_05136_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  and _28172_ (_05137_, _05136_, _04503_);
  and _28173_ (_05138_, _05137_, _05135_);
  or _28174_ (_05139_, _05138_, _05134_);
  and _28175_ (_05140_, _05139_, _05049_);
  and _28176_ (_05141_, _05013_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _28177_ (_05142_, _05004_, _04503_);
  or _28178_ (_05143_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or _28179_ (_05144_, _05001_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and _28180_ (_05145_, _05144_, _05143_);
  or _28181_ (_05146_, _05145_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _28182_ (_05147_, _05146_, _05142_);
  and _28183_ (_05148_, _05147_, _05141_);
  or _28184_ (_05149_, _05148_, _05140_);
  and _28185_ (_05150_, _05139_, _05013_);
  or _28186_ (_05151_, _05150_, _05012_);
  and _28187_ (_05152_, _05151_, _05149_);
  and _28188_ (_05153_, _05152_, _05131_);
  and _28189_ (_05154_, _05153_, _05121_);
  and _28190_ (_05155_, _05154_, _05111_);
  or _28191_ (_05156_, _05155_, _05092_);
  nor _28192_ (_05157_, _04307_, _01231_);
  and _28193_ (_05158_, _04795_, _13921_);
  nor _28194_ (_05159_, _05158_, _05157_);
  and _28195_ (_05160_, _05157_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _28196_ (_05161_, _05157_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _28197_ (_05162_, _05161_, _05160_);
  and _28198_ (_05163_, _05162_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _28199_ (_05164_, _05162_, _08967_);
  or _28200_ (_05165_, _05164_, _05163_);
  and _28201_ (_05166_, _05165_, _04327_);
  or _28202_ (_05167_, _05166_, _05159_);
  and _28203_ (_05168_, _05162_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not _28204_ (_05169_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor _28205_ (_05170_, _05162_, _05169_);
  or _28206_ (_05171_, _05170_, _05168_);
  and _28207_ (_05172_, _05171_, _04309_);
  and _28208_ (_05173_, _05162_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor _28209_ (_05174_, _05162_, _08608_);
  or _28210_ (_05175_, _05174_, _05173_);
  and _28211_ (_05176_, _05175_, _04307_);
  and _28212_ (_05177_, _05162_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor _28213_ (_05178_, _05162_, _08639_);
  or _28214_ (_05179_, _05178_, _05177_);
  and _28215_ (_05180_, _05179_, _04357_);
  or _28216_ (_05181_, _05180_, _05176_);
  or _28217_ (_05182_, _05181_, _05172_);
  or _28218_ (_05183_, _05182_, _05167_);
  or _28219_ (_05184_, _05162_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor _28220_ (_05185_, _04780_, _04328_);
  nand _28221_ (_05186_, _05185_, _05184_);
  nand _28222_ (_05187_, _05186_, _05159_);
  or _28223_ (_05188_, _05162_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor _28224_ (_05189_, _04806_, _04344_);
  and _28225_ (_05190_, _05189_, _05188_);
  or _28226_ (_05191_, _05162_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor _28227_ (_05192_, _04786_, _04308_);
  and _28228_ (_05193_, _05192_, _05191_);
  or _28229_ (_05194_, _05162_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor _28230_ (_05195_, _04823_, _04358_);
  and _28231_ (_05196_, _05195_, _05194_);
  or _28232_ (_05197_, _05196_, _05193_);
  or _28233_ (_05198_, _05197_, _05190_);
  or _28234_ (_05199_, _05198_, _05187_);
  nor _28235_ (_05200_, _04793_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _28236_ (_05201_, _04846_, _04782_);
  nor _28237_ (_05202_, _05201_, _13921_);
  not _28238_ (_05203_, _05202_);
  nor _28239_ (_05204_, _05203_, _05200_);
  nor _28240_ (_05205_, _04814_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and _28241_ (_05206_, _04846_, _04825_);
  nor _28242_ (_05207_, _05206_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  not _28243_ (_05208_, _05207_);
  nor _28244_ (_05209_, _05208_, _05205_);
  nor _28245_ (_05210_, _05209_, _05204_);
  not _28246_ (_05211_, _05210_);
  or _28247_ (_05212_, _01350_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or _28248_ (_05213_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and _28249_ (_05214_, _05213_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and _28250_ (_05215_, _05214_, _05212_);
  and _28251_ (_05216_, _05215_, _04327_);
  and _28252_ (_05217_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08967_);
  nor _28253_ (_05218_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  nor _28254_ (_05219_, _05218_, _05217_);
  and _28255_ (_05220_, _05219_, _04310_);
  nor _28256_ (_05221_, _05220_, _05216_);
  and _28257_ (_05222_, _05221_, _05211_);
  not _28258_ (_05223_, _08139_);
  nor _28259_ (_05224_, _05223_, first_instr);
  nand _28260_ (_05225_, _05224_, _04830_);
  nor _28261_ (_05226_, _05225_, _05222_);
  and _28262_ (_05227_, _05226_, _05199_);
  and _28263_ (_05228_, _05227_, _05183_);
  and _28264_ (_05229_, _05228_, _04417_);
  and _28265_ (_05230_, _05229_, _05156_);
  nor _28266_ (_05231_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28267_ (_05232_, _10057_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28268_ (_05233_, _05232_, _05231_);
  and _28269_ (_05234_, _05233_, _04846_);
  nor _28270_ (_05235_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28271_ (_05236_, _10290_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28272_ (_05237_, _05236_, _05235_);
  and _28273_ (_05238_, _05237_, _04779_);
  nor _28274_ (_05239_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28275_ (_05240_, _09807_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28276_ (_05241_, _05240_, _05239_);
  and _28277_ (_05242_, _05241_, _04795_);
  nor _28278_ (_05243_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28279_ (_05244_, _10501_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28280_ (_05245_, _05244_, _05243_);
  and _28281_ (_05246_, _05245_, _04736_);
  or _28282_ (_05247_, _05246_, _05242_);
  or _28283_ (_05248_, _05247_, _05238_);
  or _28284_ (_05249_, _05248_, _05234_);
  and _28285_ (_05250_, _05249_, _01350_);
  nor _28286_ (_05251_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28287_ (_05252_, _11260_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28288_ (_05253_, _05252_, _05251_);
  and _28289_ (_05254_, _05253_, _04846_);
  nor _28290_ (_05255_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28291_ (_05256_, _12474_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28292_ (_05257_, _05256_, _05255_);
  and _28293_ (_05258_, _05257_, _04779_);
  nor _28294_ (_05259_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28295_ (_05260_, _10710_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28296_ (_05261_, _05260_, _05259_);
  and _28297_ (_05262_, _05261_, _04795_);
  nor _28298_ (_05263_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28299_ (_05264_, _12861_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28300_ (_05265_, _05264_, _05263_);
  and _28301_ (_05266_, _05265_, _04736_);
  or _28302_ (_05267_, _05266_, _05262_);
  or _28303_ (_05268_, _05267_, _05258_);
  or _28304_ (_05269_, _05268_, _05254_);
  and _28305_ (_05270_, _05269_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _28306_ (_05271_, _05270_, _05250_);
  and _28307_ (_05272_, _05271_, _04830_);
  nor _28308_ (_05273_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28309_ (_05274_, _10072_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28310_ (_05275_, _05274_, _05273_);
  and _28311_ (_05276_, _05275_, _04846_);
  nor _28312_ (_05277_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28313_ (_05278_, _10301_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28314_ (_05279_, _05278_, _05277_);
  and _28315_ (_05280_, _05279_, _04779_);
  nor _28316_ (_05281_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28317_ (_05282_, _09821_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28318_ (_05283_, _05282_, _05281_);
  and _28319_ (_05284_, _05283_, _04795_);
  nor _28320_ (_05285_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28321_ (_05286_, _10512_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28322_ (_05287_, _05286_, _05285_);
  and _28323_ (_05288_, _05287_, _04736_);
  or _28324_ (_05289_, _05288_, _05284_);
  or _28325_ (_05290_, _05289_, _05280_);
  or _28326_ (_05291_, _05290_, _05276_);
  and _28327_ (_05292_, _05291_, _01350_);
  nor _28328_ (_05293_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28329_ (_05294_, _12185_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28330_ (_05295_, _05294_, _05293_);
  and _28331_ (_05296_, _05295_, _04846_);
  nor _28332_ (_05297_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28333_ (_05298_, _12488_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28334_ (_05299_, _05298_, _05297_);
  and _28335_ (_05300_, _05299_, _04779_);
  nor _28336_ (_05301_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28337_ (_05302_, _10727_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28338_ (_05303_, _05302_, _05301_);
  and _28339_ (_05304_, _05303_, _04795_);
  nor _28340_ (_05305_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28341_ (_05306_, _12874_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28342_ (_05307_, _05306_, _05305_);
  and _28343_ (_05308_, _05307_, _04736_);
  or _28344_ (_05309_, _05308_, _05304_);
  or _28345_ (_05310_, _05309_, _05300_);
  or _28346_ (_05311_, _05310_, _05296_);
  and _28347_ (_05312_, _05311_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _28348_ (_05313_, _05312_, _05292_);
  and _28349_ (_05314_, _05313_, _04830_);
  nor _28350_ (_05315_, _05314_, _05272_);
  nor _28351_ (_05316_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28352_ (_05317_, _10474_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28353_ (_05318_, _05317_, _05316_);
  and _28354_ (_05319_, _05318_, _04736_);
  nor _28355_ (_05320_, _05319_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor _28356_ (_05321_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28357_ (_05322_, _09771_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28358_ (_05323_, _05322_, _05321_);
  and _28359_ (_05324_, _05323_, _04795_);
  not _28360_ (_05325_, _05324_);
  nor _28361_ (_05326_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28362_ (_05327_, _10016_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28363_ (_05328_, _05327_, _05326_);
  and _28364_ (_05329_, _05328_, _04846_);
  nor _28365_ (_05330_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28366_ (_05331_, _10263_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28367_ (_05332_, _05331_, _05330_);
  and _28368_ (_05333_, _05332_, _04779_);
  nor _28369_ (_05334_, _05333_, _05329_);
  and _28370_ (_05335_, _05334_, _05325_);
  and _28371_ (_05336_, _05335_, _05320_);
  nor _28372_ (_05337_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28373_ (_05338_, _12833_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28374_ (_05339_, _05338_, _05337_);
  and _28375_ (_05340_, _05339_, _04736_);
  nor _28376_ (_05341_, _05340_, _01350_);
  nor _28377_ (_05342_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28378_ (_05343_, _10685_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28379_ (_05344_, _05343_, _05342_);
  and _28380_ (_05345_, _05344_, _04795_);
  not _28381_ (_05346_, _05345_);
  nor _28382_ (_05347_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28383_ (_05348_, _11230_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28384_ (_05349_, _05348_, _05347_);
  and _28385_ (_05350_, _05349_, _04846_);
  nor _28386_ (_05351_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28387_ (_05352_, _12448_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28388_ (_05353_, _05352_, _05351_);
  and _28389_ (_05354_, _05353_, _04779_);
  nor _28390_ (_05355_, _05354_, _05350_);
  and _28391_ (_05356_, _05355_, _05346_);
  and _28392_ (_05357_, _05356_, _05341_);
  nor _28393_ (_05358_, _05357_, _05336_);
  and _28394_ (_05359_, _05358_, _04830_);
  not _28395_ (_05360_, _05359_);
  nor _28396_ (_05361_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28397_ (_05362_, _10037_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28398_ (_05363_, _05362_, _05361_);
  and _28399_ (_05364_, _05363_, _04846_);
  nor _28400_ (_05365_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28401_ (_05366_, _10276_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28402_ (_05367_, _05366_, _05365_);
  and _28403_ (_05368_, _05367_, _04779_);
  nor _28404_ (_05369_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28405_ (_05370_, _09792_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28406_ (_05371_, _05370_, _05369_);
  and _28407_ (_05372_, _05371_, _04795_);
  nor _28408_ (_05373_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28409_ (_05374_, _10489_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28410_ (_05375_, _05374_, _05373_);
  and _28411_ (_05376_, _05375_, _04736_);
  or _28412_ (_05377_, _05376_, _05372_);
  or _28413_ (_05378_, _05377_, _05368_);
  or _28414_ (_05379_, _05378_, _05364_);
  and _28415_ (_05380_, _05379_, _01350_);
  nor _28416_ (_05381_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28417_ (_05382_, _11247_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28418_ (_05383_, _05382_, _05381_);
  and _28419_ (_05384_, _05383_, _04846_);
  nor _28420_ (_05385_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28421_ (_05386_, _12463_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28422_ (_05387_, _05386_, _05385_);
  and _28423_ (_05388_, _05387_, _04779_);
  nor _28424_ (_05389_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28425_ (_05390_, _10699_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28426_ (_05391_, _05390_, _05389_);
  and _28427_ (_05392_, _05391_, _04795_);
  nor _28428_ (_05393_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28429_ (_05394_, _12848_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28430_ (_05395_, _05394_, _05393_);
  and _28431_ (_05396_, _05395_, _04736_);
  or _28432_ (_05397_, _05396_, _05392_);
  or _28433_ (_05398_, _05397_, _05388_);
  or _28434_ (_05399_, _05398_, _05384_);
  and _28435_ (_05400_, _05399_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or _28436_ (_05401_, _05400_, _05380_);
  nor _28437_ (_05402_, _05401_, _05360_);
  and _28438_ (_05403_, _05402_, _05315_);
  and _28439_ (_05404_, _05403_, _05230_);
  and _28440_ (property_invalid_ajmp, _05404_, _04999_);
  and _28441_ (_05405_, _04736_, _01350_);
  nor _28442_ (_05406_, _04736_, _01350_);
  nor _28443_ (_05407_, _05406_, _05405_);
  not _28444_ (_05408_, _05407_);
  and _28445_ (_05409_, _04846_, _04839_);
  or _28446_ (_05410_, _05409_, _05408_);
  and _28447_ (_05411_, _04833_, _04736_);
  and _28448_ (_05412_, _04845_, _04795_);
  and _28449_ (_05413_, _04851_, _04779_);
  or _28450_ (_05414_, _05413_, _05412_);
  or _28451_ (_05415_, _05414_, _05411_);
  or _28452_ (_05416_, _05415_, _05410_);
  and _28453_ (_05417_, _04863_, _04846_);
  or _28454_ (_05418_, _05417_, _05407_);
  and _28455_ (_05419_, _04858_, _04736_);
  and _28456_ (_05420_, _04868_, _04795_);
  and _28457_ (_05421_, _04873_, _04779_);
  or _28458_ (_05422_, _05421_, _05420_);
  or _28459_ (_05423_, _05422_, _05419_);
  or _28460_ (_05424_, _05423_, _05418_);
  nand _28461_ (_05425_, _05424_, _05416_);
  nor _28462_ (_05426_, _05425_, _05222_);
  nand _28463_ (_05427_, _05426_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  or _28464_ (_05428_, _05426_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and _28465_ (_05429_, _05428_, _05427_);
  nor _28466_ (_05430_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28467_ (_05431_, _10315_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28468_ (_05432_, _05431_, _05430_);
  and _28469_ (_05433_, _05432_, _04846_);
  or _28470_ (_05434_, _05433_, _05408_);
  nor _28471_ (_05435_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28472_ (_05436_, _09834_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28473_ (_05437_, _05436_, _05435_);
  and _28474_ (_05438_, _05437_, _04736_);
  nor _28475_ (_05439_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28476_ (_05440_, _10086_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28477_ (_05441_, _05440_, _05439_);
  and _28478_ (_05442_, _05441_, _04795_);
  nor _28479_ (_05443_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28480_ (_05444_, _10525_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28481_ (_05445_, _05444_, _05443_);
  and _28482_ (_05446_, _05445_, _04779_);
  or _28483_ (_05447_, _05446_, _05442_);
  or _28484_ (_05448_, _05447_, _05438_);
  or _28485_ (_05449_, _05448_, _05434_);
  nor _28486_ (_05450_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28487_ (_05451_, _12501_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28488_ (_05452_, _05451_, _05450_);
  and _28489_ (_05453_, _05452_, _04846_);
  or _28490_ (_05454_, _05453_, _05407_);
  nor _28491_ (_05455_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28492_ (_05456_, _10743_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28493_ (_05457_, _05456_, _05455_);
  and _28494_ (_05458_, _05457_, _04736_);
  nor _28495_ (_05459_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28496_ (_05460_, _12196_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28497_ (_05461_, _05460_, _05459_);
  and _28498_ (_05462_, _05461_, _04795_);
  nor _28499_ (_05463_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28500_ (_05464_, _12887_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28501_ (_05465_, _05464_, _05463_);
  and _28502_ (_05466_, _05465_, _04779_);
  or _28503_ (_05467_, _05466_, _05462_);
  or _28504_ (_05468_, _05467_, _05458_);
  or _28505_ (_05469_, _05468_, _05454_);
  nand _28506_ (_05470_, _05469_, _05449_);
  nor _28507_ (_05471_, _05470_, _05222_);
  nand _28508_ (_05472_, _05471_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or _28509_ (_05473_, _05471_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and _28510_ (_05474_, _05473_, _05472_);
  or _28511_ (_05475_, _05474_, _05429_);
  and _28512_ (_05476_, _04958_, _04846_);
  or _28513_ (_05477_, _05476_, _05408_);
  and _28514_ (_05478_, _04962_, _04736_);
  and _28515_ (_05479_, _04949_, _04795_);
  and _28516_ (_05480_, _04953_, _04779_);
  or _28517_ (_05481_, _05480_, _05479_);
  or _28518_ (_05482_, _05481_, _05478_);
  or _28519_ (_05483_, _05482_, _05477_);
  and _28520_ (_05484_, _04974_, _04846_);
  or _28521_ (_05485_, _05484_, _05407_);
  and _28522_ (_05486_, _04979_, _04736_);
  and _28523_ (_05487_, _04970_, _04795_);
  and _28524_ (_05488_, _04983_, _04779_);
  or _28525_ (_05489_, _05488_, _05487_);
  or _28526_ (_05490_, _05489_, _05486_);
  or _28527_ (_05491_, _05490_, _05485_);
  nand _28528_ (_05492_, _05491_, _05483_);
  nor _28529_ (_05493_, _05492_, _05222_);
  nor _28530_ (_05494_, _05493_, _01149_);
  and _28531_ (_05495_, _05493_, _01149_);
  or _28532_ (_05496_, _05495_, _05494_);
  not _28533_ (_05497_, _05222_);
  and _28534_ (_05498_, _04907_, _04795_);
  and _28535_ (_05499_, _04923_, _04779_);
  and _28536_ (_05500_, _04912_, _04846_);
  and _28537_ (_05501_, _04917_, _04736_);
  or _28538_ (_05502_, _05501_, _05500_);
  or _28539_ (_05503_, _05502_, _05499_);
  or _28540_ (_05504_, _05503_, _05498_);
  and _28541_ (_05505_, _05504_, _05408_);
  and _28542_ (_05506_, _04885_, _04795_);
  and _28543_ (_05507_, _04899_, _04779_);
  and _28544_ (_05508_, _04894_, _04736_);
  and _28545_ (_05509_, _04890_, _04846_);
  or _28546_ (_05510_, _05509_, _05508_);
  or _28547_ (_05511_, _05510_, _05507_);
  or _28548_ (_05512_, _05511_, _05506_);
  and _28549_ (_05513_, _05512_, _05407_);
  or _28550_ (_05514_, _05513_, _05505_);
  and _28551_ (_05515_, _05514_, _05497_);
  and _28552_ (_05516_, _05515_, _01188_);
  nor _28553_ (_05517_, _05515_, _01188_);
  or _28554_ (_05518_, _05517_, _05516_);
  or _28555_ (_05519_, _05518_, _05496_);
  or _28556_ (_05520_, _05519_, _05475_);
  and _28557_ (_05521_, _05349_, _04795_);
  and _28558_ (_05522_, _05339_, _04779_);
  and _28559_ (_05523_, _05344_, _04736_);
  and _28560_ (_05524_, _05353_, _04846_);
  or _28561_ (_05525_, _05524_, _05523_);
  or _28562_ (_05526_, _05525_, _05522_);
  or _28563_ (_05527_, _05526_, _05521_);
  and _28564_ (_05528_, _05527_, _05408_);
  and _28565_ (_05529_, _05328_, _04795_);
  and _28566_ (_05530_, _05318_, _04779_);
  and _28567_ (_05531_, _05323_, _04736_);
  and _28568_ (_05532_, _05332_, _04846_);
  or _28569_ (_05533_, _05532_, _05531_);
  or _28570_ (_05534_, _05533_, _05530_);
  or _28571_ (_05535_, _05534_, _05529_);
  and _28572_ (_05536_, _05535_, _05407_);
  or _28573_ (_05537_, _05536_, _05528_);
  and _28574_ (_05538_, _05537_, _05497_);
  nand _28575_ (_05539_, _05538_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or _28576_ (_05540_, _05538_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  and _28577_ (_05541_, _05540_, _05539_);
  and _28578_ (_05542_, _05367_, _04846_);
  and _28579_ (_05543_, _05375_, _04779_);
  and _28580_ (_05544_, _05371_, _04736_);
  or _28581_ (_05545_, _05544_, _05543_);
  or _28582_ (_05546_, _05545_, _05542_);
  and _28583_ (_05547_, _05363_, _04795_);
  or _28584_ (_05548_, _05547_, _05408_);
  or _28585_ (_05549_, _05548_, _05546_);
  and _28586_ (_05550_, _05387_, _04846_);
  or _28587_ (_05551_, _05550_, _05407_);
  and _28588_ (_05552_, _05391_, _04736_);
  and _28589_ (_05553_, _05383_, _04795_);
  and _28590_ (_05554_, _05395_, _04779_);
  or _28591_ (_05555_, _05554_, _05553_);
  or _28592_ (_05556_, _05555_, _05552_);
  or _28593_ (_05557_, _05556_, _05551_);
  nand _28594_ (_05558_, _05557_, _05549_);
  nor _28595_ (_05559_, _05558_, _05222_);
  nor _28596_ (_05560_, _05559_, _05013_);
  and _28597_ (_05561_, _05559_, _05013_);
  or _28598_ (_05562_, _05561_, _05560_);
  or _28599_ (_05563_, _05562_, _05541_);
  and _28600_ (_05564_, _05253_, _04795_);
  and _28601_ (_05565_, _05265_, _04779_);
  and _28602_ (_05566_, _05261_, _04736_);
  and _28603_ (_05567_, _05257_, _04846_);
  or _28604_ (_05568_, _05567_, _05566_);
  or _28605_ (_05569_, _05568_, _05565_);
  or _28606_ (_05570_, _05569_, _05564_);
  and _28607_ (_05571_, _05570_, _05408_);
  and _28608_ (_05572_, _05233_, _04795_);
  and _28609_ (_05573_, _05245_, _04779_);
  and _28610_ (_05574_, _05237_, _04846_);
  and _28611_ (_05575_, _05241_, _04736_);
  or _28612_ (_05576_, _05575_, _05574_);
  or _28613_ (_05577_, _05576_, _05573_);
  or _28614_ (_05578_, _05577_, _05572_);
  and _28615_ (_05579_, _05578_, _05407_);
  or _28616_ (_05580_, _05579_, _05571_);
  and _28617_ (_05581_, _05580_, _05497_);
  nand _28618_ (_05582_, _05581_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _28619_ (_05583_, _05581_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _28620_ (_05584_, _05583_, _05582_);
  and _28621_ (_05585_, _05279_, _04846_);
  or _28622_ (_05586_, _05585_, _05408_);
  and _28623_ (_05587_, _05283_, _04736_);
  and _28624_ (_05588_, _05275_, _04795_);
  and _28625_ (_05589_, _05287_, _04779_);
  or _28626_ (_05590_, _05589_, _05588_);
  or _28627_ (_05591_, _05590_, _05587_);
  or _28628_ (_05592_, _05591_, _05586_);
  and _28629_ (_05593_, _05295_, _04795_);
  and _28630_ (_05594_, _05299_, _04846_);
  or _28631_ (_05595_, _05594_, _05593_);
  and _28632_ (_05596_, _05303_, _04736_);
  and _28633_ (_05597_, _05307_, _04779_);
  or _28634_ (_05598_, _05597_, _05407_);
  or _28635_ (_05599_, _05598_, _05596_);
  or _28636_ (_05600_, _05599_, _05595_);
  nand _28637_ (_05601_, _05600_, _05592_);
  nor _28638_ (_05602_, _05601_, _05222_);
  nand _28639_ (_05603_, _05602_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _28640_ (_05604_, _05602_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _28641_ (_05605_, _05604_, _05603_);
  or _28642_ (_05606_, _05605_, _05584_);
  or _28643_ (_05607_, _05606_, _05563_);
  or _28644_ (_05608_, _05607_, _05520_);
  or _28645_ (_05609_, _04412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _28646_ (_05610_, _04412_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _28647_ (_05611_, _05610_, _05609_);
  and _28648_ (_05612_, _04455_, _01144_);
  nor _28649_ (_05613_, _04455_, _01144_);
  or _28650_ (_05614_, _05613_, _05612_);
  or _28651_ (_05615_, _05614_, _05611_);
  or _28652_ (_05616_, _04499_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand _28653_ (_05617_, _04499_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and _28654_ (_05618_, _05617_, _05616_);
  nor _28655_ (_05619_, _04548_, _01220_);
  and _28656_ (_05620_, _04548_, _01220_);
  or _28657_ (_05621_, _05620_, _05619_);
  or _28658_ (_05622_, _05621_, _05618_);
  or _28659_ (_05623_, _05622_, _05615_);
  or _28660_ (_05624_, _04604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand _28661_ (_05625_, _04604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and _28662_ (_05626_, _05625_, _05624_);
  nor _28663_ (_05627_, _04646_, _00687_);
  and _28664_ (_05628_, _04646_, _00687_);
  or _28665_ (_05629_, _05628_, _05627_);
  or _28666_ (_05630_, _05629_, _05626_);
  and _28667_ (_05631_, _04729_, _00659_);
  nor _28668_ (_05632_, _04729_, _00659_);
  or _28669_ (_05633_, _05632_, _05631_);
  and _28670_ (_05634_, _04688_, _00619_);
  nor _28671_ (_05635_, _04688_, _00619_);
  or _28672_ (_05636_, _05635_, _05634_);
  or _28673_ (_05637_, _05636_, _05633_);
  or _28674_ (_05638_, _05637_, _05630_);
  or _28675_ (_05639_, _05638_, _05623_);
  or _28676_ (_05640_, _05639_, _05608_);
  nor _28677_ (_05641_, _04992_, _04931_);
  not _28678_ (_05642_, _04879_);
  and _28679_ (_05643_, _05401_, _04830_);
  and _28680_ (_05644_, _05360_, _05315_);
  and _28681_ (_05645_, _05644_, _05643_);
  and _28682_ (_05646_, _05645_, _05642_);
  and _28683_ (_05647_, _05646_, _05641_);
  and _28684_ (_05648_, _05647_, _05230_);
  and _28685_ (property_invalid_ljmp, _05648_, _05640_);
  and _28686_ (_05649_, _04688_, _04773_);
  nor _28687_ (_05650_, _04688_, _04773_);
  nor _28688_ (_05651_, _05650_, _05649_);
  and _28689_ (_05652_, _04688_, _04762_);
  nor _28690_ (_05653_, _04688_, _04762_);
  and _28691_ (_05654_, _04688_, _04767_);
  and _28692_ (_05655_, _04940_, _04688_);
  nor _28693_ (_05656_, _04940_, _04688_);
  nor _28694_ (_05657_, _04936_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _28695_ (_05658_, _05657_, _04937_);
  and _28696_ (_05659_, _05658_, _04688_);
  nor _28697_ (_05660_, _05658_, _04688_);
  nor _28698_ (_05661_, _05660_, _05659_);
  and _28699_ (_05662_, _04741_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _28700_ (_05663_, _05662_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _28701_ (_05664_, _05663_, _04936_);
  and _28702_ (_05665_, _05664_, _04688_);
  nor _28703_ (_05666_, _05664_, _04688_);
  nor _28704_ (_05667_, _04741_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _28705_ (_05668_, _05667_, _05662_);
  and _28706_ (_05669_, _05668_, _04688_);
  nor _28707_ (_05670_, _04740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _28708_ (_05671_, _05670_, _04741_);
  and _28709_ (_05672_, _05671_, _04688_);
  nor _28710_ (_05673_, _05671_, _04688_);
  nor _28711_ (_05674_, _04739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _28712_ (_05675_, _05674_, _04740_);
  and _28713_ (_05676_, _05675_, _04729_);
  nor _28714_ (_05677_, _05675_, _04729_);
  nor _28715_ (_05678_, _05677_, _05676_);
  not _28716_ (_05679_, _05678_);
  and _28717_ (_05680_, _04737_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _28718_ (_05681_, _05680_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _28719_ (_05682_, _05681_, _04739_);
  and _28720_ (_05683_, _05682_, _04604_);
  nor _28721_ (_05684_, _05682_, _04604_);
  nor _28722_ (_05685_, _05684_, _05683_);
  not _28723_ (_05686_, _05685_);
  nor _28724_ (_05687_, _04737_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _28725_ (_05688_, _05687_, _05680_);
  and _28726_ (_05689_, _05688_, _04646_);
  and _28727_ (_05690_, _04499_, _05408_);
  nor _28728_ (_05691_, _04499_, _05408_);
  nor _28729_ (_05692_, _04846_, _04779_);
  not _28730_ (_05693_, _05692_);
  and _28731_ (_05694_, _05693_, _04548_);
  and _28732_ (_05695_, _04412_, _12949_);
  and _28733_ (_05696_, _04455_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28734_ (_05697_, _04412_, _12949_);
  nor _28735_ (_05698_, _05697_, _05695_);
  and _28736_ (_05699_, _05698_, _05696_);
  nor _28737_ (_05700_, _05699_, _05695_);
  nor _28738_ (_05701_, _05693_, _04548_);
  nor _28739_ (_05702_, _05701_, _05694_);
  not _28740_ (_05703_, _05702_);
  nor _28741_ (_05704_, _05703_, _05700_);
  nor _28742_ (_05705_, _05704_, _05694_);
  nor _28743_ (_05706_, _05705_, _05691_);
  nor _28744_ (_05707_, _05706_, _05690_);
  nor _28745_ (_05708_, _05688_, _04646_);
  nor _28746_ (_05709_, _05708_, _05689_);
  not _28747_ (_05710_, _05709_);
  nor _28748_ (_05711_, _05710_, _05707_);
  nor _28749_ (_05712_, _05711_, _05689_);
  nor _28750_ (_05713_, _05712_, _05686_);
  nor _28751_ (_05714_, _05713_, _05683_);
  nor _28752_ (_05715_, _05714_, _05679_);
  nor _28753_ (_05716_, _05715_, _05676_);
  nor _28754_ (_05717_, _05716_, _05673_);
  or _28755_ (_05718_, _05717_, _05672_);
  nor _28756_ (_05719_, _05668_, _04688_);
  nor _28757_ (_05720_, _05719_, _05669_);
  and _28758_ (_05721_, _05720_, _05718_);
  nor _28759_ (_05722_, _05721_, _05669_);
  nor _28760_ (_05723_, _05722_, _05666_);
  or _28761_ (_05724_, _05723_, _05665_);
  and _28762_ (_05725_, _05724_, _05661_);
  nor _28763_ (_05726_, _05725_, _05659_);
  nor _28764_ (_05727_, _05726_, _05656_);
  or _28765_ (_05728_, _05727_, _05655_);
  nor _28766_ (_05729_, _04688_, _04767_);
  nor _28767_ (_05730_, _05729_, _05654_);
  and _28768_ (_05731_, _05730_, _05728_);
  nor _28769_ (_05732_, _05731_, _05654_);
  nor _28770_ (_05733_, _05732_, _05653_);
  or _28771_ (_05734_, _05733_, _05652_);
  and _28772_ (_05735_, _05734_, _05651_);
  nor _28773_ (_05736_, _05735_, _05649_);
  and _28774_ (_05737_, _04688_, _04751_);
  nor _28775_ (_05738_, _04688_, _04751_);
  or _28776_ (_05739_, _05738_, _05737_);
  and _28777_ (_05740_, _05739_, _05736_);
  nor _28778_ (_05741_, _05739_, _05736_);
  or _28779_ (_05742_, _05741_, _05740_);
  nor _28780_ (_05743_, _05742_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  and _28781_ (_05744_, _05742_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor _28782_ (_05745_, _05734_, _05651_);
  nor _28783_ (_05746_, _05745_, _05735_);
  nor _28784_ (_05747_, _05746_, _00659_);
  and _28785_ (_05748_, _05746_, _00659_);
  not _28786_ (_05749_, _05732_);
  not _28787_ (_05750_, _04688_);
  nand _28788_ (_05751_, _05750_, _04765_);
  or _28789_ (_05752_, _05750_, _04765_);
  and _28790_ (_05753_, _05752_, _05751_);
  nor _28791_ (_05754_, _05753_, _05749_);
  not _28792_ (_05755_, _04946_);
  and _28793_ (_05756_, _05755_, _04688_);
  nor _28794_ (_05757_, _05755_, _04688_);
  nor _28795_ (_05758_, _05757_, _05756_);
  or _28796_ (_05759_, _05758_, _05726_);
  nand _28797_ (_05760_, _05758_, _05726_);
  and _28798_ (_05761_, _05760_, _05759_);
  nor _28799_ (_05762_, _05724_, _05661_);
  nor _28800_ (_05763_, _05762_, _05725_);
  nor _28801_ (_05764_, _05763_, _01220_);
  and _28802_ (_05765_, _05763_, _01220_);
  nor _28803_ (_05766_, _05720_, _05718_);
  nor _28804_ (_05767_, _05766_, _05721_);
  and _28805_ (_05768_, _05767_, _01144_);
  nor _28806_ (_05769_, _05672_, _05673_);
  nor _28807_ (_05770_, _05769_, _05716_);
  and _28808_ (_05771_, _05769_, _05716_);
  nor _28809_ (_05772_, _05771_, _05770_);
  and _28810_ (_05773_, _05772_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor _28811_ (_05774_, _05772_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and _28812_ (_05775_, _05714_, _05679_);
  nor _28813_ (_05776_, _05775_, _05715_);
  and _28814_ (_05777_, _05776_, _01188_);
  nor _28815_ (_05778_, _05776_, _01188_);
  and _28816_ (_05779_, _05712_, _05686_);
  nor _28817_ (_05780_, _05779_, _05713_);
  nor _28818_ (_05781_, _05780_, _01192_);
  and _28819_ (_05782_, _05780_, _01192_);
  and _28820_ (_05783_, _05710_, _05707_);
  nor _28821_ (_05784_, _05783_, _05711_);
  nor _28822_ (_05785_, _05784_, _04608_);
  nor _28823_ (_05786_, _05691_, _05690_);
  and _28824_ (_05787_, _05786_, _05705_);
  nor _28825_ (_05788_, _05786_, _05705_);
  nor _28826_ (_05789_, _05788_, _05787_);
  and _28827_ (_05790_, _05789_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _28828_ (_05791_, _05789_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _28829_ (_05792_, _05703_, _05700_);
  nor _28830_ (_05793_, _05792_, _05704_);
  and _28831_ (_05794_, _05793_, _04503_);
  nor _28832_ (_05795_, _05698_, _05696_);
  nor _28833_ (_05796_, _05795_, _05699_);
  nor _28834_ (_05797_, _05796_, _05013_);
  and _28835_ (_05798_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _28836_ (_05799_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _28837_ (_05800_, _05799_, _05798_);
  not _28838_ (_05801_, _05800_);
  nand _28839_ (_05802_, _05801_, _04455_);
  or _28840_ (_05803_, _05801_, _04455_);
  and _28841_ (_05804_, _05803_, _05802_);
  and _28842_ (_05805_, _05796_, _05013_);
  or _28843_ (_05806_, _05805_, _05804_);
  or _28844_ (_05807_, _05806_, _05797_);
  nor _28845_ (_05808_, _05793_, _04503_);
  or _28846_ (_05809_, _05808_, _05807_);
  or _28847_ (_05810_, _05809_, _05794_);
  or _28848_ (_05811_, _05810_, _05791_);
  or _28849_ (_05812_, _05811_, _05790_);
  and _28850_ (_05813_, _05784_, _04608_);
  or _28851_ (_05814_, _05813_, _05812_);
  or _28852_ (_05815_, _05814_, _05785_);
  or _28853_ (_05816_, _05815_, _05782_);
  or _28854_ (_05817_, _05816_, _05781_);
  or _28855_ (_05818_, _05817_, _05778_);
  or _28856_ (_05819_, _05818_, _05777_);
  or _28857_ (_05820_, _05819_, _05774_);
  or _28858_ (_05821_, _05820_, _05773_);
  or _28859_ (_05822_, _05821_, _05768_);
  or _28860_ (_05823_, _05664_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _28861_ (_05824_, _05664_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _28862_ (_05825_, _05824_, _05823_);
  or _28863_ (_05826_, _05825_, _04688_);
  nand _28864_ (_05827_, _05825_, _04688_);
  and _28865_ (_05828_, _05827_, _05826_);
  and _28866_ (_05829_, _05828_, _05722_);
  nor _28867_ (_05830_, _05767_, _01144_);
  nor _28868_ (_05831_, _05828_, _05722_);
  or _28869_ (_05832_, _05831_, _05830_);
  or _28870_ (_05833_, _05832_, _05829_);
  or _28871_ (_05834_, _05833_, _05822_);
  or _28872_ (_05835_, _05834_, _05765_);
  or _28873_ (_05836_, _05835_, _05764_);
  or _28874_ (_05837_, _05836_, _05761_);
  or _28875_ (_05838_, _05837_, _05754_);
  nor _28876_ (_05839_, _05730_, _05728_);
  nor _28877_ (_05840_, _05839_, _05731_);
  nor _28878_ (_05841_, _05840_, _00687_);
  and _28879_ (_05842_, _05753_, _05749_);
  and _28880_ (_05843_, _05840_, _00687_);
  or _28881_ (_05844_, _05843_, _05842_);
  or _28882_ (_05845_, _05844_, _05841_);
  or _28883_ (_05846_, _05845_, _05838_);
  or _28884_ (_05847_, _05846_, _05748_);
  or _28885_ (_05848_, _05847_, _05747_);
  or _28886_ (_05849_, _05848_, _05744_);
  or _28887_ (_05850_, _05849_, _05743_);
  not _28888_ (_05851_, _04931_);
  and _28889_ (_05852_, _04992_, _05851_);
  and _28890_ (_05853_, _05445_, _04736_);
  nor _28891_ (_05854_, _05853_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and _28892_ (_05855_, _05437_, _04795_);
  not _28893_ (_05856_, _05855_);
  and _28894_ (_05857_, _05441_, _04846_);
  and _28895_ (_05858_, _05432_, _04779_);
  nor _28896_ (_05859_, _05858_, _05857_);
  and _28897_ (_05860_, _05859_, _05856_);
  and _28898_ (_05861_, _05860_, _05854_);
  and _28899_ (_05862_, _05465_, _04736_);
  nor _28900_ (_05863_, _05862_, _01350_);
  and _28901_ (_05864_, _05461_, _04846_);
  not _28902_ (_05865_, _05864_);
  and _28903_ (_05866_, _05452_, _04779_);
  and _28904_ (_05867_, _05457_, _04795_);
  nor _28905_ (_05868_, _05867_, _05866_);
  and _28906_ (_05869_, _05868_, _05865_);
  and _28907_ (_05870_, _05869_, _05863_);
  or _28908_ (_05871_, _05870_, _05861_);
  not _28909_ (_05872_, _05871_);
  and _28910_ (_05873_, _05872_, _04830_);
  nor _28911_ (_05874_, _05873_, _04879_);
  nor _28912_ (_05875_, _05643_, _05359_);
  and _28913_ (_05876_, _05875_, _05315_);
  and _28914_ (_05877_, _05876_, _05874_);
  and _28915_ (_05878_, _05877_, _05852_);
  and _28916_ (_05879_, _05878_, _05230_);
  and _28917_ (property_invalid_sjmp, _05879_, _05850_);
  and _28918_ (_05880_, _07455_, _07454_);
  nand _28919_ (_05881_, _05880_, _08436_);
  nor _28920_ (_05882_, _05881_, _06968_);
  and _28921_ (_05883_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand _28922_ (_05884_, _07467_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor _28923_ (_05885_, _07475_, _07165_);
  not _28924_ (_05886_, _05885_);
  or _28925_ (_05887_, _05886_, _07472_);
  or _28926_ (_05888_, _05887_, _05884_);
  and _28927_ (_05889_, _05888_, _05883_);
  and _28928_ (_05890_, _05889_, _05881_);
  or _28929_ (_05891_, _05890_, _07459_);
  or _28930_ (_05892_, _05891_, _05882_);
  nand _28931_ (_05893_, _07459_, _07317_);
  and _28932_ (_05894_, _05893_, _06989_);
  and _28933_ (_04835_, _05894_, _05892_);
  not _28934_ (_05895_, _04992_);
  nor _28935_ (_05896_, _05401_, _05313_);
  and _28936_ (_05897_, _05896_, _05272_);
  and _28937_ (_05898_, _05897_, _05359_);
  and _28938_ (_05899_, _04930_, _04878_);
  and _28939_ (_05900_, _05899_, _05898_);
  and _28940_ (_05901_, _05900_, _05873_);
  and _28941_ (_05902_, _05643_, _05359_);
  and _28942_ (_05903_, _05902_, _05315_);
  not _28943_ (_05904_, _04878_);
  or _28944_ (_05905_, _05871_, _05904_);
  and _28945_ (_05906_, _05905_, _04931_);
  and _28946_ (_05907_, _05906_, _05903_);
  or _28947_ (_05908_, _05907_, _05901_);
  and _28948_ (_05909_, _05908_, _05895_);
  and _28949_ (_05910_, _05876_, _05873_);
  not _28950_ (_05911_, _05873_);
  and _28951_ (_05912_, _05898_, _05911_);
  or _28952_ (_05913_, _05912_, _05910_);
  and _28953_ (_05914_, _05852_, _05904_);
  and _28954_ (_05915_, _05914_, _05913_);
  or _28955_ (_05916_, _05915_, _05909_);
  and _28956_ (_05917_, _05160_, _04756_);
  and _28957_ (_05918_, _05917_, _04742_);
  and _28958_ (_05919_, _05918_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _28959_ (_05920_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and _28960_ (_05921_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor _28961_ (_05922_, _05921_, _05920_);
  or _28962_ (_05923_, _05922_, _05919_);
  nand _28963_ (_05924_, _05922_, _05919_);
  and _28964_ (_05925_, _05924_, _05923_);
  and _28965_ (_05926_, _05160_, _04738_);
  and _28966_ (_05927_, _05926_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _28967_ (_05928_, _05926_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _28968_ (_05929_, _05928_, _05927_);
  nor _28969_ (_05930_, _05929_, _01188_);
  nor _28970_ (_05931_, _05918_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _28971_ (_05932_, _05931_, _05919_);
  nor _28972_ (_05933_, _05932_, _01220_);
  or _28973_ (_05934_, _05933_, _05930_);
  or _28974_ (_05935_, _05934_, _05925_);
  and _28975_ (_05936_, _05917_, _04744_);
  and _28976_ (_05937_, _05936_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _28977_ (_05938_, _05936_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _28978_ (_05939_, _05938_, _05937_);
  and _28979_ (_05940_, _05939_, _00687_);
  and _28980_ (_05941_, _05929_, _01188_);
  or _28981_ (_05942_, _05941_, _05940_);
  and _28982_ (_05943_, _05917_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and _28983_ (_05944_, _05943_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _28984_ (_05945_, _05943_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _28985_ (_05946_, _05945_, _05944_);
  and _28986_ (_05947_, _05946_, _01227_);
  and _28987_ (_05948_, _05932_, _01220_);
  or _28988_ (_05949_, _05948_, _05947_);
  or _28989_ (_05950_, _05949_, _05942_);
  nor _28990_ (_05951_, _05162_, _05001_);
  and _28991_ (_05952_, _05162_, _05001_);
  or _28992_ (_05953_, _05952_, _05951_);
  and _28993_ (_05954_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _28994_ (_05955_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor _28995_ (_05956_, _05955_, _05954_);
  nand _28996_ (_05957_, _05956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or _28997_ (_05958_, _05956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and _28998_ (_05959_, _05958_, _05957_);
  nand _28999_ (_05960_, _05959_, _05801_);
  or _29000_ (_05961_, _05159_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand _29001_ (_05962_, _05159_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and _29002_ (_05963_, _05962_, _05961_);
  or _29003_ (_05964_, _05963_, _05960_);
  or _29004_ (_05965_, _05964_, _05953_);
  and _29005_ (_05966_, _05160_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _29006_ (_05967_, _05160_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor _29007_ (_05968_, _05967_, _05966_);
  and _29008_ (_05969_, _05968_, _04608_);
  nor _29009_ (_05970_, _05968_, _04608_);
  or _29010_ (_05971_, _05970_, _05969_);
  or _29011_ (_05972_, _05971_, _05965_);
  nor _29012_ (_05973_, _05917_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _29013_ (_05974_, _05973_, _05943_);
  nor _29014_ (_05975_, _05974_, _01144_);
  and _29015_ (_05976_, _05974_, _01144_);
  or _29016_ (_05977_, _05976_, _05975_);
  or _29017_ (_05978_, _05977_, _05972_);
  nor _29018_ (_05979_, _05946_, _01227_);
  nor _29019_ (_05980_, _05939_, _00687_);
  or _29020_ (_05981_, _05980_, _05979_);
  or _29021_ (_05982_, _05981_, _05978_);
  or _29022_ (_05983_, _05982_, _05950_);
  or _29023_ (_05984_, _05983_, _05935_);
  and _29024_ (_05985_, _05937_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _29025_ (_05986_, _05985_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _29026_ (_05987_, _05985_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _29027_ (_05988_, _05987_, _05986_);
  nand _29028_ (_05989_, _05988_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or _29029_ (_05990_, _05988_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _29030_ (_05991_, _05990_, _05989_);
  nor _29031_ (_05992_, _05937_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _29032_ (_05993_, _05992_, _05985_);
  and _29033_ (_05994_, _05993_, _01686_);
  nor _29034_ (_05995_, _05993_, _01686_);
  nor _29035_ (_05996_, _05966_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _29036_ (_05997_, _05996_, _05926_);
  nor _29037_ (_05998_, _05997_, _01192_);
  and _29038_ (_05999_, _05997_, _01192_);
  or _29039_ (_06000_, _05999_, _05998_);
  nor _29040_ (_06001_, _05927_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _29041_ (_06002_, _06001_, _05917_);
  nor _29042_ (_06003_, _06002_, _01149_);
  and _29043_ (_06004_, _06002_, _01149_);
  or _29044_ (_06005_, _06004_, _06003_);
  or _29045_ (_06006_, _06005_, _06000_);
  or _29046_ (_06007_, _06006_, _05995_);
  or _29047_ (_06008_, _06007_, _05994_);
  or _29048_ (_06009_, _06008_, _05991_);
  and _29049_ (_06010_, _05986_, _00655_);
  nor _29050_ (_06011_, _05986_, _00655_);
  or _29051_ (_06012_, _06011_, _06010_);
  nor _29052_ (_06013_, _06012_, _00619_);
  and _29053_ (_06014_, _06012_, _00619_);
  or _29054_ (_06015_, _06014_, _06013_);
  or _29055_ (_06016_, _06015_, _06009_);
  or _29056_ (_06017_, _06016_, _05984_);
  and _29057_ (_06018_, _06017_, _05230_);
  and _29058_ (property_invalid_pcp3, _06018_, _05916_);
  or _29059_ (_06019_, _05658_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand _29060_ (_06020_, _05658_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and _29061_ (_06021_, _06020_, _06019_);
  or _29062_ (_06022_, _05668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand _29063_ (_06023_, _05668_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and _29064_ (_06024_, _06023_, _06022_);
  and _29065_ (_06025_, _05671_, _01149_);
  nor _29066_ (_06026_, _05671_, _01149_);
  or _29067_ (_06027_, _06026_, _06025_);
  nor _29068_ (_06028_, _05675_, _01188_);
  and _29069_ (_06029_, _05675_, _01188_);
  or _29070_ (_06030_, _06029_, _06028_);
  nor _29071_ (_06031_, _05682_, _01192_);
  and _29072_ (_06032_, _05682_, _01192_);
  or _29073_ (_06033_, _06032_, _06031_);
  and _29074_ (_06034_, _05407_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor _29075_ (_06035_, _05407_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _29076_ (_06036_, _06035_, _06034_);
  and _29077_ (_06037_, _05692_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nand _29078_ (_06038_, _05956_, _05800_);
  nor _29079_ (_06039_, _05692_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or _29080_ (_06040_, _06039_, _06038_);
  or _29081_ (_06041_, _06040_, _06037_);
  or _29082_ (_06042_, _06041_, _06036_);
  nor _29083_ (_06043_, _05688_, _04608_);
  and _29084_ (_06044_, _05688_, _04608_);
  or _29085_ (_06045_, _06044_, _06043_);
  or _29086_ (_06046_, _06045_, _06042_);
  or _29087_ (_06047_, _06046_, _06033_);
  or _29088_ (_06048_, _06047_, _06030_);
  or _29089_ (_06049_, _06048_, _06027_);
  or _29090_ (_06050_, _06049_, _06024_);
  or _29091_ (_06051_, _06050_, _05825_);
  or _29092_ (_06052_, _06051_, _06021_);
  or _29093_ (_06053_, _06052_, _04946_);
  or _29094_ (_06054_, _06053_, _04778_);
  and _29095_ (_06055_, _04931_, _05642_);
  and _29096_ (_06056_, _06055_, _05644_);
  or _29097_ (_06057_, _05900_, _05895_);
  or _29098_ (_06058_, _06057_, _06056_);
  and _29099_ (_06059_, _05871_, _05314_);
  and _29100_ (_06060_, _05873_, _05904_);
  and _29101_ (_06061_, _06060_, _05897_);
  or _29102_ (_06062_, _06061_, _06059_);
  and _29103_ (_06063_, _06062_, _05851_);
  or _29104_ (_06064_, _06063_, _05646_);
  or _29105_ (_06065_, _06064_, _06058_);
  and _29106_ (_06066_, _05643_, _05272_);
  and _29107_ (_06067_, _06066_, _05873_);
  and _29108_ (_06068_, _06067_, _04879_);
  not _29109_ (_06069_, _05358_);
  and _29110_ (_06070_, _05897_, _06069_);
  or _29111_ (_06071_, _06070_, _05645_);
  or _29112_ (_06072_, _06071_, _06068_);
  and _29113_ (_06073_, _06072_, _04931_);
  and _29114_ (_06074_, _05898_, _05642_);
  and _29115_ (_06075_, _05899_, _05314_);
  and _29116_ (_06076_, _06075_, _05872_);
  or _29117_ (_06077_, _06076_, _04992_);
  or _29118_ (_06078_, _06077_, _06074_);
  or _29119_ (_06079_, _06078_, _06073_);
  and _29120_ (_06080_, _06079_, _06065_);
  and _29121_ (_06081_, _06066_, _05911_);
  and _29122_ (_06082_, _05644_, _04878_);
  or _29123_ (_06083_, _06082_, _06081_);
  and _29124_ (_06084_, _06083_, _05852_);
  and _29125_ (_06085_, _05912_, _04931_);
  and _29126_ (_06086_, _05897_, _04879_);
  and _29127_ (_06087_, _06086_, _05641_);
  or _29128_ (_06088_, _06087_, _06085_);
  or _29129_ (_06089_, _06088_, _06084_);
  or _29130_ (_06090_, _06089_, _06080_);
  and _29131_ (_06091_, _06090_, _05230_);
  and _29132_ (property_invalid_pcp2, _06091_, _06054_);
  and _29133_ (_06092_, _03503_, _09009_);
  and _29134_ (_06093_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and _29135_ (_06094_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor _29136_ (_06095_, _06094_, _06093_);
  nor _29137_ (_06096_, _06095_, _13986_);
  and _29138_ (_06097_, _04006_, _11821_);
  or _29139_ (_06098_, _06097_, _06096_);
  or _29140_ (_06099_, _06098_, _06092_);
  and _29141_ (_04843_, _06099_, _06989_);
  and _29142_ (_06100_, _05875_, _05895_);
  or _29143_ (_06101_, _06100_, _06070_);
  and _29144_ (_06102_, _06101_, _05874_);
  and _29145_ (_06103_, _06069_, _05272_);
  nor _29146_ (_06104_, _04992_, _04878_);
  and _29147_ (_06105_, _06104_, _06103_);
  and _29148_ (_06106_, _05314_, _05904_);
  and _29149_ (_06107_, _06106_, _05873_);
  or _29150_ (_06108_, _06107_, _05903_);
  or _29151_ (_06109_, _06108_, _06105_);
  or _29152_ (_06110_, _06109_, _06102_);
  and _29153_ (_06111_, _06110_, _05851_);
  and _29154_ (_06112_, _06067_, _05642_);
  or _29155_ (_06113_, _06103_, _05902_);
  and _29156_ (_06114_, _04991_, _04931_);
  and _29157_ (_06115_, _06114_, _06113_);
  nor _29158_ (_06116_, _06115_, _06112_);
  nor _29159_ (_06117_, _06116_, _05314_);
  and _29160_ (_06118_, _06069_, _04878_);
  and _29161_ (_06119_, _06118_, _04992_);
  or _29162_ (_06120_, _06119_, _06059_);
  or _29163_ (_06121_, _06120_, _06081_);
  and _29164_ (_06122_, _06121_, _04931_);
  or _29165_ (_06123_, _06106_, _04991_);
  or _29166_ (_06124_, _06075_, _04989_);
  and _29167_ (_06125_, _06124_, _06123_);
  or _29168_ (_06126_, _06066_, _05314_);
  and _29169_ (_06127_, _06126_, _05641_);
  and _29170_ (_06128_, _05871_, _04878_);
  and _29171_ (_06129_, _06128_, _05897_);
  and _29172_ (_06130_, _06129_, _05852_);
  or _29173_ (_06131_, _06130_, _06127_);
  or _29174_ (_06132_, _06131_, _06125_);
  or _29175_ (_06133_, _06132_, _06122_);
  or _29176_ (_06134_, _06133_, _06117_);
  or _29177_ (_06135_, _06134_, _06111_);
  not _29178_ (_06136_, _04756_);
  nand _29179_ (_06137_, _04737_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _29180_ (_06138_, _06137_, _06136_);
  and _29181_ (_06139_, _06138_, _04744_);
  and _29182_ (_06140_, _06139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and _29183_ (_06141_, _06140_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and _29184_ (_06142_, _06141_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _29185_ (_06143_, _06142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and _29186_ (_06144_, _06142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor _29187_ (_06145_, _06144_, _06143_);
  and _29188_ (_06146_, _06145_, _00619_);
  nor _29189_ (_06147_, _06141_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor _29190_ (_06148_, _06147_, _06142_);
  nand _29191_ (_06149_, _06148_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  or _29192_ (_06150_, _06148_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  and _29193_ (_06151_, _06150_, _06149_);
  nor _29194_ (_06152_, _06145_, _00619_);
  or _29195_ (_06153_, _06152_, _06151_);
  or _29196_ (_06154_, _06153_, _06146_);
  and _29197_ (_06155_, _04740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _29198_ (_06156_, _06155_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and _29199_ (_06157_, _06155_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor _29200_ (_06158_, _06157_, _06156_);
  and _29201_ (_06159_, _06158_, _01149_);
  nor _29202_ (_06160_, _06158_, _01149_);
  and _29203_ (_06161_, _06138_, _04742_);
  nor _29204_ (_06162_, _06161_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and _29205_ (_06163_, _06161_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor _29206_ (_06164_, _06163_, _06162_);
  nor _29207_ (_06165_, _06164_, _01220_);
  and _29208_ (_06166_, _06164_, _01220_);
  or _29209_ (_06167_, _06166_, _06165_);
  nor _29210_ (_06168_, _06139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor _29211_ (_06169_, _06168_, _06140_);
  nor _29212_ (_06170_, _06169_, _00687_);
  and _29213_ (_06171_, _06169_, _00687_);
  or _29214_ (_06172_, _06171_, _06170_);
  or _29215_ (_06173_, _06172_, _06167_);
  or _29216_ (_06174_, _06173_, _06160_);
  or _29217_ (_06175_, _06174_, _06159_);
  nor _29218_ (_06176_, _06140_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor _29219_ (_06177_, _06176_, _06141_);
  nor _29220_ (_06178_, _06177_, _01686_);
  and _29221_ (_06179_, _04739_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor _29222_ (_06180_, _06179_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor _29223_ (_06181_, _06180_, _06155_);
  and _29224_ (_06182_, _06181_, _01188_);
  nor _29225_ (_06183_, _06181_, _01188_);
  or _29226_ (_06184_, _06183_, _06182_);
  or _29227_ (_06185_, _06184_, _06178_);
  and _29228_ (_06186_, _06138_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _29229_ (_06187_, _06138_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor _29230_ (_06188_, _06187_, _06186_);
  nor _29231_ (_06189_, _06188_, _01144_);
  and _29232_ (_06190_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _04608_);
  nor _29233_ (_06191_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and _29234_ (_06192_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor _29235_ (_06193_, _06192_, _06191_);
  nor _29236_ (_06194_, _06193_, _06137_);
  nor _29237_ (_06195_, _06194_, _06190_);
  and _29238_ (_06196_, _01346_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nor _29239_ (_06197_, _06196_, _06193_);
  or _29240_ (_06198_, _06197_, _06137_);
  or _29241_ (_06199_, _06198_, _06195_);
  nand _29242_ (_06200_, _06197_, _06195_);
  and _29243_ (_06201_, _06200_, _06199_);
  and _29244_ (_06202_, _06188_, _01144_);
  or _29245_ (_06203_, _06202_, _06201_);
  or _29246_ (_06204_, _06203_, _06189_);
  or _29247_ (_06205_, _06163_, _05922_);
  nand _29248_ (_06206_, _06163_, _05922_);
  and _29249_ (_06207_, _06206_, _06205_);
  nor _29250_ (_06208_, _04316_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and _29251_ (_06209_, _04316_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or _29252_ (_06210_, _06209_, _06208_);
  or _29253_ (_06211_, _05959_, _05800_);
  nor _29254_ (_06212_, _04312_, _04503_);
  and _29255_ (_06213_, _04312_, _04503_);
  or _29256_ (_06214_, _06213_, _06212_);
  or _29257_ (_06215_, _06214_, _06211_);
  or _29258_ (_06216_, _06215_, _06210_);
  or _29259_ (_06217_, _06216_, _06207_);
  or _29260_ (_06218_, _06217_, _06204_);
  and _29261_ (_06219_, _06177_, _01686_);
  and _29262_ (_06220_, _06186_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _29263_ (_06221_, _06186_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor _29264_ (_06222_, _06221_, _06220_);
  or _29265_ (_06223_, _06222_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand _29266_ (_06224_, _06222_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and _29267_ (_06225_, _06224_, _06223_);
  or _29268_ (_06226_, _06225_, _06219_);
  or _29269_ (_06227_, _06226_, _06218_);
  or _29270_ (_06228_, _06227_, _06185_);
  or _29271_ (_06229_, _06228_, _06175_);
  or _29272_ (_06230_, _06229_, _06154_);
  and _29273_ (_06231_, _06230_, _05230_);
  and _29274_ (property_invalid_pcp1, _06231_, _06135_);
  and _29275_ (_06232_, _03503_, _09599_);
  and _29276_ (_06233_, _03498_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and _29277_ (_06234_, _00919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor _29278_ (_06235_, _06234_, _06233_);
  nor _29279_ (_06236_, _06235_, _13986_);
  and _29280_ (_06237_, _04006_, _09009_);
  or _29281_ (_06238_, _06237_, _06236_);
  or _29282_ (_06239_, _06238_, _06232_);
  and _29283_ (_04848_, _06239_, _06989_);
  and _29284_ (_06240_, _05223_, first_instr);
  or _29285_ (_00000_, _06240_, rst);
  or _29286_ (_06241_, _13959_, _13969_);
  nor _29287_ (_06242_, _06241_, _00918_);
  and _29288_ (_06243_, _00918_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or _29289_ (_06244_, _06243_, _06242_);
  and _29290_ (_06245_, _13968_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or _29291_ (_06246_, _06245_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and _29292_ (_06247_, _06246_, _13959_);
  nor _29293_ (_06248_, _06247_, _06244_);
  nor _29294_ (_06249_, _06248_, _13986_);
  and _29295_ (_06250_, _04181_, _09599_);
  or _29296_ (_06251_, _06250_, _06249_);
  and _29297_ (_04872_, _06251_, _06989_);
  nor _29298_ (_06252_, _10970_, _04286_);
  nor _29299_ (_06253_, _07145_, _03252_);
  and _29300_ (_06254_, _06253_, _09580_);
  nand _29301_ (_06255_, _07071_, _07056_);
  and _29302_ (_06256_, _06255_, _03245_);
  nor _29303_ (_06257_, _06256_, _09575_);
  or _29304_ (_06258_, _06257_, _07077_);
  or _29305_ (_06259_, _06258_, _06254_);
  and _29306_ (_06260_, _07077_, _03252_);
  nor _29307_ (_06261_, _06260_, _07046_);
  and _29308_ (_06262_, _06261_, _06259_);
  or _29309_ (_06263_, _06262_, _07050_);
  or _29310_ (_06264_, _06263_, _06252_);
  nand _29311_ (_06265_, _07050_, _03245_);
  and _29312_ (_06266_, _06265_, _06989_);
  and _29313_ (_04889_, _06266_, _06264_);
  and _29314_ (_06267_, _07077_, _03256_);
  nor _29315_ (_06268_, _07145_, _03256_);
  and _29316_ (_06269_, _06268_, _09580_);
  not _29317_ (_06270_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand _29318_ (_06271_, _02808_, _06270_);
  and _29319_ (_06272_, _06271_, _06255_);
  or _29320_ (_06273_, _06272_, _07077_);
  nor _29321_ (_06274_, _06273_, _06269_);
  or _29322_ (_06275_, _06274_, _06267_);
  nand _29323_ (_06276_, _06275_, _04286_);
  nand _29324_ (_06277_, _07118_, _07046_);
  and _29325_ (_06278_, _06277_, _06276_);
  or _29326_ (_06279_, _06278_, _07050_);
  nand _29327_ (_06280_, _07050_, _06270_);
  and _29328_ (_06281_, _06280_, _06989_);
  and _29329_ (_04896_, _06281_, _06279_);
  and _29330_ (_06282_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and _29331_ (_06283_, _06282_, _09580_);
  and _29332_ (_06284_, _07071_, _07062_);
  nor _29333_ (_06285_, _06284_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor _29334_ (_06286_, _06285_, _04293_);
  or _29335_ (_06287_, _06286_, _07077_);
  or _29336_ (_06288_, _06287_, _06283_);
  nor _29337_ (_06289_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor _29338_ (_06290_, _06289_, _07046_);
  and _29339_ (_06291_, _06290_, _06288_);
  and _29340_ (_06292_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or _29341_ (_06293_, _06292_, _07050_);
  or _29342_ (_06294_, _06293_, _06291_);
  nand _29343_ (_06295_, _07260_, _07050_);
  and _29344_ (_06296_, _06295_, _06989_);
  and _29345_ (_04909_, _06296_, _06294_);
  and _29346_ (_06297_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and _29347_ (_06298_, _06297_, _09580_);
  nand _29348_ (_06299_, _07071_, _07061_);
  and _29349_ (_06300_, _06299_, _03049_);
  nor _29350_ (_06301_, _06300_, _06284_);
  or _29351_ (_06302_, _06301_, _07077_);
  or _29352_ (_06303_, _06302_, _06298_);
  nor _29353_ (_06304_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor _29354_ (_06305_, _06304_, _07046_);
  and _29355_ (_06306_, _06305_, _06303_);
  and _29356_ (_06307_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or _29357_ (_06308_, _06307_, _07050_);
  or _29358_ (_06309_, _06308_, _06306_);
  nand _29359_ (_06310_, _07317_, _07050_);
  and _29360_ (_06311_, _06310_, _06989_);
  and _29361_ (_04916_, _06311_, _06309_);
  and _29362_ (_06312_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and _29363_ (_06313_, _06312_, _09580_);
  and _29364_ (_06314_, _07071_, _07060_);
  or _29365_ (_06315_, _06314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and _29366_ (_06316_, _06315_, _06299_);
  or _29367_ (_06317_, _06316_, _07077_);
  or _29368_ (_06318_, _06317_, _06313_);
  nor _29369_ (_06319_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor _29370_ (_06320_, _06319_, _07046_);
  and _29371_ (_06321_, _06320_, _06318_);
  and _29372_ (_06322_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or _29373_ (_06323_, _06322_, _07050_);
  or _29374_ (_06324_, _06323_, _06321_);
  nand _29375_ (_06325_, _11529_, _07050_);
  and _29376_ (_06326_, _06325_, _06989_);
  and _29377_ (_04920_, _06326_, _06324_);
  nor _29378_ (_06327_, _10970_, _14146_);
  and _29379_ (_06328_, _08999_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and _29380_ (_06329_, _06981_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  and _29381_ (_06330_, _06329_, _09002_);
  or _29382_ (_06331_, _06330_, _06328_);
  or _29383_ (_06332_, _06331_, _06327_);
  and _29384_ (_04922_, _06332_, _06989_);
  and _29385_ (_06333_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and _29386_ (_06334_, _06333_, _09580_);
  and _29387_ (_06335_, _07071_, _07059_);
  nor _29388_ (_06336_, _06335_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor _29389_ (_06337_, _06336_, _06314_);
  or _29390_ (_06338_, _06337_, _07077_);
  or _29391_ (_06339_, _06338_, _06334_);
  nor _29392_ (_06340_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor _29393_ (_06341_, _06340_, _07046_);
  and _29394_ (_06342_, _06341_, _06339_);
  and _29395_ (_06343_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or _29396_ (_06344_, _06343_, _07050_);
  or _29397_ (_06345_, _06344_, _06342_);
  nand _29398_ (_06346_, _09008_, _07050_);
  and _29399_ (_06347_, _06346_, _06989_);
  and _29400_ (_04924_, _06347_, _06345_);
  and _29401_ (_06348_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor _29402_ (_06349_, _08139_, _04608_);
  or _29403_ (_06350_, _06349_, _06348_);
  and _29404_ (_04941_, _06350_, _06989_);
  and _29405_ (_06351_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor _29406_ (_06352_, _08139_, _05001_);
  or _29407_ (_06353_, _06352_, _06351_);
  and _29408_ (_04943_, _06353_, _06989_);
  and _29409_ (_06354_, _07146_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and _29410_ (_06355_, _06354_, _09580_);
  and _29411_ (_06356_, _09577_, _03143_);
  nor _29412_ (_06357_, _06356_, _06335_);
  or _29413_ (_06358_, _06357_, _07077_);
  or _29414_ (_06359_, _06358_, _06355_);
  nor _29415_ (_06360_, _09574_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor _29416_ (_06361_, _06360_, _07046_);
  and _29417_ (_06362_, _06361_, _06359_);
  and _29418_ (_06363_, _07046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or _29419_ (_06364_, _06363_, _07050_);
  or _29420_ (_06365_, _06364_, _06362_);
  nand _29421_ (_06366_, _09598_, _07050_);
  and _29422_ (_06367_, _06366_, _06989_);
  and _29423_ (_04945_, _06367_, _06365_);
  nand _29424_ (_06368_, _05880_, _07089_);
  nor _29425_ (_06369_, _06368_, _06968_);
  or _29426_ (_06370_, _05885_, _07472_);
  or _29427_ (_06371_, _06370_, _05884_);
  nand _29428_ (_06372_, _06371_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand _29429_ (_06373_, _06372_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and _29430_ (_06374_, _06373_, _06368_);
  or _29431_ (_06375_, _06374_, _07459_);
  or _29432_ (_06376_, _06375_, _06369_);
  nand _29433_ (_06377_, _09008_, _07459_);
  and _29434_ (_06378_, _06377_, _06989_);
  and _29435_ (_04978_, _06378_, _06376_);
  and _29436_ (_06379_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor _29437_ (_06380_, _08139_, _04503_);
  or _29438_ (_06381_, _06380_, _06379_);
  and _29439_ (_04990_, _06381_, _06989_);
  nor _29440_ (_06382_, _01811_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  or _29441_ (_06383_, _05887_, _07468_);
  and _29442_ (_06384_, _06383_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or _29443_ (_06385_, _06384_, _06382_);
  and _29444_ (_06386_, _05880_, _07048_);
  or _29445_ (_06387_, _06386_, _06385_);
  nand _29446_ (_06388_, _06386_, _06968_);
  and _29447_ (_06389_, _06388_, _06387_);
  or _29448_ (_06390_, _06389_, _07459_);
  nand _29449_ (_06391_, _07459_, _07118_);
  and _29450_ (_06392_, _06391_, _06989_);
  and _29451_ (_05002_, _06392_, _06390_);
  and _29452_ (_06393_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor _29453_ (_06394_, _08139_, _05013_);
  or _29454_ (_06395_, _06394_, _06393_);
  and _29455_ (_05018_, _06395_, _06989_);
  and _29456_ (_06396_, _08139_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor _29457_ (_06397_, _08139_, _04416_);
  or _29458_ (_06398_, _06397_, _06396_);
  and _29459_ (_05033_, _06398_, _06989_);
  dff _29460_ (first_instr, _00000_, clk);
  dff _29461_ (\oc8051_symbolic_cxrom1.regarray[10] [0], _14649_, clk);
  dff _29462_ (\oc8051_symbolic_cxrom1.regarray[10] [1], _14650_, clk);
  dff _29463_ (\oc8051_symbolic_cxrom1.regarray[10] [2], _14651_, clk);
  dff _29464_ (\oc8051_symbolic_cxrom1.regarray[10] [3], _14652_, clk);
  dff _29465_ (\oc8051_symbolic_cxrom1.regarray[10] [4], _14653_, clk);
  dff _29466_ (\oc8051_symbolic_cxrom1.regarray[10] [5], _14654_, clk);
  dff _29467_ (\oc8051_symbolic_cxrom1.regarray[10] [6], _09711_, clk);
  dff _29468_ (\oc8051_symbolic_cxrom1.regarray[10] [7], _14655_, clk);
  dff _29469_ (\oc8051_symbolic_cxrom1.regarray[9] [0], _14707_, clk);
  dff _29470_ (\oc8051_symbolic_cxrom1.regarray[9] [1], _09612_, clk);
  dff _29471_ (\oc8051_symbolic_cxrom1.regarray[9] [2], _09617_, clk);
  dff _29472_ (\oc8051_symbolic_cxrom1.regarray[9] [3], _09622_, clk);
  dff _29473_ (\oc8051_symbolic_cxrom1.regarray[9] [4], _14708_, clk);
  dff _29474_ (\oc8051_symbolic_cxrom1.regarray[9] [5], _14709_, clk);
  dff _29475_ (\oc8051_symbolic_cxrom1.regarray[9] [6], _14710_, clk);
  dff _29476_ (\oc8051_symbolic_cxrom1.regarray[9] [7], _09635_, clk);
  dff _29477_ (\oc8051_symbolic_cxrom1.regarray[8] [0], _09522_, clk);
  dff _29478_ (\oc8051_symbolic_cxrom1.regarray[8] [1], _14702_, clk);
  dff _29479_ (\oc8051_symbolic_cxrom1.regarray[8] [2], _09526_, clk);
  dff _29480_ (\oc8051_symbolic_cxrom1.regarray[8] [3], _14703_, clk);
  dff _29481_ (\oc8051_symbolic_cxrom1.regarray[8] [4], _14704_, clk);
  dff _29482_ (\oc8051_symbolic_cxrom1.regarray[8] [5], _14705_, clk);
  dff _29483_ (\oc8051_symbolic_cxrom1.regarray[8] [6], _09540_, clk);
  dff _29484_ (\oc8051_symbolic_cxrom1.regarray[8] [7], _14706_, clk);
  dff _29485_ (\oc8051_symbolic_cxrom1.regarray[7] [0], _14694_, clk);
  dff _29486_ (\oc8051_symbolic_cxrom1.regarray[7] [1], _14695_, clk);
  dff _29487_ (\oc8051_symbolic_cxrom1.regarray[7] [2], _14696_, clk);
  dff _29488_ (\oc8051_symbolic_cxrom1.regarray[7] [3], _14697_, clk);
  dff _29489_ (\oc8051_symbolic_cxrom1.regarray[7] [4], _14698_, clk);
  dff _29490_ (\oc8051_symbolic_cxrom1.regarray[7] [5], _14699_, clk);
  dff _29491_ (\oc8051_symbolic_cxrom1.regarray[7] [6], _14700_, clk);
  dff _29492_ (\oc8051_symbolic_cxrom1.regarray[7] [7], _14701_, clk);
  dff _29493_ (\oc8051_symbolic_cxrom1.regarray[6] [0], _09328_, clk);
  dff _29494_ (\oc8051_symbolic_cxrom1.regarray[6] [1], _14691_, clk);
  dff _29495_ (\oc8051_symbolic_cxrom1.regarray[6] [2], _09335_, clk);
  dff _29496_ (\oc8051_symbolic_cxrom1.regarray[6] [3], _14692_, clk);
  dff _29497_ (\oc8051_symbolic_cxrom1.regarray[6] [4], _14693_, clk);
  dff _29498_ (\oc8051_symbolic_cxrom1.regarray[6] [5], _09346_, clk);
  dff _29499_ (\oc8051_symbolic_cxrom1.regarray[6] [6], _09351_, clk);
  dff _29500_ (\oc8051_symbolic_cxrom1.regarray[6] [7], _09354_, clk);
  dff _29501_ (\oc8051_symbolic_cxrom1.regarray[5] [0], _09235_, clk);
  dff _29502_ (\oc8051_symbolic_cxrom1.regarray[5] [1], _09238_, clk);
  dff _29503_ (\oc8051_symbolic_cxrom1.regarray[5] [2], _14690_, clk);
  dff _29504_ (\oc8051_symbolic_cxrom1.regarray[5] [3], _09243_, clk);
  dff _29505_ (\oc8051_symbolic_cxrom1.regarray[5] [4], _09247_, clk);
  dff _29506_ (\oc8051_symbolic_cxrom1.regarray[5] [5], _09251_, clk);
  dff _29507_ (\oc8051_symbolic_cxrom1.regarray[5] [6], _09254_, clk);
  dff _29508_ (\oc8051_symbolic_cxrom1.regarray[5] [7], _09257_, clk);
  dff _29509_ (\oc8051_symbolic_cxrom1.regarray[1] [0], _08840_, clk);
  dff _29510_ (\oc8051_symbolic_cxrom1.regarray[1] [1], _14666_, clk);
  dff _29511_ (\oc8051_symbolic_cxrom1.regarray[1] [2], _14667_, clk);
  dff _29512_ (\oc8051_symbolic_cxrom1.regarray[1] [3], _14668_, clk);
  dff _29513_ (\oc8051_symbolic_cxrom1.regarray[1] [4], _14669_, clk);
  dff _29514_ (\oc8051_symbolic_cxrom1.regarray[1] [5], _14670_, clk);
  dff _29515_ (\oc8051_symbolic_cxrom1.regarray[1] [6], _14671_, clk);
  dff _29516_ (\oc8051_symbolic_cxrom1.regarray[1] [7], _14672_, clk);
  dff _29517_ (\oc8051_symbolic_cxrom1.regarray[0] [0], _14642_, clk);
  dff _29518_ (\oc8051_symbolic_cxrom1.regarray[0] [1], _14643_, clk);
  dff _29519_ (\oc8051_symbolic_cxrom1.regarray[0] [2], _14644_, clk);
  dff _29520_ (\oc8051_symbolic_cxrom1.regarray[0] [3], _14645_, clk);
  dff _29521_ (\oc8051_symbolic_cxrom1.regarray[0] [4], _08749_, clk);
  dff _29522_ (\oc8051_symbolic_cxrom1.regarray[0] [5], _14646_, clk);
  dff _29523_ (\oc8051_symbolic_cxrom1.regarray[0] [6], _14647_, clk);
  dff _29524_ (\oc8051_symbolic_cxrom1.regarray[0] [7], _14648_, clk);
  dff _29525_ (\oc8051_symbolic_cxrom1.regarray[3] [0], _14680_, clk);
  dff _29526_ (\oc8051_symbolic_cxrom1.regarray[3] [1], _14681_, clk);
  dff _29527_ (\oc8051_symbolic_cxrom1.regarray[3] [2], _14682_, clk);
  dff _29528_ (\oc8051_symbolic_cxrom1.regarray[3] [3], _14683_, clk);
  dff _29529_ (\oc8051_symbolic_cxrom1.regarray[3] [4], _14684_, clk);
  dff _29530_ (\oc8051_symbolic_cxrom1.regarray[3] [5], _14685_, clk);
  dff _29531_ (\oc8051_symbolic_cxrom1.regarray[3] [6], _14686_, clk);
  dff _29532_ (\oc8051_symbolic_cxrom1.regarray[3] [7], _09047_, clk);
  dff _29533_ (\oc8051_symbolic_cxrom1.regarray[2] [0], _14673_, clk);
  dff _29534_ (\oc8051_symbolic_cxrom1.regarray[2] [1], _14674_, clk);
  dff _29535_ (\oc8051_symbolic_cxrom1.regarray[2] [2], _14675_, clk);
  dff _29536_ (\oc8051_symbolic_cxrom1.regarray[2] [3], _14676_, clk);
  dff _29537_ (\oc8051_symbolic_cxrom1.regarray[2] [4], _14677_, clk);
  dff _29538_ (\oc8051_symbolic_cxrom1.regarray[2] [5], _08962_, clk);
  dff _29539_ (\oc8051_symbolic_cxrom1.regarray[2] [6], _14678_, clk);
  dff _29540_ (\oc8051_symbolic_cxrom1.regarray[2] [7], _14679_, clk);
  dff _29541_ (\oc8051_symbolic_cxrom1.regarray[4] [0], _09135_, clk);
  dff _29542_ (\oc8051_symbolic_cxrom1.regarray[4] [1], _09137_, clk);
  dff _29543_ (\oc8051_symbolic_cxrom1.regarray[4] [2], _09141_, clk);
  dff _29544_ (\oc8051_symbolic_cxrom1.regarray[4] [3], _14687_, clk);
  dff _29545_ (\oc8051_symbolic_cxrom1.regarray[4] [4], _14688_, clk);
  dff _29546_ (\oc8051_symbolic_cxrom1.regarray[4] [5], _14689_, clk);
  dff _29547_ (\oc8051_symbolic_cxrom1.regarray[4] [6], _09152_, clk);
  dff _29548_ (\oc8051_symbolic_cxrom1.regarray[4] [7], _09154_, clk);
  dff _29549_ (\oc8051_symbolic_cxrom1.regvalid [0], _07214_, clk);
  dff _29550_ (\oc8051_symbolic_cxrom1.regvalid [1], _07241_, clk);
  dff _29551_ (\oc8051_symbolic_cxrom1.regvalid [2], _07280_, clk);
  dff _29552_ (\oc8051_symbolic_cxrom1.regvalid [3], _07329_, clk);
  dff _29553_ (\oc8051_symbolic_cxrom1.regvalid [4], _07388_, clk);
  dff _29554_ (\oc8051_symbolic_cxrom1.regvalid [5], _07451_, clk);
  dff _29555_ (\oc8051_symbolic_cxrom1.regvalid [6], _07503_, clk);
  dff _29556_ (\oc8051_symbolic_cxrom1.regvalid [7], _07599_, clk);
  dff _29557_ (\oc8051_symbolic_cxrom1.regvalid [8], _07673_, clk);
  dff _29558_ (\oc8051_symbolic_cxrom1.regvalid [9], _07773_, clk);
  dff _29559_ (\oc8051_symbolic_cxrom1.regvalid [10], _07869_, clk);
  dff _29560_ (\oc8051_symbolic_cxrom1.regvalid [11], _07980_, clk);
  dff _29561_ (\oc8051_symbolic_cxrom1.regvalid [12], _08081_, clk);
  dff _29562_ (\oc8051_symbolic_cxrom1.regvalid [13], _08217_, clk);
  dff _29563_ (\oc8051_symbolic_cxrom1.regvalid [14], _08347_, clk);
  dff _29564_ (\oc8051_symbolic_cxrom1.regvalid [15], _07163_, clk);
  dff _29565_ (\oc8051_symbolic_cxrom1.regarray[15] [0], _10126_, clk);
  dff _29566_ (\oc8051_symbolic_cxrom1.regarray[15] [1], _10131_, clk);
  dff _29567_ (\oc8051_symbolic_cxrom1.regarray[15] [2], _10133_, clk);
  dff _29568_ (\oc8051_symbolic_cxrom1.regarray[15] [3], _10135_, clk);
  dff _29569_ (\oc8051_symbolic_cxrom1.regarray[15] [4], _10137_, clk);
  dff _29570_ (\oc8051_symbolic_cxrom1.regarray[15] [5], _10139_, clk);
  dff _29571_ (\oc8051_symbolic_cxrom1.regarray[15] [6], _10144_, clk);
  dff _29572_ (\oc8051_symbolic_cxrom1.regarray[15] [7], _07192_, clk);
  dff _29573_ (\oc8051_symbolic_cxrom1.regarray[13] [0], _14665_, clk);
  dff _29574_ (\oc8051_symbolic_cxrom1.regarray[13] [1], _09956_, clk);
  dff _29575_ (\oc8051_symbolic_cxrom1.regarray[13] [2], _09961_, clk);
  dff _29576_ (\oc8051_symbolic_cxrom1.regarray[13] [3], _09963_, clk);
  dff _29577_ (\oc8051_symbolic_cxrom1.regarray[13] [4], _09967_, clk);
  dff _29578_ (\oc8051_symbolic_cxrom1.regarray[13] [5], _09971_, clk);
  dff _29579_ (\oc8051_symbolic_cxrom1.regarray[13] [6], _09973_, clk);
  dff _29580_ (\oc8051_symbolic_cxrom1.regarray[13] [7], _09978_, clk);
  dff _29581_ (\oc8051_symbolic_cxrom1.regarray[14] [0], _10042_, clk);
  dff _29582_ (\oc8051_symbolic_cxrom1.regarray[14] [1], _10047_, clk);
  dff _29583_ (\oc8051_symbolic_cxrom1.regarray[14] [2], _10049_, clk);
  dff _29584_ (\oc8051_symbolic_cxrom1.regarray[14] [3], _10051_, clk);
  dff _29585_ (\oc8051_symbolic_cxrom1.regarray[14] [4], _10053_, clk);
  dff _29586_ (\oc8051_symbolic_cxrom1.regarray[14] [5], _10055_, clk);
  dff _29587_ (\oc8051_symbolic_cxrom1.regarray[14] [6], _10058_, clk);
  dff _29588_ (\oc8051_symbolic_cxrom1.regarray[14] [7], _10062_, clk);
  dff _29589_ (\oc8051_symbolic_cxrom1.regarray[12] [0], _09864_, clk);
  dff _29590_ (\oc8051_symbolic_cxrom1.regarray[12] [1], _09867_, clk);
  dff _29591_ (\oc8051_symbolic_cxrom1.regarray[12] [2], _09869_, clk);
  dff _29592_ (\oc8051_symbolic_cxrom1.regarray[12] [3], _09874_, clk);
  dff _29593_ (\oc8051_symbolic_cxrom1.regarray[12] [4], _09877_, clk);
  dff _29594_ (\oc8051_symbolic_cxrom1.regarray[12] [5], _09880_, clk);
  dff _29595_ (\oc8051_symbolic_cxrom1.regarray[12] [6], _14664_, clk);
  dff _29596_ (\oc8051_symbolic_cxrom1.regarray[12] [7], _09885_, clk);
  dff _29597_ (\oc8051_symbolic_cxrom1.regarray[11] [0], _14656_, clk);
  dff _29598_ (\oc8051_symbolic_cxrom1.regarray[11] [1], _14657_, clk);
  dff _29599_ (\oc8051_symbolic_cxrom1.regarray[11] [2], _14658_, clk);
  dff _29600_ (\oc8051_symbolic_cxrom1.regarray[11] [3], _14659_, clk);
  dff _29601_ (\oc8051_symbolic_cxrom1.regarray[11] [4], _14660_, clk);
  dff _29602_ (\oc8051_symbolic_cxrom1.regarray[11] [5], _14661_, clk);
  dff _29603_ (\oc8051_symbolic_cxrom1.regarray[11] [6], _14662_, clk);
  dff _29604_ (\oc8051_symbolic_cxrom1.regarray[11] [7], _14663_, clk);
  dff _29605_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _13463_, clk);
  dff _29606_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _13118_, clk);
  dff _29607_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _13114_, clk);
  dff _29608_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _12965_, clk);
  dff _29609_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _04086_, clk);
  dff _29610_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _04206_, clk);
  dff _29611_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _04099_, clk);
  dff _29612_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _04196_, clk);
  dff _29613_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03313_, clk);
  dff _29614_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _11967_, clk);
  dff _29615_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _12000_, clk);
  dff _29616_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _11997_, clk);
  dff _29617_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _04104_, clk);
  dff _29618_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _12133_, clk);
  dff _29619_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _12387_, clk);
  dff _29620_ (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _04199_, clk);
  dff _29621_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11307_, clk);
  dff _29622_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _12373_, clk);
  dff _29623_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _11323_, clk);
  dff _29624_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _11318_, clk);
  dff _29625_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _11487_, clk);
  dff _29626_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _11384_, clk);
  dff _29627_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _11362_, clk);
  dff _29628_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11357_, clk);
  dff _29629_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _11434_, clk);
  dff _29630_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _08135_, clk);
  dff _29631_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _11200_, clk);
  dff _29632_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _11228_, clk);
  dff _29633_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _11222_, clk);
  dff _29634_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _11633_, clk);
  dff _29635_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _11268_, clk);
  dff _29636_ (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _11259_, clk);
  dff _29637_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _06825_, clk);
  dff _29638_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _06827_, clk);
  dff _29639_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _06829_, clk);
  dff _29640_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _06831_, clk);
  dff _29641_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _06833_, clk);
  dff _29642_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _06836_, clk);
  dff _29643_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _06838_, clk);
  dff _29644_ (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _06671_, clk);
  dff _29645_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _04487_, clk);
  dff _29646_ (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _06674_, clk);
  dff _29647_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _09999_, clk);
  dff _29648_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _03758_, clk);
  dff _29649_ (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _00258_, clk);
  dff _29650_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _03795_, clk);
  dff _29651_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _03766_, clk);
  dff _29652_ (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _03634_, clk);
  dff _29653_ (\oc8051_top_1.oc8051_decoder1.mem_act [0], _03693_, clk);
  dff _29654_ (\oc8051_top_1.oc8051_decoder1.mem_act [1], _03715_, clk);
  dff _29655_ (\oc8051_top_1.oc8051_decoder1.mem_act [2], _03636_, clk);
  dff _29656_ (\oc8051_top_1.oc8051_decoder1.state [0], _03721_, clk);
  dff _29657_ (\oc8051_top_1.oc8051_decoder1.state [1], _03638_, clk);
  dff _29658_ (\oc8051_top_1.oc8051_decoder1.op [0], _03829_, clk);
  dff _29659_ (\oc8051_top_1.oc8051_decoder1.op [1], _03833_, clk);
  dff _29660_ (\oc8051_top_1.oc8051_decoder1.op [2], _03835_, clk);
  dff _29661_ (\oc8051_top_1.oc8051_decoder1.op [3], _03837_, clk);
  dff _29662_ (\oc8051_top_1.oc8051_decoder1.op [4], _03839_, clk);
  dff _29663_ (\oc8051_top_1.oc8051_decoder1.op [5], _03841_, clk);
  dff _29664_ (\oc8051_top_1.oc8051_decoder1.op [6], _03854_, clk);
  dff _29665_ (\oc8051_top_1.oc8051_decoder1.op [7], _03641_, clk);
  dff _29666_ (\oc8051_top_1.oc8051_decoder1.src_sel3 , _03643_, clk);
  dff _29667_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _03518_, clk);
  dff _29668_ (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _03645_, clk);
  dff _29669_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _03541_, clk);
  dff _29670_ (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _03648_, clk);
  dff _29671_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _03557_, clk);
  dff _29672_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _03566_, clk);
  dff _29673_ (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _03655_, clk);
  dff _29674_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _03579_, clk);
  dff _29675_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _03598_, clk);
  dff _29676_ (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _03657_, clk);
  dff _29677_ (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _03719_, clk);
  dff _29678_ (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _03659_, clk);
  dff _29679_ (\oc8051_top_1.oc8051_decoder1.alu_op [0], _03815_, clk);
  dff _29680_ (\oc8051_top_1.oc8051_decoder1.alu_op [1], _03869_, clk);
  dff _29681_ (\oc8051_top_1.oc8051_decoder1.alu_op [2], _03879_, clk);
  dff _29682_ (\oc8051_top_1.oc8051_decoder1.alu_op [3], _03662_, clk);
  dff _29683_ (\oc8051_top_1.oc8051_decoder1.psw_set [0], _03995_, clk);
  dff _29684_ (\oc8051_top_1.oc8051_decoder1.psw_set [1], _03664_, clk);
  dff _29685_ (\oc8051_top_1.oc8051_decoder1.wr , _03666_, clk);
  dff _29686_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _03764_, clk);
  dff _29687_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _14572_, clk);
  dff _29688_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _11893_, clk);
  dff _29689_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _09305_, clk);
  dff _29690_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _13146_, clk);
  dff _29691_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _09122_, clk);
  dff _29692_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _04117_, clk);
  dff _29693_ (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _14014_, clk);
  dff _29694_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _01250_, clk);
  dff _29695_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _04211_, clk);
  dff _29696_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _13157_, clk);
  dff _29697_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _04214_, clk);
  dff _29698_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _02297_, clk);
  dff _29699_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _04524_, clk);
  dff _29700_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _04216_, clk);
  dff _29701_ (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _04034_, clk);
  dff _29702_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _03072_, clk);
  dff _29703_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _00442_, clk);
  dff _29704_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _10877_, clk);
  dff _29705_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _00494_, clk);
  dff _29706_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _03327_, clk);
  dff _29707_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _12693_, clk);
  dff _29708_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _12672_, clk);
  dff _29709_ (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _02737_, clk);
  dff _29710_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _03345_, clk);
  dff _29711_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _03364_, clk);
  dff _29712_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _13272_, clk);
  dff _29713_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _01662_, clk);
  dff _29714_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _00529_, clk);
  dff _29715_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _03439_, clk);
  dff _29716_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _01770_, clk);
  dff _29717_ (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _03992_, clk);
  dff _29718_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _08521_, clk);
  dff _29719_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _08660_, clk);
  dff _29720_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _04112_, clk);
  dff _29721_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _01526_, clk);
  dff _29722_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _12548_, clk);
  dff _29723_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _12655_, clk);
  dff _29724_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _03447_, clk);
  dff _29725_ (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _01800_, clk);
  dff _29726_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _11031_, clk);
  dff _29727_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _07336_, clk);
  dff _29728_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _03957_, clk);
  dff _29729_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _12976_, clk);
  dff _29730_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _03354_, clk);
  dff _29731_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _04003_, clk);
  dff _29732_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _04922_, clk);
  dff _29733_ (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _04207_, clk);
  dff _29734_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _02650_, clk);
  dff _29735_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _13446_, clk);
  dff _29736_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _01208_, clk);
  dff _29737_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _09596_, clk);
  dff _29738_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _13225_, clk);
  dff _29739_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _12039_, clk);
  dff _29740_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _09662_, clk);
  dff _29741_ (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _12810_, clk);
  dff _29742_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _01240_, clk);
  dff _29743_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _12941_, clk);
  dff _29744_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _11005_, clk);
  dff _29745_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _13597_, clk);
  dff _29746_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _08073_, clk);
  dff _29747_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _06571_, clk);
  dff _29748_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _02294_, clk);
  dff _29749_ (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _13343_, clk);
  dff _29750_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _08194_, clk);
  dff _29751_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _08111_, clk);
  dff _29752_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _07933_, clk);
  dff _29753_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _08088_, clk);
  dff _29754_ (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _03549_, clk);
  dff _29755_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _05033_, clk);
  dff _29756_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _05018_, clk);
  dff _29757_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _04990_, clk);
  dff _29758_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _04943_, clk);
  dff _29759_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _04941_, clk);
  dff _29760_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _00638_, clk);
  dff _29761_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _04566_, clk);
  dff _29762_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _02965_, clk);
  dff _29763_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _02962_, clk);
  dff _29764_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _02922_, clk);
  dff _29765_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _00667_, clk);
  dff _29766_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _02100_, clk);
  dff _29767_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _01835_, clk);
  dff _29768_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _02058_, clk);
  dff _29769_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _02001_, clk);
  dff _29770_ (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _14123_, clk);
  dff _29771_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _11677_, clk);
  dff _29772_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _10989_, clk);
  dff _29773_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _00681_, clk);
  dff _29774_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _01629_, clk);
  dff _29775_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _01627_, clk);
  dff _29776_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _00588_, clk);
  dff _29777_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _00575_, clk);
  dff _29778_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _00457_, clk);
  dff _29779_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _00445_, clk);
  dff _29780_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _00679_, clk);
  dff _29781_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _00663_, clk);
  dff _29782_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _06580_, clk);
  dff _29783_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _14585_, clk);
  dff _29784_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _14583_, clk);
  dff _29785_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _14403_, clk);
  dff _29786_ (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _14264_, clk);
  dff _29787_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _04306_, clk);
  dff _29788_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _04532_, clk);
  dff _29789_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _04360_, clk);
  dff _29790_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _10020_, clk);
  dff _29791_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _09691_, clk);
  dff _29792_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _09812_, clk);
  dff _29793_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _03712_, clk);
  dff _29794_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _03706_, clk);
  dff _29795_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _10029_, clk);
  dff _29796_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _04068_, clk);
  dff _29797_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _04061_, clk);
  dff _29798_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _04059_, clk);
  dff _29799_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _10025_, clk);
  dff _29800_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _03150_, clk);
  dff _29801_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _00705_, clk);
  dff _29802_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _02578_, clk);
  dff _29803_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _01817_, clk);
  dff _29804_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _01721_, clk);
  dff _29805_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _10036_, clk);
  dff _29806_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _03489_, clk);
  dff _29807_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _03521_, clk);
  dff _29808_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _03512_, clk);
  dff _29809_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _10033_, clk);
  dff _29810_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _09687_, clk);
  dff _29811_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _14024_, clk);
  dff _29812_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _13822_, clk);
  dff _29813_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _13954_, clk);
  dff _29814_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _13872_, clk);
  dff _29815_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _10045_, clk);
  dff _29816_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _00387_, clk);
  dff _29817_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _00055_, clk);
  dff _29818_ (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _14019_, clk);
  dff _29819_ (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _14216_, clk);
  dff _29820_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _10056_, clk);
  dff _29821_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _09677_, clk);
  dff _29822_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _09795_, clk);
  dff _29823_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _14142_, clk);
  dff _29824_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _14393_, clk);
  dff _29825_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _01178_, clk);
  dff _29826_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _09919_, clk);
  dff _29827_ (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _03539_, clk);
  dff _29828_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _09922_, clk);
  dff _29829_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _09747_, clk);
  dff _29830_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _00596_, clk);
  dff _29831_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _09929_, clk);
  dff _29832_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _10114_, clk);
  dff _29833_ (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _09651_, clk);
  dff _29834_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _09936_, clk);
  dff _29835_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _09733_, clk);
  dff _29836_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _04007_, clk);
  dff _29837_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _03810_, clk);
  dff _29838_ (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _03808_, clk);
  dff _29839_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _00250_, clk);
  dff _29840_ (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _03755_, clk);
  dff _29841_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _10079_, clk);
  dff _29842_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _04585_, clk);
  dff _29843_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _04582_, clk);
  dff _29844_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _04572_, clk);
  dff _29845_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _04568_, clk);
  dff _29846_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _10074_, clk);
  dff _29847_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _09791_, clk);
  dff _29848_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _04137_, clk);
  dff _29849_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _04134_, clk);
  dff _29850_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _04130_, clk);
  dff _29851_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _04122_, clk);
  dff _29852_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _04114_, clk);
  dff _29853_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _10092_, clk);
  dff _29854_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _04236_, clk);
  dff _29855_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _04233_, clk);
  dff _29856_ (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _03742_, clk);
  dff _29857_ (\oc8051_top_1.oc8051_memory_interface1.pc [0], _03399_, clk);
  dff _29858_ (\oc8051_top_1.oc8051_memory_interface1.pc [1], _03374_, clk);
  dff _29859_ (\oc8051_top_1.oc8051_memory_interface1.pc [2], _03372_, clk);
  dff _29860_ (\oc8051_top_1.oc8051_memory_interface1.pc [3], _10101_, clk);
  dff _29861_ (\oc8051_top_1.oc8051_memory_interface1.pc [4], _03831_, clk);
  dff _29862_ (\oc8051_top_1.oc8051_memory_interface1.pc [5], _03723_, clk);
  dff _29863_ (\oc8051_top_1.oc8051_memory_interface1.pc [6], _03682_, clk);
  dff _29864_ (\oc8051_top_1.oc8051_memory_interface1.pc [7], _03651_, clk);
  dff _29865_ (\oc8051_top_1.oc8051_memory_interface1.pc [8], _10098_, clk);
  dff _29866_ (\oc8051_top_1.oc8051_memory_interface1.pc [9], _09669_, clk);
  dff _29867_ (\oc8051_top_1.oc8051_memory_interface1.pc [10], _02056_, clk);
  dff _29868_ (\oc8051_top_1.oc8051_memory_interface1.pc [11], _01860_, clk);
  dff _29869_ (\oc8051_top_1.oc8051_memory_interface1.pc [12], _02024_, clk);
  dff _29870_ (\oc8051_top_1.oc8051_memory_interface1.pc [13], _01870_, clk);
  dff _29871_ (\oc8051_top_1.oc8051_memory_interface1.pc [14], _01865_, clk);
  dff _29872_ (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03726_, clk);
  dff _29873_ (\oc8051_top_1.oc8051_memory_interface1.int_ack , _14022_, clk);
  dff _29874_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _03331_, clk);
  dff _29875_ (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _03350_, clk);
  dff _29876_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _01023_, clk);
  dff _29877_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _01000_, clk);
  dff _29878_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _10112_, clk);
  dff _29879_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _01734_, clk);
  dff _29880_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _01732_, clk);
  dff _29881_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _01697_, clk);
  dff _29882_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _01695_, clk);
  dff _29883_ (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _03329_, clk);
  dff _29884_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _09655_, clk);
  dff _29885_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _00647_, clk);
  dff _29886_ (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _03315_, clk);
  dff _29887_ (\oc8051_top_1.oc8051_memory_interface1.reti , _03444_, clk);
  dff _29888_ (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _10129_, clk);
  dff _29889_ (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _00160_, clk);
  dff _29890_ (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _00121_, clk);
  dff _29891_ (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _00148_, clk);
  dff _29892_ (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _00136_, clk);
  dff _29893_ (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _00130_, clk);
  dff _29894_ (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _00128_, clk);
  dff _29895_ (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03428_, clk);
  dff _29896_ (\oc8051_top_1.oc8051_memory_interface1.cdone , _03420_, clk);
  dff _29897_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _03413_, clk);
  dff _29898_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _14255_, clk);
  dff _29899_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _14227_, clk);
  dff _29900_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _14225_, clk);
  dff _29901_ (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _00256_, clk);
  dff _29902_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _13207_, clk);
  dff _29903_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _13154_, clk);
  dff _29904_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _13137_, clk);
  dff _29905_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _13103_, clk);
  dff _29906_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _10142_, clk);
  dff _29907_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _09628_, clk);
  dff _29908_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _12121_, clk);
  dff _29909_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _12104_, clk);
  dff _29910_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _12057_, clk);
  dff _29911_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _10446_, clk);
  dff _29912_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _12478_, clk);
  dff _29913_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _12405_, clk);
  dff _29914_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _12475_, clk);
  dff _29915_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _12445_, clk);
  dff _29916_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _12441_, clk);
  dff _29917_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _12423_, clk);
  dff _29918_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _12414_, clk);
  dff _29919_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _10400_, clk);
  dff _29920_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _09624_, clk);
  dff _29921_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _09779_, clk);
  dff _29922_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11592_, clk);
  dff _29923_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _11544_, clk);
  dff _29924_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _10452_, clk);
  dff _29925_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _11826_, clk);
  dff _29926_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _11854_, clk);
  dff _29927_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _11847_, clk);
  dff _29928_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _11831_, clk);
  dff _29929_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _10449_, clk);
  dff _29930_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _09620_, clk);
  dff _29931_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _08105_, clk);
  dff _29932_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _03985_, clk);
  dff _29933_ (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _02597_, clk);
  dff _29934_ (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _03156_, clk);
  dff _29935_ (\oc8051_top_1.oc8051_memory_interface1.istb_t , _03146_, clk);
  dff _29936_ (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _03135_, clk);
  dff _29937_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01803_, clk);
  dff _29938_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01762_, clk);
  dff _29939_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01711_, clk);
  dff _29940_ (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01669_, clk);
  dff _29941_ (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _00261_, clk);
  dff _29942_ (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0], clk);
  dff _29943_ (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1], clk);
  dff _29944_ (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2], clk);
  dff _29945_ (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3], clk);
  dff _29946_ (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4], clk);
  dff _29947_ (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5], clk);
  dff _29948_ (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6], clk);
  dff _29949_ (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7], clk);
  dff _29950_ (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8], clk);
  dff _29951_ (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9], clk);
  dff _29952_ (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10], clk);
  dff _29953_ (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11], clk);
  dff _29954_ (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12], clk);
  dff _29955_ (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13], clk);
  dff _29956_ (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14], clk);
  dff _29957_ (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15], clk);
  dff _29958_ (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16], clk);
  dff _29959_ (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17], clk);
  dff _29960_ (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18], clk);
  dff _29961_ (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19], clk);
  dff _29962_ (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20], clk);
  dff _29963_ (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21], clk);
  dff _29964_ (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22], clk);
  dff _29965_ (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23], clk);
  dff _29966_ (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24], clk);
  dff _29967_ (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25], clk);
  dff _29968_ (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26], clk);
  dff _29969_ (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27], clk);
  dff _29970_ (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28], clk);
  dff _29971_ (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29], clk);
  dff _29972_ (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30], clk);
  dff _29973_ (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31], clk);
  dff _29974_ (\oc8051_top_1.oc8051_sfr1.pres_ow , _04227_, clk);
  dff _29975_ (\oc8051_top_1.oc8051_sfr1.prescaler [0], _01821_, clk);
  dff _29976_ (\oc8051_top_1.oc8051_sfr1.prescaler [1], _14087_, clk);
  dff _29977_ (\oc8051_top_1.oc8051_sfr1.prescaler [2], _14082_, clk);
  dff _29978_ (\oc8051_top_1.oc8051_sfr1.prescaler [3], _04224_, clk);
  dff _29979_ (\oc8051_top_1.oc8051_sfr1.bit_out , _04219_, clk);
  dff _29980_ (\oc8051_top_1.oc8051_sfr1.wait_data , _04570_, clk);
  dff _29981_ (\oc8051_top_1.oc8051_sfr1.dat0 [0], _01825_, clk);
  dff _29982_ (\oc8051_top_1.oc8051_sfr1.dat0 [1], _13592_, clk);
  dff _29983_ (\oc8051_top_1.oc8051_sfr1.dat0 [2], _13580_, clk);
  dff _29984_ (\oc8051_top_1.oc8051_sfr1.dat0 [3], _13573_, clk);
  dff _29985_ (\oc8051_top_1.oc8051_sfr1.dat0 [4], _01823_, clk);
  dff _29986_ (\oc8051_top_1.oc8051_sfr1.dat0 [5], _01187_, clk);
  dff _29987_ (\oc8051_top_1.oc8051_sfr1.dat0 [6], _13423_, clk);
  dff _29988_ (\oc8051_top_1.oc8051_sfr1.dat0 [7], _04355_, clk);
  dff _29989_ (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _04353_, clk);
  dff _29990_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _06542_, clk);
  dff _29991_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _06536_, clk);
  dff _29992_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _03047_, clk);
  dff _29993_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _06641_, clk);
  dff _29994_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _06638_, clk);
  dff _29995_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _06626_, clk);
  dff _29996_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _02542_, clk);
  dff _29997_ (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _09804_, clk);
  dff _29998_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _03687_, clk);
  dff _29999_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _02805_, clk);
  dff _30000_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _02759_, clk);
  dff _30001_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _02563_, clk);
  dff _30002_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _02622_, clk);
  dff _30003_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _01201_, clk);
  dff _30004_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _02756_, clk);
  dff _30005_ (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _04485_, clk);
  dff _30006_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _07834_, clk);
  dff _30007_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _07829_, clk);
  dff _30008_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _07820_, clk);
  dff _30009_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _07806_, clk);
  dff _30010_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _07785_, clk);
  dff _30011_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _07767_, clk);
  dff _30012_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _07764_, clk);
  dff _30013_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _13651_, clk);
  dff _30014_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _07578_, clk);
  dff _30015_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _07635_, clk);
  dff _30016_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _07620_, clk);
  dff _30017_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _07616_, clk);
  dff _30018_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _07592_, clk);
  dff _30019_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _07584_, clk);
  dff _30020_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _07581_, clk);
  dff _30021_ (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _13649_, clk);
  dff _30022_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _02576_, clk);
  dff _30023_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00348_, clk);
  dff _30024_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00345_, clk);
  dff _30025_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00327_, clk);
  dff _30026_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00325_, clk);
  dff _30027_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00321_, clk);
  dff _30028_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00318_, clk);
  dff _30029_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00310_, clk);
  dff _30030_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _12565_, clk);
  dff _30031_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00289_, clk);
  dff _30032_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _12832_, clk);
  dff _30033_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _12851_, clk);
  dff _30034_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00275_, clk);
  dff _30035_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00272_, clk);
  dff _30036_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _03486_, clk);
  dff _30037_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00254_, clk);
  dff _30038_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00252_, clk);
  dff _30039_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _13415_, clk);
  dff _30040_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00228_, clk);
  dff _30041_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00222_, clk);
  dff _30042_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _04835_, clk);
  dff _30043_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _04978_, clk);
  dff _30044_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _05002_, clk);
  dff _30045_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _01362_, clk);
  dff _30046_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00181_, clk);
  dff _30047_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00179_, clk);
  dff _30048_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00162_, clk);
  dff _30049_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _04527_, clk);
  dff _30050_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00140_, clk);
  dff _30051_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00138_, clk);
  dff _30052_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00123_, clk);
  dff _30053_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00111_, clk);
  dff _30054_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00119_, clk);
  dff _30055_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00117_, clk);
  dff _30056_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00113_, clk);
  dff _30057_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _04529_, clk);
  dff _30058_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00050_, clk);
  dff _30059_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00048_, clk);
  dff _30060_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00031_, clk);
  dff _30061_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00028_, clk);
  dff _30062_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00026_, clk);
  dff _30063_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00024_, clk);
  dff _30064_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00009_, clk);
  dff _30065_ (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _04539_, clk);
  dff _30066_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _02937_, clk);
  dff _30067_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _02911_, clk);
  dff _30068_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _03081_, clk);
  dff _30069_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _02939_, clk);
  dff _30070_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _03079_, clk);
  dff _30071_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _02909_, clk);
  dff _30072_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _03077_, clk);
  dff _30073_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _00018_, clk);
  dff _30074_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _02935_, clk);
  dff _30075_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _03087_, clk);
  dff _30076_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _02907_, clk);
  dff _30077_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _03083_, clk);
  dff _30078_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _03055_, clk);
  dff _30079_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _03053_, clk);
  dff _30080_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _02933_, clk);
  dff _30081_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _14607_, clk);
  dff _30082_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _03091_, clk);
  dff _30083_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _02903_, clk);
  dff _30084_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _03089_, clk);
  dff _30085_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _03058_, clk);
  dff _30086_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _03057_, clk);
  dff _30087_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _02905_, clk);
  dff _30088_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _03085_, clk);
  dff _30089_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _07448_, clk);
  dff _30090_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _02928_, clk);
  dff _30091_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _02899_, clk);
  dff _30092_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _03098_, clk);
  dff _30093_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _02930_, clk);
  dff _30094_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _03095_, clk);
  dff _30095_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _02900_, clk);
  dff _30096_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _03093_, clk);
  dff _30097_ (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _00502_, clk);
  dff _30098_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _03873_, clk);
  dff _30099_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _03864_, clk);
  dff _30100_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _03825_, clk);
  dff _30101_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _03793_, clk);
  dff _30102_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _03127_, clk);
  dff _30103_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _03561_, clk);
  dff _30104_ (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _03209_, clk);
  dff _30105_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _03456_, clk);
  dff _30106_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _04799_, clk);
  dff _30107_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _04801_, clk);
  dff _30108_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _04805_, clk);
  dff _30109_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _04813_, clk);
  dff _30110_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _04815_, clk);
  dff _30111_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _04817_, clk);
  dff _30112_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _04819_, clk);
  dff _30113_ (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _03475_, clk);
  dff _30114_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _02689_, clk);
  dff _30115_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _02698_, clk);
  dff _30116_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _14456_, clk);
  dff _30117_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _14121_, clk);
  dff _30118_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _14115_, clk);
  dff _30119_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _14118_, clk);
  dff _30120_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _14111_, clk);
  dff _30121_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _14105_, clk);
  dff _30122_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _14108_, clk);
  dff _30123_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _02695_, clk);
  dff _30124_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _14127_, clk);
  dff _30125_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _14085_, clk);
  dff _30126_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _14090_, clk);
  dff _30127_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _14072_, clk);
  dff _30128_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _14075_, clk);
  dff _30129_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _14064_, clk);
  dff _30130_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _14059_, clk);
  dff _30131_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _02692_, clk);
  dff _30132_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _02684_, clk);
  dff _30133_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _02683_, clk);
  dff _30134_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _14006_, clk);
  dff _30135_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _14009_, clk);
  dff _30136_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _13910_, clk);
  dff _30137_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _13907_, clk);
  dff _30138_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _13908_, clk);
  dff _30139_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _13802_, clk);
  dff _30140_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _13798_, clk);
  dff _30141_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _02680_, clk);
  dff _30142_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _13788_, clk);
  dff _30143_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _13817_, clk);
  dff _30144_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _13809_, clk);
  dff _30145_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _13815_, clk);
  dff _30146_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _13812_, clk);
  dff _30147_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _13766_, clk);
  dff _30148_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _13768_, clk);
  dff _30149_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _02671_, clk);
  dff _30150_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _02677_, clk);
  dff _30151_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _13745_, clk);
  dff _30152_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _13710_, clk);
  dff _30153_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _13707_, clk);
  dff _30154_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _13729_, clk);
  dff _30155_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _13735_, clk);
  dff _30156_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _13919_, clk);
  dff _30157_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _13914_, clk);
  dff _30158_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _02668_, clk);
  dff _30159_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _09976_, clk);
  dff _30160_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _08250_, clk);
  dff _30161_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _08297_, clk);
  dff _30162_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _08321_, clk);
  dff _30163_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _03971_, clk);
  dff _30164_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _03966_, clk);
  dff _30165_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _03942_, clk);
  dff _30166_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _03917_, clk);
  dff _30167_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _03929_, clk);
  dff _30168_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _03926_, clk);
  dff _30169_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _03920_, clk);
  dff _30170_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _08181_, clk);
  dff _30171_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _03862_, clk);
  dff _30172_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _03791_, clk);
  dff _30173_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _03821_, clk);
  dff _30174_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _03805_, clk);
  dff _30175_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _03802_, clk);
  dff _30176_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _03799_, clk);
  dff _30177_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _03761_, clk);
  dff _30178_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _08108_, clk);
  dff _30179_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _08266_, clk);
  dff _30180_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _03698_, clk);
  dff _30181_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _03679_, clk);
  dff _30182_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _03675_, clk);
  dff _30183_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _03672_, clk);
  dff _30184_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _03669_, clk);
  dff _30185_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _04896_, clk);
  dff _30186_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _04889_, clk);
  dff _30187_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _08330_, clk);
  dff _30188_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _04945_, clk);
  dff _30189_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _04924_, clk);
  dff _30190_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _04920_, clk);
  dff _30191_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _04916_, clk);
  dff _30192_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _04909_, clk);
  dff _30193_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _04594_, clk);
  dff _30194_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _04592_, clk);
  dff _30195_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _10680_, clk);
  dff _30196_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _13884_, clk);
  dff _30197_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _04555_, clk);
  dff _30198_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _04550_, clk);
  dff _30199_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _04547_, clk);
  dff _30200_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _04544_, clk);
  dff _30201_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _03622_, clk);
  dff _30202_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _03619_, clk);
  dff _30203_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _03617_, clk);
  dff _30204_ (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _11486_, clk);
  dff _30205_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _08094_, clk);
  dff _30206_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _07997_, clk);
  dff _30207_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _07969_, clk);
  dff _30208_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _07992_, clk);
  dff _30209_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _07989_, clk);
  dff _30210_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _07976_, clk);
  dff _30211_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _07973_, clk);
  dff _30212_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _07959_, clk);
  dff _30213_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _08054_, clk);
  dff _30214_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _08100_, clk);
  dff _30215_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _08097_, clk);
  dff _30216_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _13093_, clk);
  dff _30217_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _12170_, clk);
  dff _30218_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _12160_, clk);
  dff _30219_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00213_, clk);
  dff _30220_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _12208_, clk);
  dff _30221_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _12229_, clk);
  dff _30222_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _12220_, clk);
  dff _30223_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _02284_, clk);
  dff _30224_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _12214_, clk);
  dff _30225_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _02225_, clk);
  dff _30226_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _08809_, clk);
  dff _30227_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _03479_, clk);
  dff _30228_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _12211_, clk);
  dff _30229_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _00465_, clk);
  dff _30230_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _00453_, clk);
  dff _30231_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _14139_, clk);
  dff _30232_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _13758_, clk);
  dff _30233_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _12863_, clk);
  dff _30234_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _12440_, clk);
  dff _30235_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _11465_, clk);
  dff _30236_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00188_, clk);
  dff _30237_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _12085_, clk);
  dff _30238_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _12082_, clk);
  dff _30239_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _12075_, clk);
  dff _30240_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _12060_, clk);
  dff _30241_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _01896_, clk);
  dff _30242_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _03422_, clk);
  dff _30243_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _00794_, clk);
  dff _30244_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _12052_, clk);
  dff _30245_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _04872_, clk);
  dff _30246_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _04848_, clk);
  dff _30247_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _04843_, clk);
  dff _30248_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _04563_, clk);
  dff _30249_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _04560_, clk);
  dff _30250_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _04557_, clk);
  dff _30251_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _04339_, clk);
  dff _30252_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _04334_, clk);
  dff _30253_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _04282_, clk);
  dff _30254_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _04187_, clk);
  dff _30255_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00230_, clk);
  dff _30256_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _02723_, clk);
  dff _30257_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _02705_, clk);
  dff _30258_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _02703_, clk);
  dff _30259_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _02300_, clk);
  dff _30260_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _02286_, clk);
  dff _30261_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _02185_, clk);
  dff _30262_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _02212_, clk);
  dff _30263_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _12115_, clk);
  dff _30264_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01673_, clk);
  dff _30265_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01649_, clk);
  dff _30266_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _00219_, clk);
  dff _30267_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _00639_, clk);
  dff _30268_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _00570_, clk);
  dff _30269_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _00334_, clk);
  dff _30270_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _13365_, clk);
  dff _30271_ (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _12128_, clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
endmodule
