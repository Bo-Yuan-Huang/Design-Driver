
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid_ajmp, ABINPUT, ABINPUT000, ABINPUT000000);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  input [8:0] ABINPUT;
  input [16:0] ABINPUT000;
  input [16:0] ABINPUT000000;
  input clk;
  wire [31:0] cxrom_data_out;
  wire cy;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [16:0] \oc8051_top_1.ABINPUT000 ;
  wire [16:0] \oc8051_top_1.ABINPUT000000 ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT ;
  wire [16:0] \oc8051_top_1.oc8051_alu1.ABINPUT000 ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire \oc8051_top_1.oc8051_alu1.divOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.mulOv ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.mulsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid_ajmp;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  not (_04856_, rst);
  not (_04857_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  not (_04858_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not (_04859_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_04860_, \oc8051_top_1.oc8051_decoder1.wr , _04859_);
  and (_04861_, _04860_, _04858_);
  and (_04862_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_04863_, _04862_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_04864_, _04863_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_04865_, _04864_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_04866_, _04865_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  and (_04867_, _04866_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_04868_, _04867_);
  not (_04869_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_04870_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _04859_);
  and (_04871_, _04870_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_04872_, _04871_, _04869_);
  or (_04873_, _04866_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  and (_04874_, _04873_, _04872_);
  nand (_04875_, _04874_, _04868_);
  and (_04876_, _04871_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_04877_, _04876_);
  not (_04878_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_04879_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _04859_);
  and (_04880_, _04879_, _04878_);
  and (_04881_, _04880_, _04869_);
  nand (_04882_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  and (_04883_, _04882_, _04877_);
  and (_04884_, _04870_, _04869_);
  not (_04885_, _04884_);
  nor (_04886_, _04885_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  nand (_04887_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_04888_, _04880_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  nand (_04889_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  and (_04890_, _04889_, _04887_);
  and (_04892_, _04890_, _04883_);
  and (_04893_, _04892_, _04875_);
  nand (_04894_, _04867_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  or (_04895_, _04867_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  and (_04896_, _04895_, _04894_);
  nand (_04897_, _04896_, _04872_);
  nand (_04898_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_04899_, _04898_, _04877_);
  nand (_04900_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nand (_04901_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_04902_, _04901_, _04900_);
  and (_04903_, _04902_, _04899_);
  and (_04904_, _04903_, _04897_);
  and (_04905_, _04904_, _04893_);
  not (_04906_, _04865_);
  or (_04907_, _04864_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  and (_04908_, _04907_, _04872_);
  and (_04909_, _04908_, _04906_);
  not (_04910_, _04909_);
  nand (_04911_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  and (_04912_, _04911_, _04877_);
  nor (_04913_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  nor (_04914_, _04913_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_04915_, _04914_, _04879_);
  nand (_04916_, _04915_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nand (_04917_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  and (_04918_, _04917_, _04916_);
  nand (_04919_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_04920_, _04919_, _04918_);
  and (_04921_, _04920_, _04912_);
  and (_04922_, _04921_, _04910_);
  or (_04923_, _04865_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nand (_04924_, _04923_, _04872_);
  or (_04925_, _04924_, _04866_);
  nand (_04926_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nand (_04927_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_04928_, _04927_, _04926_);
  nand (_04929_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_04930_, _04929_, _04877_);
  and (_04931_, _04930_, _04928_);
  and (_04932_, _04931_, _04925_);
  not (_04933_, _04932_);
  nor (_04934_, _04933_, _04922_);
  and (_04935_, _04934_, _04905_);
  and (_04936_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  and (_04937_, _04881_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_04938_, _04937_, _04936_);
  nor (_04939_, _04863_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_04940_, _04939_, _04864_);
  and (_04941_, _04940_, _04872_);
  not (_04942_, _04941_);
  nand (_04943_, _04915_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nand (_04944_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  and (_04945_, _04944_, _04943_);
  and (_04946_, _04945_, _04942_);
  and (_04947_, _04946_, _04938_);
  not (_04948_, _04947_);
  nand (_04949_, _04888_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  nand (_04950_, _04915_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  and (_04951_, _04950_, _04949_);
  not (_04952_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nand (_04953_, _04872_, _04952_);
  nand (_04954_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nand (_04955_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  and (_04956_, _04955_, _04954_);
  and (_04957_, _04956_, _04953_);
  and (_04958_, _04957_, _04951_);
  not (_04959_, _04958_);
  nor (_04960_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_04961_, _04960_, _04862_);
  nand (_04962_, _04961_, _04872_);
  nand (_04963_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  and (_04964_, _04963_, _04962_);
  nand (_04965_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand (_04966_, _04888_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  nand (_04967_, _04915_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  and (_04968_, _04967_, _04966_);
  and (_04969_, _04968_, _04965_);
  and (_04971_, _04969_, _04964_);
  not (_04972_, _04872_);
  nor (_04973_, _04862_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  or (_04974_, _04973_, _04863_);
  or (_04975_, _04974_, _04972_);
  nand (_04976_, _04886_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  and (_04977_, _04976_, _04975_);
  nand (_04978_, _04881_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  nand (_04979_, _04888_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  nand (_04980_, _04915_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  and (_04981_, _04980_, _04979_);
  and (_04982_, _04981_, _04978_);
  and (_04984_, _04982_, _04977_);
  and (_04985_, _04984_, _04971_);
  and (_04986_, _04985_, _04959_);
  and (_04987_, _04986_, _04948_);
  and (_04988_, _04987_, _04935_);
  and (_04989_, _04971_, _04958_);
  and (_04990_, _04989_, _04984_);
  and (_04991_, _04990_, _04948_);
  and (_04992_, _04991_, _04935_);
  and (_04993_, _04932_, _04922_);
  and (_04994_, _04993_, _04905_);
  and (_04995_, _04994_, _04985_);
  not (_04996_, _04971_);
  nor (_04997_, _04996_, _04958_);
  and (_04998_, _04984_, _04947_);
  and (_04999_, _04998_, _04997_);
  and (_05000_, _04999_, _04935_);
  and (_05001_, _04998_, _04989_);
  and (_05002_, _05001_, _04935_);
  or (_05003_, _05002_, _05000_);
  or (_05004_, _05003_, _04995_);
  or (_05005_, _05004_, _04992_);
  or (_05006_, _05005_, _04988_);
  nand (_05007_, _05006_, _04861_);
  and (_05008_, _05005_, _04861_);
  nor (_05009_, _05008_, _05007_);
  nor (_05010_, _05009_, _04857_);
  not (_05011_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  not (_05012_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  not (_05013_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_05014_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], _05013_);
  nand (_05015_, _05014_, _05012_);
  nor (_05016_, _05015_, _05011_);
  not (_05017_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  or (_05018_, _05012_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or (_05019_, _05018_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nor (_05020_, _05019_, _05017_);
  nor (_05021_, _05020_, _05016_);
  not (_05022_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  or (_05023_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  or (_05024_, _05023_, _05013_);
  nor (_05025_, _05024_, _05022_);
  not (_05026_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  or (_05027_, _05018_, _05013_);
  nor (_05028_, _05027_, _05026_);
  nor (_05029_, _05028_, _05025_);
  and (_05030_, _05029_, _05021_);
  not (_05031_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_05032_, _05031_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  nor (_05033_, _05032_, ABINPUT[7]);
  nand (_05034_, _05031_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  nor (_05035_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nor (_05036_, _05035_, _05033_);
  nor (_05037_, _05023_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_05038_, _05037_, _05036_);
  and (_05039_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_05040_, _05039_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_05041_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  not (_05042_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nand (_05043_, _05039_, _05013_);
  nor (_05044_, _05043_, _05042_);
  nor (_05045_, _05044_, _05041_);
  not (_05046_, _05045_);
  nor (_05047_, _05046_, _05038_);
  and (_05048_, _05047_, _05030_);
  not (_05049_, _05048_);
  or (_05050_, _05032_, ABINPUT[0]);
  or (_05051_, _05034_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nand (_05052_, _05051_, _05050_);
  not (_05053_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  nand (_05054_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  and (_05055_, _05054_, _05053_);
  or (_05056_, _05055_, _05052_);
  not (_05057_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_05058_, _05055_, _05057_);
  nand (_05059_, _05058_, _05056_);
  not (_05060_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  nor (_05061_, _05015_, _05060_);
  not (_05062_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  nor (_05063_, _05019_, _05062_);
  nor (_05064_, _05063_, _05061_);
  not (_05065_, _05027_);
  and (_05066_, _05065_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_05067_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_05068_, _05024_, _05067_);
  nor (_05069_, _05068_, _05066_);
  and (_05070_, _05069_, _05064_);
  nor (_05071_, _05032_, ABINPUT[5]);
  nor (_05072_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nor (_05073_, _05072_, _05071_);
  and (_05074_, _05073_, _05037_);
  not (_05075_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_05076_, _05043_, _05075_);
  and (_05077_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nor (_05078_, _05077_, _05076_);
  not (_05079_, _05078_);
  nor (_05080_, _05079_, _05074_);
  and (_05081_, _05080_, _05070_);
  not (_05082_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  or (_05083_, _05015_, _05082_);
  not (_05084_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  or (_05085_, _05019_, _05084_);
  and (_05086_, _05085_, _05083_);
  not (_05087_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_05088_, _05027_, _05087_);
  not (_05089_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_05090_, _05024_, _05089_);
  nor (_05091_, _05090_, _05088_);
  and (_05092_, _05091_, _05086_);
  not (_05093_, _05037_);
  or (_05094_, _05032_, ABINPUT[4]);
  or (_05095_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_05096_, _05095_, _05094_);
  or (_05097_, _05096_, _05093_);
  and (_05098_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  not (_05099_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_05100_, _05043_, _05099_);
  nor (_05101_, _05100_, _05098_);
  and (_05102_, _05101_, _05097_);
  and (_05103_, _05102_, _05092_);
  not (_05104_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  or (_05105_, _05019_, _05104_);
  not (_05106_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  or (_05107_, _05015_, _05106_);
  and (_05108_, _05107_, _05105_);
  not (_05109_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_05110_, _05027_, _05109_);
  not (_05111_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_05112_, _05024_, _05111_);
  and (_05114_, _05112_, _05110_);
  and (_05115_, _05114_, _05108_);
  or (_05117_, _05032_, ABINPUT[1]);
  or (_05118_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  nand (_05119_, _05118_, _05117_);
  or (_05120_, _05119_, _05093_);
  nand (_05121_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  not (_05122_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_05123_, _05043_, _05122_);
  and (_05124_, _05123_, _05121_);
  and (_05125_, _05124_, _05120_);
  and (_05126_, _05125_, _05115_);
  or (_05128_, _05032_, ABINPUT[2]);
  or (_05129_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_05130_, _05129_, _05128_);
  or (_05131_, _05130_, _05093_);
  not (_05132_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  or (_05134_, _05019_, _05132_);
  not (_05135_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  or (_05137_, _05015_, _05135_);
  and (_05138_, _05137_, _05134_);
  and (_05139_, _05138_, _05131_);
  not (_05140_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_05141_, _05027_, _05140_);
  not (_05142_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_05144_, _05024_, _05142_);
  and (_05145_, _05144_, _05141_);
  nand (_05146_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  not (_05147_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_05148_, _05043_, _05147_);
  and (_05149_, _05148_, _05146_);
  and (_05150_, _05149_, _05145_);
  and (_05151_, _05150_, _05139_);
  not (_05152_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_05153_, _05019_, _05152_);
  not (_05154_, \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  or (_05155_, _05015_, _05154_);
  and (_05156_, _05155_, _05153_);
  not (_05157_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_05158_, _05024_, _05157_);
  not (_05159_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_05160_, _05027_, _05159_);
  and (_05161_, _05160_, _05158_);
  and (_05162_, _05161_, _05156_);
  or (_05163_, _05032_, ABINPUT[3]);
  or (_05164_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_05165_, _05164_, _05163_);
  or (_05166_, _05165_, _05093_);
  not (_05167_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_05168_, _05043_, _05167_);
  nand (_05169_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  and (_05170_, _05169_, _05168_);
  and (_05171_, _05170_, _05166_);
  and (_05172_, _05171_, _05162_);
  and (_05173_, _05172_, _05151_);
  and (_05174_, _05173_, _05126_);
  and (_05175_, _05174_, _05103_);
  and (_05176_, _05175_, _05081_);
  not (_05177_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  nor (_05178_, _05015_, _05177_);
  not (_05179_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  nor (_05180_, _05019_, _05179_);
  nor (_05181_, _05180_, _05178_);
  not (_05183_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  nor (_05184_, _05027_, _05183_);
  not (_05185_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_05186_, _05024_, _05185_);
  nor (_05187_, _05186_, _05184_);
  and (_05188_, _05187_, _05181_);
  nor (_05189_, _05032_, ABINPUT[6]);
  nor (_05190_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nor (_05191_, _05190_, _05189_);
  and (_05192_, _05191_, _05037_);
  and (_05193_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  not (_05194_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_05195_, _05043_, _05194_);
  nor (_05196_, _05195_, _05193_);
  not (_05197_, _05196_);
  nor (_05198_, _05197_, _05192_);
  and (_05199_, _05198_, _05188_);
  nand (_05201_, _05199_, _05176_);
  nand (_05202_, _05201_, _05059_);
  not (_05204_, _05103_);
  not (_05205_, _05172_);
  nand (_05206_, _05125_, _05115_);
  nand (_05207_, _05150_, _05139_);
  and (_05208_, _05207_, _05206_);
  and (_05209_, _05208_, _05205_);
  and (_05210_, _05209_, _05204_);
  nor (_05211_, _05199_, _05081_);
  and (_05212_, _05211_, _05210_);
  or (_05213_, _05212_, _05059_);
  and (_05214_, _05213_, _05202_);
  nand (_05215_, _05214_, _05049_);
  not (_05216_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_05217_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _04859_);
  and (_05218_, _05217_, _05216_);
  and (_05220_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _04859_);
  and (_05221_, _05220_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_05223_, _05221_, _05218_);
  or (_05224_, _05214_, _05049_);
  and (_05225_, _05224_, _05223_);
  and (_05226_, _05225_, _05215_);
  and (_05227_, _05058_, _05056_);
  and (_05228_, _05227_, _05048_);
  not (_05229_, _05228_);
  and (_05230_, _05217_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_05231_, _05230_, _05221_);
  not (_05232_, _05231_);
  nor (_05233_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_05234_, _05233_, _05036_);
  not (_05236_, _05234_);
  and (_05237_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_05238_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  not (_05239_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_05240_, _05239_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  and (_05241_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_05242_, _05241_, _05238_);
  and (_05243_, _05242_, _05236_);
  and (_05244_, _05243_, _05059_);
  nor (_05245_, _05244_, _05232_);
  and (_05246_, _05245_, _05229_);
  nor (_05247_, _05246_, _05226_);
  and (_05248_, _05243_, _05048_);
  not (_05249_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_05250_, _04859_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_05252_, _05250_, _05249_);
  not (_05253_, _05220_);
  nor (_05254_, _05253_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_05255_, _05254_, _05252_);
  not (_05256_, _05255_);
  nor (_05257_, _05256_, _05248_);
  nor (_05258_, _05250_, _05217_);
  and (_05259_, _05258_, _05254_);
  nor (_05260_, _05243_, _05048_);
  nor (_05261_, _05260_, _05248_);
  and (_05262_, _05261_, _05259_);
  nor (_05263_, _05262_, _05257_);
  not (_05264_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_05265_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _04859_);
  and (_05266_, _05265_, _05264_);
  and (_05267_, _05266_, _05230_);
  and (_05268_, _05267_, _05260_);
  and (_05269_, _05266_, _05218_);
  and (_05270_, _05269_, _05048_);
  nor (_05271_, _05270_, _05268_);
  nor (_05272_, _05265_, _05220_);
  and (_05273_, _05272_, _05258_);
  not (_05274_, _05273_);
  nand (_05275_, _05272_, _05250_);
  nand (_05276_, _05266_, _05249_);
  and (_05277_, _05276_, _05275_);
  and (_05278_, _05277_, _05274_);
  and (_05279_, _05221_, _05249_);
  and (_05280_, _05254_, _05217_);
  nor (_05281_, _05280_, _05279_);
  and (_05282_, _05281_, _05278_);
  nor (_05283_, _05282_, _05048_);
  not (_05284_, _05283_);
  and (_05285_, _05284_, _05271_);
  and (_05286_, _05285_, _05263_);
  and (_05287_, _05286_, _05247_);
  not (_05288_, _05287_);
  and (_05289_, _05288_, _05009_);
  or (_05290_, _05289_, _05010_);
  and (_13054_, _05290_, _04856_);
  and (_05291_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _04859_);
  and (_05292_, _05291_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  not (_05293_, _05292_);
  nor (_05294_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_05295_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_05296_, _05295_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_05297_, _05296_, _05294_);
  not (_05298_, _05297_);
  nor (_05299_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_05300_, _05022_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_05301_, _05300_, _05299_);
  not (_05303_, _05301_);
  nor (_05304_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_05305_, _05185_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_05306_, _05305_, _05304_);
  not (_05307_, _05306_);
  nor (_05308_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_05309_, _05089_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_05310_, _05309_, _05308_);
  nor (_05312_, _05032_, ABINPUT[8]);
  nor (_05313_, _05034_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nor (_05314_, _05313_, _05312_);
  and (_05315_, _05314_, _05233_);
  not (_05316_, _05315_);
  and (_05317_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  and (_05318_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_05319_, _05318_, _05317_);
  and (_05320_, _05319_, _05316_);
  not (_05321_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nor (_05322_, _05019_, _05321_);
  not (_05323_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  nor (_05324_, _05015_, _05323_);
  nor (_05325_, _05324_, _05322_);
  nor (_05326_, _05024_, _05295_);
  not (_05327_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_05328_, _05027_, _05327_);
  nor (_05329_, _05328_, _05326_);
  and (_05330_, _05329_, _05325_);
  and (_05331_, _05314_, _05037_);
  not (_05332_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_05333_, _05043_, _05332_);
  and (_05334_, _05040_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  nor (_05335_, _05334_, _05333_);
  not (_05336_, _05335_);
  nor (_05337_, _05336_, _05331_);
  and (_05338_, _05337_, _05330_);
  nor (_05339_, _05338_, _05320_);
  not (_05340_, _05339_);
  and (_05341_, _05233_, _05073_);
  not (_05342_, _05341_);
  and (_05343_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  and (_05344_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_05345_, _05344_, _05343_);
  and (_05346_, _05345_, _05342_);
  nor (_05347_, _05346_, _05081_);
  and (_05348_, _05346_, _05081_);
  nor (_05349_, _05348_, _05347_);
  not (_05350_, _05233_);
  nor (_05351_, _05350_, _05096_);
  not (_05352_, _05351_);
  and (_05353_, _05237_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  and (_05354_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_05355_, _05354_, _05353_);
  and (_05356_, _05355_, _05352_);
  nor (_05357_, _05356_, _05103_);
  and (_05359_, _05356_, _05103_);
  nor (_05360_, _05359_, _05357_);
  not (_05362_, _05360_);
  or (_05363_, _05350_, _05165_);
  and (_05365_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and (_05366_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_05367_, _05366_, _05365_);
  and (_05368_, _05367_, _05363_);
  nor (_05369_, _05368_, _05172_);
  not (_05370_, _05369_);
  and (_05371_, _05368_, _05172_);
  nor (_05372_, _05371_, _05369_);
  or (_05373_, _05350_, _05130_);
  nand (_05374_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  nand (_05375_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_05376_, _05375_, _05374_);
  nand (_05377_, _05376_, _05373_);
  and (_05378_, _05377_, _05207_);
  or (_05379_, _05350_, _05119_);
  nand (_05380_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  nand (_05381_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  and (_05382_, _05381_, _05380_);
  and (_05383_, _05382_, _05379_);
  not (_05384_, _05383_);
  and (_05385_, _05384_, _05206_);
  and (_05386_, _05376_, _05373_);
  and (_05387_, _05386_, _05151_);
  nor (_05388_, _05387_, _05378_);
  and (_05389_, _05388_, _05385_);
  or (_05390_, _05389_, _05378_);
  nand (_05391_, _05390_, _05372_);
  nand (_05392_, _05391_, _05370_);
  and (_05393_, _05392_, _05362_);
  nor (_05394_, _05392_, _05362_);
  or (_05395_, _05394_, _05393_);
  and (_05396_, _05383_, _05126_);
  nor (_05397_, _05396_, _05385_);
  and (_05398_, _05397_, _05059_);
  and (_05399_, _05398_, _05388_);
  or (_05400_, _05390_, _05372_);
  and (_05401_, _05400_, _05391_);
  and (_05402_, _05401_, _05399_);
  and (_05403_, _05402_, _05395_);
  not (_05404_, _05359_);
  and (_05405_, _05392_, _05404_);
  or (_05406_, _05405_, _05357_);
  or (_05407_, _05406_, _05403_);
  nand (_05408_, _05407_, _05349_);
  and (_05409_, _05233_, _05191_);
  not (_05410_, _05409_);
  and (_05411_, _05237_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  and (_05412_, _05240_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nor (_05413_, _05412_, _05411_);
  and (_05414_, _05413_, _05410_);
  nor (_05415_, _05414_, _05199_);
  and (_05416_, _05414_, _05199_);
  nor (_05417_, _05416_, _05415_);
  and (_05418_, _05417_, _05347_);
  nor (_05419_, _05417_, _05347_);
  nor (_05420_, _05419_, _05418_);
  not (_05421_, _05420_);
  or (_05422_, _05421_, _05408_);
  not (_05423_, _05261_);
  nor (_05424_, _05418_, _05415_);
  nor (_05425_, _05424_, _05423_);
  and (_05426_, _05424_, _05423_);
  nor (_05427_, _05426_, _05425_);
  not (_05428_, _05427_);
  or (_05429_, _05428_, _05422_);
  nor (_05430_, _05425_, _05260_);
  and (_05431_, _05430_, _05429_);
  and (_05432_, _05338_, _05320_);
  or (_05433_, _05432_, _05431_);
  nand (_05434_, _05433_, _05340_);
  nor (_05435_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_05436_, _05111_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_05437_, _05436_, _05435_);
  and (_05438_, _05437_, _05434_);
  nor (_05439_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_05440_, _05142_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_05441_, _05440_, _05439_);
  and (_05442_, _05441_, _05438_);
  nor (_05443_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_05444_, _05157_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_05445_, _05444_, _05443_);
  and (_05446_, _05445_, _05442_);
  and (_05447_, _05446_, _05310_);
  nor (_05448_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_05449_, _05067_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_05450_, _05449_, _05448_);
  nand (_05451_, _05450_, _05447_);
  or (_05452_, _05451_, _05307_);
  or (_05453_, _05452_, _05303_);
  or (_05454_, _05453_, _05298_);
  and (_05455_, _05272_, _05252_);
  nand (_05456_, _05453_, _05298_);
  and (_05457_, _05456_, _05455_);
  and (_05458_, _05457_, _05454_);
  not (_05459_, _05320_);
  nor (_05460_, _05243_, _05059_);
  nor (_05461_, _05460_, _05244_);
  and (_05462_, _05199_, _05048_);
  and (_05463_, _05338_, _05462_);
  and (_05464_, _05463_, _05176_);
  and (_05465_, _05464_, _05383_);
  and (_05466_, _05465_, _05386_);
  and (_05467_, _05466_, _05368_);
  and (_05468_, _05467_, _05356_);
  and (_05469_, _05468_, _05346_);
  and (_05470_, _05414_, _05059_);
  nand (_05471_, _05470_, _05469_);
  not (_05472_, _05368_);
  nor (_05473_, _05338_, _05048_);
  and (_05474_, _05473_, _05211_);
  and (_05475_, _05474_, _05210_);
  and (_05476_, _05475_, _05384_);
  and (_05477_, _05476_, _05377_);
  and (_05478_, _05477_, _05472_);
  nor (_05479_, _05414_, _05059_);
  nor (_05480_, _05356_, _05346_);
  and (_05481_, _05480_, _05479_);
  nand (_05482_, _05481_, _05478_);
  and (_05483_, _05482_, _05471_);
  nor (_05484_, _05483_, _05461_);
  nand (_05485_, _05484_, _05459_);
  or (_05486_, _05484_, _05459_);
  and (_05487_, _05486_, _05485_);
  and (_05488_, _05487_, _05223_);
  and (_05489_, _05254_, _05230_);
  not (_05490_, _05489_);
  nor (_05491_, _05490_, _05103_);
  and (_05492_, _05231_, _05227_);
  or (_05493_, _05492_, _05273_);
  and (_05494_, _05493_, _05459_);
  or (_05495_, _05232_, _05227_);
  nor (_05496_, _05495_, _05338_);
  and (_05497_, _05266_, _05258_);
  and (_05498_, _05497_, ABINPUT000000[16]);
  and (_05499_, _05272_, _05230_);
  and (_05500_, _05499_, ABINPUT000[16]);
  or (_05501_, _05500_, _05498_);
  or (_05502_, _05501_, _05496_);
  or (_05503_, _05502_, _05494_);
  or (_05504_, _05503_, _05491_);
  or (_05506_, _05504_, _05488_);
  or (_05507_, _05506_, _05458_);
  or (_05509_, _05507_, _05293_);
  and (_05510_, _04861_, _04885_);
  and (_05512_, _05510_, _04947_);
  not (_05513_, _04893_);
  nor (_05515_, _04904_, _05513_);
  and (_05517_, _05515_, _04993_);
  nor (_05519_, _04971_, _04958_);
  and (_05520_, _05519_, _04984_);
  and (_05522_, _05520_, _05517_);
  and (_05524_, _05522_, _05512_);
  nor (_05525_, _05338_, _05274_);
  nor (_05526_, _05338_, _05059_);
  nor (_05527_, _05320_, _05227_);
  or (_05528_, _05527_, _05526_);
  and (_05529_, _05528_, _05231_);
  not (_05530_, _05338_);
  nor (_05531_, _05227_, _05048_);
  nor (_05532_, _05531_, _05228_);
  and (_05533_, _05532_, _05214_);
  nor (_05534_, _05533_, _05530_);
  and (_05535_, _05533_, _05530_);
  nor (_05536_, _05535_, _05534_);
  and (_05537_, _05536_, _05223_);
  nor (_05538_, _05537_, _05529_);
  and (_05540_, _05252_, _05221_);
  and (_05541_, _05540_, _05059_);
  and (_05542_, _05258_, _05221_);
  and (_05543_, _05542_, _05206_);
  nor (_05544_, _05543_, _05541_);
  nand (_05545_, _05544_, _05538_);
  and (_05546_, _05280_, _05049_);
  not (_05547_, _05546_);
  nor (_05548_, _05432_, _05256_);
  nor (_05549_, _05432_, _05339_);
  and (_05550_, _05549_, _05259_);
  nor (_05551_, _05550_, _05548_);
  nand (_05552_, _05551_, _05547_);
  or (_05553_, _05552_, _05545_);
  and (_05554_, _05339_, _05267_);
  and (_05555_, _05338_, _05269_);
  nor (_05556_, _05555_, _05554_);
  and (_05557_, _05266_, _05252_);
  not (_05558_, _05557_);
  nor (_05559_, _05173_, _05103_);
  and (_05560_, _05559_, _05557_);
  not (_05561_, _05560_);
  or (_05562_, _05338_, _05462_);
  and (_05563_, _05562_, _05227_);
  and (_05564_, _05563_, _05561_);
  not (_05565_, _05081_);
  and (_05567_, _05560_, _05565_);
  nor (_05568_, _05567_, _05564_);
  and (_05569_, _05568_, _05462_);
  or (_05570_, _05569_, _05564_);
  and (_05571_, _05570_, _05338_);
  nor (_05572_, _05570_, _05338_);
  or (_05573_, _05572_, _05571_);
  nor (_05574_, _05573_, _05558_);
  and (_05576_, _05497_, ABINPUT000000[8]);
  nor (_05577_, _05576_, _05574_);
  nand (_05578_, _05577_, _05556_);
  and (_05579_, _05549_, _05431_);
  nor (_05580_, _05549_, _05431_);
  or (_05581_, _05580_, _05579_);
  and (_05582_, _05581_, _05455_);
  and (_05583_, _05272_, _05218_);
  not (_05584_, _05583_);
  not (_05585_, _05549_);
  and (_05586_, _05243_, _05049_);
  not (_05587_, _05199_);
  and (_05588_, _05414_, _05587_);
  not (_05589_, _05346_);
  and (_05590_, _05589_, _05081_);
  nor (_05591_, _05417_, _05590_);
  nor (_05592_, _05591_, _05588_);
  nor (_05593_, _05592_, _05261_);
  nor (_05594_, _05593_, _05586_);
  and (_05595_, _05592_, _05261_);
  nor (_05596_, _05595_, _05593_);
  not (_05597_, _05596_);
  and (_05598_, _05417_, _05590_);
  nor (_05599_, _05598_, _05591_);
  not (_05600_, _05599_);
  not (_05601_, _05349_);
  nor (_05602_, _05472_, _05172_);
  or (_05603_, _05377_, _05151_);
  and (_05604_, _05384_, _05126_);
  or (_05605_, _05604_, _05388_);
  nand (_05606_, _05605_, _05603_);
  not (_05607_, _05606_);
  nor (_05608_, _05607_, _05372_);
  nor (_05609_, _05608_, _05602_);
  nor (_05610_, _05609_, _05360_);
  and (_05611_, _05609_, _05360_);
  or (_05612_, _05611_, _05610_);
  and (_05613_, _05607_, _05372_);
  or (_05614_, _05613_, _05608_);
  and (_05615_, _05604_, _05388_);
  not (_05616_, _05615_);
  nand (_05617_, _05616_, _05605_);
  nor (_05618_, _05397_, _05227_);
  and (_05619_, _05618_, _05617_);
  and (_05620_, _05619_, _05614_);
  and (_05621_, _05620_, _05612_);
  not (_05622_, _05356_);
  or (_05623_, _05622_, _05103_);
  and (_05624_, _05622_, _05103_);
  or (_05625_, _05609_, _05624_);
  and (_05626_, _05625_, _05623_);
  or (_05627_, _05626_, _05621_);
  and (_05628_, _05627_, _05601_);
  and (_05629_, _05628_, _05600_);
  and (_05630_, _05629_, _05597_);
  or (_05631_, _05630_, _05594_);
  and (_05632_, _05631_, _05585_);
  nor (_05633_, _05631_, _05585_);
  nor (_05634_, _05633_, _05632_);
  nor (_05635_, _05634_, _05584_);
  and (_05636_, _05499_, ABINPUT000[8]);
  or (_05637_, _05636_, _05635_);
  or (_05638_, _05637_, _05582_);
  or (_05639_, _05638_, _05578_);
  or (_05640_, _05639_, _05553_);
  or (_05641_, _05640_, _05525_);
  and (_05642_, _05641_, _05524_);
  not (_05643_, _05524_);
  and (_05644_, _05643_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_05645_, _05644_, _05292_);
  or (_05646_, _05645_, _05642_);
  and (_05647_, _05646_, _04856_);
  and (_03221_, _05647_, _05509_);
  nor (_05648_, _05356_, _05232_);
  nand (_05649_, _05209_, _05227_);
  nand (_05650_, _05174_, _05059_);
  and (_05651_, _05650_, _05649_);
  nand (_05652_, _05651_, _05103_);
  or (_05653_, _05651_, _05103_);
  and (_05654_, _05653_, _05223_);
  and (_05655_, _05654_, _05652_);
  nor (_05656_, _05655_, _05648_);
  nor (_05657_, _05282_, _05103_);
  not (_05658_, _05657_);
  and (_05659_, _05360_, _05259_);
  not (_05660_, _05659_);
  nor (_05661_, _05359_, _05256_);
  not (_05662_, _05661_);
  and (_05663_, _05357_, _05267_);
  and (_05664_, _05269_, _05103_);
  nor (_05665_, _05664_, _05663_);
  and (_05666_, _05665_, _05662_);
  and (_05667_, _05666_, _05660_);
  and (_05668_, _05667_, _05658_);
  and (_05669_, _05668_, _05656_);
  not (_05670_, _05669_);
  and (_05671_, _05002_, _04861_);
  and (_05672_, _05671_, _05670_);
  not (_05673_, _04861_);
  and (_05674_, _04991_, _04994_);
  and (_05675_, _04999_, _04994_);
  and (_05676_, _05001_, _04994_);
  or (_05677_, _05676_, _05675_);
  nor (_05678_, _05677_, _05674_);
  and (_05679_, _04994_, _04987_);
  nor (_05680_, _05002_, _05679_);
  and (_05681_, _05680_, _05678_);
  or (_05682_, _05681_, _05673_);
  or (_05683_, _05682_, _04995_);
  and (_05684_, _05683_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  or (_05685_, _05684_, _05672_);
  and (_04850_, _05685_, _04856_);
  and (_05686_, _05199_, _05227_);
  not (_05687_, _05686_);
  nor (_05688_, _05470_, _05232_);
  and (_05689_, _05688_, _05687_);
  and (_05690_, _05081_, _05227_);
  not (_05692_, _05690_);
  and (_05693_, _05210_, _05227_);
  or (_05694_, _05693_, _05176_);
  and (_05696_, _05694_, _05692_);
  or (_05698_, _05587_, _05696_);
  nand (_05699_, _05587_, _05696_);
  and (_05700_, _05699_, _05223_);
  and (_05701_, _05700_, _05698_);
  nor (_05702_, _05701_, _05689_);
  nor (_05703_, _05282_, _05199_);
  not (_05704_, _05703_);
  and (_05705_, _05417_, _05259_);
  not (_05707_, _05705_);
  nor (_05708_, _05416_, _05256_);
  not (_05710_, _05708_);
  and (_05711_, _05415_, _05267_);
  and (_05713_, _05269_, _05199_);
  nor (_05714_, _05713_, _05711_);
  and (_05715_, _05714_, _05710_);
  and (_05716_, _05715_, _05707_);
  and (_05717_, _05716_, _05704_);
  nand (_05718_, _05717_, _05702_);
  and (_05719_, _05000_, _04861_);
  and (_05720_, _05719_, _05718_);
  nand (_05721_, _05004_, _04861_);
  not (_05722_, _05721_);
  nand (_05723_, _05722_, _05682_);
  and (_05724_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  or (_05725_, _05724_, _05720_);
  and (_04852_, _05725_, _04856_);
  not (_05726_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor (_05727_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_05728_, _05727_, _05726_);
  nor (_05729_, \oc8051_top_1.oc8051_decoder1.state [0], \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_05730_, _05729_, _04859_);
  and (_05731_, _05730_, _05728_);
  not (_05732_, _05731_);
  not (_05733_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05734_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_05735_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  not (_05736_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not (_05737_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_05738_, _05737_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_05739_, _05738_, _05736_);
  or (_05740_, _05739_, _05735_);
  and (_05741_, _05737_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_05742_, _05741_, _05736_);
  nand (_05743_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_05744_, _05743_, _05740_);
  not (_05745_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nand (_05746_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_05747_, _05746_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  or (_05748_, _05747_, _05745_);
  not (_05749_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  or (_05750_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_05751_, _05750_, _05736_);
  or (_05752_, _05751_, _05749_);
  and (_05753_, _05752_, _05748_);
  not (_05754_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_05755_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_05756_, _05755_, _05736_);
  or (_05757_, _05756_, _05754_);
  and (_05758_, _05755_, _05736_);
  nand (_05759_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_05760_, _05759_, _05757_);
  and (_05761_, _05760_, _05753_);
  nand (_05762_, _05761_, _05744_);
  nand (_05763_, _05762_, _05734_);
  nand (_05764_, _05763_, _05733_);
  nor (_05765_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _05733_);
  not (_05766_, _05765_);
  and (_05767_, _05766_, _05764_);
  or (_05768_, _05767_, _05732_);
  not (_05769_, _05728_);
  nor (_05770_, _05730_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_05771_, _05770_, _05769_);
  and (_05772_, _05771_, _05768_);
  not (_05773_, _05772_);
  not (_05774_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  or (_05775_, _05747_, _05774_);
  nand (_05776_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_05777_, _05776_, _05775_);
  not (_05778_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  or (_05779_, _05756_, _05778_);
  nand (_05780_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_05781_, _05780_, _05779_);
  not (_05782_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  or (_05783_, _05751_, _05782_);
  not (_05784_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  or (_05785_, _05739_, _05784_);
  and (_05786_, _05785_, _05783_);
  and (_05787_, _05786_, _05781_);
  nand (_05788_, _05787_, _05777_);
  nand (_05789_, _05788_, _05734_);
  nand (_05790_, _05789_, _05733_);
  nor (_05791_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _05733_);
  not (_05792_, _05791_);
  and (_05793_, _05792_, _05790_);
  or (_05794_, _05793_, _05732_);
  nor (_05795_, _05730_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_05796_, _05795_, _05769_);
  nand (_05797_, _05796_, _05794_);
  and (_05798_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_05799_, _05798_);
  nand (_05800_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_05801_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_05802_, _05801_, _05800_);
  not (_05803_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  or (_05804_, _05756_, _05803_);
  not (_05805_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  or (_05806_, _05751_, _05805_);
  and (_05807_, _05806_, _05804_);
  not (_05808_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  or (_05810_, _05747_, _05808_);
  not (_05811_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  or (_05812_, _05739_, _05811_);
  and (_05813_, _05812_, _05810_);
  and (_05814_, _05813_, _05807_);
  and (_05815_, _05814_, _05802_);
  or (_05816_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_05817_, _05816_, _05815_);
  nand (_05818_, _05817_, _05799_);
  or (_05819_, _05818_, _05732_);
  nor (_05820_, _05730_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_05821_, _05820_, _05769_);
  nand (_05822_, _05821_, _05819_);
  and (_05823_, _05822_, _05797_);
  not (_05824_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  or (_05825_, _05751_, _05824_);
  not (_05826_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  or (_05827_, _05747_, _05826_);
  and (_05828_, _05827_, _05825_);
  not (_05829_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  or (_05830_, _05739_, _05829_);
  and (_05831_, _05830_, _05828_);
  nand (_05832_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_05833_, _05832_, _05734_);
  not (_05834_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  or (_05835_, _05756_, _05834_);
  nand (_05836_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_05837_, _05836_, _05835_);
  and (_05838_, _05837_, _05833_);
  nand (_05839_, _05838_, _05831_);
  or (_05840_, _05839_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_05841_, _05733_, \oc8051_top_1.oc8051_memory_interface1.cdata [1]);
  not (_05842_, _05841_);
  and (_05843_, _05842_, _05840_);
  or (_05844_, _05843_, _05732_);
  nor (_05845_, _05730_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_05846_, _05845_, _05769_);
  and (_05847_, _05846_, _05844_);
  and (_05848_, _05847_, _05823_);
  and (_05849_, _05848_, _05773_);
  not (_05850_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_05851_, _05751_, _05850_);
  not (_05852_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_05853_, _05747_, _05852_);
  and (_05854_, _05853_, _05851_);
  not (_05855_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  or (_05856_, _05739_, _05855_);
  and (_05857_, _05856_, _05854_);
  nand (_05858_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_05860_, _05858_, _05734_);
  not (_05861_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_05862_, _05756_, _05861_);
  nand (_05863_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_05864_, _05863_, _05862_);
  and (_05865_, _05864_, _05860_);
  nand (_05866_, _05865_, _05857_);
  or (_05867_, _05866_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_05868_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _05733_);
  not (_05869_, _05868_);
  and (_05870_, _05869_, _05867_);
  or (_05871_, _05870_, _05732_);
  nor (_05872_, _05730_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_05873_, _05872_, _05769_);
  and (_05874_, _05873_, _05871_);
  not (_05875_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  or (_05876_, _05739_, _05875_);
  nand (_05877_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_05878_, _05877_, _05876_);
  not (_05879_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  or (_05880_, _05747_, _05879_);
  not (_05881_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  or (_05882_, _05751_, _05881_);
  and (_05883_, _05882_, _05880_);
  not (_05884_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  or (_05885_, _05756_, _05884_);
  nand (_05886_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  and (_05888_, _05886_, _05885_);
  and (_05889_, _05888_, _05883_);
  nand (_05890_, _05889_, _05878_);
  and (_05891_, _05890_, _05734_);
  or (_05892_, _05891_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_05893_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _05733_);
  not (_05894_, _05893_);
  and (_05895_, _05894_, _05892_);
  or (_05896_, _05895_, _05732_);
  nor (_05897_, _05730_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_05898_, _05897_, _05769_);
  and (_05899_, _05898_, _05896_);
  not (_05900_, _05899_);
  nand (_05901_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_05902_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_05903_, _05902_, _05901_);
  not (_05904_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  or (_05905_, _05756_, _05904_);
  not (_05906_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  or (_05907_, _05747_, _05906_);
  and (_05908_, _05907_, _05905_);
  not (_05909_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  or (_05910_, _05751_, _05909_);
  not (_05911_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  or (_05912_, _05739_, _05911_);
  and (_05913_, _05912_, _05910_);
  and (_05914_, _05913_, _05908_);
  and (_05915_, _05914_, _05903_);
  or (_05916_, _05915_, _05816_);
  and (_05917_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.cdata [7]);
  not (_05918_, _05917_);
  nand (_05919_, _05918_, _05916_);
  or (_05920_, _05919_, _05732_);
  nor (_05921_, _05730_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_05922_, _05921_, _05769_);
  nand (_05923_, _05922_, _05920_);
  and (_05924_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_05925_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  or (_05926_, _05925_, _05924_);
  and (_05927_, _05750_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_05928_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_05929_, _05746_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_05930_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_05932_, _05930_, _05928_);
  and (_05933_, _05755_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_05934_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_05935_, _05738_, _05736_);
  and (_05936_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  or (_05937_, _05936_, _05934_);
  or (_05938_, _05937_, _05932_);
  or (_05939_, _05938_, _05926_);
  not (_05940_, _05939_);
  nor (_05941_, _05940_, _05816_);
  and (_05942_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  or (_05943_, _05942_, _05941_);
  or (_05944_, _05943_, _05732_);
  nor (_05945_, _05730_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_05946_, _05945_, _05769_);
  nand (_05947_, _05946_, _05944_);
  and (_05948_, _05947_, _05923_);
  and (_05949_, _05948_, _05900_);
  and (_05950_, _05949_, _05874_);
  and (_05951_, _05950_, _05849_);
  not (_05952_, _05847_);
  and (_05953_, _05772_, _05952_);
  and (_05954_, _05953_, _05823_);
  and (_05955_, _05954_, _05874_);
  or (_05956_, _05955_, _05951_);
  not (_05957_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_05958_, \oc8051_top_1.oc8051_decoder1.state [1], _04859_);
  and (_05959_, _05958_, _05957_);
  and (_05960_, _05959_, _05956_);
  or (_05961_, _05960_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_05962_, _05729_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_05963_, _05796_, _05794_);
  and (_05964_, _05847_, _05963_);
  and (_05965_, _05964_, _05822_);
  and (_05966_, _05965_, _05949_);
  and (_05967_, _05946_, _05944_);
  and (_05968_, _05967_, _05899_);
  and (_05969_, _05968_, _05874_);
  and (_05970_, _05969_, _05965_);
  or (_05971_, _05970_, _05966_);
  not (_05972_, _05874_);
  and (_05973_, _05822_, _05972_);
  and (_05974_, _05973_, _05964_);
  and (_05976_, _05922_, _05920_);
  and (_05977_, _05947_, _05976_);
  and (_05978_, _05977_, _05899_);
  and (_05979_, _05978_, _05974_);
  or (_05980_, _05979_, _05971_);
  nor (_05982_, _05772_, _05847_);
  and (_05983_, _05982_, _05823_);
  and (_05984_, _05967_, _05900_);
  and (_05985_, _05984_, _05976_);
  and (_05986_, _05985_, _05972_);
  and (_05987_, _05986_, _05983_);
  and (_05988_, _05985_, _05965_);
  or (_05989_, _05988_, _05987_);
  or (_05990_, _05989_, _05980_);
  or (_05991_, _05990_, _05956_);
  and (_05992_, _05991_, _05962_);
  not (_05993_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_05994_, \oc8051_top_1.oc8051_decoder1.state [0], _04859_);
  and (_05995_, _05994_, _05993_);
  and (_05996_, _05978_, _05972_);
  and (_05997_, _05822_, _05963_);
  and (_05998_, _05982_, _05997_);
  and (_05999_, _05998_, _05996_);
  and (_06000_, _05977_, _05900_);
  and (_06001_, _06000_, _05972_);
  and (_06002_, _06001_, _05998_);
  nor (_06003_, _06002_, _05999_);
  not (_06004_, _06003_);
  and (_06005_, _06004_, _05995_);
  or (_06006_, _06005_, _05992_);
  or (_06007_, _06006_, _05961_);
  or (_06008_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _04859_);
  and (_06009_, _06008_, _04856_);
  and (_04891_, _06009_, _06007_);
  nor (_06010_, _05282_, _05151_);
  not (_06011_, _06010_);
  and (_06012_, _05151_, _05059_);
  and (_06013_, _05207_, _05227_);
  nor (_06014_, _06013_, _06012_);
  or (_06015_, _06014_, _05126_);
  nand (_06016_, _06014_, _05126_);
  and (_06017_, _06016_, _05223_);
  nand (_06018_, _06017_, _06015_);
  not (_06019_, _05259_);
  or (_06020_, _05387_, _05378_);
  or (_06021_, _06020_, _06019_);
  or (_06022_, _05387_, _05256_);
  nand (_06023_, _05378_, _05267_);
  and (_06024_, _05377_, _05231_);
  and (_06025_, _05269_, _05151_);
  nor (_06026_, _06025_, _06024_);
  and (_06027_, _06026_, _06023_);
  and (_06028_, _06027_, _06022_);
  and (_06029_, _06028_, _06021_);
  and (_06030_, _06029_, _06018_);
  and (_06032_, _06030_, _06011_);
  not (_06033_, _06032_);
  and (_06034_, _06033_, _05009_);
  not (_06035_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  nor (_06036_, _05009_, _06035_);
  or (_06037_, _06036_, _06034_);
  and (_04983_, _06037_, _04856_);
  nand (_06038_, _05008_, _05678_);
  or (_06039_, _05003_, _05679_);
  and (_06040_, _06039_, _04861_);
  or (_06041_, _06040_, _06038_);
  and (_06042_, _06041_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  and (_06043_, _04992_, _04861_);
  and (_06044_, _06043_, _06033_);
  or (_06045_, _06044_, _06042_);
  and (_05235_, _06045_, _04856_);
  not (_06046_, _05675_);
  and (_06047_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_06048_, _06032_, _06046_);
  or (_06049_, _06048_, _05673_);
  or (_06050_, _06049_, _06047_);
  or (_06051_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_06052_, _06051_, _04856_);
  and (_06640_, _06052_, _06050_);
  and (_06053_, _05338_, _05459_);
  nor (_06054_, _05632_, _06053_);
  or (_06055_, _06054_, _05584_);
  nand (_06056_, _05434_, _05455_);
  nor (_06057_, _05572_, _05059_);
  nand (_06058_, _05572_, _05059_);
  nand (_06059_, _06058_, _05557_);
  or (_06060_, _06059_, _06057_);
  nor (_06061_, _05338_, _05490_);
  not (_06062_, _05052_);
  and (_06063_, _05055_, _06062_);
  and (_06064_, _05254_, _05218_);
  and (_06065_, _05267_, _06062_);
  nor (_06066_, _06065_, _06064_);
  nor (_06067_, _06066_, _06063_);
  nor (_06068_, _06067_, _06061_);
  and (_06069_, _05058_, _05052_);
  and (_06070_, _05259_, _05056_);
  nor (_06071_, _06070_, _05255_);
  nor (_06072_, _06071_, _06069_);
  not (_06073_, _06072_);
  and (_06074_, _05540_, _05206_);
  not (_06075_, _05269_);
  and (_06076_, _06075_, _05227_);
  and (_06077_, _05542_, _05052_);
  nor (_06078_, _06077_, _05273_);
  and (_06079_, _06078_, _05059_);
  nor (_06080_, _06079_, _06076_);
  nor (_06081_, _06080_, _06074_);
  and (_06082_, _06081_, _06073_);
  and (_06083_, _06082_, _06068_);
  and (_06084_, _06083_, _05561_);
  and (_06086_, _06084_, _06060_);
  and (_06087_, _06086_, _06056_);
  and (_06088_, _06087_, _06055_);
  not (_06089_, _05517_);
  not (_06090_, _04984_);
  and (_06091_, _04997_, _06090_);
  and (_06092_, _04860_, _04885_);
  and (_06093_, _06092_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not (_06094_, _06093_);
  nor (_06095_, _06094_, _04947_);
  nand (_06096_, _06095_, _06091_);
  nor (_06097_, _06096_, _06089_);
  nand (_06098_, _06097_, _06088_);
  not (_06099_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_06100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _06099_);
  not (_06101_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  not (_06102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_06103_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  not (_06104_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_06105_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _06104_);
  nor (_06106_, _06105_, _06103_);
  nor (_06107_, _06106_, _06102_);
  or (_06108_, _06107_, _06101_);
  and (_06109_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_06110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _06104_);
  nor (_06112_, _06110_, _06109_);
  nor (_06113_, _06112_, _06102_);
  and (_06114_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_06115_, _06104_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  or (_06116_, _06115_, _06114_);
  not (_06117_, _06116_);
  nand (_06118_, _06117_, _06113_);
  or (_06119_, _06118_, _06108_);
  and (_06120_, _06119_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_06121_, _06120_, _06100_);
  or (_06122_, _06121_, _06097_);
  and (_06123_, _06122_, _06098_);
  not (_06124_, _05510_);
  nor (_06125_, _06124_, _04947_);
  and (_06126_, _06125_, _04990_);
  and (_06127_, _06126_, _05517_);
  or (_06128_, _06127_, _06123_);
  not (_06129_, _06127_);
  or (_06130_, _06129_, _05718_);
  and (_06131_, _06130_, _04856_);
  and (_08562_, _06131_, _06128_);
  and (_06132_, _04932_, _04893_);
  not (_06133_, _04904_);
  and (_06134_, _06095_, _04922_);
  and (_06135_, _06134_, _06133_);
  and (_06136_, _06135_, _06132_);
  nand (_06137_, _06136_, _04958_);
  and (_06138_, _06137_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_06139_, _06138_, _06127_);
  and (_06140_, _04948_, _04922_);
  nor (_06141_, _06094_, _04904_);
  and (_06142_, _06141_, _06140_);
  and (_06143_, _06142_, _06132_);
  nand (_06144_, _06087_, _06055_);
  and (_06145_, _04996_, _04958_);
  and (_06146_, _06145_, _06090_);
  and (_06147_, _06146_, _06144_);
  and (_06148_, _04984_, _04958_);
  or (_06149_, _04989_, _06148_);
  and (_06150_, _06149_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_06151_, _06150_, _06147_);
  and (_06152_, _06151_, _06143_);
  or (_06153_, _06152_, _06139_);
  nand (_06154_, _06127_, _05287_);
  and (_06155_, _06154_, _04856_);
  and (_08584_, _06155_, _06153_);
  nand (_06156_, _06107_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and (_06157_, _06116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  or (_06159_, _06157_, _06113_);
  or (_06160_, _06159_, _06156_);
  nand (_06161_, _06160_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand (_06162_, _06161_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_06163_, _05517_, _04987_);
  and (_06164_, _06163_, _06093_);
  or (_06165_, _06164_, _06162_);
  and (_06166_, _06165_, _06129_);
  nand (_06168_, _06164_, _06088_);
  and (_06169_, _06168_, _06166_);
  nor (_06170_, _06129_, _06032_);
  or (_06171_, _06170_, _06169_);
  and (_08683_, _06171_, _04856_);
  and (_06172_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_06173_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _06104_);
  and (_06174_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_06175_, _06174_, _06173_);
  and (_06176_, _06175_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_06177_, _06176_, _06102_);
  and (_06178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_06179_, _06178_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_06180_, _06179_);
  and (_06181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_06182_, _06181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_06183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_06184_, _06183_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_06185_, _06184_, _06182_);
  and (_06186_, _06185_, _06180_);
  not (_06187_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_06188_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nor (_06189_, _06188_, _06187_);
  nand (_06190_, _06189_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  not (_06191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_06192_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_06193_, _06192_, _06191_);
  and (_06194_, _06193_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_06195_, _06194_);
  and (_06196_, _06195_, _06190_);
  and (_06197_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_06198_, _06197_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_06199_, _06198_);
  and (_06200_, _06199_, _06196_);
  and (_06201_, _06200_, _06186_);
  nor (_06202_, _06201_, _06177_);
  and (_06203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _06102_);
  not (_06204_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_06205_, _06178_, _06204_);
  not (_06206_, _06205_);
  not (_06207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_06208_, _06181_, _06207_);
  not (_06209_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_06210_, _06183_, _06209_);
  nor (_06211_, _06210_, _06208_);
  and (_06212_, _06211_, _06206_);
  not (_06213_, _06212_);
  and (_06214_, _06213_, _06203_);
  not (_06215_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_06216_, _06189_, _06215_);
  not (_06217_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_06218_, _06193_, _06217_);
  nor (_06219_, _06218_, _06216_);
  not (_06220_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_06221_, _06197_, _06220_);
  not (_06222_, _06221_);
  nand (_06223_, _06222_, _06219_);
  and (_06224_, _06223_, _06203_);
  or (_06225_, _06224_, _06214_);
  nor (_06226_, _06225_, _06202_);
  and (_06227_, _06226_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  not (_06228_, _06202_);
  nor (_06229_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _06104_);
  and (_06230_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _06104_);
  nor (_06231_, _06230_, _06229_);
  nor (_06232_, _06231_, _06228_);
  or (_06233_, _06232_, _06227_);
  or (_06234_, _06233_, _06172_);
  not (_06235_, _06172_);
  or (_06236_, _06231_, _06235_);
  and (_06237_, _06236_, _04856_);
  and (_09163_, _06237_, _06234_);
  and (_06238_, _05731_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_06240_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_06241_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_06242_, _06238_, _06241_);
  or (_06243_, _06242_, _06240_);
  and (_09192_, _06243_, _04856_);
  nand (_06244_, _06228_, _06214_);
  or (_06245_, _06186_, _06177_);
  and (_06246_, _06245_, _06235_);
  and (_06248_, _06246_, _06244_);
  nor (_06249_, _06172_, _06104_);
  nor (_06250_, _06235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  nor (_06251_, _06250_, _06249_);
  or (_06252_, _06251_, _06248_);
  or (_06253_, _06224_, _06202_);
  not (_06254_, _06200_);
  or (_06255_, _06245_, _06254_);
  and (_06256_, _06255_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_06257_, _06256_, _06253_);
  or (_06258_, _06257_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_06259_, _06258_, _04856_);
  and (_09318_, _06259_, _06252_);
  and (_06260_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_06261_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_06262_, _06238_, _06261_);
  or (_06263_, _06262_, _06260_);
  and (_09528_, _06263_, _04856_);
  nand (_06264_, _06201_, _06102_);
  or (_06265_, _06264_, _06225_);
  nand (_06266_, _06229_, _06172_);
  and (_06267_, _06266_, _04856_);
  and (_10162_, _06267_, _06265_);
  and (_06268_, _05519_, _06090_);
  and (_06269_, _04933_, _04893_);
  and (_06270_, _06269_, _06142_);
  and (_06271_, _06270_, _06268_);
  or (_06272_, _06271_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_06273_, _04933_, _04922_);
  and (_06274_, _06273_, _05515_);
  and (_06275_, _06274_, _06126_);
  not (_06276_, _06275_);
  and (_06277_, _06276_, _06272_);
  nand (_06278_, _06271_, _06088_);
  and (_06279_, _06278_, _06277_);
  nor (_06280_, _05338_, _05282_);
  not (_06281_, _06280_);
  and (_06282_, _06281_, _05556_);
  and (_06283_, _06282_, _05551_);
  and (_06284_, _06283_, _05538_);
  nor (_06285_, _06284_, _06276_);
  or (_06286_, _06285_, _06279_);
  and (_10217_, _06286_, _04856_);
  not (_06287_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_06288_, _06172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_06289_, _06288_, _06287_);
  or (_06290_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _06104_);
  or (_06291_, _06253_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_06292_, _06291_, _06290_);
  and (_06293_, _06292_, _06248_);
  or (_06294_, _06293_, _06289_);
  and (_10318_, _06294_, _04856_);
  nor (_06295_, _04947_, _04922_);
  and (_06296_, _06295_, _06141_);
  and (_06297_, _06296_, _06269_);
  and (_06298_, _06297_, _06268_);
  nand (_06299_, _06298_, _06088_);
  or (_06300_, _06298_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_06301_, _06268_, _05512_);
  nor (_06302_, _04932_, _04922_);
  and (_06303_, _06302_, _05515_);
  and (_06304_, _06303_, _06301_);
  not (_06305_, _06304_);
  and (_06306_, _06305_, _06300_);
  and (_06307_, _06306_, _06299_);
  nor (_06308_, _06305_, _06284_);
  or (_06309_, _06308_, _06307_);
  and (_10339_, _06309_, _04856_);
  and (_06310_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _04856_);
  and (_10459_, _06310_, _06172_);
  and (_06311_, _06268_, _06095_);
  and (_06312_, _06311_, _05517_);
  nand (_06313_, _06312_, _06088_);
  nor (_06314_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_06316_, _06314_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  nand (_06317_, _06157_, _06112_);
  or (_06318_, _06317_, _06108_);
  and (_06319_, _06318_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_06320_, _06319_, _06316_);
  or (_06321_, _06320_, _06312_);
  and (_06322_, _06321_, _06129_);
  and (_06323_, _06322_, _06313_);
  nor (_06324_, _06284_, _06129_);
  or (_06325_, _06324_, _06323_);
  and (_10480_, _06325_, _04856_);
  and (_10675_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _04856_);
  and (_06326_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  or (_06327_, _06156_, _06118_);
  and (_06328_, _06327_, _06326_);
  and (_06329_, _05520_, _04948_);
  and (_06330_, _06329_, _05517_);
  and (_06331_, _06330_, _06093_);
  or (_06332_, _06331_, _06328_);
  and (_06333_, _06332_, _06129_);
  nand (_06334_, _06331_, _06088_);
  and (_06335_, _06334_, _06333_);
  nor (_06336_, _06129_, _05669_);
  or (_06337_, _06336_, _06335_);
  and (_10816_, _06337_, _04856_);
  and (_06338_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  or (_06339_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nand (_06340_, _06339_, _04856_);
  nor (_11292_, _06340_, _06338_);
  nor (_11844_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  or (_06341_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not (_06342_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_06343_, _06238_, _06342_);
  and (_06344_, _06343_, _04856_);
  and (_12295_, _06344_, _06341_);
  not (_06345_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_06346_, _06338_, _06345_);
  and (_06347_, _06346_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor (_06348_, _06338_, _06345_);
  or (_06349_, _06348_, _06346_);
  nand (_06350_, _06349_, _04856_);
  nor (_12580_, _06350_, _06347_);
  or (_06351_, _04992_, _05003_);
  and (_06352_, _06351_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_06353_, _06352_, _04861_);
  or (_06354_, _05007_, _04995_);
  and (_06355_, _06354_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  or (_06356_, _05385_, _06019_);
  and (_06357_, _06356_, _05256_);
  or (_06358_, _06357_, _05396_);
  nand (_06359_, _05385_, _05267_);
  or (_06360_, _06075_, _05206_);
  and (_06361_, _06360_, _06359_);
  or (_06362_, _05383_, _05232_);
  not (_06363_, _05223_);
  or (_06364_, _06363_, _05206_);
  and (_06365_, _06364_, _06362_);
  or (_06366_, _05282_, _05126_);
  and (_06367_, _06366_, _06365_);
  and (_06368_, _06367_, _06361_);
  and (_06369_, _06368_, _06358_);
  nor (_06370_, _06369_, _05673_);
  and (_06371_, _06370_, _04988_);
  or (_06372_, _06371_, _06355_);
  or (_06373_, _06372_, _06353_);
  and (_13213_, _06373_, _04856_);
  and (_06374_, _06354_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_06375_, _05718_, _04988_);
  and (_06376_, _06351_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  or (_06377_, _06376_, _06375_);
  and (_06378_, _06377_, _04861_);
  or (_06379_, _06378_, _06374_);
  and (_01164_, _06379_, _04856_);
  and (_06380_, _06038_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_06381_, _06370_, _04992_);
  and (_06382_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_06383_, _06382_, _06039_);
  or (_06384_, _06383_, _06381_);
  or (_06385_, _06384_, _06380_);
  and (_01432_, _06385_, _04856_);
  nand (_06386_, _05721_, _05008_);
  and (_06387_, _06386_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nor (_06388_, _05282_, _05081_);
  not (_06389_, _06388_);
  not (_06390_, _05693_);
  nand (_06391_, _05175_, _05059_);
  nand (_06392_, _06391_, _06390_);
  nand (_06393_, _06392_, _05565_);
  or (_06395_, _06392_, _05565_);
  and (_06396_, _06395_, _05223_);
  nand (_06397_, _06396_, _06393_);
  nand (_06398_, _05349_, _05259_);
  and (_06399_, _05347_, _05267_);
  and (_06400_, _05269_, _05081_);
  nor (_06401_, _06400_, _06399_);
  and (_06402_, _05346_, _05059_);
  nor (_06403_, _06402_, _05232_);
  and (_06404_, _06403_, _05692_);
  nor (_06405_, _05348_, _05256_);
  nor (_06406_, _06405_, _06404_);
  and (_06407_, _06406_, _06401_);
  and (_06408_, _06407_, _06398_);
  and (_06409_, _06408_, _06397_);
  nand (_06410_, _06409_, _06389_);
  and (_06411_, _06410_, _06043_);
  or (_06412_, _06411_, _06387_);
  and (_01517_, _06412_, _04856_);
  and (_06413_, _06354_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_06414_, _06410_, _04988_);
  and (_06415_, _06351_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or (_06416_, _06415_, _06414_);
  and (_06417_, _06416_, _04861_);
  or (_06418_, _06417_, _06413_);
  and (_01547_, _06418_, _04856_);
  and (_06419_, _05719_, _05670_);
  and (_06420_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  or (_06421_, _06420_, _06419_);
  and (_01669_, _06421_, _04856_);
  and (_06422_, _06041_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_06423_, _06043_, _05670_);
  or (_06424_, _06423_, _06422_);
  and (_01710_, _06424_, _04856_);
  and (_06425_, _06041_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_06426_, _06043_, _05288_);
  or (_06427_, _06426_, _06425_);
  and (_01955_, _06427_, _04856_);
  nand (_06428_, _05452_, _05303_);
  and (_06429_, _06428_, _05453_);
  nand (_06430_, _06429_, _05455_);
  and (_06431_, _05483_, _05243_);
  not (_06432_, _06431_);
  nor (_06433_, _05483_, _05243_);
  nor (_06434_, _06433_, _06363_);
  and (_06435_, _06434_, _06432_);
  nor (_06436_, _05531_, _05460_);
  nor (_06437_, _06436_, _05232_);
  not (_06438_, _06437_);
  nor (_06439_, _05490_, _05172_);
  not (_06440_, _06439_);
  nor (_06441_, _05274_, _05243_);
  and (_06442_, _05497_, ABINPUT000000[15]);
  and (_06443_, _05499_, ABINPUT000[15]);
  nor (_06444_, _06443_, _06442_);
  not (_06445_, _06444_);
  nor (_06446_, _06445_, _06441_);
  and (_06448_, _06446_, _06440_);
  and (_06449_, _06448_, _06438_);
  not (_06450_, _06449_);
  nor (_06451_, _06450_, _06435_);
  nand (_06452_, _06451_, _06430_);
  or (_06453_, _06452_, _05293_);
  not (_06454_, _05455_);
  and (_06455_, _05428_, _05422_);
  nor (_06456_, _06455_, _06454_);
  and (_06457_, _06456_, _05429_);
  not (_06458_, _06457_);
  nor (_06459_, _05629_, _05597_);
  nor (_06460_, _06459_, _05630_);
  nor (_06461_, _06460_, _05584_);
  and (_06462_, _05568_, _05199_);
  nor (_06463_, _06462_, _05048_);
  nor (_06464_, _06463_, _05569_);
  nor (_06466_, _06464_, _05558_);
  not (_06468_, _05279_);
  or (_06469_, _05338_, _06468_);
  and (_06470_, _05499_, ABINPUT000[7]);
  not (_06471_, _06470_);
  and (_06473_, _06471_, _06469_);
  and (_06474_, _05280_, _05587_);
  nor (_06475_, _05274_, _05048_);
  and (_06476_, _05497_, ABINPUT000000[7]);
  or (_06477_, _06476_, _06475_);
  nor (_06478_, _06477_, _06474_);
  and (_06479_, _06478_, _05271_);
  and (_06480_, _06479_, _06473_);
  and (_06481_, _06480_, _05263_);
  not (_06482_, _06481_);
  nor (_06483_, _06482_, _06466_);
  and (_06485_, _06483_, _05247_);
  not (_06486_, _06485_);
  nor (_06487_, _06486_, _06461_);
  and (_06488_, _06487_, _06458_);
  nor (_06489_, _06488_, _05643_);
  and (_06490_, _05643_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_06491_, _06490_, _05292_);
  or (_06492_, _06491_, _06489_);
  and (_06493_, _06492_, _04856_);
  and (_02380_, _06493_, _06453_);
  and (_06494_, _06145_, _04984_);
  and (_06495_, _06494_, _05512_);
  and (_06496_, _06495_, _05517_);
  nor (_06497_, _06496_, _05292_);
  not (_06498_, _06497_);
  nand (_06499_, _06498_, _06488_);
  or (_06500_, _06498_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_06501_, _06500_, _04856_);
  and (_02512_, _06501_, _06499_);
  nor (_06502_, _05401_, _05399_);
  not (_06503_, _06502_);
  nor (_06504_, _05402_, _06454_);
  and (_06505_, _06504_, _06503_);
  not (_06506_, _06505_);
  nor (_06507_, _05619_, _05614_);
  nor (_06508_, _06507_, _05620_);
  nor (_06509_, _06508_, _05584_);
  not (_06510_, _06509_);
  and (_06511_, _05173_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_06512_, _05559_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_06513_, _06512_, _05207_);
  nor (_06514_, _06513_, _05172_);
  nor (_06515_, _06514_, _06511_);
  nor (_06516_, _06515_, _05558_);
  nor (_06517_, _05371_, _05256_);
  and (_06518_, _05372_, _05259_);
  or (_06519_, _06518_, _06517_);
  not (_06520_, _06519_);
  and (_06521_, _05280_, _05207_);
  and (_06522_, _05497_, ABINPUT000000[3]);
  and (_06523_, _05499_, ABINPUT000[3]);
  nor (_06524_, _06523_, _06522_);
  not (_06525_, _06524_);
  nor (_06526_, _06525_, _06521_);
  or (_06527_, _06468_, _05103_);
  nor (_06528_, _05274_, _05172_);
  not (_06529_, _06528_);
  and (_06530_, _06529_, _06527_);
  and (_06531_, _06530_, _06526_);
  and (_06532_, _06531_, _06520_);
  not (_06533_, _06532_);
  nor (_06534_, _06533_, _06516_);
  not (_06535_, _06534_);
  or (_06536_, _06012_, _05206_);
  or (_06537_, _06013_, _05126_);
  nand (_06538_, _06537_, _06536_);
  or (_06539_, _06538_, _05172_);
  nand (_06540_, _06538_, _05172_);
  and (_06541_, _06540_, _05223_);
  and (_06542_, _06541_, _06539_);
  nor (_06543_, _05368_, _05232_);
  or (_06544_, _06543_, _06542_);
  not (_06545_, _06544_);
  and (_06546_, _05369_, _05267_);
  and (_06547_, _05269_, _05172_);
  nor (_06548_, _06547_, _06546_);
  nand (_06549_, _06548_, _06545_);
  nor (_06550_, _06549_, _06535_);
  and (_06551_, _06550_, _06510_);
  and (_06552_, _06551_, _06506_);
  nand (_06553_, _06552_, _06498_);
  or (_06554_, _06498_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_06555_, _06554_, _04856_);
  and (_02954_, _06555_, _06553_);
  nor (_06556_, _05402_, _05395_);
  or (_06557_, _06556_, _06454_);
  nor (_06558_, _06557_, _05403_);
  not (_06559_, _06558_);
  nor (_06560_, _05620_, _05612_);
  nor (_06561_, _06560_, _05621_);
  nor (_06562_, _06561_, _05584_);
  not (_06563_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_06564_, _05173_, _06563_);
  nor (_06565_, _06564_, _05204_);
  or (_06566_, _06565_, _05558_);
  nor (_06567_, _06566_, _05559_);
  and (_06568_, _05280_, _05205_);
  and (_06569_, _05497_, ABINPUT000000[4]);
  and (_06570_, _05499_, ABINPUT000[4]);
  nor (_06571_, _06570_, _06569_);
  not (_06572_, _06571_);
  nor (_06573_, _06572_, _06568_);
  nor (_06574_, _05274_, _05103_);
  not (_06575_, _06574_);
  or (_06576_, _06468_, _05081_);
  and (_06578_, _06576_, _06575_);
  and (_06579_, _06578_, _06573_);
  not (_06580_, _06579_);
  nor (_06581_, _06580_, _06567_);
  and (_06582_, _06581_, _05667_);
  and (_06583_, _06582_, _05656_);
  not (_06584_, _06583_);
  nor (_06585_, _06584_, _06562_);
  and (_06586_, _06585_, _06559_);
  nand (_06587_, _06586_, _06498_);
  not (_06588_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  nand (_06589_, _06497_, _06588_);
  and (_06590_, _06589_, _04856_);
  and (_03036_, _06590_, _06587_);
  and (_06591_, _05683_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_06592_, _05671_, _05288_);
  or (_06593_, _06592_, _06591_);
  and (_03190_, _06593_, _04856_);
  and (_06594_, _05985_, _05874_);
  and (_06595_, _06594_, _05849_);
  and (_06596_, _05968_, _05923_);
  and (_06597_, _06596_, _05972_);
  and (_06598_, _05848_, _05772_);
  and (_06599_, _06598_, _06597_);
  and (_06600_, _06597_, _05849_);
  or (_06601_, _06600_, _06599_);
  nor (_06602_, _06601_, _06595_);
  and (_06603_, _05985_, _05983_);
  nor (_06604_, _06603_, _05951_);
  nand (_06605_, _06604_, _06602_);
  and (_06606_, _05997_, _05953_);
  and (_06607_, _06606_, _05969_);
  and (_06608_, _05949_, _05972_);
  and (_06609_, _06606_, _06608_);
  and (_06610_, _06594_, _06606_);
  or (_06611_, _06610_, _06609_);
  and (_06612_, _05978_, _05874_);
  and (_06613_, _06612_, _05849_);
  and (_06614_, _05986_, _05849_);
  nor (_06615_, _06614_, _06613_);
  not (_06616_, _06615_);
  or (_06617_, _06616_, _06611_);
  or (_06618_, _06617_, _06607_);
  and (_06619_, _05984_, _05923_);
  and (_06620_, _06619_, _05972_);
  and (_06621_, _06598_, _06620_);
  and (_06622_, _06620_, _05849_);
  or (_06623_, _06622_, _06621_);
  and (_06624_, _06000_, _05874_);
  and (_06625_, _06624_, _05849_);
  and (_06626_, _06606_, _06001_);
  or (_06627_, _06626_, _06625_);
  and (_06628_, _06606_, _05986_);
  and (_06629_, _06606_, _05950_);
  or (_06630_, _06629_, _06628_);
  or (_06631_, _06630_, _06627_);
  or (_06632_, _06631_, _06623_);
  or (_06633_, _06632_, _06618_);
  or (_06634_, _06633_, _06605_);
  and (_06635_, _06619_, _05874_);
  and (_06636_, _06635_, _05848_);
  not (_06637_, _05822_);
  or (_06638_, _05964_, _06637_);
  and (_06639_, _06638_, _06001_);
  or (_06641_, _06639_, _06636_);
  or (_06642_, _06641_, _05955_);
  or (_06643_, _06642_, _06634_);
  and (_06644_, _06643_, _05730_);
  and (_06645_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_06646_, _06005_, _05960_);
  not (_06647_, _05959_);
  nand (_06648_, _05983_, _05950_);
  nor (_06649_, _06648_, _06647_);
  or (_06650_, _06649_, _06646_);
  or (_06651_, _06650_, _06645_);
  or (_06652_, _06651_, _06644_);
  and (_03594_, _06652_, _04856_);
  not (_06653_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_06654_, _05291_, _06653_);
  and (_06655_, _06654_, _05507_);
  not (_06656_, _06654_);
  and (_06657_, _06268_, _06144_);
  nor (_06658_, _06268_, _05332_);
  or (_06659_, _06658_, _06657_);
  nor (_06660_, _06653_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_06661_, _06660_, _04859_);
  nor (_06662_, _04904_, _04893_);
  and (_06663_, _06662_, _06273_);
  and (_06664_, _06663_, _05001_);
  and (_06665_, _06664_, _05510_);
  nor (_06666_, _06665_, _06661_);
  and (_06667_, _06666_, _06656_);
  nor (_06668_, _04948_, _04904_);
  and (_06669_, _06668_, _04922_);
  nor (_06670_, _04932_, _04893_);
  and (_06671_, _06670_, _06093_);
  and (_06672_, _06671_, _06669_);
  and (_06673_, _06672_, _06667_);
  nand (_06674_, _06673_, _06659_);
  not (_06675_, _06666_);
  and (_06676_, _06675_, _05641_);
  not (_06677_, _06672_);
  and (_06678_, _06677_, _06667_);
  and (_06679_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_06680_, _06679_, _06676_);
  nand (_06681_, _06680_, _06674_);
  and (_06682_, _06681_, _06656_);
  or (_06684_, _06682_, _06655_);
  and (_04014_, _06684_, _04856_);
  not (_06685_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_06686_, _05679_, _04861_);
  nor (_06687_, _06686_, _06685_);
  not (_06688_, _06686_);
  nor (_06689_, _06688_, _05287_);
  or (_06690_, _06689_, _06687_);
  and (_04065_, _06690_, _04856_);
  or (_06691_, _06497_, _05641_);
  or (_06692_, _06498_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_06693_, _06692_, _04856_);
  and (_04848_, _06693_, _06691_);
  and (_06694_, _06033_, _05671_);
  and (_06695_, _04995_, _04861_);
  or (_06696_, _06695_, _05682_);
  and (_06697_, _06696_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  or (_06698_, _06697_, _06694_);
  and (_04849_, _06698_, _04856_);
  or (_06699_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_06700_, _06238_, _05185_);
  and (_06701_, _06700_, _04856_);
  and (_04851_, _06701_, _06699_);
  and (_06702_, _06386_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor (_06703_, _05282_, _05172_);
  or (_06704_, _06703_, _06519_);
  or (_06705_, _06704_, _06549_);
  and (_06706_, _06705_, _06043_);
  or (_06707_, _06706_, _06702_);
  and (_04853_, _06707_, _04856_);
  not (_06708_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_06709_, _05675_, _06708_);
  and (_06710_, _06705_, _05675_);
  or (_06711_, _06710_, _06709_);
  or (_06712_, _06711_, _05673_);
  or (_06713_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_06714_, _06713_, _04856_);
  and (_04854_, _06714_, _06712_);
  and (_06715_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_06716_, _06705_, _05719_);
  or (_06717_, _06716_, _06715_);
  and (_04855_, _06717_, _04856_);
  and (_06718_, _06033_, _05719_);
  and (_06719_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  or (_06720_, _06719_, _06718_);
  and (_04970_, _06720_, _04856_);
  and (_06721_, _04856_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06722_, _06721_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_06723_, _05998_, _06608_);
  or (_06724_, _06723_, _06611_);
  and (_06725_, _05998_, _05950_);
  or (_06726_, _06725_, _06629_);
  or (_06727_, _06726_, _06724_);
  nand (_06728_, _06612_, _05983_);
  not (_06729_, _06728_);
  or (_06730_, _05847_, _06637_);
  nor (_06731_, _06730_, _05797_);
  and (_06732_, _06620_, _06731_);
  and (_06733_, _06732_, _05772_);
  or (_06734_, _06733_, _06729_);
  and (_06735_, _06732_, _05773_);
  and (_06736_, _06620_, _05848_);
  and (_06737_, _05969_, _05923_);
  and (_06738_, _06737_, _05849_);
  or (_06739_, _06738_, _06736_);
  or (_06740_, _06739_, _06735_);
  or (_06741_, _06740_, _06734_);
  or (_06742_, _06741_, _06727_);
  nor (_06743_, _05822_, _05874_);
  and (_06744_, _06743_, _05949_);
  or (_06745_, _06594_, _05950_);
  and (_06746_, _06745_, _06637_);
  or (_06747_, _06746_, _06744_);
  nor (_06748_, _06601_, _05966_);
  not (_06749_, _06748_);
  and (_06750_, _06743_, _06596_);
  and (_06751_, _06598_, _05948_);
  or (_06752_, _06751_, _06750_);
  or (_06753_, _06752_, _06749_);
  or (_06754_, _06753_, _06747_);
  and (_06755_, _06597_, _05965_);
  and (_06756_, _06620_, _05965_);
  or (_06757_, _06756_, _06755_);
  or (_06758_, _06757_, _05988_);
  and (_06759_, _05998_, _05986_);
  or (_06760_, _06759_, _06628_);
  and (_06761_, _06597_, _06731_);
  and (_06762_, _05983_, _05996_);
  and (_06763_, _06743_, _05984_);
  or (_06764_, _06763_, _06762_);
  or (_06765_, _06764_, _06761_);
  or (_06766_, _06765_, _06760_);
  or (_06767_, _06766_, _06758_);
  or (_06768_, _06767_, _06754_);
  or (_06769_, _06768_, _06742_);
  and (_06770_, _05730_, _04856_);
  and (_06771_, _06770_, _06769_);
  or (_05113_, _06771_, _06722_);
  and (_06772_, _05968_, _05976_);
  and (_06773_, _06772_, _05874_);
  nand (_06774_, _06773_, _05848_);
  nand (_06775_, _06773_, _05983_);
  and (_06776_, _06775_, _06774_);
  and (_06777_, _06772_, _05972_);
  and (_06778_, _06777_, _05983_);
  and (_06779_, _06777_, _05848_);
  nor (_06780_, _06779_, _06778_);
  and (_06781_, _06780_, _06776_);
  not (_06782_, _06770_);
  and (_06783_, _06598_, _06000_);
  or (_06784_, _06783_, _06782_);
  or (_05116_, _06784_, _06781_);
  and (_06786_, _06598_, _05996_);
  and (_06787_, _06624_, _05983_);
  or (_06788_, _06787_, _06786_);
  and (_06789_, _06763_, _05976_);
  or (_06790_, _06789_, _05988_);
  or (_06791_, _06790_, _06760_);
  or (_06792_, _06791_, _06788_);
  and (_06793_, _06792_, _05730_);
  and (_06794_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_06795_, _06794_, _06005_);
  or (_06796_, _06795_, _06793_);
  and (_05127_, _06796_, _04856_);
  and (_06797_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_06798_, _06797_);
  not (_06799_, _05962_);
  or (_06800_, _06737_, _06624_);
  and (_06801_, _06800_, _06598_);
  nor (_06802_, _06801_, _06786_);
  and (_06803_, _06802_, _06003_);
  nor (_06804_, _06803_, _06799_);
  not (_06805_, _06804_);
  and (_06806_, _05983_, _06596_);
  and (_06807_, _06806_, _05959_);
  and (_06808_, _06619_, _05983_);
  and (_06809_, _06808_, _05959_);
  nor (_06810_, _06809_, _06807_);
  not (_06811_, _06810_);
  not (_06812_, _05729_);
  nor (_06813_, _06003_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06814_, _06813_, _06812_);
  nor (_06815_, _06814_, _06811_);
  nand (_06816_, _06815_, _06805_);
  nand (_06817_, _06816_, _04859_);
  and (_06818_, _06817_, _06798_);
  not (_06819_, _06818_);
  and (_06820_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_06821_, _06820_);
  and (_06822_, _05948_, _05899_);
  and (_06823_, _06822_, _05849_);
  not (_06824_, _06823_);
  nand (_06825_, _06001_, _05965_);
  and (_06826_, _06825_, _06824_);
  nand (_06827_, _06594_, _05983_);
  nand (_06828_, _06777_, _05965_);
  and (_06829_, _06828_, _06827_);
  and (_06830_, _06829_, _06826_);
  and (_06831_, _05965_, _05874_);
  and (_06832_, _06619_, _06831_);
  and (_06833_, _06822_, _05965_);
  or (_06834_, _06833_, _06832_);
  and (_06835_, _06000_, _06831_);
  and (_06836_, _06612_, _05965_);
  nor (_06837_, _06836_, _05966_);
  not (_06838_, _06837_);
  or (_06839_, _06838_, _06835_);
  nor (_06840_, _06839_, _06834_);
  and (_06841_, _06840_, _06830_);
  not (_06842_, _06802_);
  nor (_06843_, _06842_, _06758_);
  nand (_06844_, _06843_, _06841_);
  nand (_06845_, _06844_, _05962_);
  and (_06846_, _05994_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_06847_, _06823_, _06846_);
  nor (_06848_, _06847_, _06807_);
  nand (_06849_, _06848_, _06845_);
  nand (_06850_, _06849_, _04859_);
  nand (_06851_, _06850_, _06821_);
  and (_06852_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_06853_, _06852_);
  and (_06854_, _06822_, _05972_);
  nand (_06855_, _06854_, _05983_);
  not (_06856_, _06855_);
  and (_06857_, _06822_, _05874_);
  nand (_06858_, _06857_, _05983_);
  nand (_06859_, _06858_, _06648_);
  nor (_06860_, _06859_, _06856_);
  and (_06861_, _06612_, _06606_);
  and (_06862_, _06624_, _06606_);
  nor (_06863_, _06862_, _06861_);
  and (_06864_, _06863_, _06860_);
  and (_06865_, _06001_, _05849_);
  or (_06866_, _06865_, _06636_);
  nand (_06867_, _06635_, _06606_);
  nand (_06868_, _06822_, _06606_);
  nand (_06869_, _06868_, _06867_);
  nor (_06870_, _06869_, _06866_);
  and (_06871_, _06777_, _06606_);
  and (_06872_, _05996_, _05849_);
  nor (_06873_, _06872_, _06871_);
  and (_06875_, _06873_, _06870_);
  and (_06876_, _06875_, _06864_);
  nor (_06877_, _06609_, _05979_);
  or (_06878_, _06762_, _06738_);
  nor (_06879_, _06878_, _06623_);
  nand (_06880_, _06620_, _06606_);
  and (_06882_, _06880_, _06728_);
  nor (_06883_, _06610_, _06629_);
  and (_06885_, _06883_, _06615_);
  and (_06886_, _06885_, _06882_);
  and (_06887_, _06886_, _06879_);
  and (_06888_, _06597_, _06606_);
  or (_06889_, _06888_, _06628_);
  nor (_06890_, _06889_, _06603_);
  and (_06891_, _06890_, _06824_);
  and (_06892_, _06743_, _05978_);
  nor (_06893_, _06892_, _06627_);
  and (_06894_, _06893_, _06602_);
  and (_06895_, _06894_, _06891_);
  and (_06897_, _06895_, _06887_);
  and (_06898_, _06897_, _06877_);
  nand (_06899_, _06898_, _06876_);
  nand (_06900_, _06899_, _05962_);
  not (_06901_, _06847_);
  and (_06902_, _06901_, _06810_);
  nand (_06903_, _06902_, _06900_);
  nand (_06904_, _06903_, _04859_);
  and (_06905_, _06904_, _06853_);
  or (_06906_, _06905_, _06851_);
  or (_06907_, _06906_, _06819_);
  nor (_06908_, _05730_, _05104_);
  and (_06910_, _05730_, _05734_);
  not (_06911_, _06910_);
  and (_06912_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_06913_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_06915_, _06913_, _06912_);
  and (_06916_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_06917_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_06918_, _06917_, _06916_);
  and (_06919_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_06920_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_06921_, _06920_, _06919_);
  and (_06922_, _06921_, _06918_);
  and (_06923_, _06922_, _06915_);
  nor (_06924_, _06923_, _06911_);
  nor (_06925_, _06924_, _06908_);
  or (_06926_, _06925_, _06907_);
  and (_06928_, _06905_, _06851_);
  and (_06929_, _06928_, _06818_);
  not (_06930_, _04922_);
  and (_06931_, _05510_, _05001_);
  and (_06932_, _06931_, _04934_);
  and (_06934_, _06932_, _06662_);
  not (_06935_, _06934_);
  and (_06936_, _06935_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_06937_, _06934_, _06410_);
  nor (_06938_, _06937_, _06936_);
  nor (_06940_, _06938_, _06930_);
  and (_06941_, _06938_, _06930_);
  nor (_06943_, _06941_, _06940_);
  and (_06944_, _06935_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_06946_, _06935_, _05669_);
  nor (_06947_, _06946_, _06944_);
  and (_06948_, _06947_, _04948_);
  or (_06949_, _06947_, _04948_);
  nor (_06950_, _05772_, _04958_);
  and (_06951_, _05772_, _04958_);
  or (_06952_, _06951_, _05007_);
  nor (_06953_, _06952_, _06950_);
  nand (_06955_, _06953_, _06949_);
  nor (_06956_, _06955_, _06948_);
  and (_06957_, _06956_, _06943_);
  and (_06958_, _06957_, _06369_);
  not (_06959_, _06938_);
  nor (_06960_, _06947_, _05773_);
  and (_06961_, _06960_, _06959_);
  and (_06962_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_06963_, _06947_, _05773_);
  and (_06964_, _06963_, _06938_);
  and (_06965_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  nor (_06966_, _06965_, _06962_);
  nor (_06967_, _06947_, _05772_);
  and (_06968_, _06967_, _06959_);
  and (_06969_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_06970_, _06960_, _06938_);
  and (_06971_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_06972_, _06971_, _06969_);
  and (_06973_, _06972_, _06966_);
  not (_06974_, _06957_);
  and (_06976_, _06963_, _06959_);
  nand (_06977_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_06978_, _06947_, _05772_);
  and (_06979_, _06978_, _06938_);
  nand (_06980_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  and (_06981_, _06980_, _06977_);
  not (_06982_, _06978_);
  nor (_06983_, _06982_, _06938_);
  nand (_06984_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_06985_, _06967_, _06938_);
  nand (_06986_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_06987_, _06986_, _06984_);
  and (_06988_, _06987_, _06981_);
  and (_06989_, _06988_, _06974_);
  and (_06990_, _06989_, _06973_);
  nor (_06991_, _06990_, _06958_);
  nand (_06992_, _06991_, _06929_);
  and (_06993_, _06992_, _06926_);
  nand (_06994_, _06904_, _06853_);
  and (_06995_, _06994_, _06851_);
  nand (_06996_, _06995_, _06818_);
  not (_06997_, _06369_);
  and (_06998_, _05510_, _04999_);
  and (_06999_, _06998_, _05517_);
  nand (_07000_, _06999_, _06997_);
  or (_07001_, _06999_, _04952_);
  and (_07002_, _07001_, _07000_);
  and (_07003_, _07002_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_07004_, _07002_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_07005_, _07004_, _07003_);
  nor (_07006_, _07005_, _04872_);
  not (_07007_, _07006_);
  and (_07008_, _07007_, _04953_);
  nor (_07009_, _07008_, _06999_);
  not (_07010_, _07009_);
  and (_07011_, _07010_, _07000_);
  or (_07012_, _07011_, _06996_);
  and (_07013_, _06850_, _06821_);
  and (_07014_, _06905_, _07013_);
  nand (_07015_, _07014_, _06818_);
  or (_07016_, _07015_, _05773_);
  and (_07017_, _07016_, _07012_);
  and (_07018_, _07017_, _06993_);
  nor (_07019_, _05730_, _05132_);
  and (_07020_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_07021_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_07022_, _07021_, _07020_);
  and (_07023_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_07024_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_07025_, _07024_, _07023_);
  and (_07026_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_07027_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_07028_, _07027_, _07026_);
  and (_07029_, _07028_, _07025_);
  and (_07030_, _07029_, _07022_);
  nor (_07031_, _07030_, _06911_);
  nor (_07032_, _07031_, _07019_);
  or (_07033_, _07032_, _06907_);
  or (_07034_, _07015_, _05952_);
  and (_07035_, _07034_, _07033_);
  and (_07036_, _06957_, _06032_);
  and (_07037_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_07038_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_07039_, _07038_, _07037_);
  and (_07040_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_07041_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nor (_07042_, _07041_, _07040_);
  and (_07043_, _07042_, _07039_);
  nand (_07044_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nand (_07045_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_07046_, _07045_, _07044_);
  nand (_07047_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nand (_07048_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_07049_, _07048_, _07047_);
  and (_07050_, _07049_, _07046_);
  and (_07051_, _07050_, _06974_);
  and (_07052_, _07051_, _07043_);
  nor (_07053_, _07052_, _07036_);
  nand (_07054_, _07053_, _06929_);
  not (_07055_, _06999_);
  or (_07056_, _07055_, _06032_);
  not (_07057_, _04962_);
  nand (_07058_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  and (_07059_, _07058_, _07056_);
  and (_07060_, _07059_, _07003_);
  nor (_07061_, _07059_, _07003_);
  nor (_07062_, _07061_, _07060_);
  nor (_07063_, _07062_, _04872_);
  nor (_07064_, _07063_, _07057_);
  nor (_07065_, _07064_, _06999_);
  not (_07066_, _07065_);
  and (_07067_, _07066_, _07056_);
  or (_07068_, _07067_, _06996_);
  or (_07069_, _06994_, _07013_);
  or (_07070_, _07069_, _06818_);
  and (_07071_, _07070_, _07068_);
  and (_07072_, _07071_, _07054_);
  nand (_07073_, _07072_, _07035_);
  and (_07074_, _07073_, _07018_);
  or (_07075_, _07015_, _05797_);
  nor (_07076_, _05730_, _05152_);
  and (_07077_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_07078_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_07079_, _07078_, _07077_);
  and (_07080_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_07081_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_07082_, _07081_, _07080_);
  and (_07083_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_07084_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_07085_, _07084_, _07083_);
  and (_07086_, _07085_, _07082_);
  and (_07087_, _07086_, _07079_);
  nor (_07088_, _07087_, _06911_);
  nor (_07089_, _07088_, _07076_);
  or (_07090_, _07089_, _06907_);
  and (_07091_, _07090_, _07075_);
  and (_07092_, _06995_, _06818_);
  nand (_07093_, _06999_, _06705_);
  nand (_07094_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_07095_, _07094_, _07093_);
  and (_07096_, _07095_, _07060_);
  nor (_07097_, _07095_, _07060_);
  or (_07098_, _07097_, _07096_);
  nand (_07099_, _07098_, _04972_);
  nand (_07100_, _07099_, _04975_);
  nand (_07101_, _07100_, _07055_);
  nand (_07102_, _07101_, _07093_);
  nand (_07103_, _07102_, _07092_);
  or (_07104_, _06974_, _06705_);
  nand (_07105_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nand (_07106_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_07108_, _07106_, _07105_);
  nand (_07109_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nand (_07110_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_07111_, _07110_, _07109_);
  and (_07112_, _07111_, _07108_);
  not (_07113_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  nand (_07114_, _06960_, _06959_);
  or (_07115_, _07114_, _07113_);
  nand (_07116_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_07117_, _07116_, _07115_);
  nand (_07118_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nand (_07119_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_07120_, _07119_, _07118_);
  and (_07121_, _07120_, _07117_);
  and (_07122_, _07121_, _06974_);
  nand (_07123_, _07122_, _07112_);
  and (_07124_, _07123_, _07104_);
  nand (_07125_, _07124_, _06929_);
  and (_07126_, _07125_, _07103_);
  and (_07127_, _07126_, _07091_);
  or (_07128_, _07015_, _06947_);
  nor (_07129_, _05730_, _05084_);
  and (_07130_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_07131_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_07132_, _07131_, _07130_);
  and (_07133_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_07134_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_07135_, _07134_, _07133_);
  and (_07136_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_07137_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_07138_, _07137_, _07136_);
  and (_07139_, _07138_, _07135_);
  and (_07140_, _07139_, _07132_);
  nor (_07141_, _07140_, _06911_);
  nor (_07142_, _07141_, _07129_);
  or (_07143_, _07142_, _06907_);
  and (_07144_, _07143_, _07128_);
  nor (_07145_, _07055_, _05669_);
  and (_07146_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_07147_, _07146_, _07145_);
  and (_07148_, _07147_, _07096_);
  nor (_07149_, _07147_, _07096_);
  or (_07150_, _07149_, _07148_);
  nand (_07151_, _07150_, _04972_);
  nand (_07152_, _07151_, _04942_);
  and (_07153_, _07152_, _07055_);
  nor (_07154_, _07153_, _07145_);
  or (_07155_, _07154_, _06996_);
  and (_07156_, _06957_, _05669_);
  and (_07157_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_07158_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  nor (_07159_, _07158_, _07157_);
  and (_07160_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_07161_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_07162_, _07161_, _07160_);
  and (_07163_, _07162_, _07159_);
  nand (_07164_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nand (_07165_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_07166_, _07165_, _07164_);
  nand (_07167_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  nand (_07168_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_07169_, _07168_, _07167_);
  and (_07170_, _07169_, _07166_);
  and (_07171_, _07170_, _06974_);
  and (_07172_, _07171_, _07163_);
  nor (_07173_, _07172_, _07156_);
  nand (_07174_, _07173_, _06929_);
  and (_07175_, _07174_, _07155_);
  and (_07176_, _07175_, _07144_);
  and (_07177_, _07176_, _07127_);
  nor (_07178_, _05730_, _05062_);
  and (_07179_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_07180_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_07181_, _07180_, _07179_);
  and (_07182_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_07183_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_07184_, _07183_, _07182_);
  and (_07185_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_07186_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_07187_, _07186_, _07185_);
  and (_07188_, _07187_, _07184_);
  and (_07189_, _07188_, _07181_);
  nor (_07190_, _06911_, _07189_);
  nor (_07191_, _07190_, _07178_);
  or (_07192_, _07191_, _06907_);
  or (_07193_, _07015_, _06938_);
  and (_07194_, _07193_, _07192_);
  nor (_07195_, _06974_, _06410_);
  and (_07196_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_07197_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  nor (_07198_, _07197_, _07196_);
  and (_07199_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  and (_07200_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_07201_, _07200_, _07199_);
  and (_07202_, _07201_, _07198_);
  nand (_07203_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nand (_07204_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_07205_, _07204_, _07203_);
  nand (_07206_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  nand (_07207_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_07208_, _07207_, _07206_);
  and (_07209_, _07208_, _07205_);
  and (_07210_, _07209_, _06974_);
  and (_07211_, _07210_, _07202_);
  nor (_07212_, _07211_, _07195_);
  nand (_07213_, _07212_, _06929_);
  and (_07214_, _06999_, _06410_);
  and (_07215_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_07216_, _07215_, _07214_);
  nand (_07217_, _07216_, _07148_);
  or (_07218_, _07216_, _07148_);
  nand (_07219_, _07218_, _07217_);
  nand (_07220_, _07219_, _04972_);
  nand (_07221_, _07220_, _04910_);
  and (_07222_, _07221_, _07055_);
  or (_07223_, _07222_, _07214_);
  nand (_07224_, _07223_, _07092_);
  or (_07225_, _06851_, _06818_);
  and (_07226_, _07225_, _07224_);
  and (_07227_, _07226_, _07213_);
  and (_07228_, _07227_, _07194_);
  or (_07229_, _06974_, _05718_);
  nand (_07230_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  nand (_07231_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_07232_, _07231_, _07230_);
  nand (_07233_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nand (_07234_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_07235_, _07234_, _07233_);
  and (_07236_, _07235_, _07232_);
  nand (_07237_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nand (_07238_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_07239_, _07238_, _07237_);
  nand (_07240_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  nand (_07241_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_07242_, _07241_, _07240_);
  and (_07243_, _07242_, _07239_);
  and (_07244_, _07243_, _06974_);
  nand (_07245_, _07244_, _07236_);
  and (_07246_, _07245_, _07229_);
  nand (_07247_, _07246_, _06929_);
  nor (_07248_, _05730_, _05179_);
  and (_07249_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_07250_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_07251_, _07250_, _07249_);
  and (_07252_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_07253_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_07254_, _07253_, _07252_);
  and (_07255_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_07256_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_07257_, _07256_, _07255_);
  and (_07258_, _07257_, _07254_);
  and (_07259_, _07258_, _07251_);
  nor (_07260_, _07259_, _06911_);
  nor (_07261_, _07260_, _07248_);
  or (_07262_, _07261_, _06907_);
  and (_07263_, _07262_, _07247_);
  and (_07264_, _06999_, _05718_);
  and (_07265_, _07216_, _07148_);
  and (_07266_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_07267_, _07266_, _07264_);
  nand (_07268_, _07267_, _07265_);
  or (_07269_, _07267_, _07265_);
  nand (_07270_, _07269_, _07268_);
  nand (_07271_, _07270_, _04972_);
  nand (_07272_, _07271_, _04925_);
  and (_07273_, _07272_, _07055_);
  nor (_07274_, _07273_, _07264_);
  or (_07275_, _07274_, _07013_);
  nand (_07276_, _07275_, _06818_);
  and (_07277_, _07069_, _06906_);
  nand (_07278_, _07277_, _07276_);
  and (_07279_, _07278_, _07263_);
  or (_07280_, _06928_, _06818_);
  nor (_07281_, _05730_, _05017_);
  and (_07282_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_07283_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_07284_, _07283_, _07282_);
  and (_07285_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_07286_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_07287_, _07286_, _07285_);
  and (_07288_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_07289_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_07290_, _07289_, _07288_);
  and (_07291_, _07290_, _07287_);
  and (_07292_, _07291_, _07284_);
  nor (_07293_, _07292_, _06911_);
  nor (_07294_, _07293_, _07281_);
  or (_07295_, _07294_, _06907_);
  and (_07296_, _07295_, _07280_);
  nor (_07297_, _07055_, _05287_);
  and (_07299_, _07267_, _07265_);
  and (_07300_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_07301_, _07300_, _07297_);
  or (_07303_, _07301_, _07299_);
  nand (_07304_, _07301_, _07299_);
  nand (_07305_, _07304_, _07303_);
  nand (_07306_, _07305_, _04972_);
  nand (_07308_, _07306_, _04875_);
  and (_07309_, _07308_, _07055_);
  or (_07310_, _07309_, _07297_);
  nand (_07311_, _07310_, _07092_);
  nand (_07312_, _06957_, _05287_);
  or (_07314_, _07114_, _04857_);
  nand (_07315_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_07316_, _07315_, _07314_);
  nand (_07317_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  nand (_07319_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  and (_07320_, _07319_, _07317_);
  and (_07321_, _07320_, _07316_);
  nand (_07322_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nand (_07323_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_07325_, _07323_, _07322_);
  nand (_07326_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  nand (_07327_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_07328_, _07327_, _07326_);
  and (_07330_, _07328_, _07325_);
  and (_07331_, _07330_, _06974_);
  nand (_07333_, _07331_, _07321_);
  and (_07334_, _07333_, _07312_);
  nand (_07335_, _07334_, _06929_);
  and (_07336_, _07335_, _07311_);
  and (_07337_, _07336_, _07296_);
  and (_07338_, _06999_, _06284_);
  and (_07339_, _07055_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  or (_07340_, _07339_, _07304_);
  nand (_07341_, _07339_, _07304_);
  nand (_07342_, _07341_, _07340_);
  nand (_07343_, _07342_, _04972_);
  and (_07344_, _07055_, _04897_);
  and (_07345_, _07344_, _07343_);
  nor (_07346_, _07345_, _07338_);
  nand (_07347_, _07346_, _06995_);
  nand (_07348_, _06957_, _06284_);
  and (_07349_, _06968_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_07350_, _06979_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_07351_, _07350_, _07349_);
  and (_07352_, _06961_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_07353_, _06983_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  or (_07354_, _07353_, _07352_);
  or (_07355_, _07354_, _07351_);
  nand (_07356_, _06970_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nand (_07357_, _06964_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_07358_, _07357_, _07356_);
  nand (_07359_, _06976_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nand (_07360_, _06985_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_07361_, _07360_, _07359_);
  and (_07362_, _07361_, _07358_);
  nand (_07363_, _07362_, _06974_);
  or (_07364_, _07363_, _07355_);
  and (_07365_, _07364_, _07348_);
  nand (_07366_, _07365_, _06929_);
  nor (_07367_, _05730_, _05321_);
  and (_07368_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_07369_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_07370_, _07369_, _07368_);
  and (_07371_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_07372_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_07373_, _07372_, _07371_);
  and (_07374_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  and (_07375_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_07376_, _07375_, _07374_);
  and (_07377_, _07376_, _07373_);
  and (_07378_, _07377_, _07370_);
  nor (_07379_, _07378_, _06911_);
  nor (_07380_, _07379_, _07367_);
  or (_07381_, _07380_, _06906_);
  and (_07382_, _07381_, _06818_);
  and (_07383_, _07382_, _07366_);
  nand (_07384_, _07383_, _07347_);
  and (_07385_, _07384_, _07337_);
  and (_07386_, _07385_, _07279_);
  and (_07387_, _07386_, _07228_);
  and (_07388_, _07387_, _07177_);
  and (_07389_, _07388_, _07074_);
  and (_07390_, _07389_, _05292_);
  not (_07391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  nand (_07392_, _07017_, _06993_);
  or (_07393_, _07073_, _07392_);
  nand (_07394_, _07175_, _07144_);
  and (_07395_, _07394_, _07127_);
  not (_07396_, _07395_);
  or (_07397_, _07396_, _07393_);
  nand (_07398_, _07227_, _07194_);
  nand (_07399_, _07278_, _07263_);
  and (_07400_, _07383_, _07347_);
  or (_07401_, _07400_, _07337_);
  or (_07402_, _07401_, _07399_);
  or (_07403_, _07402_, _07398_);
  or (_07404_, _07403_, _07397_);
  nor (_07405_, _07404_, _07391_);
  nand (_07406_, _07126_, _07091_);
  and (_07407_, _07394_, _07406_);
  not (_07408_, _07407_);
  or (_07409_, _07408_, _07393_);
  or (_07410_, _07409_, _07403_);
  not (_07411_, _07410_);
  and (_07412_, _07411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_07414_, _07412_, _07405_);
  and (_07415_, _07072_, _07035_);
  or (_07417_, _07415_, _07392_);
  or (_07418_, _07417_, _07396_);
  or (_07420_, _07418_, _07403_);
  not (_07422_, _07420_);
  and (_07424_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_07425_, _07073_, _07018_);
  or (_07426_, _07408_, _07425_);
  or (_07428_, _07426_, _07403_);
  not (_07429_, _07428_);
  and (_07430_, _07429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_07432_, _07430_, _07424_);
  or (_07433_, _07432_, _07414_);
  nand (_07435_, _07386_, _07228_);
  or (_07436_, _07397_, _07435_);
  not (_07437_, _07436_);
  and (_07438_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_07439_, _07415_, _07018_);
  or (_07440_, _07439_, _07396_);
  or (_07441_, _07403_, _07440_);
  not (_07442_, _07441_);
  and (_07443_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or (_07444_, _07443_, _07438_);
  and (_07445_, _07415_, _07018_);
  and (_07446_, _07395_, _07445_);
  and (_07447_, _07385_, _07399_);
  and (_07448_, _07447_, _07228_);
  and (_07449_, _07448_, _07446_);
  and (_07450_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_07451_, _07447_, _07398_);
  and (_07452_, _07073_, _07392_);
  and (_07453_, _07452_, _07406_);
  and (_07454_, _07453_, _07176_);
  and (_07455_, _07454_, _07451_);
  and (_07456_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_07457_, _07456_, _07450_);
  or (_07458_, _07457_, _07444_);
  or (_07459_, _07458_, _07433_);
  not (_07460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_07461_, _07415_, _07392_);
  and (_07462_, _07461_, _07395_);
  nand (_07463_, _07462_, _07387_);
  nor (_07464_, _07463_, _07460_);
  or (_07465_, _07440_, _07435_);
  not (_07466_, _07465_);
  and (_07467_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or (_07468_, _07467_, _07464_);
  or (_07469_, _07418_, _07435_);
  not (_07470_, _07469_);
  and (_07471_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or (_07472_, _07426_, _07435_);
  not (_07473_, _07472_);
  and (_07474_, _07473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or (_07475_, _07474_, _07471_);
  or (_07476_, _07475_, _07468_);
  nor (_07477_, _07409_, _07435_);
  and (_07478_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_07479_, _07454_, _07387_);
  and (_07480_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  or (_07481_, _07480_, _07478_);
  and (_07482_, _07386_, _07398_);
  nand (_07483_, _07482_, _07462_);
  not (_07484_, _07483_);
  and (_07485_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  nand (_07486_, _07482_, _07446_);
  not (_07487_, _07486_);
  and (_07488_, _07487_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_07489_, _07488_, _07485_);
  or (_07490_, _07489_, _07481_);
  or (_07491_, _07490_, _07476_);
  or (_07492_, _07491_, _07459_);
  and (_07493_, _07389_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_07494_, _07388_, _07452_);
  and (_07495_, _07494_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_07496_, _07495_, _07493_);
  and (_07497_, _07445_, _07177_);
  and (_07498_, _07497_, _07398_);
  nor (_07499_, _07401_, _07279_);
  and (_07500_, _07499_, _07498_);
  and (_07501_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_07502_, _07387_, _07177_);
  or (_07503_, _07502_, _07425_);
  nor (_07504_, _07503_, _07011_);
  or (_07505_, _07504_, _07501_);
  or (_07506_, _07505_, _07496_);
  and (_07507_, _07448_, _07497_);
  and (_07508_, _06635_, _06731_);
  nor (_07509_, _07508_, _06866_);
  and (_07510_, _06637_, _05874_);
  and (_07511_, _07510_, _05985_);
  nor (_07512_, _07511_, _06744_);
  and (_07513_, _06635_, _05965_);
  nor (_07514_, _06619_, _05950_);
  nor (_07515_, _07514_, _05822_);
  nor (_07516_, _07515_, _07513_);
  nor (_07518_, _06756_, _06750_);
  and (_07519_, _07518_, _07516_);
  and (_07521_, _07519_, _07512_);
  nor (_07522_, _06888_, _06609_);
  nor (_07523_, _06755_, _06595_);
  and (_07525_, _07523_, _07522_);
  and (_07526_, _07525_, _06748_);
  and (_07527_, _07526_, _07521_);
  and (_07528_, _07527_, _06887_);
  and (_07530_, _07528_, _07509_);
  nor (_07531_, _07530_, _06799_);
  or (_07532_, _07531_, p2_in[0]);
  not (_07533_, _07531_);
  or (_07535_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_07536_, _07535_, _07532_);
  and (_07538_, _07536_, _07507_);
  and (_07539_, _07451_, _07497_);
  or (_07541_, _07531_, p3_in[0]);
  or (_07542_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_07544_, _07542_, _07541_);
  and (_07545_, _07544_, _07539_);
  or (_07546_, _07545_, _07538_);
  and (_07547_, _07387_, _07497_);
  or (_07548_, _07531_, p0_in[0]);
  or (_07549_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_07550_, _07549_, _07548_);
  and (_07551_, _07550_, _07547_);
  and (_07552_, _07482_, _07497_);
  or (_07553_, _07531_, p1_in[0]);
  or (_07554_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_07555_, _07554_, _07553_);
  and (_07556_, _07555_, _07552_);
  or (_07557_, _07556_, _07551_);
  or (_07558_, _07557_, _07546_);
  or (_07559_, _07558_, _07506_);
  not (_07560_, _07402_);
  and (_07561_, _07560_, _07498_);
  nor (_07562_, _06666_, _06488_);
  and (_07563_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_07564_, _07563_, _07562_);
  nor (_07565_, _07564_, _06654_);
  not (_07566_, _07565_);
  and (_07567_, _06654_, _06452_);
  not (_07568_, _06673_);
  nor (_07569_, _06146_, _05042_);
  nor (_07570_, _07569_, _06147_);
  nor (_07571_, _07570_, _07568_);
  nor (_07572_, _07571_, _07567_);
  nand (_07573_, _07572_, _07566_);
  nand (_07574_, _07573_, _06684_);
  or (_07575_, _07573_, _06684_);
  and (_07576_, _07575_, _07574_);
  or (_07577_, _05445_, _05442_);
  nor (_07578_, _05446_, _06454_);
  nand (_07579_, _07578_, _07577_);
  nor (_07580_, _05466_, _05227_);
  nor (_07581_, _05477_, _05059_);
  nor (_07582_, _07581_, _07580_);
  and (_07583_, _07582_, _05368_);
  nor (_07584_, _07582_, _05368_);
  or (_07585_, _07584_, _07583_);
  and (_07586_, _07585_, _05223_);
  nor (_07587_, _05490_, _05048_);
  nor (_07588_, _05368_, _05274_);
  and (_07589_, _05497_, ABINPUT000000[11]);
  or (_07590_, _07589_, _07588_);
  nor (_07591_, _07590_, _07587_);
  nor (_07592_, _05232_, _05172_);
  and (_07593_, _05499_, ABINPUT000[11]);
  nor (_07594_, _07593_, _07592_);
  and (_07595_, _07594_, _07591_);
  not (_07596_, _07595_);
  nor (_07597_, _07596_, _07586_);
  nand (_07598_, _07597_, _07579_);
  nand (_07599_, _07598_, _06654_);
  nor (_07600_, _06672_, _05167_);
  nor (_07601_, _07600_, _06675_);
  and (_07602_, _06494_, _06144_);
  nor (_07603_, _06494_, _05167_);
  or (_07604_, _07603_, _07602_);
  nand (_07605_, _07604_, _06672_);
  and (_07606_, _07605_, _07601_);
  nor (_07607_, _06654_, _06552_);
  nor (_07609_, _07607_, _06667_);
  or (_07610_, _07609_, _07606_);
  nand (_07612_, _07610_, _07599_);
  or (_07613_, _05446_, _05310_);
  nor (_07614_, _05447_, _06454_);
  nand (_07616_, _07614_, _07613_);
  and (_07617_, _05478_, _05227_);
  and (_07619_, _05467_, _05059_);
  nor (_07620_, _07619_, _07617_);
  and (_07621_, _07620_, _05356_);
  not (_07622_, _07621_);
  nor (_07624_, _07620_, _05356_);
  nor (_07625_, _07624_, _06363_);
  and (_07626_, _07625_, _07622_);
  nor (_07628_, _05356_, _05274_);
  and (_07629_, _05497_, ABINPUT000000[12]);
  or (_07631_, _07629_, _07628_);
  nor (_07632_, _07631_, _06061_);
  nor (_07633_, _05232_, _05103_);
  and (_07634_, _05499_, ABINPUT000[12]);
  nor (_07636_, _07634_, _07633_);
  and (_07637_, _07636_, _07632_);
  not (_07638_, _07637_);
  nor (_07639_, _07638_, _07626_);
  nand (_07640_, _07639_, _07616_);
  or (_07641_, _07640_, _06656_);
  and (_07642_, _06144_, _05520_);
  nor (_07643_, _05520_, _05099_);
  or (_07644_, _07643_, _07642_);
  nand (_07645_, _07644_, _06673_);
  nor (_07646_, _06666_, _06586_);
  and (_07647_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_07648_, _07647_, _07646_);
  and (_07649_, _07648_, _07645_);
  nand (_07650_, _07649_, _06656_);
  nand (_07651_, _07650_, _07641_);
  nand (_07652_, _07651_, _07612_);
  or (_07653_, _07651_, _07612_);
  and (_07654_, _07653_, _07652_);
  or (_07655_, _05437_, _05434_);
  nor (_07656_, _05438_, _06454_);
  nand (_07657_, _07656_, _07655_);
  and (_07658_, _05464_, _05059_);
  and (_07659_, _05475_, _05227_);
  nor (_07660_, _07659_, _07658_);
  and (_07661_, _07660_, _05383_);
  nor (_07662_, _07660_, _05383_);
  nor (_07663_, _07662_, _07661_);
  and (_07664_, _07663_, _05223_);
  nor (_07665_, _05490_, _05081_);
  nor (_07666_, _05383_, _05274_);
  and (_07667_, _05497_, ABINPUT000000[9]);
  or (_07668_, _07667_, _07666_);
  nor (_07669_, _07668_, _07665_);
  and (_07670_, _05231_, _05206_);
  and (_07671_, _05499_, ABINPUT000[9]);
  nor (_07672_, _07671_, _07670_);
  and (_07673_, _07672_, _07669_);
  not (_07674_, _07673_);
  nor (_07675_, _07674_, _07664_);
  nand (_07676_, _07675_, _07657_);
  and (_07677_, _07676_, _06654_);
  nor (_07678_, _05397_, _05059_);
  nor (_07679_, _07678_, _05398_);
  not (_07680_, _07679_);
  nor (_07681_, _05455_, _05583_);
  nor (_07682_, _07681_, _07680_);
  not (_07683_, _07682_);
  and (_07684_, _05530_, _06064_);
  and (_07685_, _05489_, _05059_);
  and (_07686_, _05497_, ABINPUT000000[1]);
  and (_07687_, _05499_, ABINPUT000[1]);
  nor (_07688_, _07687_, _07686_);
  not (_07689_, _07688_);
  nor (_07690_, _07689_, _07685_);
  not (_07691_, _07690_);
  nor (_07692_, _07691_, _07684_);
  or (_07693_, _06468_, _05151_);
  nor (_07694_, _05557_, _05273_);
  nor (_07695_, _07694_, _05126_);
  not (_07696_, _07695_);
  and (_07697_, _07696_, _07693_);
  and (_07698_, _07697_, _07692_);
  and (_07699_, _07698_, _06365_);
  and (_07700_, _07699_, _06361_);
  and (_07701_, _07700_, _06358_);
  and (_07702_, _07701_, _07683_);
  nor (_07703_, _07702_, _06666_);
  and (_07704_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_07705_, _07704_, _07703_);
  nor (_07706_, _07705_, _06654_);
  nor (_07707_, _07706_, _07677_);
  and (_07708_, _06144_, _04990_);
  nor (_07709_, _04990_, _05122_);
  or (_07710_, _07709_, _07708_);
  nand (_07711_, _07710_, _06673_);
  and (_07712_, _07711_, _07707_);
  and (_07713_, _06144_, _04986_);
  nor (_07714_, _04986_, _05147_);
  or (_07715_, _07714_, _07713_);
  nand (_07716_, _07715_, _06673_);
  or (_07717_, _05441_, _05438_);
  nor (_07718_, _05442_, _06454_);
  nand (_07719_, _07718_, _07717_);
  and (_07720_, _05476_, _05227_);
  and (_07721_, _05465_, _05059_);
  nor (_07722_, _07721_, _07720_);
  nor (_07723_, _07722_, _05377_);
  and (_07724_, _07722_, _05377_);
  nor (_07725_, _07724_, _07723_);
  nor (_07726_, _07725_, _06363_);
  nor (_07727_, _05490_, _05199_);
  and (_07729_, _05377_, _05273_);
  and (_07730_, _05497_, ABINPUT000000[10]);
  or (_07732_, _07730_, _07729_);
  nor (_07733_, _07732_, _07727_);
  and (_07735_, _05231_, _05207_);
  and (_07736_, _05499_, ABINPUT000[10]);
  nor (_07737_, _07736_, _07735_);
  and (_07739_, _07737_, _07733_);
  not (_07740_, _07739_);
  nor (_07741_, _07740_, _07726_);
  nand (_07743_, _07741_, _07719_);
  and (_07744_, _07743_, _06654_);
  nor (_07746_, _05618_, _05617_);
  nor (_07748_, _07746_, _05619_);
  nor (_07749_, _07748_, _05584_);
  not (_07751_, _07749_);
  or (_07752_, _06468_, _05172_);
  and (_07753_, _05497_, ABINPUT000000[2]);
  and (_07754_, _05499_, ABINPUT000[2]);
  nor (_07755_, _07754_, _07753_);
  and (_07756_, _07755_, _07752_);
  and (_07757_, _05273_, _05207_);
  and (_07758_, _05280_, _05206_);
  nor (_07759_, _07758_, _07757_);
  and (_07760_, _07759_, _07756_);
  and (_07761_, _07760_, _06030_);
  and (_07762_, _06512_, _05207_);
  nor (_07763_, _07762_, _06513_);
  nor (_07764_, _07763_, _05558_);
  not (_07765_, _05385_);
  and (_07766_, _06020_, _07765_);
  or (_07767_, _07766_, _05389_);
  and (_07768_, _07767_, _05398_);
  nor (_07769_, _07767_, _05398_);
  or (_07770_, _07769_, _07768_);
  and (_07771_, _07770_, _05455_);
  nor (_07772_, _07771_, _07764_);
  and (_07773_, _07772_, _07761_);
  and (_07774_, _07773_, _07751_);
  nor (_07775_, _07774_, _06666_);
  and (_07776_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  nor (_07777_, _07776_, _07775_);
  nor (_07778_, _07777_, _06654_);
  nor (_07779_, _07778_, _07744_);
  nand (_07780_, _07779_, _07716_);
  nand (_07781_, _07780_, _07712_);
  or (_07782_, _07780_, _07712_);
  nand (_07783_, _07782_, _07781_);
  nand (_07784_, _07783_, _07654_);
  or (_07785_, _07783_, _07654_);
  nand (_07786_, _07785_, _07784_);
  nor (_07787_, _05627_, _05349_);
  and (_07788_, _05627_, _05349_);
  nor (_07789_, _07788_, _07787_);
  and (_07790_, _07789_, _05583_);
  not (_07791_, _07790_);
  nor (_07792_, _05407_, _05349_);
  nor (_07793_, _07792_, _06454_);
  and (_07794_, _07793_, _05408_);
  nor (_07795_, _05560_, _05565_);
  not (_07796_, _07795_);
  nor (_07797_, _05567_, _05558_);
  and (_07798_, _07797_, _07796_);
  and (_07799_, _05280_, _05204_);
  and (_07800_, _05497_, ABINPUT000000[5]);
  and (_07801_, _05499_, ABINPUT000[5]);
  nor (_07802_, _07801_, _07800_);
  not (_07803_, _07802_);
  nor (_07804_, _07803_, _07799_);
  or (_07805_, _06468_, _05199_);
  not (_07806_, _07805_);
  nor (_07807_, _05274_, _05081_);
  nor (_07808_, _07807_, _07806_);
  and (_07809_, _07808_, _07804_);
  not (_07810_, _07809_);
  nor (_07811_, _07810_, _07798_);
  and (_07812_, _07811_, _06409_);
  not (_07813_, _07812_);
  nor (_07814_, _07813_, _07794_);
  and (_07815_, _07814_, _07791_);
  nor (_07816_, _07815_, _06666_);
  and (_07817_, _06678_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_07818_, _07817_, _07816_);
  nor (_07819_, _07818_, _06654_);
  not (_07820_, _07819_);
  or (_07821_, _05450_, _05447_);
  and (_07822_, _05451_, _05455_);
  and (_07823_, _07822_, _07821_);
  and (_07824_, _05468_, _05059_);
  and (_07825_, _07617_, _05622_);
  nor (_07826_, _07825_, _07824_);
  nand (_07828_, _07826_, _05346_);
  or (_07829_, _07826_, _05346_);
  and (_07831_, _07829_, _07828_);
  and (_07832_, _07831_, _05223_);
  and (_07833_, _05489_, _05206_);
  nand (_07835_, _05081_, _05059_);
  and (_07836_, _05346_, _05227_);
  nor (_07838_, _07836_, _05232_);
  and (_07840_, _07838_, _07835_);
  nor (_07841_, _05346_, _05274_);
  and (_07843_, _05497_, ABINPUT000000[13]);
  and (_07845_, _05499_, ABINPUT000[13]);
  or (_07846_, _07845_, _07843_);
  or (_07847_, _07846_, _07841_);
  or (_07848_, _07847_, _07840_);
  or (_07850_, _07848_, _07833_);
  or (_07851_, _07850_, _07832_);
  or (_07853_, _07851_, _07823_);
  nand (_07854_, _07853_, _06654_);
  and (_07855_, _04989_, _06090_);
  and (_07857_, _07855_, _06144_);
  nor (_07858_, _07855_, _05075_);
  or (_07859_, _07858_, _07857_);
  nand (_07860_, _07859_, _06673_);
  and (_07861_, _07860_, _07854_);
  nand (_07862_, _07861_, _07820_);
  nor (_07863_, _06672_, _05194_);
  nor (_07864_, _07863_, _06675_);
  and (_07865_, _06091_, _06144_);
  nor (_07866_, _06091_, _05194_);
  or (_07867_, _07866_, _07865_);
  nand (_07868_, _07867_, _06673_);
  and (_07869_, _07868_, _07864_);
  nor (_07870_, _05628_, _05600_);
  nor (_07871_, _07870_, _05629_);
  nor (_07872_, _07871_, _05584_);
  not (_07873_, _07872_);
  and (_07874_, _05421_, _05408_);
  nor (_07875_, _07874_, _06454_);
  and (_07876_, _07875_, _05422_);
  nor (_07877_, _05568_, _05199_);
  nor (_07878_, _07877_, _06462_);
  nor (_07879_, _07878_, _05558_);
  and (_07880_, _05280_, _05565_);
  and (_07881_, _05497_, ABINPUT000000[6]);
  and (_07882_, _05499_, ABINPUT000[6]);
  nor (_07883_, _07882_, _07881_);
  not (_07884_, _07883_);
  nor (_07885_, _07884_, _07880_);
  or (_07886_, _06468_, _05048_);
  nor (_07887_, _05274_, _05199_);
  not (_07888_, _07887_);
  and (_07889_, _07888_, _07886_);
  and (_07890_, _07889_, _07885_);
  and (_07891_, _07890_, _05716_);
  not (_07892_, _07891_);
  nor (_07893_, _07892_, _07879_);
  and (_07894_, _07893_, _05702_);
  not (_07895_, _07894_);
  nor (_07896_, _07895_, _07876_);
  and (_07897_, _07896_, _07873_);
  and (_07898_, _07897_, _06675_);
  or (_07899_, _07898_, _07869_);
  nand (_07900_, _07899_, _06656_);
  nand (_07901_, _05451_, _05307_);
  and (_07902_, _05452_, _05455_);
  and (_07903_, _07902_, _07901_);
  not (_07904_, _05414_);
  nor (_07905_, _07825_, _05469_);
  nor (_07906_, _07905_, _07836_);
  or (_07907_, _07906_, _07904_);
  nand (_07908_, _07906_, _07904_);
  and (_07909_, _07908_, _07907_);
  and (_07910_, _07909_, _05223_);
  and (_07911_, _05489_, _05207_);
  nor (_07912_, _05199_, _05227_);
  or (_07913_, _07912_, _05479_);
  and (_07914_, _07913_, _05231_);
  nor (_07915_, _05414_, _05274_);
  and (_07916_, _05497_, ABINPUT000000[14]);
  and (_07917_, _05499_, ABINPUT000[14]);
  or (_07918_, _07917_, _07916_);
  or (_07919_, _07918_, _07915_);
  or (_07920_, _07919_, _07914_);
  or (_07921_, _07920_, _07911_);
  or (_07922_, _07921_, _07910_);
  or (_07924_, _07922_, _07903_);
  or (_07925_, _07924_, _06656_);
  nand (_07927_, _07925_, _07900_);
  nand (_07928_, _07927_, _07862_);
  or (_07929_, _07927_, _07862_);
  nand (_07931_, _07929_, _07928_);
  nand (_07932_, _07931_, _07786_);
  or (_07933_, _07931_, _07786_);
  nand (_07935_, _07933_, _07932_);
  nor (_07936_, _07935_, _07576_);
  and (_07937_, _07935_, _07576_);
  or (_07939_, _07937_, _07936_);
  and (_07940_, _07939_, _07561_);
  and (_07942_, _07499_, _07228_);
  and (_07943_, _07942_, _07497_);
  and (_07944_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_07945_, _07944_, _07940_);
  or (_07947_, _07945_, _07559_);
  or (_07948_, _07947_, _07492_);
  nor (_07949_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  not (_07951_, _07949_);
  nand (_07952_, _07951_, _07561_);
  or (_07953_, _07502_, _07439_);
  or (_07954_, _07953_, _05293_);
  nand (_07955_, _07943_, _06654_);
  and (_07956_, _07955_, _07954_);
  nand (_07957_, _07956_, _07952_);
  nand (_07958_, _07957_, _04859_);
  or (_07959_, _07228_, _06930_);
  or (_07960_, _07398_, _04922_);
  nand (_07961_, _07960_, _07959_);
  or (_07962_, _07392_, _04958_);
  or (_07963_, _07018_, _04959_);
  nand (_07964_, _07963_, _07962_);
  nor (_07965_, _07964_, _07961_);
  or (_07966_, _07073_, _04971_);
  or (_07967_, _07279_, _04932_);
  or (_07968_, _07399_, _04933_);
  and (_07969_, _07968_, _07967_);
  or (_07970_, _07337_, _04893_);
  nand (_07971_, _07336_, _07296_);
  or (_07972_, _07971_, _05513_);
  and (_07973_, _07972_, _07970_);
  nor (_07974_, _07973_, _07969_);
  and (_07975_, _07974_, _07966_);
  and (_07976_, _07975_, _07965_);
  or (_07977_, _07176_, _04947_);
  or (_07978_, _07394_, _04948_);
  and (_07979_, _07978_, _07977_);
  or (_07980_, _07400_, _04904_);
  or (_07981_, _07384_, _06133_);
  and (_07982_, _07981_, _07980_);
  nor (_07983_, _07982_, _07979_);
  or (_07984_, _07127_, _06090_);
  or (_07985_, _07406_, _04984_);
  nand (_07986_, _07985_, _07984_);
  or (_07987_, _07415_, _04996_);
  nand (_07988_, _07987_, _06092_);
  nor (_07989_, _07988_, _07986_);
  and (_07990_, _07989_, _07983_);
  nand (_07991_, _07990_, _07976_);
  or (_07992_, _04904_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  or (_07993_, _07992_, _07991_);
  not (_07994_, _07961_);
  and (_07995_, _07974_, _07994_);
  and (_07996_, _07995_, _07983_);
  not (_07997_, _07453_);
  and (_07998_, _07997_, _06141_);
  nand (_07999_, _07998_, _07996_);
  nand (_08000_, _07943_, _06660_);
  and (_08001_, _08000_, _07999_);
  nand (_08002_, _08001_, _07993_);
  nand (_08003_, _08002_, _04859_);
  and (_08004_, _08003_, _07958_);
  and (_08005_, _08004_, _07948_);
  and (_08006_, _07410_, _07404_);
  and (_08007_, _07428_, _07420_);
  and (_08008_, _08007_, _08006_);
  and (_08009_, _07441_, _07436_);
  nor (_08010_, _07455_, _07449_);
  and (_08011_, _08010_, _08009_);
  and (_08012_, _08011_, _08008_);
  and (_08013_, _07465_, _07463_);
  and (_08014_, _07472_, _07469_);
  and (_08015_, _08014_, _08013_);
  nor (_08016_, _07479_, _07477_);
  and (_08017_, _07486_, _07483_);
  and (_08018_, _08017_, _08016_);
  and (_08019_, _08018_, _08015_);
  and (_08021_, _08019_, _08012_);
  nor (_08022_, _07943_, _07561_);
  nand (_08024_, _07385_, _07497_);
  or (_08025_, _07502_, _07417_);
  and (_08027_, _07953_, _08025_);
  and (_08028_, _07388_, _07461_);
  nor (_08029_, _08028_, _07500_);
  and (_08031_, _08029_, _08027_);
  and (_08032_, _08031_, _08024_);
  and (_08033_, _08032_, _08022_);
  nand (_08034_, _08033_, _08021_);
  and (_08036_, _08034_, _07958_);
  nand (_08037_, _08036_, _08003_);
  and (_08038_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or (_08040_, _08038_, _08005_);
  or (_08041_, _08040_, _07390_);
  nand (_08043_, _07390_, _07702_);
  and (_08044_, _08043_, _04856_);
  and (_05133_, _08044_, _08041_);
  and (_08046_, _06721_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_08047_, _06624_, _05998_);
  or (_08048_, _08047_, _06838_);
  or (_08049_, _08048_, _06727_);
  and (_08050_, _07510_, _05978_);
  or (_08051_, _08050_, _06747_);
  and (_08052_, _06612_, _05998_);
  or (_08053_, _08052_, _06788_);
  or (_08054_, _08053_, _08051_);
  or (_08055_, _08054_, _08049_);
  and (_08056_, _08055_, _06770_);
  or (_05136_, _08056_, _08046_);
  nor (_08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , rst);
  and (_08058_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  not (_08059_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor (_08060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_08061_, _08060_, _08059_);
  and (_08062_, _08061_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_08063_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_08064_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _08063_);
  not (_08065_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_08066_, _08065_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_08067_, _08066_, _08064_);
  not (_08068_, _08067_);
  and (_08069_, _08068_, _08062_);
  not (_08070_, _08060_);
  and (_08071_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_08072_, _08071_, _08070_);
  not (_08073_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_08074_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _08073_);
  and (_08075_, _08074_, _08059_);
  and (_08076_, _08075_, _08060_);
  nor (_08077_, _08076_, _08062_);
  not (_08078_, _08077_);
  nor (_08079_, _08078_, _08072_);
  nor (_08080_, _08079_, _08069_);
  and (_08081_, _08060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_08082_, _08081_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  or (_08083_, _08082_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_08084_, _08083_, _08080_);
  and (_08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _04856_);
  and (_08086_, _08067_, _08062_);
  nor (_08087_, _08086_, _08082_);
  or (_08088_, _08087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_08089_, _08088_, _08085_);
  and (_08090_, _08089_, _08084_);
  or (_05143_, _08090_, _08058_);
  not (_08091_, _05843_);
  not (_08092_, _05818_);
  and (_08093_, _08092_, _05793_);
  and (_08094_, _08093_, _08091_);
  and (_08095_, _08094_, _05767_);
  not (_08096_, _05895_);
  and (_08097_, _08096_, _05870_);
  and (_08098_, _05943_, _05919_);
  and (_08099_, _08098_, _08097_);
  and (_08100_, _08099_, _08095_);
  not (_08101_, _05919_);
  nor (_08102_, _05943_, _08101_);
  and (_08103_, _05895_, _05870_);
  and (_08104_, _08103_, _08102_);
  and (_08105_, _08104_, _08094_);
  nor (_08106_, _08105_, _08100_);
  nor (_08107_, _05818_, _05793_);
  nor (_08108_, _05767_, _05843_);
  and (_08109_, _08108_, _08107_);
  nor (_08110_, _05943_, _05919_);
  and (_08111_, _08110_, _08097_);
  not (_08112_, _05870_);
  and (_08113_, _05895_, _08112_);
  and (_08114_, _08113_, _08110_);
  or (_08115_, _08114_, _08111_);
  and (_08116_, _08115_, _08109_);
  not (_08117_, _05767_);
  and (_08119_, _08107_, _05843_);
  and (_08120_, _08119_, _08117_);
  and (_08121_, _08110_, _08096_);
  and (_08122_, _08121_, _08120_);
  nor (_08123_, _08122_, _08116_);
  nand (_08124_, _08123_, _08106_);
  and (_08125_, _05943_, _08101_);
  and (_08126_, _08125_, _08103_);
  and (_08127_, _08126_, _08109_);
  and (_08128_, _08107_, _08091_);
  not (_08130_, _08128_);
  and (_08131_, _08125_, _08113_);
  nor (_08132_, _08131_, _05767_);
  nor (_08133_, _08132_, _08130_);
  nor (_08134_, _08133_, _08127_);
  nor (_08135_, _05895_, _05870_);
  and (_08136_, _08135_, _08102_);
  and (_08137_, _08136_, _08109_);
  and (_08138_, _08098_, _08096_);
  and (_08139_, _05818_, _05870_);
  and (_08140_, _08139_, _08138_);
  nor (_08142_, _08140_, _08137_);
  nand (_08143_, _08142_, _08134_);
  or (_08144_, _08143_, _08124_);
  or (_08145_, _08119_, _08109_);
  and (_08146_, _08125_, _08097_);
  and (_08147_, _08146_, _08109_);
  and (_08149_, _08098_, _05895_);
  or (_08150_, _08149_, _08147_);
  and (_08151_, _08150_, _08145_);
  not (_08152_, _08109_);
  and (_08153_, _08110_, _08103_);
  and (_08154_, _08125_, _08135_);
  nor (_08155_, _08154_, _08153_);
  nor (_08156_, _08155_, _08152_);
  and (_08157_, _08108_, _08093_);
  and (_08158_, _08102_, _08112_);
  and (_08159_, _08158_, _08157_);
  and (_08160_, _08119_, _05767_);
  and (_08161_, _08160_, _08126_);
  or (_08162_, _08161_, _08159_);
  or (_08163_, _08162_, _08156_);
  and (_08164_, _08153_, _08120_);
  and (_08165_, _08102_, _08096_);
  and (_08166_, _08160_, _08165_);
  or (_08167_, _08166_, _08164_);
  and (_08168_, _08120_, _08114_);
  and (_08169_, _08102_, _05895_);
  and (_08170_, _05843_, _05870_);
  and (_08171_, _08170_, _08093_);
  or (_08172_, _08171_, _08139_);
  and (_08173_, _08172_, _08169_);
  or (_08174_, _08173_, _08168_);
  or (_08175_, _08174_, _08167_);
  or (_08176_, _08175_, _08163_);
  or (_08177_, _08176_, _08151_);
  or (_08178_, _08177_, _08144_);
  and (_08179_, _08178_, _05731_);
  and (_08180_, _05728_, _04859_);
  and (_08181_, _08180_, _05957_);
  nor (_08182_, _08181_, _05993_);
  or (_08183_, _08182_, rst);
  or (_05182_, _08183_, _08179_);
  and (_08184_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_08185_, _06626_, _05730_);
  or (_08186_, _08185_, _08184_);
  or (_08187_, _08186_, _06005_);
  and (_05200_, _08187_, _04856_);
  and (_08188_, _06410_, _05719_);
  and (_08189_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  or (_08190_, _08189_, _08188_);
  and (_05203_, _08190_, _04856_);
  and (_08191_, _06721_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_08192_, _05986_, _05950_);
  and (_08193_, _08192_, _05965_);
  or (_08194_, _06789_, _06628_);
  or (_08195_, _08194_, _06872_);
  or (_08196_, _08195_, _08193_);
  or (_08197_, _06786_, _06610_);
  and (_08198_, _06594_, _05848_);
  or (_08199_, _06613_, _08198_);
  or (_08200_, _06746_, _06726_);
  or (_08201_, _08200_, _08199_);
  or (_08202_, _08201_, _08197_);
  or (_08203_, _08202_, _08196_);
  and (_08204_, _08203_, _06770_);
  or (_05219_, _08204_, _08191_);
  and (_08205_, _06721_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_08206_, _06808_, _06806_);
  not (_08207_, _08206_);
  and (_08208_, _06777_, _05998_);
  and (_08209_, _06598_, _05986_);
  or (_08210_, _08209_, _08208_);
  or (_08211_, _08210_, _08207_);
  and (_08212_, _06783_, _05972_);
  and (_08213_, _06001_, _05983_);
  not (_08214_, _06858_);
  or (_08215_, _08214_, _08198_);
  or (_08216_, _08215_, _08213_);
  and (_08217_, _06855_, _06648_);
  not (_08218_, _08217_);
  or (_08219_, _08218_, _06614_);
  or (_08220_, _08219_, _08216_);
  or (_08221_, _08220_, _08212_);
  or (_08222_, _08221_, _08211_);
  and (_08223_, _08222_, _06770_);
  or (_05222_, _08223_, _08205_);
  and (_08224_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_08225_, _06686_, _06410_);
  or (_08226_, _08225_, _08224_);
  and (_05251_, _08226_, _04856_);
  and (_08228_, _05969_, _06637_);
  or (_08229_, _08228_, _05955_);
  or (_08231_, _06892_, _06790_);
  or (_08232_, _08231_, _08229_);
  or (_08233_, _06641_, _05980_);
  or (_08235_, _08233_, _06747_);
  or (_08236_, _08235_, _08232_);
  or (_08237_, _08236_, _06634_);
  and (_08238_, _08237_, _05730_);
  and (_08239_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_08240_, _08239_, _06650_);
  or (_08241_, _08240_, _08238_);
  and (_05302_, _08241_, _04856_);
  and (_08242_, _06822_, _06731_);
  and (_08243_, _06822_, _06637_);
  or (_08244_, _08243_, _08242_);
  and (_08245_, _06624_, _05965_);
  and (_08246_, _07510_, _06000_);
  or (_08247_, _08246_, _06833_);
  or (_08248_, _08247_, _08245_);
  or (_08249_, _08248_, _08244_);
  or (_08250_, _08047_, _06862_);
  or (_08251_, _08250_, _08249_);
  and (_08252_, _08251_, _05730_);
  and (_08253_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_08254_, _08253_, _06813_);
  or (_08255_, _08254_, _08252_);
  and (_05311_, _08255_, _04856_);
  and (_05358_, _05919_, _04856_);
  nor (_05361_, _07380_, rst);
  nor (_08256_, _05730_, _05323_);
  not (_08257_, _05730_);
  and (_08258_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_08259_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_08260_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_08261_, _08260_, _08259_);
  and (_08262_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_08263_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_08264_, _08263_, _08262_);
  and (_08265_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_08266_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_08267_, _08266_, _08265_);
  and (_08268_, _08267_, _08264_);
  and (_08269_, _08268_, _08261_);
  nor (_08270_, _08269_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_08271_, _08270_, _08258_);
  nor (_08272_, _08271_, _08257_);
  nor (_08273_, _08272_, _08256_);
  nor (_05364_, _08273_, rst);
  nor (_08274_, _04948_, _04922_);
  and (_08275_, _04932_, _05513_);
  and (_08276_, _08275_, _08274_);
  and (_08277_, _08276_, _06141_);
  and (_08278_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_08280_, _08278_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_08281_, _05627_, _05583_);
  and (_08282_, _05407_, _05455_);
  nand (_08284_, _05273_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_08285_, _08284_, _08278_);
  or (_08286_, _08285_, _08282_);
  or (_08287_, _08286_, _08281_);
  and (_08288_, _08287_, _08280_);
  or (_08289_, _08288_, _08277_);
  or (_08290_, _06146_, _06563_);
  nand (_08291_, _08290_, _08277_);
  or (_08292_, _08291_, _06147_);
  and (_08294_, _08292_, _08289_);
  or (_08295_, _08294_, _06934_);
  nand (_08296_, _06934_, _05287_);
  and (_08298_, _08296_, _04856_);
  and (_05505_, _08298_, _08295_);
  and (_05508_, _05767_, _04856_);
  and (_05511_, _05843_, _04856_);
  and (_05514_, _05793_, _04856_);
  and (_05516_, _05818_, _04856_);
  and (_05518_, _05870_, _04856_);
  and (_05521_, _05895_, _04856_);
  and (_05523_, _05943_, _04856_);
  and (_08304_, _08277_, _06091_);
  nand (_08305_, _08304_, _06088_);
  or (_08306_, _08304_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_08308_, _08306_, _06935_);
  and (_08309_, _08308_, _08305_);
  and (_08310_, _06934_, _05718_);
  or (_08311_, _08310_, _08309_);
  and (_05539_, _08311_, _04856_);
  nand (_08312_, _07897_, _06498_);
  not (_08313_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  nand (_08314_, _06497_, _08313_);
  and (_08315_, _08314_, _04856_);
  and (_05566_, _08315_, _08312_);
  nand (_08316_, _07815_, _06498_);
  or (_08317_, _06498_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_08318_, _08317_, _04856_);
  and (_05575_, _08318_, _08316_);
  or (_08319_, _07676_, _05293_);
  or (_08320_, _05524_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  nand (_08321_, _07702_, _05524_);
  and (_08322_, _08321_, _08320_);
  or (_08323_, _08322_, _05292_);
  and (_08324_, _08323_, _04856_);
  and (_05691_, _08324_, _08319_);
  or (_08325_, _07924_, _05293_);
  nor (_08326_, _07897_, _05643_);
  not (_08327_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  nor (_08328_, _05524_, _08327_);
  or (_08329_, _08328_, _05292_);
  or (_08330_, _08329_, _08326_);
  and (_08331_, _08330_, _04856_);
  and (_05695_, _08331_, _08325_);
  or (_08332_, _07853_, _05293_);
  nor (_08333_, _07815_, _05643_);
  and (_08334_, _05643_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_08335_, _08334_, _05292_);
  or (_08336_, _08335_, _08333_);
  and (_08337_, _08336_, _04856_);
  and (_05697_, _08337_, _08332_);
  or (_08338_, _07743_, _05293_);
  nor (_08339_, _07774_, _05643_);
  not (_08340_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  nor (_08341_, _05524_, _08340_);
  or (_08342_, _08341_, _05292_);
  or (_08343_, _08342_, _08339_);
  and (_08344_, _08343_, _04856_);
  and (_05706_, _08344_, _08338_);
  or (_08345_, _07640_, _05293_);
  nor (_08346_, _06586_, _05643_);
  not (_08347_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  nor (_08348_, _05524_, _08347_);
  or (_08349_, _08348_, _05292_);
  or (_08350_, _08349_, _08346_);
  and (_08351_, _08350_, _04856_);
  and (_05709_, _08351_, _08345_);
  or (_08352_, _07598_, _05293_);
  nor (_08353_, _06552_, _05643_);
  and (_08354_, _05643_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_08355_, _08354_, _05292_);
  or (_08356_, _08355_, _08353_);
  and (_08357_, _08356_, _04856_);
  and (_05712_, _08357_, _08352_);
  nor (_08358_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_08359_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08360_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _08359_);
  nor (_08361_, _08360_, _08358_);
  not (_08363_, \oc8051_symbolic_cxrom1.regvalid [13]);
  not (_08364_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_08365_, _05746_, _05736_);
  nor (_08366_, _08365_, _08257_);
  nor (_08367_, _08366_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_08368_, _08367_, _08364_);
  and (_08369_, _08368_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_08370_, _08368_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_08371_, _08370_, _08369_);
  nor (_08372_, _08371_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08373_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _08359_);
  nor (_08375_, _08373_, _08372_);
  and (_08376_, _08375_, _08363_);
  nor (_08377_, _08375_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08378_, _08377_, _08376_);
  not (_08380_, _08378_);
  nor (_08381_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08382_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _08359_);
  nor (_08383_, _08382_, _08381_);
  not (_08385_, _08383_);
  and (_08386_, _08367_, _08364_);
  nor (_08387_, _08386_, _08368_);
  nor (_08389_, _08387_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08390_, _08359_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor (_08392_, _08390_, _08389_);
  and (_08393_, _08392_, _08385_);
  nand (_08394_, _08393_, _08380_);
  and (_08396_, _08394_, _08361_);
  nor (_08397_, _08392_, _08385_);
  not (_08398_, _08397_);
  not (_08399_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_08401_, _08375_, _08399_);
  and (_08403_, _08375_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08404_, _08403_, _08401_);
  nor (_08405_, _08404_, _08398_);
  and (_08406_, _08392_, _08383_);
  not (_08407_, _08406_);
  not (_08408_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_08409_, _08375_, _08408_);
  nor (_08410_, _08375_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_08411_, _08410_, _08409_);
  nor (_08412_, _08411_, _08407_);
  nor (_08413_, _08412_, _08405_);
  not (_08414_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08415_, _08375_, _08414_);
  nor (_08416_, _08392_, _08383_);
  not (_08417_, _08416_);
  nor (_08418_, _08375_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08419_, _08418_, _08417_);
  or (_08420_, _08419_, _08415_);
  and (_08421_, _08420_, _08413_);
  and (_08422_, _08421_, _08396_);
  not (_08423_, _08392_);
  and (_08424_, _08375_, \oc8051_symbolic_cxrom1.regvalid [12]);
  not (_08425_, _08375_);
  and (_08426_, _08425_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_08427_, _08426_, _08424_);
  nor (_08428_, _08427_, _08423_);
  nor (_08429_, _08392_, _08375_);
  and (_08430_, _08429_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_08431_, _08423_, _08375_);
  and (_08432_, _08431_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_08433_, _08432_, _08430_);
  not (_08434_, _08433_);
  nor (_08435_, _08434_, _08428_);
  nor (_08436_, _08435_, _08383_);
  and (_08437_, _08429_, _08383_);
  and (_08438_, _08437_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not (_08439_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_08440_, _08375_, _08439_);
  nor (_08441_, _08375_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08442_, _08441_, _08440_);
  nor (_08443_, _08442_, _08407_);
  and (_08444_, _08375_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08445_, _08444_, _08397_);
  or (_08446_, _08445_, _08361_);
  or (_08447_, _08446_, _08443_);
  or (_08448_, _08447_, _08438_);
  nor (_08449_, _08448_, _08436_);
  nor (_08450_, _08449_, _08422_);
  not (_08451_, _08450_);
  and (_08452_, _08451_, word_in[7]);
  not (_08453_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_08454_, _08361_, _08453_);
  or (_08455_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_08456_, _08455_, _08454_);
  and (_08457_, _08456_, _08406_);
  not (_08458_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_08459_, _08361_, _08458_);
  or (_08460_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_08461_, _08460_, _08459_);
  and (_08462_, _08461_, _08397_);
  or (_08463_, _08462_, _08457_);
  not (_08464_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_08465_, _08361_, _08464_);
  or (_08466_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_08467_, _08466_, _08465_);
  and (_08468_, _08467_, _08393_);
  not (_08469_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_08470_, _08361_, _08469_);
  or (_08471_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_08472_, _08471_, _08470_);
  and (_08473_, _08472_, _08416_);
  or (_08474_, _08473_, _08468_);
  or (_08475_, _08474_, _08463_);
  and (_08476_, _08475_, _08375_);
  not (_08477_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_08478_, _08361_, _08477_);
  or (_08479_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_08480_, _08479_, _08478_);
  and (_08481_, _08480_, _08437_);
  and (_08482_, _08406_, _08425_);
  not (_08483_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_08484_, _08361_, _08483_);
  or (_08485_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_08486_, _08485_, _08484_);
  and (_08487_, _08486_, _08482_);
  not (_08488_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_08489_, _08361_, _08488_);
  or (_08490_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_08491_, _08490_, _08489_);
  and (_08493_, _08491_, _08393_);
  not (_08494_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_08495_, _08361_, _08494_);
  or (_08496_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_08498_, _08496_, _08495_);
  and (_08500_, _08498_, _08416_);
  or (_08502_, _08500_, _08493_);
  and (_08503_, _08502_, _08425_);
  or (_08505_, _08503_, _08487_);
  or (_08506_, _08505_, _08481_);
  or (_08507_, _08506_, _08476_);
  and (_08509_, _08507_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _08509_, _08452_);
  and (_08511_, _08385_, _08361_);
  not (_08512_, _08511_);
  and (_08514_, _08383_, _08361_);
  nor (_08515_, _08514_, _08392_);
  and (_08516_, _08514_, _08392_);
  nor (_08517_, _08516_, _08515_);
  not (_08518_, _08517_);
  nor (_08519_, _08518_, _08442_);
  nor (_08520_, _08516_, _08425_);
  and (_08521_, _08516_, _08425_);
  nor (_08522_, _08521_, _08520_);
  nor (_08523_, _08522_, _08517_);
  and (_08524_, _08523_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08525_, _08522_, _08518_);
  and (_08526_, _08525_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08527_, _08526_, _08524_);
  nor (_08528_, _08527_, _08519_);
  nor (_08529_, _08528_, _08512_);
  not (_08530_, _08529_);
  not (_08531_, _08514_);
  nor (_08532_, _08518_, _08427_);
  and (_08533_, _08525_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_08534_, _08533_, _08532_);
  or (_08535_, _08534_, _08531_);
  nand (_08536_, _08521_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08537_, _08536_, _08535_);
  and (_08538_, _08537_, _08530_);
  not (_08539_, _08361_);
  and (_08540_, _08383_, _08539_);
  not (_08541_, _08540_);
  nor (_08542_, _08518_, _08411_);
  and (_08543_, _08523_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08544_, _08525_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_08545_, _08544_, _08543_);
  nor (_08546_, _08545_, _08542_);
  nor (_08547_, _08546_, _08541_);
  nor (_08548_, _08383_, _08361_);
  not (_08549_, _08548_);
  nor (_08550_, _08518_, _08378_);
  and (_08551_, _08523_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08552_, _08525_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08553_, _08552_, _08551_);
  nor (_08554_, _08553_, _08550_);
  nor (_08555_, _08554_, _08549_);
  nor (_08556_, _08555_, _08547_);
  and (_08557_, _08556_, _08538_);
  or (_08558_, _08514_, _08548_);
  not (_08559_, _08558_);
  not (_08560_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_08561_, _08361_, _08560_);
  or (_08563_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_08564_, _08563_, _08561_);
  and (_08565_, _08564_, _08559_);
  not (_08566_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_08567_, _08361_, _08566_);
  or (_08568_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_08569_, _08568_, _08567_);
  and (_08570_, _08569_, _08558_);
  or (_08571_, _08570_, _08565_);
  and (_08572_, _08571_, _08523_);
  and (_08573_, _08517_, _08375_);
  not (_08574_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_08575_, _08361_, _08574_);
  or (_08576_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_08577_, _08576_, _08575_);
  and (_08578_, _08577_, _08559_);
  not (_08579_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_08580_, _08361_, _08579_);
  or (_08581_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_08583_, _08581_, _08580_);
  and (_08585_, _08583_, _08558_);
  or (_08586_, _08585_, _08578_);
  and (_08587_, _08586_, _08573_);
  or (_08588_, _08587_, _08572_);
  and (_08589_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_08590_, _08361_, _08494_);
  or (_08591_, _08590_, _08589_);
  and (_08592_, _08591_, _08558_);
  not (_08593_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_08594_, _08361_, _08593_);
  or (_08595_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_08596_, _08595_, _08594_);
  and (_08597_, _08596_, _08559_);
  or (_08598_, _08597_, _08592_);
  and (_08599_, _08598_, _08525_);
  and (_08600_, _08517_, _08425_);
  not (_08601_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_08602_, _08361_, _08601_);
  or (_08603_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_08604_, _08603_, _08602_);
  and (_08605_, _08604_, _08558_);
  not (_08606_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_08607_, _08361_, _08606_);
  or (_08608_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_08609_, _08608_, _08607_);
  and (_08610_, _08609_, _08559_);
  or (_08611_, _08610_, _08605_);
  and (_08612_, _08611_, _08600_);
  or (_08613_, _08612_, _08599_);
  nor (_08614_, _08613_, _08588_);
  nor (_08615_, _08614_, _08557_);
  and (_08616_, _08557_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _08616_, _08615_);
  nor (_08617_, _08406_, _08416_);
  and (_08618_, _08407_, _08375_);
  or (_08619_, _08618_, _08482_);
  nor (_08620_, _08619_, _08617_);
  and (_08621_, _08620_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not (_08622_, _08621_);
  not (_08623_, _08617_);
  nor (_08624_, _08623_, _08442_);
  and (_08625_, _08619_, _08623_);
  and (_08626_, _08625_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_08627_, _08626_, _08624_);
  and (_08628_, _08627_, _08622_);
  nor (_08629_, _08628_, _08549_);
  not (_08630_, _08629_);
  nor (_08631_, _08623_, _08427_);
  and (_08632_, _08620_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_08633_, _08632_, _08631_);
  or (_08634_, _08633_, _08541_);
  or (_08635_, _08375_, _08361_);
  nor (_08636_, _08635_, _08407_);
  nand (_08637_, _08636_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08638_, _08637_, _08634_);
  and (_08639_, _08638_, _08630_);
  nor (_08640_, _08623_, _08378_);
  and (_08641_, _08620_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_08642_, _08625_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_08643_, _08642_, _08641_);
  nor (_08644_, _08643_, _08640_);
  nor (_08645_, _08644_, _08531_);
  and (_08646_, _08620_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_08647_, _08646_);
  nor (_08648_, _08623_, _08411_);
  and (_08649_, _08625_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08650_, _08649_, _08648_);
  and (_08651_, _08650_, _08647_);
  nor (_08652_, _08651_, _08512_);
  nor (_08653_, _08652_, _08645_);
  and (_08654_, _08653_, _08639_);
  and (_08655_, _08486_, _08393_);
  and (_08656_, _08498_, _08375_);
  or (_08657_, _08656_, _08655_);
  and (_08658_, _08491_, _08397_);
  and (_08659_, _08480_, _08416_);
  or (_08660_, _08659_, _08658_);
  nor (_08661_, _08660_, _08657_);
  nor (_08662_, _08661_, _08619_);
  and (_08663_, _08467_, _08397_);
  and (_08664_, _08461_, _08416_);
  or (_08665_, _08664_, _08663_);
  and (_08666_, _08456_, _08393_);
  and (_08667_, _08472_, _08406_);
  or (_08668_, _08667_, _08666_);
  or (_08669_, _08668_, _08665_);
  and (_08670_, _08669_, _08619_);
  nor (_08671_, _08670_, _08662_);
  nor (_08672_, _08671_, _08654_);
  and (_08673_, _08654_, word_in[23]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _08673_, _08672_);
  and (_08674_, _08516_, _08375_);
  and (_08675_, _08674_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_08676_, _08549_, _08392_);
  nor (_08677_, _08549_, _08392_);
  nor (_08678_, _08677_, _08676_);
  not (_08679_, _08678_);
  nor (_08680_, _08442_, _08679_);
  and (_08681_, _08676_, _08375_);
  nor (_08682_, _08676_, _08375_);
  nor (_08684_, _08682_, _08681_);
  and (_08685_, _08684_, _08679_);
  and (_08686_, _08685_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_08687_, _08686_, _08680_);
  nor (_08688_, _08687_, _08531_);
  nor (_08689_, _08679_, _08427_);
  nor (_08690_, _08684_, _08678_);
  and (_08692_, _08690_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_08693_, _08685_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_08695_, _08693_, _08692_);
  nor (_08696_, _08695_, _08689_);
  nor (_08698_, _08696_, _08512_);
  or (_08699_, _08698_, _08688_);
  nor (_08700_, _08699_, _08675_);
  nor (_08701_, _08679_, _08378_);
  and (_08703_, _08685_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08704_, _08690_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08706_, _08704_, _08703_);
  nor (_08707_, _08706_, _08701_);
  nor (_08708_, _08707_, _08541_);
  nor (_08710_, _08679_, _08411_);
  and (_08711_, _08685_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08712_, _08711_, _08710_);
  nor (_08713_, _08712_, _08549_);
  and (_08714_, _08677_, _08401_);
  or (_08715_, _08714_, _08713_);
  nor (_08716_, _08715_, _08708_);
  and (_08717_, _08716_, _08700_);
  and (_08718_, _08569_, _08559_);
  and (_08719_, _08564_, _08558_);
  or (_08720_, _08719_, _08718_);
  and (_08721_, _08720_, _08685_);
  and (_08722_, _08591_, _08559_);
  and (_08723_, _08596_, _08558_);
  or (_08724_, _08723_, _08722_);
  and (_08725_, _08724_, _08690_);
  and (_08726_, _08678_, _08425_);
  and (_08727_, _08604_, _08559_);
  and (_08728_, _08609_, _08558_);
  or (_08729_, _08728_, _08727_);
  and (_08730_, _08729_, _08726_);
  and (_08731_, _08678_, _08375_);
  and (_08732_, _08583_, _08559_);
  and (_08733_, _08577_, _08558_);
  or (_08734_, _08733_, _08732_);
  and (_08735_, _08734_, _08731_);
  or (_08736_, _08735_, _08730_);
  or (_08737_, _08736_, _08725_);
  nor (_08738_, _08737_, _08721_);
  nor (_08739_, _08738_, _08717_);
  and (_08740_, _08717_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08740_, _08739_);
  and (_08741_, _08392_, _08375_);
  or (_08742_, _08741_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_05809_, _08742_, _04856_);
  and (_08743_, _08717_, _04856_);
  and (_08744_, _08743_, _08678_);
  and (_08745_, _08744_, _08684_);
  and (_08746_, _08745_, _08548_);
  and (_08747_, _08654_, _04856_);
  and (_08748_, _08747_, _08617_);
  and (_08749_, _08748_, _08619_);
  and (_08750_, _08749_, _08511_);
  and (_08751_, _08557_, _04856_);
  and (_08752_, _08751_, _08540_);
  and (_08753_, _08752_, _08573_);
  and (_08754_, _08422_, _04856_);
  and (_08755_, _08754_, _08383_);
  nor (_08756_, _08450_, rst);
  and (_08757_, _08756_, _08741_);
  and (_08758_, _08757_, _08755_);
  nor (_08759_, _08758_, _08453_);
  and (_08760_, _08756_, word_in[7]);
  and (_08761_, _08760_, _08758_);
  or (_08762_, _08761_, _08759_);
  or (_08763_, _08762_, _08753_);
  not (_08764_, word_in[15]);
  nand (_08765_, _08753_, _08764_);
  and (_08766_, _08765_, _08763_);
  or (_08767_, _08766_, _08750_);
  not (_08768_, _08750_);
  and (_08769_, _08747_, word_in[23]);
  or (_08770_, _08769_, _08768_);
  and (_08771_, _08770_, _08767_);
  or (_08772_, _08771_, _08746_);
  not (_08773_, _08746_);
  and (_08774_, _08743_, word_in[31]);
  or (_08775_, _08774_, _08773_);
  and (_13255_, _08775_, _08772_);
  or (_08776_, _08690_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_05859_, _08776_, _04856_);
  and (_08777_, _08690_, _08540_);
  and (_08778_, _08416_, _08425_);
  or (_08779_, _08778_, _08674_);
  or (_08780_, _08779_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08781_, _08780_, _08777_);
  and (_05887_, _08781_, _04856_);
  and (_08782_, _08726_, _08540_);
  or (_08783_, _08782_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08784_, _08779_, _08783_);
  and (_05931_, _08784_, _04856_);
  and (_08785_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  not (_08786_, _07390_);
  nand (_08787_, _08003_, _07958_);
  not (_08788_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_08789_, _07410_, _08788_);
  not (_08790_, _07404_);
  nand (_08791_, _08790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_08792_, _08791_, _08789_);
  nand (_08793_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  not (_08794_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_08795_, _07428_, _08794_);
  and (_08796_, _08795_, _08793_);
  and (_08797_, _08796_, _08792_);
  nand (_08798_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  nand (_08799_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_08800_, _08799_, _08798_);
  nand (_08801_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  nand (_08802_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_08803_, _08802_, _08801_);
  and (_08804_, _08803_, _08800_);
  and (_08805_, _08804_, _08797_);
  not (_08806_, _07463_);
  nand (_08807_, _08806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  not (_08808_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  or (_08809_, _07465_, _08808_);
  and (_08810_, _08809_, _08807_);
  nand (_08811_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  not (_08812_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_08813_, _07472_, _08812_);
  and (_08814_, _08813_, _08811_);
  and (_08815_, _08814_, _08810_);
  not (_08816_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_08817_, _07486_, _08816_);
  nand (_08818_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  and (_08819_, _08818_, _08817_);
  nand (_08820_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nand (_08821_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_08822_, _08821_, _08820_);
  and (_08823_, _08822_, _08819_);
  and (_08824_, _08823_, _08815_);
  and (_08825_, _08824_, _08805_);
  or (_08826_, _07503_, _07154_);
  nand (_08827_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_08828_, _08827_, _08826_);
  or (_08829_, _08025_, _06588_);
  or (_08830_, _07953_, _08347_);
  and (_08831_, _08830_, _08829_);
  and (_08832_, _08831_, _08828_);
  nor (_08833_, _07531_, p0_in[3]);
  not (_08834_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_08835_, _07531_, _08834_);
  nor (_08836_, _08835_, _08833_);
  nand (_08837_, _08836_, _07547_);
  nor (_08838_, _07531_, p1_in[3]);
  not (_08839_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_08840_, _07531_, _08839_);
  nor (_08841_, _08840_, _08838_);
  nand (_08842_, _08841_, _07552_);
  and (_08843_, _08842_, _08837_);
  nor (_08844_, _07531_, p2_in[3]);
  not (_08845_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_08846_, _07531_, _08845_);
  nor (_08847_, _08846_, _08844_);
  nand (_08848_, _08847_, _07507_);
  nor (_08849_, _07531_, p3_in[3]);
  not (_08850_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_08851_, _07531_, _08850_);
  nor (_08852_, _08851_, _08849_);
  nand (_08853_, _08852_, _07539_);
  and (_08854_, _08853_, _08848_);
  and (_08855_, _08854_, _08843_);
  and (_08856_, _08855_, _08832_);
  nand (_08857_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nand (_08858_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_08859_, _08858_, _08857_);
  and (_08860_, _08859_, _08856_);
  and (_08861_, _08860_, _08825_);
  or (_08862_, _08861_, _08787_);
  nand (_08863_, _08862_, _08786_);
  or (_08864_, _08863_, _08785_);
  nand (_08865_, _07390_, _06586_);
  and (_08866_, _08865_, _04856_);
  and (_05975_, _08866_, _08864_);
  or (_08867_, _08429_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_05981_, _08867_, _04856_);
  not (_08868_, _08429_);
  nor (_08869_, _08423_, _08375_);
  and (_08870_, _08869_, _08548_);
  or (_08871_, _08870_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_08872_, _08871_, _08868_);
  or (_08873_, _08512_, _08392_);
  nor (_08874_, _08873_, _08375_);
  and (_08875_, _08677_, _08426_);
  or (_08876_, _08875_, _08437_);
  or (_08877_, _08876_, _08874_);
  or (_08878_, _08877_, _08872_);
  and (_06031_, _08878_, _04856_);
  and (_08880_, _08514_, _08429_);
  or (_08882_, _08870_, _08880_);
  or (_08883_, _08406_, _08375_);
  or (_08884_, _08883_, _08882_);
  and (_08885_, _08884_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08886_, _08869_, _08511_);
  and (_08887_, _08782_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08888_, _08887_, _08886_);
  nor (_08889_, _08888_, _08885_);
  nor (_08890_, _08889_, _08682_);
  and (_08891_, _08778_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08892_, _08891_, _08782_);
  or (_08893_, _08892_, _08870_);
  or (_08894_, _08893_, _08880_);
  or (_08895_, _08894_, _08890_);
  and (_06085_, _08895_, _04856_);
  and (_08896_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_08897_, _08790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  not (_08898_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_08899_, _07410_, _08898_);
  or (_08900_, _08899_, _08897_);
  not (_08901_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  nor (_08902_, _07428_, _08901_);
  and (_08903_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_08904_, _08903_, _08902_);
  or (_08905_, _08904_, _08900_);
  and (_08906_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_08907_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_08908_, _08907_, _08906_);
  and (_08909_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_08910_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_08911_, _08910_, _08909_);
  or (_08912_, _08911_, _08908_);
  or (_08913_, _08912_, _08905_);
  and (_08914_, _08806_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_08915_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_08916_, _08915_, _08914_);
  and (_08917_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_08918_, _07473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_08919_, _08918_, _08917_);
  or (_08920_, _08919_, _08916_);
  and (_08921_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  not (_08922_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor (_08923_, _07486_, _08922_);
  or (_08924_, _08923_, _08921_);
  and (_08925_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_08926_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_08927_, _08926_, _08925_);
  or (_08928_, _08927_, _08924_);
  or (_08929_, _08928_, _08920_);
  or (_08930_, _08929_, _08913_);
  and (_08931_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_08932_, _08028_, _07102_);
  or (_08933_, _08932_, _08931_);
  and (_08934_, _07494_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  and (_08935_, _07389_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  or (_08936_, _08935_, _08934_);
  or (_08937_, _08936_, _08933_);
  or (_08938_, _07531_, p1_in[2]);
  or (_08939_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_08940_, _08939_, _08938_);
  and (_08941_, _08940_, _07552_);
  or (_08942_, _07531_, p0_in[2]);
  or (_08943_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_08944_, _08943_, _08942_);
  and (_08945_, _08944_, _07547_);
  or (_08946_, _08945_, _08941_);
  or (_08947_, _07531_, p3_in[2]);
  or (_08948_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_08949_, _08948_, _08947_);
  and (_08950_, _08949_, _07539_);
  or (_08951_, _07531_, p2_in[2]);
  or (_08952_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_08953_, _08952_, _08951_);
  and (_08954_, _08953_, _07507_);
  or (_08955_, _08954_, _08950_);
  or (_08956_, _08955_, _08946_);
  or (_08957_, _08956_, _08937_);
  and (_08958_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_08959_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_08960_, _08959_, _08958_);
  or (_08961_, _08960_, _08957_);
  or (_08962_, _08961_, _08930_);
  and (_08963_, _08962_, _08004_);
  or (_08964_, _08963_, _07390_);
  or (_08965_, _08964_, _08896_);
  nand (_08966_, _07390_, _06552_);
  and (_08967_, _08966_, _04856_);
  and (_06111_, _08967_, _08965_);
  and (_08968_, _08676_, _08425_);
  or (_08969_, _08520_, _08968_);
  and (_08970_, _08868_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08971_, _08970_, _08635_);
  or (_08972_, _08971_, _08636_);
  and (_08973_, _08972_, _08883_);
  and (_08974_, _08882_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08975_, _08974_, _08886_);
  or (_08976_, _08975_, _08973_);
  and (_08977_, _08976_, _08969_);
  or (_08978_, _08974_, _08972_);
  and (_08979_, _08978_, _08674_);
  and (_08980_, _08782_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08981_, _08778_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08982_, _08981_, _08880_);
  or (_08983_, _08982_, _08980_);
  or (_08984_, _08983_, _08870_);
  or (_08985_, _08984_, _08979_);
  or (_08986_, _08985_, _08977_);
  and (_06158_, _08986_, _04856_);
  and (_08987_, _06668_, _06132_);
  and (_08988_, _08987_, _04922_);
  and (_08989_, _08988_, _06268_);
  nand (_08990_, _08989_, _06088_);
  or (_08991_, _08989_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_08992_, _08991_, _06093_);
  and (_08993_, _08992_, _08990_);
  and (_08994_, _05517_, _05001_);
  nand (_08995_, _08994_, _06284_);
  or (_08996_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_08997_, _08996_, _05510_);
  and (_08998_, _08997_, _08995_);
  not (_08999_, _06092_);
  and (_09000_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_09001_, _09000_, rst);
  or (_09002_, _09001_, _08998_);
  or (_06167_, _09002_, _08993_);
  or (_09003_, _08516_, _08375_);
  and (_09004_, _08429_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_09005_, _08636_, _08375_);
  and (_09006_, _09005_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_09007_, _08385_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_09008_, _09007_, _08869_);
  or (_09009_, _09008_, _08521_);
  or (_09010_, _09009_, _09006_);
  or (_09011_, _09010_, _09004_);
  and (_09012_, _09011_, _09003_);
  or (_09013_, _09004_, _08870_);
  or (_09014_, _09013_, _08886_);
  or (_09015_, _09014_, _08636_);
  or (_09016_, _09015_, _09012_);
  and (_06239_, _09016_, _04856_);
  and (_09017_, _08987_, _06930_);
  and (_09018_, _09017_, _06268_);
  nand (_09019_, _09018_, _06088_);
  or (_09020_, _09018_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_09021_, _09020_, _06093_);
  and (_09022_, _09021_, _09019_);
  and (_09023_, _05515_, _04934_);
  and (_09024_, _09023_, _05001_);
  nand (_09025_, _09024_, _06284_);
  or (_09026_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_09027_, _09026_, _05510_);
  and (_09028_, _09027_, _09025_);
  and (_09029_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_09030_, _09029_, rst);
  or (_09031_, _09030_, _09028_);
  or (_06247_, _09031_, _09022_);
  nor (_09032_, _08726_, _08685_);
  and (_09033_, _09032_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_09034_, _08559_, _08869_);
  and (_09035_, _09034_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_09037_, _08677_, _08375_);
  and (_09038_, _08726_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_09039_, _09038_, _09037_);
  or (_09040_, _09039_, _09035_);
  or (_09041_, _09040_, _09033_);
  and (_09042_, _09041_, _08375_);
  and (_09043_, _08429_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_09044_, _08870_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_09045_, _08886_, _08521_);
  or (_09046_, _09045_, _09044_);
  or (_09047_, _09046_, _09043_);
  or (_09048_, _09047_, _08636_);
  or (_09049_, _09048_, _09042_);
  and (_06315_, _09049_, _04856_);
  not (_09050_, _08677_);
  and (_09051_, _08520_, _09050_);
  or (_09052_, _09051_, _08674_);
  nor (_09053_, _08873_, _08425_);
  and (_09054_, _08883_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_09055_, _09054_, _09053_);
  and (_09056_, _09055_, _09052_);
  or (_09057_, _08886_, _08726_);
  and (_09058_, _09057_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_09059_, _08635_, _08417_);
  and (_09060_, _09059_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_09061_, _09060_, _08636_);
  or (_09062_, _09061_, _09058_);
  or (_09063_, _09062_, _08521_);
  or (_09064_, _09063_, _09037_);
  or (_09065_, _09064_, _09056_);
  and (_06394_, _09065_, _04856_);
  and (_09066_, _06612_, _06731_);
  or (_09067_, _08208_, _09066_);
  and (_09068_, _06773_, _05998_);
  or (_09069_, _09068_, _06002_);
  or (_09070_, _06594_, _05949_);
  and (_09071_, _09070_, _05998_);
  or (_09072_, _09071_, _09069_);
  or (_09074_, _09072_, _09067_);
  and (_09075_, _06857_, _06731_);
  or (_09076_, _09075_, _05999_);
  or (_09077_, _09076_, _06783_);
  and (_09078_, _07510_, _06619_);
  or (_09079_, _09078_, _08243_);
  or (_09080_, _09079_, _07508_);
  or (_09081_, _09080_, _09077_);
  and (_09082_, _06635_, _05849_);
  and (_09083_, _06597_, _05998_);
  or (_09084_, _09083_, _09082_);
  or (_09085_, _09084_, _08245_);
  or (_09086_, _06759_, _06751_);
  or (_09087_, _09086_, _08250_);
  and (_09088_, _06737_, _06598_);
  and (_09089_, _06737_, _05998_);
  or (_09090_, _09089_, _09088_);
  and (_09091_, _06773_, _06606_);
  and (_09092_, _06620_, _05998_);
  or (_09093_, _09092_, _09091_);
  or (_09094_, _09093_, _09090_);
  or (_09095_, _09094_, _09087_);
  or (_09096_, _09095_, _09085_);
  and (_09097_, _08242_, _05972_);
  or (_09098_, _09097_, _05970_);
  or (_09099_, _08247_, _07513_);
  or (_09100_, _09099_, _09098_);
  or (_09101_, _09100_, _08229_);
  or (_09102_, _09101_, _05951_);
  or (_09103_, _09102_, _09096_);
  or (_09104_, _09103_, _09081_);
  or (_09105_, _09104_, _09074_);
  and (_09106_, _09105_, _05730_);
  and (_09107_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_09108_, _06003_, _05962_);
  not (_09109_, _06783_);
  nand (_09110_, _09109_, _06780_);
  and (_09111_, _09110_, _05995_);
  or (_09112_, _09111_, _09108_);
  or (_09113_, _09112_, _09107_);
  or (_09114_, _09113_, _09106_);
  and (_06447_, _09114_, _04856_);
  and (_06465_, _07612_, _04856_);
  and (_09115_, _05515_, _04947_);
  and (_09116_, _09115_, _06302_);
  and (_09117_, _09116_, _06268_);
  or (_09118_, _09117_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_09119_, _09118_, _06093_);
  nand (_09120_, _09117_, _06088_);
  and (_09121_, _09120_, _09119_);
  and (_09122_, _06302_, _05001_);
  and (_09123_, _09122_, _05515_);
  not (_09124_, _09123_);
  nor (_09125_, _09124_, _06284_);
  and (_09126_, _09124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_09127_, _09126_, _09125_);
  and (_09128_, _09127_, _05510_);
  and (_09129_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_09130_, _09129_, rst);
  or (_09131_, _09130_, _09128_);
  or (_06467_, _09131_, _09121_);
  and (_09132_, _09115_, _06273_);
  and (_09133_, _09132_, _06268_);
  nand (_09134_, _09133_, _06088_);
  or (_09135_, _09133_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_09136_, _09135_, _06093_);
  and (_09137_, _09136_, _09134_);
  and (_09138_, _06274_, _05001_);
  not (_09139_, _09138_);
  nor (_09140_, _09139_, _06284_);
  and (_09141_, _09139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_09142_, _09141_, _09140_);
  and (_09143_, _09142_, _05510_);
  and (_09144_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_09145_, _09144_, rst);
  or (_09146_, _09145_, _09143_);
  or (_06472_, _09146_, _09137_);
  and (_09147_, _08540_, _08731_);
  not (_09148_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_09149_, _08558_, _09148_);
  and (_09150_, _09149_, _08726_);
  or (_09151_, _09150_, _09147_);
  and (_09152_, _08600_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nand (_09153_, _08515_, _08873_);
  and (_09154_, _09153_, _08444_);
  or (_09155_, _09154_, _09152_);
  or (_09156_, _09155_, _09151_);
  or (_09157_, _08521_, _09037_);
  and (_09158_, _09157_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_09159_, _09059_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_09160_, _09159_, _09158_);
  or (_09161_, _09160_, _09156_);
  and (_09162_, _08520_, _08417_);
  and (_09164_, _09162_, _09161_);
  or (_09165_, _09158_, _09053_);
  or (_09166_, _09165_, _09164_);
  and (_09167_, _09166_, _09051_);
  and (_09168_, _09161_, _08674_);
  and (_09169_, _08617_, _08425_);
  and (_09170_, _09169_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_09171_, _08636_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_09172_, _08778_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_09173_, _09172_, _08521_);
  or (_09174_, _09173_, _09171_);
  or (_09175_, _09174_, _09037_);
  or (_09176_, _09175_, _09170_);
  or (_09177_, _09176_, _09168_);
  or (_09178_, _09177_, _09167_);
  and (_06484_, _09178_, _04856_);
  and (_09179_, _08514_, _08731_);
  and (_09180_, _08741_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_09181_, _09180_, _09179_);
  and (_09182_, _08559_, _08429_);
  or (_09183_, _09059_, _08521_);
  or (_09184_, _09183_, _09182_);
  and (_09185_, _09184_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_09186_, _08600_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_09187_, _09186_, _09037_);
  or (_09188_, _09187_, _09147_);
  or (_09189_, _09188_, _09185_);
  or (_09190_, _09189_, _09181_);
  or (_09191_, _09190_, _09053_);
  and (_06577_, _09191_, _04856_);
  not (_09193_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_09194_, _09052_, _09193_);
  and (_09195_, _08681_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_09196_, _09195_, _08731_);
  or (_09197_, _09196_, _09194_);
  and (_06683_, _09197_, _04856_);
  and (_09198_, _08619_, _08617_);
  or (_09199_, _09198_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_06785_, _09199_, _04856_);
  and (_09200_, _06301_, _05517_);
  or (_09201_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_09202_, _09201_, _04856_);
  not (_09203_, _09200_);
  or (_09204_, _09203_, _06705_);
  and (_06874_, _09204_, _09202_);
  and (_09205_, _05510_, _04987_);
  and (_09206_, _09205_, _09023_);
  and (_09207_, _09206_, _08060_);
  and (_09208_, _09207_, _06410_);
  and (_09209_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_09210_, _09209_, _08060_);
  and (_09211_, _08070_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_09212_, _09211_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_09213_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_09214_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  and (_09215_, _09214_, _09213_);
  and (_09216_, _09215_, _09212_);
  nor (_09217_, _09216_, _09210_);
  not (_09218_, _09217_);
  and (_09219_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_09220_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_09221_, _09220_, _09219_);
  nor (_09222_, _09221_, _09206_);
  and (_09223_, _09206_, _08070_);
  and (_09224_, _09223_, _05670_);
  or (_09225_, _09224_, _09222_);
  or (_09226_, _09225_, _09208_);
  and (_06881_, _09226_, _04856_);
  and (_09227_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nor (_09228_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_09229_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_09230_, _09229_, _09228_);
  nor (_09231_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_09232_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_09233_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_09234_, _09233_, _09232_);
  and (_09235_, _09234_, _09231_);
  and (_09236_, _09235_, _09230_);
  and (_09237_, _09236_, _09210_);
  or (_09238_, _09237_, _09217_);
  and (_09239_, _09238_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nor (_09240_, _09239_, _09227_);
  nor (_09241_, _09240_, _09206_);
  nor (_09242_, _08070_, _06369_);
  and (_09243_, _09242_, _09206_);
  or (_09244_, _09243_, _09241_);
  and (_06884_, _09244_, _04856_);
  or (_09245_, _08573_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_06896_, _09245_, _04856_);
  and (_09246_, _05719_, _05288_);
  and (_09247_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  or (_09248_, _09247_, _09246_);
  and (_06909_, _09248_, _04856_);
  not (_09249_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_09250_, _08072_, _08062_);
  or (_09251_, _09250_, _09249_);
  and (_09252_, _09251_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_09253_, _08062_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_09254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_09255_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_09256_, _09255_, _09254_);
  and (_09257_, _09256_, _09253_);
  or (_09258_, _09257_, _09252_);
  and (_06914_, _09258_, _04856_);
  and (_09259_, _06296_, _06132_);
  and (_09260_, _09259_, _06146_);
  nand (_09261_, _09260_, _06088_);
  or (_09262_, _09260_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_09263_, _09023_, _06126_);
  not (_09264_, _09263_);
  and (_09265_, _09264_, _09262_);
  and (_09266_, _09265_, _09261_);
  nor (_09267_, _09264_, _05287_);
  or (_09268_, _09267_, _09266_);
  and (_06927_, _09268_, _04856_);
  or (_09269_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  or (_09270_, _09269_, _09259_);
  not (_09271_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_09272_, _04986_, _09271_);
  nand (_09273_, _09272_, _09259_);
  or (_09274_, _09273_, _07713_);
  and (_09275_, _09274_, _09270_);
  or (_09276_, _09275_, _09263_);
  nand (_09277_, _09263_, _06032_);
  and (_09278_, _09277_, _04856_);
  and (_06933_, _09278_, _09276_);
  or (_09279_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_09280_, _09279_, _04856_);
  nand (_09281_, _09200_, _05669_);
  and (_06939_, _09281_, _09280_);
  not (_09282_, _06284_);
  and (_09283_, _09207_, _09282_);
  and (_09284_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_09285_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_09286_, _09285_, _09284_);
  nor (_09287_, _09286_, _09206_);
  and (_09288_, _09223_, _05288_);
  or (_09289_, _09288_, _09287_);
  or (_09290_, _09289_, _09283_);
  and (_06942_, _09290_, _04856_);
  nand (_09291_, _09223_, _06369_);
  nand (_09292_, _09207_, _06032_);
  and (_09293_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  and (_09294_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  or (_09295_, _09294_, _09293_);
  or (_09296_, _09295_, _09206_);
  and (_09297_, _09296_, _04856_);
  and (_09298_, _09297_, _09292_);
  and (_06945_, _09298_, _09291_);
  and (_09299_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_09300_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_06954_, _09300_, _09299_);
  or (_09301_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  or (_09302_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  and (_09303_, _09302_, _09301_);
  or (_09304_, _09303_, _09206_);
  and (_09305_, _09304_, _04856_);
  nand (_09306_, _09223_, _06284_);
  and (_06975_, _09306_, _09305_);
  or (_09307_, _06607_, _05999_);
  or (_09308_, _06636_, _06599_);
  or (_09309_, _09308_, _09307_);
  and (_09310_, _08228_, _05976_);
  or (_09311_, _09310_, _08245_);
  or (_09312_, _09088_, _06621_);
  or (_09313_, _09312_, _09311_);
  or (_09314_, _09313_, _09309_);
  and (_09315_, _06772_, _06831_);
  and (_09316_, _06598_, _06624_);
  or (_09317_, _06787_, _09316_);
  or (_09319_, _09317_, _09315_);
  or (_09320_, _09319_, _09099_);
  or (_09321_, _09079_, _06869_);
  or (_09322_, _09321_, _09087_);
  or (_09323_, _09322_, _09320_);
  or (_09324_, _09323_, _09314_);
  or (_09325_, _09324_, _09074_);
  and (_09326_, _09325_, _05730_);
  and (_09327_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_09328_, _09327_, _09112_);
  or (_09329_, _09328_, _09326_);
  and (_07107_, _09329_, _04856_);
  and (_09330_, _08751_, _08674_);
  not (_09331_, _09330_);
  not (_09332_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_09333_, _08756_, _08383_);
  not (_09334_, _09333_);
  not (_09335_, _08754_);
  and (_09336_, _08756_, _09335_);
  and (_09337_, _09336_, _09334_);
  and (_09338_, _09337_, _08429_);
  nor (_09339_, _09338_, _09332_);
  and (_09340_, _09338_, word_in[0]);
  or (_09341_, _09340_, _09339_);
  and (_09342_, _09341_, _09331_);
  and (_09343_, _09330_, word_in[8]);
  or (_09344_, _09343_, _09342_);
  nand (_09345_, _08747_, _08777_);
  and (_09346_, _09345_, _09344_);
  and (_09347_, _08511_, _08741_);
  and (_09348_, _09347_, _08743_);
  and (_09349_, _08747_, word_in[16]);
  and (_09350_, _09349_, _08777_);
  or (_09351_, _09350_, _09348_);
  or (_09352_, _09351_, _09346_);
  not (_09353_, _09348_);
  or (_09354_, _09353_, word_in[24]);
  and (_07298_, _09354_, _09352_);
  not (_09355_, _09338_);
  or (_09356_, _09355_, word_in[1]);
  or (_09357_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_09358_, _09357_, _09331_);
  and (_09359_, _09358_, _09356_);
  and (_09360_, _09330_, word_in[9]);
  nor (_09361_, _09360_, _09359_);
  nand (_09362_, _09361_, _09345_);
  or (_09363_, _09345_, word_in[17]);
  and (_09364_, _09363_, _09353_);
  and (_09365_, _09364_, _09362_);
  and (_09366_, _08743_, word_in[25]);
  and (_09367_, _09366_, _09348_);
  or (_07302_, _09367_, _09365_);
  and (_09368_, _08743_, word_in[26]);
  and (_09369_, _09368_, _09348_);
  or (_09370_, _09355_, word_in[2]);
  or (_09371_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_09372_, _09371_, _09331_);
  and (_09373_, _09372_, _09370_);
  and (_09374_, _09330_, word_in[10]);
  nor (_09375_, _09374_, _09373_);
  nand (_09376_, _09375_, _09345_);
  or (_09377_, _09345_, word_in[18]);
  and (_09378_, _09377_, _09353_);
  and (_09379_, _09378_, _09376_);
  or (_07307_, _09379_, _09369_);
  and (_09380_, _08743_, word_in[27]);
  and (_09381_, _09380_, _09348_);
  or (_09382_, _09355_, word_in[3]);
  or (_09383_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_09384_, _09383_, _09331_);
  and (_09385_, _09384_, _09382_);
  and (_09386_, _09330_, word_in[11]);
  nor (_09387_, _09386_, _09385_);
  nand (_09388_, _09387_, _09345_);
  or (_09389_, _09345_, word_in[19]);
  and (_09390_, _09389_, _09353_);
  and (_09391_, _09390_, _09388_);
  or (_07313_, _09391_, _09381_);
  or (_09392_, _09355_, word_in[4]);
  or (_09393_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_09394_, _09393_, _09331_);
  and (_09395_, _09394_, _09392_);
  and (_09396_, _09330_, word_in[12]);
  nor (_09397_, _09396_, _09395_);
  nand (_09398_, _09397_, _09345_);
  or (_09399_, _09345_, word_in[20]);
  and (_09400_, _09399_, _09353_);
  and (_09401_, _09400_, _09398_);
  and (_09402_, _08743_, word_in[28]);
  and (_09403_, _09402_, _09348_);
  or (_07318_, _09403_, _09401_);
  or (_09404_, _09355_, word_in[5]);
  or (_09405_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_09406_, _09405_, _09331_);
  and (_09407_, _09406_, _09404_);
  and (_09408_, _09330_, word_in[13]);
  nor (_09409_, _09408_, _09407_);
  nand (_09410_, _09409_, _09345_);
  or (_09411_, _09345_, word_in[21]);
  and (_09412_, _09411_, _09353_);
  and (_09413_, _09412_, _09410_);
  and (_09414_, _08743_, word_in[29]);
  and (_09415_, _09414_, _09348_);
  or (_07324_, _09415_, _09413_);
  or (_09416_, _09355_, word_in[6]);
  or (_09417_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_09418_, _09417_, _09331_);
  and (_09419_, _09418_, _09416_);
  and (_09420_, _09330_, word_in[14]);
  nor (_09421_, _09420_, _09419_);
  nand (_09422_, _09421_, _09345_);
  or (_09423_, _09345_, word_in[22]);
  and (_09424_, _09423_, _09353_);
  and (_09425_, _09424_, _09422_);
  and (_09426_, _08743_, word_in[30]);
  and (_09427_, _09426_, _09348_);
  or (_07329_, _09427_, _09425_);
  and (_09428_, _09348_, word_in[31]);
  or (_09429_, _09355_, word_in[7]);
  or (_09430_, _09338_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_09431_, _09430_, _09331_);
  and (_09432_, _09431_, _09429_);
  and (_09433_, _09330_, word_in[15]);
  nor (_09434_, _09433_, _09432_);
  nand (_09435_, _09434_, _09345_);
  or (_09436_, _09345_, word_in[23]);
  and (_09437_, _09436_, _09353_);
  and (_09438_, _09437_, _09435_);
  or (_07332_, _09438_, _09428_);
  and (_09439_, _08747_, _08514_);
  and (_09440_, _09439_, _08620_);
  and (_09441_, _08751_, _08548_);
  and (_09442_, _09441_, _08525_);
  not (_09443_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_09444_, _08756_, _08868_);
  and (_09445_, _08754_, _08385_);
  not (_09446_, _09445_);
  nor (_09447_, _09446_, _09444_);
  nor (_09448_, _09447_, _09443_);
  and (_09449_, _08756_, word_in[0]);
  and (_09450_, _09447_, _09449_);
  or (_09451_, _09450_, _09448_);
  or (_09452_, _09451_, _09442_);
  not (_09453_, _09442_);
  or (_09454_, _09453_, word_in[8]);
  and (_09455_, _09454_, _09452_);
  or (_09456_, _09455_, _09440_);
  and (_09457_, _08743_, _08777_);
  not (_09458_, _09457_);
  not (_09459_, _09440_);
  or (_09460_, _09459_, _09349_);
  and (_09461_, _09460_, _09458_);
  and (_09462_, _09461_, _09456_);
  and (_09463_, _09457_, word_in[24]);
  or (_07413_, _09463_, _09462_);
  and (_09464_, _08747_, word_in[17]);
  and (_09465_, _09440_, _09464_);
  and (_09466_, _08756_, word_in[1]);
  and (_09467_, _09447_, _09466_);
  not (_09468_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_09469_, _09447_, _09468_);
  nor (_09470_, _09469_, _09467_);
  nor (_09471_, _09470_, _09442_);
  and (_09472_, _09442_, word_in[9]);
  or (_09473_, _09472_, _09471_);
  and (_09474_, _09473_, _09459_);
  or (_09475_, _09474_, _09465_);
  and (_09476_, _09475_, _09458_);
  and (_09477_, _09457_, word_in[25]);
  or (_07416_, _09477_, _09476_);
  and (_09478_, _08747_, word_in[18]);
  and (_09479_, _09440_, _09478_);
  and (_09480_, _08756_, word_in[2]);
  and (_09481_, _09447_, _09480_);
  not (_09482_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_09483_, _09447_, _09482_);
  nor (_09484_, _09483_, _09481_);
  nor (_09485_, _09484_, _09442_);
  and (_09486_, _09442_, word_in[10]);
  or (_09487_, _09486_, _09485_);
  and (_09488_, _09487_, _09459_);
  or (_09489_, _09488_, _09479_);
  and (_09490_, _09489_, _09458_);
  and (_09491_, _09457_, word_in[26]);
  or (_07419_, _09491_, _09490_);
  and (_09493_, _08747_, word_in[19]);
  and (_09494_, _09440_, _09493_);
  and (_09495_, _08756_, word_in[3]);
  and (_09496_, _09447_, _09495_);
  not (_09497_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_09498_, _09447_, _09497_);
  nor (_09499_, _09498_, _09496_);
  nor (_09500_, _09499_, _09442_);
  and (_09501_, _09442_, word_in[11]);
  or (_09502_, _09501_, _09500_);
  and (_09503_, _09502_, _09459_);
  or (_09504_, _09503_, _09494_);
  and (_09505_, _09504_, _09458_);
  and (_09506_, _09457_, word_in[27]);
  or (_07421_, _09506_, _09505_);
  and (_09507_, _09457_, word_in[28]);
  not (_09508_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_09509_, _09447_, _09508_);
  and (_09510_, _08756_, word_in[4]);
  and (_09511_, _09447_, _09510_);
  or (_09512_, _09511_, _09509_);
  or (_09514_, _09512_, _09442_);
  or (_09515_, _09453_, word_in[12]);
  and (_09516_, _09515_, _09514_);
  or (_09517_, _09516_, _09440_);
  and (_09518_, _08747_, word_in[20]);
  or (_09519_, _09459_, _09518_);
  and (_09520_, _09519_, _09458_);
  and (_09522_, _09520_, _09517_);
  or (_07423_, _09522_, _09507_);
  and (_09523_, _08747_, word_in[21]);
  and (_09524_, _09440_, _09523_);
  and (_09525_, _08756_, word_in[5]);
  and (_09526_, _09447_, _09525_);
  not (_09527_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_09530_, _09447_, _09527_);
  nor (_09531_, _09530_, _09526_);
  nor (_09532_, _09531_, _09442_);
  and (_09533_, _09442_, word_in[13]);
  or (_09534_, _09533_, _09532_);
  and (_09535_, _09534_, _09459_);
  or (_09536_, _09535_, _09524_);
  and (_09537_, _09536_, _09458_);
  and (_09538_, _09457_, word_in[29]);
  or (_07427_, _09538_, _09537_);
  not (_09539_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_09540_, _09447_, _09539_);
  and (_09541_, _08756_, word_in[6]);
  and (_09542_, _09447_, _09541_);
  or (_09543_, _09542_, _09540_);
  or (_09544_, _09543_, _09442_);
  or (_09545_, _09453_, word_in[14]);
  and (_09546_, _09545_, _09544_);
  or (_09547_, _09546_, _09440_);
  and (_09548_, _08747_, word_in[22]);
  or (_09549_, _09459_, _09548_);
  and (_09550_, _09549_, _09458_);
  and (_09551_, _09550_, _09547_);
  and (_09552_, _09457_, word_in[30]);
  or (_07431_, _09552_, _09551_);
  and (_09553_, _09440_, _08769_);
  and (_09554_, _09447_, _08760_);
  nor (_09555_, _09447_, _08494_);
  or (_09556_, _09555_, _09554_);
  or (_09557_, _09556_, _09442_);
  nand (_09558_, _09442_, _08764_);
  and (_09559_, _09558_, _09459_);
  and (_09560_, _09559_, _09557_);
  or (_09561_, _09560_, _09553_);
  and (_09562_, _09561_, _09458_);
  and (_09563_, _09457_, word_in[31]);
  or (_07434_, _09563_, _09562_);
  and (_09564_, _08743_, _08674_);
  and (_09565_, _08747_, _08548_);
  and (_09566_, _09565_, _08620_);
  not (_09567_, _09566_);
  or (_09568_, _09567_, _09349_);
  and (_09569_, _08751_, _08511_);
  and (_09570_, _09569_, _08525_);
  not (_09571_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_09572_, _09333_, _09335_);
  and (_09573_, _09572_, _08429_);
  nor (_09574_, _09573_, _09571_);
  and (_09575_, _09573_, _09449_);
  or (_09576_, _09575_, _09574_);
  or (_09577_, _09576_, _09570_);
  not (_09578_, _09570_);
  or (_09579_, _09578_, word_in[8]);
  and (_09580_, _09579_, _09577_);
  or (_09581_, _09580_, _09566_);
  and (_09582_, _09581_, _09568_);
  or (_09583_, _09582_, _09564_);
  not (_09584_, _09564_);
  or (_09585_, _09584_, word_in[24]);
  and (_07517_, _09585_, _09583_);
  not (_09586_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_09587_, _09573_, _09586_);
  and (_09588_, _09573_, _09466_);
  or (_09589_, _09588_, _09587_);
  or (_09590_, _09589_, _09570_);
  or (_09591_, _09578_, word_in[9]);
  and (_09592_, _09591_, _09590_);
  or (_09593_, _09592_, _09566_);
  or (_09594_, _09567_, _09464_);
  and (_09595_, _09594_, _09584_);
  and (_09596_, _09595_, _09593_);
  and (_09597_, _09564_, word_in[25]);
  or (_07520_, _09597_, _09596_);
  or (_09598_, _09567_, _09478_);
  not (_09599_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_09600_, _09573_, _09599_);
  and (_09601_, _09573_, _09480_);
  or (_09602_, _09601_, _09600_);
  or (_09603_, _09602_, _09570_);
  or (_09604_, _09578_, word_in[10]);
  and (_09605_, _09604_, _09603_);
  or (_09606_, _09605_, _09566_);
  and (_09607_, _09606_, _09598_);
  or (_09608_, _09607_, _09564_);
  or (_09609_, _09584_, word_in[26]);
  and (_07524_, _09609_, _09608_);
  not (_09610_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_09611_, _09573_, _09610_);
  and (_09612_, _09573_, _09495_);
  or (_09613_, _09612_, _09611_);
  or (_09614_, _09613_, _09570_);
  or (_09615_, _09578_, word_in[11]);
  and (_09616_, _09615_, _09614_);
  or (_09617_, _09616_, _09566_);
  or (_09618_, _09567_, _09493_);
  and (_09619_, _09618_, _09584_);
  and (_09620_, _09619_, _09617_);
  and (_09621_, _09564_, word_in[27]);
  or (_07529_, _09621_, _09620_);
  not (_09622_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_09623_, _09573_, _09622_);
  and (_09624_, _09573_, _09510_);
  or (_09625_, _09624_, _09623_);
  or (_09626_, _09625_, _09570_);
  or (_09627_, _09578_, word_in[12]);
  and (_09628_, _09627_, _09626_);
  or (_09629_, _09628_, _09566_);
  or (_09630_, _09567_, _09518_);
  and (_09631_, _09630_, _09584_);
  and (_09632_, _09631_, _09629_);
  and (_09633_, _09564_, word_in[28]);
  or (_07534_, _09633_, _09632_);
  or (_09634_, _09567_, _09523_);
  not (_09635_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_09636_, _09573_, _09635_);
  and (_09637_, _09573_, _09525_);
  or (_09638_, _09637_, _09636_);
  or (_09639_, _09638_, _09570_);
  or (_09640_, _09578_, word_in[13]);
  and (_09641_, _09640_, _09639_);
  or (_09642_, _09641_, _09566_);
  and (_09643_, _09642_, _09634_);
  or (_09644_, _09643_, _09564_);
  or (_09645_, _09584_, word_in[29]);
  and (_07537_, _09645_, _09644_);
  or (_09646_, _09567_, _09548_);
  not (_09647_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_09648_, _09573_, _09647_);
  and (_09649_, _09573_, _09541_);
  or (_09650_, _09649_, _09648_);
  or (_09651_, _09650_, _09570_);
  or (_09652_, _09578_, word_in[14]);
  and (_09653_, _09652_, _09651_);
  or (_09654_, _09653_, _09566_);
  and (_09655_, _09654_, _09646_);
  or (_09656_, _09655_, _09564_);
  or (_09657_, _09584_, word_in[30]);
  and (_07540_, _09657_, _09656_);
  nor (_09658_, _09573_, _08593_);
  and (_09659_, _09573_, _08760_);
  or (_09660_, _09659_, _09658_);
  or (_09661_, _09660_, _09570_);
  nand (_09662_, _09570_, _08764_);
  and (_09663_, _09662_, _09661_);
  or (_09664_, _09663_, _09566_);
  or (_09665_, _09567_, _08769_);
  and (_09666_, _09665_, _09584_);
  and (_09667_, _09666_, _09664_);
  and (_09668_, _09564_, word_in[31]);
  or (_07543_, _09668_, _09667_);
  and (_09669_, _08747_, _08511_);
  and (_09670_, _09669_, _08620_);
  not (_09671_, _09670_);
  and (_09672_, _08752_, _08525_);
  not (_09673_, _08755_);
  nor (_09674_, _09444_, _09673_);
  and (_09675_, _09674_, _09449_);
  not (_09676_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  nor (_09677_, _09674_, _09676_);
  nor (_09678_, _09677_, _09675_);
  nor (_09679_, _09678_, _09672_);
  and (_09680_, _09672_, word_in[8]);
  or (_09681_, _09680_, _09679_);
  and (_09682_, _09681_, _09671_);
  and (_09683_, _08743_, _09059_);
  and (_09684_, _09670_, _09349_);
  or (_09685_, _09684_, _09683_);
  or (_09686_, _09685_, _09682_);
  not (_09687_, _09683_);
  or (_09688_, _09687_, word_in[24]);
  and (_07608_, _09688_, _09686_);
  and (_09689_, _09670_, _09464_);
  and (_09690_, _09674_, _09466_);
  not (_09691_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_09692_, _09674_, _09691_);
  nor (_09693_, _09692_, _09690_);
  nor (_09694_, _09693_, _09672_);
  and (_09695_, _09672_, word_in[9]);
  or (_09696_, _09695_, _09694_);
  and (_09697_, _09696_, _09671_);
  or (_09698_, _09697_, _09689_);
  and (_09699_, _09698_, _09687_);
  and (_09700_, _09683_, word_in[25]);
  or (_07611_, _09700_, _09699_);
  and (_09701_, _09683_, word_in[26]);
  not (_09702_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_09703_, _09674_, _09702_);
  and (_09704_, _09674_, _09480_);
  or (_09705_, _09704_, _09703_);
  or (_09706_, _09705_, _09672_);
  not (_09707_, _09672_);
  or (_09708_, _09707_, word_in[10]);
  and (_09709_, _09708_, _09706_);
  or (_09710_, _09709_, _09670_);
  or (_09711_, _09671_, _09478_);
  and (_09712_, _09711_, _09687_);
  and (_09713_, _09712_, _09710_);
  or (_07615_, _09713_, _09701_);
  and (_09714_, _09683_, word_in[27]);
  not (_09715_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_09716_, _09674_, _09715_);
  and (_09717_, _09674_, _09495_);
  or (_09718_, _09717_, _09716_);
  or (_09719_, _09718_, _09672_);
  or (_09720_, _09707_, word_in[11]);
  and (_09721_, _09720_, _09719_);
  or (_09722_, _09721_, _09670_);
  or (_09723_, _09671_, _09493_);
  and (_09724_, _09723_, _09687_);
  and (_09725_, _09724_, _09722_);
  or (_07618_, _09725_, _09714_);
  and (_09726_, _09670_, _09518_);
  and (_09727_, _09674_, _09510_);
  not (_09728_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_09729_, _09674_, _09728_);
  nor (_09730_, _09729_, _09727_);
  nor (_09731_, _09730_, _09672_);
  and (_09732_, _09672_, word_in[12]);
  or (_09733_, _09732_, _09731_);
  and (_09734_, _09733_, _09671_);
  or (_09735_, _09734_, _09726_);
  and (_09736_, _09735_, _09687_);
  and (_09737_, _09683_, word_in[28]);
  or (_07623_, _09737_, _09736_);
  and (_09738_, _09683_, word_in[29]);
  and (_09739_, _09674_, _09525_);
  not (_09740_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_09741_, _09674_, _09740_);
  nor (_09742_, _09741_, _09739_);
  nor (_09743_, _09742_, _09672_);
  and (_09744_, _09672_, word_in[13]);
  or (_09745_, _09744_, _09743_);
  or (_09746_, _09745_, _09670_);
  or (_09747_, _09671_, _09523_);
  and (_09748_, _09747_, _09687_);
  and (_09749_, _09748_, _09746_);
  or (_07627_, _09749_, _09738_);
  and (_09750_, _09683_, word_in[30]);
  and (_09751_, _09674_, _09541_);
  not (_09752_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_09753_, _09674_, _09752_);
  nor (_09754_, _09753_, _09751_);
  nor (_09755_, _09754_, _09672_);
  and (_09756_, _09672_, word_in[14]);
  or (_09757_, _09756_, _09755_);
  and (_09758_, _09757_, _09671_);
  and (_09759_, _09670_, _09548_);
  or (_09760_, _09759_, _09758_);
  and (_09761_, _09760_, _09687_);
  or (_07630_, _09761_, _09750_);
  and (_09762_, _09670_, _08769_);
  and (_09763_, _09674_, _08760_);
  nor (_09764_, _09674_, _08477_);
  or (_09765_, _09764_, _09763_);
  or (_09766_, _09765_, _09672_);
  nand (_09767_, _09672_, _08764_);
  and (_09768_, _09767_, _09671_);
  and (_09769_, _09768_, _09766_);
  or (_09770_, _09769_, _09762_);
  and (_09771_, _09770_, _09687_);
  and (_09772_, _09683_, word_in[31]);
  or (_07635_, _09772_, _09771_);
  not (_09773_, _08684_);
  and (_09774_, _08744_, _09773_);
  and (_09775_, _09774_, _08511_);
  not (_09776_, _09775_);
  not (_09777_, _08619_);
  and (_09778_, _08748_, _09777_);
  and (_09779_, _09778_, _08540_);
  and (_09780_, _09779_, _09349_);
  not (_09781_, _09779_);
  and (_09783_, _08751_, _08880_);
  not (_09784_, _09783_);
  nor (_09785_, _09333_, _08754_);
  and (_09786_, _08756_, _08869_);
  and (_09787_, _09786_, _09785_);
  and (_09789_, _09787_, word_in[0]);
  not (_09790_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_09792_, _09787_, _09790_);
  or (_09793_, _09792_, _09789_);
  and (_09795_, _09793_, _09784_);
  and (_09796_, _09783_, word_in[8]);
  or (_09797_, _09796_, _09795_);
  and (_09798_, _09797_, _09781_);
  or (_09799_, _09798_, _09780_);
  and (_09800_, _09799_, _09776_);
  and (_09801_, _08743_, word_in[24]);
  and (_09802_, _09775_, _09801_);
  or (_07728_, _09802_, _09800_);
  or (_09803_, _09784_, word_in[9]);
  not (_09804_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_09805_, _09787_, _09804_);
  and (_09807_, _09787_, word_in[1]);
  or (_09808_, _09807_, _09805_);
  or (_09809_, _09808_, _09783_);
  and (_09811_, _09809_, _09803_);
  or (_09812_, _09811_, _09779_);
  or (_09814_, _09781_, _09464_);
  and (_09815_, _09814_, _09812_);
  or (_09816_, _09815_, _09775_);
  or (_09817_, _09776_, _09366_);
  and (_07731_, _09817_, _09816_);
  not (_09818_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_09819_, _09787_, _09818_);
  and (_09821_, _09787_, word_in[2]);
  or (_09823_, _09821_, _09819_);
  and (_09824_, _09823_, _09784_);
  and (_09825_, _09783_, word_in[10]);
  or (_09826_, _09825_, _09824_);
  and (_09827_, _09826_, _09781_);
  and (_09828_, _09779_, _09478_);
  or (_09829_, _09828_, _09775_);
  or (_09830_, _09829_, _09827_);
  or (_09832_, _09776_, _09368_);
  and (_07734_, _09832_, _09830_);
  and (_09833_, _09779_, _09493_);
  not (_09834_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_09835_, _09787_, _09834_);
  and (_09836_, _09787_, word_in[3]);
  or (_09837_, _09836_, _09835_);
  and (_09838_, _09837_, _09784_);
  and (_09839_, _09783_, word_in[11]);
  or (_09840_, _09839_, _09838_);
  and (_09841_, _09840_, _09781_);
  or (_09842_, _09841_, _09833_);
  and (_09843_, _09842_, _09776_);
  and (_09844_, _09775_, _09380_);
  or (_07738_, _09844_, _09843_);
  and (_09845_, _09779_, _09518_);
  not (_09846_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_09847_, _09787_, _09846_);
  and (_09848_, _09787_, word_in[4]);
  or (_09849_, _09848_, _09847_);
  and (_09850_, _09849_, _09784_);
  and (_09851_, _09783_, word_in[12]);
  or (_09852_, _09851_, _09850_);
  and (_09853_, _09852_, _09781_);
  or (_09854_, _09853_, _09845_);
  and (_09855_, _09854_, _09776_);
  and (_09856_, _09775_, _09402_);
  or (_07742_, _09856_, _09855_);
  and (_09857_, _09779_, _09523_);
  not (_09858_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_09859_, _09787_, _09858_);
  and (_09860_, _09787_, word_in[5]);
  or (_09861_, _09860_, _09859_);
  and (_09862_, _09861_, _09784_);
  and (_09863_, _09783_, word_in[13]);
  or (_09864_, _09863_, _09862_);
  and (_09865_, _09864_, _09781_);
  or (_09866_, _09865_, _09857_);
  and (_09867_, _09866_, _09776_);
  and (_09868_, _09775_, _09414_);
  or (_07745_, _09868_, _09867_);
  and (_09869_, _09779_, _09548_);
  not (_09870_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_09871_, _09787_, _09870_);
  and (_09872_, _09787_, word_in[6]);
  or (_09873_, _09872_, _09871_);
  and (_09874_, _09873_, _09784_);
  and (_09875_, _09783_, word_in[14]);
  or (_09876_, _09875_, _09874_);
  and (_09877_, _09876_, _09781_);
  or (_09878_, _09877_, _09869_);
  and (_09879_, _09878_, _09776_);
  and (_09880_, _09775_, _09426_);
  or (_07747_, _09880_, _09879_);
  and (_09881_, _09779_, _08769_);
  nor (_09882_, _09787_, _08601_);
  and (_09883_, _09787_, word_in[7]);
  or (_09884_, _09883_, _09882_);
  and (_09885_, _09884_, _09784_);
  and (_09886_, _09783_, word_in[15]);
  or (_09887_, _09886_, _09885_);
  and (_09888_, _09887_, _09781_);
  or (_09889_, _09888_, _09881_);
  and (_09890_, _09889_, _09776_);
  and (_09891_, _09775_, _08774_);
  or (_07750_, _09891_, _09890_);
  and (_09892_, _09774_, _08540_);
  not (_09893_, _09892_);
  and (_09894_, _09778_, _08514_);
  and (_09895_, _09894_, _09349_);
  not (_09896_, _09894_);
  and (_09897_, _09441_, _08600_);
  and (_09898_, _09786_, _09445_);
  and (_09899_, _09898_, _09449_);
  not (_09900_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_09901_, _09898_, _09900_);
  nor (_09902_, _09901_, _09899_);
  nor (_09903_, _09902_, _09897_);
  and (_09904_, _09897_, word_in[8]);
  or (_09905_, _09904_, _09903_);
  and (_09906_, _09905_, _09896_);
  or (_09907_, _09906_, _09895_);
  and (_09908_, _09907_, _09893_);
  and (_09909_, _09892_, _09801_);
  or (_07827_, _09909_, _09908_);
  or (_09910_, _09896_, _09464_);
  not (_09911_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_09912_, _09898_, _09911_);
  and (_09913_, _09898_, _09466_);
  or (_09914_, _09913_, _09912_);
  or (_09915_, _09914_, _09897_);
  not (_09916_, _09897_);
  or (_09917_, _09916_, word_in[9]);
  and (_09918_, _09917_, _09915_);
  or (_09919_, _09918_, _09894_);
  and (_09920_, _09919_, _09910_);
  or (_09921_, _09920_, _09892_);
  or (_09922_, _09893_, _09366_);
  and (_07830_, _09922_, _09921_);
  and (_09923_, _09898_, _09480_);
  not (_09924_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_09925_, _09898_, _09924_);
  nor (_09926_, _09925_, _09923_);
  nor (_09927_, _09926_, _09897_);
  and (_09928_, _09897_, word_in[10]);
  or (_09929_, _09928_, _09927_);
  and (_09930_, _09929_, _09896_);
  and (_09931_, _09894_, _09478_);
  or (_09932_, _09931_, _09892_);
  or (_09933_, _09932_, _09930_);
  or (_09934_, _09893_, _09368_);
  and (_07834_, _09934_, _09933_);
  and (_09935_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  nor (_09936_, _06688_, _05669_);
  or (_09937_, _09936_, _09935_);
  and (_07837_, _09937_, _04856_);
  and (_09938_, _09898_, _09495_);
  not (_09939_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_09940_, _09898_, _09939_);
  nor (_09941_, _09940_, _09938_);
  nor (_09942_, _09941_, _09897_);
  and (_09943_, _09897_, word_in[11]);
  or (_09944_, _09943_, _09942_);
  and (_09945_, _09944_, _09896_);
  and (_09946_, _09894_, _09493_);
  or (_09947_, _09946_, _09945_);
  and (_09948_, _09947_, _09893_);
  and (_09949_, _09892_, _09380_);
  or (_07839_, _09949_, _09948_);
  or (_09950_, _05682_, _05676_);
  and (_09951_, _09950_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_09952_, _06997_, _05671_);
  or (_09953_, _05674_, _05679_);
  or (_09954_, _05675_, _09953_);
  and (_09955_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_09956_, _09955_, _09954_);
  or (_09957_, _09956_, _09952_);
  or (_09958_, _09957_, _09951_);
  and (_07842_, _09958_, _04856_);
  and (_09959_, _09894_, _09518_);
  and (_09960_, _09898_, _09510_);
  not (_09961_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_09962_, _09898_, _09961_);
  nor (_09963_, _09962_, _09960_);
  nor (_09964_, _09963_, _09897_);
  and (_09965_, _09897_, word_in[12]);
  or (_09966_, _09965_, _09964_);
  and (_09967_, _09966_, _09896_);
  or (_09968_, _09967_, _09959_);
  and (_09969_, _09968_, _09893_);
  and (_09970_, _09892_, _09402_);
  or (_07844_, _09970_, _09969_);
  not (_09971_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_09972_, _09898_, _09971_);
  and (_09973_, _09898_, _09525_);
  or (_09974_, _09973_, _09972_);
  or (_09975_, _09974_, _09897_);
  or (_09976_, _09916_, word_in[13]);
  and (_09977_, _09976_, _09975_);
  or (_09978_, _09977_, _09894_);
  or (_09979_, _09896_, _09523_);
  and (_09980_, _09979_, _09978_);
  or (_09981_, _09980_, _09892_);
  or (_09982_, _09893_, _09414_);
  and (_07849_, _09982_, _09981_);
  not (_09983_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_09985_, _09898_, _09983_);
  and (_09986_, _09898_, _09541_);
  or (_09987_, _09986_, _09985_);
  or (_09988_, _09987_, _09897_);
  or (_09989_, _09916_, word_in[14]);
  and (_09990_, _09989_, _09988_);
  and (_09991_, _09990_, _09896_);
  and (_09992_, _09894_, _09548_);
  or (_09993_, _09992_, _09892_);
  or (_09994_, _09993_, _09991_);
  or (_09995_, _09893_, _09426_);
  and (_07852_, _09995_, _09994_);
  and (_09997_, _09894_, _08769_);
  and (_09998_, _09898_, _08760_);
  nor (_09999_, _09898_, _08488_);
  nor (_10000_, _09999_, _09998_);
  nor (_10001_, _10000_, _09897_);
  and (_10002_, _09897_, word_in[15]);
  or (_10003_, _10002_, _10001_);
  and (_10004_, _10003_, _09896_);
  or (_10005_, _10004_, _09997_);
  and (_10006_, _10005_, _09893_);
  and (_10007_, _09892_, _08774_);
  or (_07856_, _10007_, _10006_);
  and (_10008_, _09774_, _08514_);
  not (_10009_, _10008_);
  and (_10010_, _09778_, _08548_);
  and (_10011_, _10010_, _09349_);
  not (_10012_, _10010_);
  and (_10013_, _09569_, _08600_);
  and (_10014_, _09572_, _08869_);
  and (_10015_, _10014_, word_in[0]);
  not (_10016_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor (_10017_, _10014_, _10016_);
  nor (_10018_, _10017_, _10015_);
  nor (_10019_, _10018_, _10013_);
  and (_10020_, _10013_, word_in[8]);
  or (_10021_, _10020_, _10019_);
  and (_10022_, _10021_, _10012_);
  or (_10023_, _10022_, _10011_);
  and (_10024_, _10023_, _10009_);
  and (_10025_, _10008_, _09801_);
  or (_07923_, _10025_, _10024_);
  not (_10026_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_10027_, _10014_, _10026_);
  and (_10028_, _10014_, word_in[1]);
  or (_10029_, _10028_, _10027_);
  or (_10030_, _10029_, _10013_);
  not (_10031_, _10013_);
  or (_10032_, _10031_, word_in[9]);
  and (_10033_, _10032_, _10030_);
  or (_10034_, _10033_, _10010_);
  or (_10035_, _10012_, _09464_);
  and (_10036_, _10035_, _10009_);
  and (_10037_, _10036_, _10034_);
  and (_10038_, _10008_, _09366_);
  or (_07926_, _10038_, _10037_);
  and (_10039_, _10010_, _09478_);
  not (_10040_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_10041_, _10014_, _10040_);
  and (_10042_, _10014_, word_in[2]);
  nor (_10043_, _10042_, _10041_);
  nor (_10044_, _10043_, _10013_);
  and (_10045_, _10013_, word_in[10]);
  or (_10046_, _10045_, _10044_);
  and (_10048_, _10046_, _10012_);
  or (_10049_, _10048_, _10039_);
  and (_10050_, _10049_, _10009_);
  and (_10051_, _10008_, _09368_);
  or (_07930_, _10051_, _10050_);
  or (_10052_, _10031_, word_in[11]);
  not (_10053_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_10054_, _10014_, _10053_);
  and (_10055_, _10014_, word_in[3]);
  or (_10056_, _10055_, _10054_);
  or (_10057_, _10056_, _10013_);
  and (_10058_, _10057_, _10052_);
  or (_10059_, _10058_, _10010_);
  or (_10061_, _10012_, _09493_);
  and (_10062_, _10061_, _10059_);
  or (_10063_, _10062_, _10008_);
  or (_10064_, _10009_, _09380_);
  and (_07934_, _10064_, _10063_);
  and (_10065_, _10010_, _09518_);
  not (_10066_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_10068_, _10014_, _10066_);
  and (_10069_, _10014_, word_in[4]);
  nor (_10070_, _10069_, _10068_);
  nor (_10071_, _10070_, _10013_);
  and (_10073_, _10013_, word_in[12]);
  or (_10074_, _10073_, _10071_);
  and (_10075_, _10074_, _10012_);
  or (_10076_, _10075_, _10065_);
  and (_10077_, _10076_, _10009_);
  and (_10078_, _10008_, _09402_);
  or (_07938_, _10078_, _10077_);
  and (_10079_, _10010_, _09523_);
  not (_10080_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_10081_, _10014_, _10080_);
  and (_10082_, _10014_, word_in[5]);
  nor (_10083_, _10082_, _10081_);
  nor (_10084_, _10083_, _10013_);
  and (_10085_, _10013_, word_in[13]);
  or (_10086_, _10085_, _10084_);
  and (_10087_, _10086_, _10012_);
  or (_10088_, _10087_, _10079_);
  and (_10089_, _10088_, _10009_);
  and (_10090_, _10008_, _09414_);
  or (_07941_, _10090_, _10089_);
  and (_10091_, _10010_, _09548_);
  not (_10092_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_10093_, _10014_, _10092_);
  and (_10094_, _10014_, word_in[6]);
  nor (_10095_, _10094_, _10093_);
  nor (_10096_, _10095_, _10013_);
  and (_10097_, _10013_, word_in[14]);
  or (_10098_, _10097_, _10096_);
  and (_10099_, _10098_, _10012_);
  or (_10100_, _10099_, _10091_);
  and (_10101_, _10100_, _10009_);
  and (_10102_, _10008_, _09426_);
  or (_07946_, _10102_, _10101_);
  and (_10103_, _10010_, _08769_);
  nor (_10104_, _10014_, _08606_);
  and (_10105_, _10014_, word_in[7]);
  nor (_10106_, _10105_, _10104_);
  nor (_10107_, _10106_, _10013_);
  and (_10108_, _10013_, word_in[15]);
  or (_10109_, _10108_, _10107_);
  and (_10110_, _10109_, _10012_);
  or (_10111_, _10110_, _10103_);
  and (_10112_, _10111_, _10009_);
  and (_10113_, _10008_, _08774_);
  or (_07950_, _10113_, _10112_);
  and (_10115_, _09774_, _08548_);
  not (_10116_, _10115_);
  and (_10117_, _09778_, _08511_);
  and (_10118_, _10117_, _09349_);
  not (_10119_, _10117_);
  and (_10120_, _08752_, _08600_);
  and (_10121_, _09786_, _08755_);
  and (_10122_, _10121_, word_in[0]);
  not (_10123_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor (_10124_, _10121_, _10123_);
  nor (_10125_, _10124_, _10122_);
  nor (_10126_, _10125_, _10120_);
  and (_10127_, _10120_, word_in[8]);
  or (_10128_, _10127_, _10126_);
  and (_10129_, _10128_, _10119_);
  or (_10130_, _10129_, _10118_);
  and (_10131_, _10130_, _10116_);
  and (_10132_, _10115_, _09801_);
  or (_08020_, _10132_, _10131_);
  and (_10133_, _10121_, word_in[1]);
  not (_10134_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_10136_, _10121_, _10134_);
  nor (_10137_, _10136_, _10133_);
  nor (_10138_, _10137_, _10120_);
  and (_10139_, _10120_, word_in[9]);
  or (_10140_, _10139_, _10138_);
  and (_10141_, _10140_, _10119_);
  and (_10142_, _10117_, _09464_);
  or (_10144_, _10142_, _10141_);
  and (_10145_, _10144_, _10116_);
  and (_10147_, _10115_, _09366_);
  or (_08023_, _10147_, _10145_);
  and (_10148_, _10121_, word_in[2]);
  not (_10149_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_10150_, _10121_, _10149_);
  nor (_10151_, _10150_, _10148_);
  nor (_10152_, _10151_, _10120_);
  and (_10153_, _10120_, word_in[10]);
  or (_10154_, _10153_, _10152_);
  and (_10155_, _10154_, _10119_);
  and (_10156_, _10117_, _09478_);
  or (_10157_, _10156_, _10155_);
  and (_10158_, _10157_, _10116_);
  and (_10159_, _10115_, _09368_);
  or (_08026_, _10159_, _10158_);
  not (_10160_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_10161_, _10121_, _10160_);
  and (_10163_, _10121_, _09495_);
  or (_10164_, _10163_, _10161_);
  or (_10165_, _10164_, _10120_);
  not (_10166_, _10120_);
  or (_10167_, _10166_, word_in[11]);
  and (_10168_, _10167_, _10165_);
  or (_10169_, _10168_, _10117_);
  or (_10170_, _10119_, _09493_);
  and (_10171_, _10170_, _10169_);
  or (_10172_, _10171_, _10115_);
  or (_10173_, _10116_, _09380_);
  and (_08030_, _10173_, _10172_);
  not (_10175_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_10176_, _10121_, _10175_);
  and (_10177_, _10121_, _09510_);
  or (_10178_, _10177_, _10176_);
  or (_10179_, _10178_, _10120_);
  or (_10180_, _10166_, word_in[12]);
  and (_10181_, _10180_, _10179_);
  or (_10182_, _10181_, _10117_);
  or (_10183_, _10119_, _09518_);
  and (_10184_, _10183_, _10182_);
  or (_10185_, _10184_, _10115_);
  or (_10186_, _10116_, _09402_);
  and (_08035_, _10186_, _10185_);
  not (_10187_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_10188_, _10121_, _10187_);
  and (_10189_, _10121_, _09525_);
  or (_10191_, _10189_, _10188_);
  or (_10192_, _10191_, _10120_);
  or (_10194_, _10166_, word_in[13]);
  and (_10195_, _10194_, _10192_);
  or (_10196_, _10195_, _10117_);
  or (_10197_, _10119_, _09523_);
  and (_10198_, _10197_, _10196_);
  or (_10200_, _10198_, _10115_);
  or (_10201_, _10116_, _09414_);
  and (_08039_, _10201_, _10200_);
  not (_10203_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_10204_, _10121_, _10203_);
  and (_10205_, _10121_, _09541_);
  or (_10206_, _10205_, _10204_);
  or (_10207_, _10206_, _10120_);
  or (_10209_, _10166_, word_in[14]);
  and (_10210_, _10209_, _10207_);
  or (_10211_, _10210_, _10117_);
  or (_10212_, _10119_, _09548_);
  and (_10213_, _10212_, _10211_);
  or (_10215_, _10213_, _10115_);
  or (_10216_, _10116_, _09426_);
  and (_08042_, _10216_, _10215_);
  nor (_10218_, _10121_, _08483_);
  and (_10219_, _10121_, _08760_);
  or (_10220_, _10219_, _10218_);
  or (_10222_, _10220_, _10120_);
  nand (_10223_, _10120_, _08764_);
  and (_10224_, _10223_, _10222_);
  or (_10225_, _10224_, _10117_);
  or (_10226_, _10119_, _08769_);
  and (_10227_, _10226_, _10225_);
  or (_10228_, _10227_, _10115_);
  or (_10229_, _10116_, _08774_);
  and (_08045_, _10229_, _10228_);
  nor (_10230_, _08076_, _08072_);
  nor (_10231_, _10230_, _08062_);
  not (_10232_, _08087_);
  or (_10233_, _10232_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_10234_, _10233_, _10231_);
  or (_10235_, _08087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_10236_, _10235_, _08085_);
  and (_10237_, _10236_, _10234_);
  or (_08118_, _10237_, _09299_);
  and (_10238_, _08743_, _08685_);
  and (_10239_, _10238_, _08511_);
  not (_10240_, _10239_);
  and (_10241_, _08747_, _08636_);
  and (_10242_, _10241_, word_in[16]);
  not (_10243_, _10241_);
  and (_10244_, _08751_, _08521_);
  not (_10245_, _10244_);
  not (_10246_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_10248_, _08756_, _08431_);
  and (_10249_, _10248_, _09785_);
  nor (_10251_, _10249_, _10246_);
  and (_10252_, _10249_, word_in[0]);
  or (_10253_, _10252_, _10251_);
  and (_10254_, _10253_, _10245_);
  and (_10255_, _10244_, word_in[8]);
  or (_10256_, _10255_, _10254_);
  and (_10258_, _10256_, _10243_);
  or (_10259_, _10258_, _10242_);
  and (_10260_, _10259_, _10240_);
  and (_10261_, _10239_, word_in[24]);
  or (_08129_, _10261_, _10260_);
  and (_10262_, _10241_, word_in[17]);
  not (_10263_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_10264_, _10249_, _10263_);
  and (_10266_, _10249_, word_in[1]);
  or (_10267_, _10266_, _10264_);
  and (_10268_, _10267_, _10245_);
  and (_10269_, _10244_, word_in[9]);
  or (_10270_, _10269_, _10268_);
  and (_10271_, _10270_, _10243_);
  or (_10272_, _10271_, _10262_);
  and (_10273_, _10272_, _10240_);
  and (_10274_, _10239_, word_in[25]);
  or (_13256_, _10274_, _10273_);
  and (_10275_, _10241_, word_in[18]);
  not (_10276_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_10277_, _10249_, _10276_);
  and (_10278_, _10249_, word_in[2]);
  or (_10279_, _10278_, _10277_);
  and (_10280_, _10279_, _10245_);
  and (_10281_, _10244_, word_in[10]);
  or (_10282_, _10281_, _10280_);
  and (_10283_, _10282_, _10243_);
  or (_10284_, _10283_, _10275_);
  and (_10285_, _10284_, _10240_);
  and (_10286_, _10239_, word_in[26]);
  or (_13257_, _10286_, _10285_);
  and (_10287_, _10241_, word_in[19]);
  not (_10288_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_10289_, _10249_, _10288_);
  and (_10290_, _10249_, word_in[3]);
  or (_10291_, _10290_, _10289_);
  and (_10292_, _10291_, _10245_);
  and (_10293_, _10244_, word_in[11]);
  or (_10294_, _10293_, _10292_);
  and (_10295_, _10294_, _10243_);
  or (_10296_, _10295_, _10287_);
  and (_10298_, _10296_, _10240_);
  and (_10299_, _10239_, word_in[27]);
  or (_08141_, _10299_, _10298_);
  and (_10300_, _10241_, word_in[20]);
  not (_10302_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_10303_, _10249_, _10302_);
  and (_10304_, _10249_, word_in[4]);
  or (_10305_, _10304_, _10303_);
  and (_10306_, _10305_, _10245_);
  and (_10307_, _10244_, word_in[12]);
  or (_10308_, _10307_, _10306_);
  and (_10309_, _10308_, _10243_);
  or (_10311_, _10309_, _10300_);
  and (_10312_, _10311_, _10240_);
  and (_10313_, _10239_, word_in[28]);
  or (_13258_, _10313_, _10312_);
  and (_10314_, _10241_, word_in[21]);
  not (_10315_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_10316_, _10249_, _10315_);
  and (_10317_, _10249_, word_in[5]);
  or (_10319_, _10317_, _10316_);
  and (_10320_, _10319_, _10245_);
  and (_10321_, _10244_, word_in[13]);
  or (_10322_, _10321_, _10320_);
  and (_10323_, _10322_, _10243_);
  or (_10324_, _10323_, _10314_);
  and (_10325_, _10324_, _10240_);
  and (_10326_, _10239_, word_in[29]);
  or (_13259_, _10326_, _10325_);
  and (_10327_, _10241_, word_in[22]);
  not (_10328_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_10329_, _10249_, _10328_);
  and (_10330_, _10249_, word_in[6]);
  or (_10331_, _10330_, _10329_);
  and (_10332_, _10331_, _10245_);
  and (_10333_, _10244_, word_in[14]);
  or (_10334_, _10333_, _10332_);
  and (_10335_, _10334_, _10243_);
  or (_10336_, _10335_, _10327_);
  and (_10338_, _10336_, _10240_);
  and (_10340_, _10239_, word_in[30]);
  or (_08148_, _10340_, _10338_);
  and (_10341_, _10241_, word_in[23]);
  nor (_10342_, _10249_, _08566_);
  and (_10343_, _10249_, word_in[7]);
  or (_10345_, _10343_, _10342_);
  and (_10346_, _10345_, _10245_);
  and (_10347_, _10244_, word_in[15]);
  or (_10348_, _10347_, _10346_);
  and (_10349_, _10348_, _10243_);
  or (_10350_, _10349_, _10341_);
  and (_10351_, _10350_, _10240_);
  and (_10352_, _10239_, word_in[31]);
  or (_13260_, _10352_, _10351_);
  and (_10353_, _08743_, _08636_);
  and (_10354_, _10353_, word_in[24]);
  and (_10355_, _09439_, _08625_);
  and (_10356_, _09441_, _08523_);
  not (_10357_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_10358_, _10248_, _09445_);
  nor (_10359_, _10358_, _10357_);
  and (_10360_, _10358_, _09449_);
  or (_10361_, _10360_, _10359_);
  or (_10362_, _10361_, _10356_);
  not (_10363_, _10356_);
  or (_10364_, _10363_, word_in[8]);
  and (_10365_, _10364_, _10362_);
  or (_10366_, _10365_, _10355_);
  not (_10367_, _10353_);
  not (_10368_, _10355_);
  or (_10369_, _10368_, _09349_);
  and (_10370_, _10369_, _10367_);
  and (_10371_, _10370_, _10366_);
  or (_13261_, _10371_, _10354_);
  or (_10372_, _10368_, _09464_);
  not (_10373_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_10375_, _10358_, _10373_);
  and (_10376_, _10358_, _09466_);
  or (_10377_, _10376_, _10375_);
  or (_10378_, _10377_, _10356_);
  or (_10379_, _10363_, word_in[9]);
  and (_10380_, _10379_, _10378_);
  or (_10381_, _10380_, _10355_);
  and (_10382_, _10381_, _10372_);
  or (_10383_, _10382_, _10353_);
  or (_10384_, _10367_, word_in[25]);
  and (_13262_, _10384_, _10383_);
  and (_10385_, _10358_, _09480_);
  not (_10386_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_10387_, _10358_, _10386_);
  nor (_10388_, _10387_, _10385_);
  nor (_10389_, _10388_, _10356_);
  and (_10390_, _10356_, word_in[10]);
  or (_10391_, _10390_, _10389_);
  and (_10392_, _10391_, _10368_);
  and (_10393_, _10355_, _09478_);
  or (_10394_, _10393_, _10353_);
  or (_10395_, _10394_, _10392_);
  or (_10396_, _10367_, word_in[26]);
  and (_13263_, _10396_, _10395_);
  and (_10397_, _10358_, _09495_);
  not (_10398_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_10399_, _10358_, _10398_);
  nor (_10400_, _10399_, _10397_);
  nor (_10401_, _10400_, _10356_);
  and (_10402_, _10356_, word_in[11]);
  or (_10403_, _10402_, _10401_);
  and (_10404_, _10403_, _10368_);
  and (_10405_, _10355_, _09493_);
  or (_10406_, _10405_, _10353_);
  or (_10407_, _10406_, _10404_);
  or (_10408_, _10367_, word_in[27]);
  and (_13264_, _10408_, _10407_);
  not (_10409_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_10410_, _10358_, _10409_);
  and (_10411_, _10358_, _09510_);
  or (_10412_, _10411_, _10410_);
  or (_10413_, _10412_, _10356_);
  or (_10414_, _10363_, word_in[12]);
  and (_10415_, _10414_, _10413_);
  or (_10417_, _10415_, _10355_);
  or (_10418_, _10368_, _09518_);
  and (_10420_, _10418_, _10367_);
  and (_10421_, _10420_, _10417_);
  and (_10422_, _10353_, word_in[28]);
  or (_13265_, _10422_, _10421_);
  and (_10423_, _10358_, _09525_);
  not (_10425_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_10426_, _10358_, _10425_);
  nor (_10428_, _10426_, _10423_);
  nor (_10429_, _10428_, _10356_);
  and (_10430_, _10356_, word_in[13]);
  or (_10431_, _10430_, _10429_);
  and (_10432_, _10431_, _10368_);
  and (_10433_, _10355_, _09523_);
  or (_10435_, _10433_, _10353_);
  or (_10436_, _10435_, _10432_);
  or (_10437_, _10367_, word_in[29]);
  and (_08227_, _10437_, _10436_);
  or (_10438_, _10368_, _09548_);
  not (_10439_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_10440_, _10358_, _10439_);
  and (_10441_, _10358_, _09541_);
  or (_10442_, _10441_, _10440_);
  or (_10444_, _10442_, _10356_);
  or (_10445_, _10363_, word_in[14]);
  and (_10446_, _10445_, _10444_);
  or (_10447_, _10446_, _10355_);
  and (_10448_, _10447_, _10438_);
  or (_10449_, _10448_, _10353_);
  or (_10450_, _10367_, word_in[30]);
  and (_08230_, _10450_, _10449_);
  nor (_10451_, _10358_, _08469_);
  and (_10452_, _10358_, _08760_);
  or (_10453_, _10452_, _10451_);
  or (_10454_, _10453_, _10356_);
  nand (_10455_, _10356_, _08764_);
  and (_10456_, _10455_, _10454_);
  or (_10457_, _10456_, _10355_);
  or (_10458_, _10368_, _08769_);
  and (_10460_, _10458_, _10367_);
  and (_10461_, _10460_, _10457_);
  and (_10462_, _10353_, word_in[31]);
  or (_08234_, _10462_, _10461_);
  and (_10463_, _05007_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  and (_10464_, _05670_, _04988_);
  and (_10465_, _05005_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  or (_10466_, _10465_, _10464_);
  and (_10467_, _10466_, _04861_);
  or (_10468_, _10467_, _10463_);
  and (_08279_, _10468_, _04856_);
  and (_10469_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  and (_10470_, _06686_, _06033_);
  or (_10472_, _10470_, _10469_);
  and (_08283_, _10472_, _04856_);
  and (_10474_, _10238_, _08514_);
  and (_10475_, _09565_, _08625_);
  not (_10476_, _10475_);
  or (_10477_, _10476_, _09349_);
  and (_10479_, _09569_, _08523_);
  not (_10481_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_10482_, _09572_, _08431_);
  nor (_10483_, _10482_, _10481_);
  and (_10484_, _10482_, word_in[0]);
  or (_10485_, _10484_, _10483_);
  or (_10486_, _10485_, _10479_);
  not (_10487_, _10479_);
  or (_10488_, _10487_, word_in[8]);
  and (_10489_, _10488_, _10486_);
  or (_10490_, _10489_, _10475_);
  and (_10491_, _10490_, _10477_);
  or (_10492_, _10491_, _10474_);
  not (_10493_, _10474_);
  or (_10494_, _10493_, word_in[24]);
  and (_08293_, _10494_, _10492_);
  not (_10495_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_10496_, _10482_, _10495_);
  and (_10497_, _10482_, word_in[1]);
  or (_10498_, _10497_, _10496_);
  or (_10500_, _10498_, _10479_);
  or (_10501_, _10487_, word_in[9]);
  and (_10502_, _10501_, _10500_);
  or (_10503_, _10502_, _10475_);
  or (_10504_, _10476_, _09464_);
  and (_10505_, _10504_, _10493_);
  and (_10506_, _10505_, _10503_);
  and (_10508_, _10474_, word_in[25]);
  or (_08297_, _10508_, _10506_);
  or (_10509_, _10476_, _09478_);
  not (_10510_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_10511_, _10482_, _10510_);
  and (_10512_, _10482_, word_in[2]);
  or (_10513_, _10512_, _10511_);
  or (_10515_, _10513_, _10479_);
  or (_10516_, _10487_, word_in[10]);
  and (_10517_, _10516_, _10515_);
  or (_10518_, _10517_, _10475_);
  and (_10519_, _10518_, _10509_);
  or (_10520_, _10519_, _10474_);
  or (_10521_, _10493_, word_in[26]);
  and (_08299_, _10521_, _10520_);
  not (_10522_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_10523_, _10482_, _10522_);
  and (_10524_, _10482_, word_in[3]);
  or (_10525_, _10524_, _10523_);
  or (_10526_, _10525_, _10479_);
  or (_10527_, _10487_, word_in[11]);
  and (_10528_, _10527_, _10526_);
  or (_10529_, _10528_, _10475_);
  or (_10530_, _10476_, _09493_);
  and (_10532_, _10530_, _10493_);
  and (_10533_, _10532_, _10529_);
  and (_10534_, _10474_, word_in[27]);
  or (_08300_, _10534_, _10533_);
  not (_10535_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_10536_, _10482_, _10535_);
  and (_10537_, _10482_, word_in[4]);
  or (_10538_, _10537_, _10536_);
  or (_10539_, _10538_, _10479_);
  or (_10540_, _10487_, word_in[12]);
  and (_10541_, _10540_, _10539_);
  or (_10542_, _10541_, _10475_);
  or (_10543_, _10476_, _09518_);
  and (_10544_, _10543_, _10493_);
  and (_10545_, _10544_, _10542_);
  and (_10546_, _10474_, word_in[28]);
  or (_08301_, _10546_, _10545_);
  not (_10548_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_10550_, _10482_, _10548_);
  and (_10551_, _10482_, word_in[5]);
  or (_10552_, _10551_, _10550_);
  or (_10554_, _10552_, _10479_);
  or (_10555_, _10487_, word_in[13]);
  and (_10556_, _10555_, _10554_);
  or (_10558_, _10556_, _10475_);
  or (_10559_, _10476_, _09523_);
  and (_10560_, _10559_, _10493_);
  and (_10561_, _10560_, _10558_);
  and (_10562_, _10474_, word_in[29]);
  or (_08302_, _10562_, _10561_);
  or (_10563_, _10476_, _09548_);
  not (_10564_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_10565_, _10482_, _10564_);
  and (_10567_, _10482_, word_in[6]);
  or (_10568_, _10567_, _10565_);
  or (_10569_, _10568_, _10479_);
  or (_10570_, _10487_, word_in[14]);
  and (_10571_, _10570_, _10569_);
  or (_10572_, _10571_, _10475_);
  and (_10573_, _10572_, _10563_);
  or (_10574_, _10573_, _10474_);
  or (_10575_, _10493_, word_in[30]);
  and (_08303_, _10575_, _10574_);
  nor (_10576_, _10482_, _08560_);
  and (_10577_, _10482_, word_in[7]);
  or (_10578_, _10577_, _10576_);
  or (_10579_, _10578_, _10479_);
  nand (_10580_, _10479_, _08764_);
  and (_10581_, _10580_, _10579_);
  or (_10582_, _10581_, _10475_);
  or (_10583_, _10476_, _08769_);
  and (_10584_, _10583_, _10493_);
  and (_10585_, _10584_, _10582_);
  and (_10586_, _10474_, word_in[31]);
  or (_08307_, _10586_, _10585_);
  and (_10587_, _05676_, _04861_);
  nand (_10588_, _10587_, _06369_);
  or (_10589_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_10590_, _10589_, _10588_);
  and (_08362_, _10590_, _04856_);
  and (_10591_, _09669_, _08625_);
  and (_10592_, _08752_, _08523_);
  not (_10593_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_10594_, _10248_, _08755_);
  nor (_10595_, _10594_, _10593_);
  and (_10596_, _10594_, _09449_);
  or (_10597_, _10596_, _10595_);
  or (_10598_, _10597_, _10592_);
  not (_10599_, _10592_);
  or (_10600_, _10599_, word_in[8]);
  and (_10601_, _10600_, _10598_);
  or (_10602_, _10601_, _10591_);
  and (_10603_, _10238_, _08548_);
  not (_10604_, _10603_);
  not (_10605_, _10591_);
  or (_10606_, _10605_, _09349_);
  and (_10607_, _10606_, _10604_);
  and (_10608_, _10607_, _10602_);
  and (_10609_, _10603_, word_in[24]);
  or (_08374_, _10609_, _10608_);
  and (_10610_, _10591_, _09464_);
  and (_10611_, _10594_, _09466_);
  not (_10612_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_10613_, _10594_, _10612_);
  nor (_10614_, _10613_, _10611_);
  nor (_10615_, _10614_, _10592_);
  and (_10616_, _10592_, word_in[9]);
  or (_10617_, _10616_, _10615_);
  and (_10618_, _10617_, _10605_);
  or (_10619_, _10618_, _10610_);
  and (_10620_, _10619_, _10604_);
  and (_10621_, _10603_, word_in[25]);
  or (_08379_, _10621_, _10620_);
  and (_10622_, _10591_, _09478_);
  and (_10623_, _10594_, _09480_);
  not (_10624_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_10625_, _10594_, _10624_);
  nor (_10626_, _10625_, _10623_);
  nor (_10627_, _10626_, _10592_);
  and (_10628_, _10592_, word_in[10]);
  or (_10629_, _10628_, _10627_);
  and (_10630_, _10629_, _10605_);
  or (_10631_, _10630_, _10622_);
  and (_10632_, _10631_, _10604_);
  and (_10633_, _10603_, word_in[26]);
  or (_08384_, _10633_, _10632_);
  and (_10634_, _10591_, _09493_);
  and (_10635_, _10594_, _09495_);
  not (_10636_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_10637_, _10594_, _10636_);
  nor (_10638_, _10637_, _10635_);
  nor (_10639_, _10638_, _10592_);
  and (_10640_, _10592_, word_in[11]);
  or (_10641_, _10640_, _10639_);
  and (_10642_, _10641_, _10605_);
  or (_10643_, _10642_, _10634_);
  and (_10644_, _10643_, _10604_);
  and (_10645_, _10603_, word_in[27]);
  or (_08388_, _10645_, _10644_);
  not (_10646_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_10647_, _10594_, _10646_);
  and (_10648_, _10594_, _09510_);
  or (_10649_, _10648_, _10647_);
  or (_10650_, _10649_, _10592_);
  or (_10651_, _10599_, word_in[12]);
  and (_10652_, _10651_, _10650_);
  or (_10653_, _10652_, _10591_);
  or (_10654_, _10605_, _09518_);
  and (_10655_, _10654_, _10604_);
  and (_10656_, _10655_, _10653_);
  and (_10657_, _10603_, word_in[28]);
  or (_08391_, _10657_, _10656_);
  and (_10658_, _10591_, _09523_);
  and (_10659_, _10594_, _09525_);
  not (_10660_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_10661_, _10594_, _10660_);
  nor (_10662_, _10661_, _10659_);
  nor (_10663_, _10662_, _10592_);
  and (_10664_, _10592_, word_in[13]);
  or (_10665_, _10664_, _10663_);
  and (_10666_, _10665_, _10605_);
  or (_10667_, _10666_, _10658_);
  and (_10668_, _10667_, _10604_);
  and (_10669_, _10603_, word_in[29]);
  or (_08395_, _10669_, _10668_);
  or (_10670_, _10605_, _09548_);
  not (_10671_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_10672_, _10594_, _10671_);
  and (_10673_, _10594_, _09541_);
  or (_10674_, _10673_, _10672_);
  or (_10676_, _10674_, _10592_);
  or (_10677_, _10599_, word_in[14]);
  and (_10678_, _10677_, _10676_);
  or (_10679_, _10678_, _10591_);
  and (_10680_, _10679_, _10670_);
  or (_10681_, _10680_, _10603_);
  or (_10682_, _10604_, word_in[30]);
  and (_08400_, _10682_, _10681_);
  nor (_10683_, _10594_, _08458_);
  and (_10684_, _10594_, _08760_);
  or (_10685_, _10684_, _10683_);
  or (_10686_, _10685_, _10592_);
  nand (_10687_, _10592_, _08764_);
  and (_10688_, _10687_, _10686_);
  or (_10689_, _10688_, _10591_);
  or (_10690_, _10605_, _08769_);
  and (_10691_, _10690_, _10604_);
  and (_10692_, _10691_, _10689_);
  and (_10693_, _10603_, word_in[31]);
  or (_08402_, _10693_, _10692_);
  and (_10694_, _08745_, _08511_);
  not (_10695_, _10694_);
  and (_10696_, _08749_, _08540_);
  and (_10697_, _10696_, _09349_);
  not (_10698_, _10696_);
  and (_10699_, _08751_, _09179_);
  not (_10700_, _10699_);
  and (_10701_, _09785_, _08757_);
  and (_10702_, _10701_, word_in[0]);
  not (_10703_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_10704_, _10701_, _10703_);
  or (_10705_, _10704_, _10702_);
  and (_10706_, _10705_, _10700_);
  and (_10707_, _10699_, word_in[8]);
  or (_10708_, _10707_, _10706_);
  and (_10709_, _10708_, _10698_);
  or (_10710_, _10709_, _10697_);
  and (_10711_, _10710_, _10695_);
  and (_10712_, _10694_, _09801_);
  or (_08492_, _10712_, _10711_);
  and (_10713_, _10696_, _09464_);
  not (_10714_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_10715_, _10701_, _10714_);
  and (_10716_, _10701_, word_in[1]);
  or (_10717_, _10716_, _10715_);
  and (_10718_, _10717_, _10700_);
  and (_10719_, _10699_, word_in[9]);
  or (_10720_, _10719_, _10718_);
  and (_10721_, _10720_, _10698_);
  or (_10722_, _10721_, _10713_);
  and (_10723_, _10722_, _10695_);
  and (_10724_, _10694_, _09366_);
  or (_08497_, _10724_, _10723_);
  and (_10725_, _10696_, _09478_);
  not (_10726_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_10727_, _10701_, _10726_);
  and (_10728_, _10701_, word_in[2]);
  or (_10729_, _10728_, _10727_);
  and (_10730_, _10729_, _10700_);
  and (_10731_, _10699_, word_in[10]);
  or (_10732_, _10731_, _10730_);
  and (_10733_, _10732_, _10698_);
  or (_10734_, _10733_, _10725_);
  and (_10735_, _10734_, _10695_);
  and (_10736_, _10694_, _09368_);
  or (_08499_, _10736_, _10735_);
  not (_10737_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_10738_, _10701_, _10737_);
  and (_10739_, _10701_, word_in[3]);
  or (_10740_, _10739_, _10738_);
  and (_10741_, _10740_, _10700_);
  and (_10742_, _10699_, word_in[11]);
  or (_10743_, _10742_, _10741_);
  and (_10744_, _10743_, _10698_);
  and (_10745_, _10696_, _09493_);
  or (_10746_, _10745_, _10694_);
  or (_10747_, _10746_, _10744_);
  or (_10748_, _10695_, _09380_);
  and (_08501_, _10748_, _10747_);
  not (_10749_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_10750_, _10701_, _10749_);
  and (_10751_, _10701_, word_in[4]);
  or (_10752_, _10751_, _10750_);
  and (_10753_, _10752_, _10700_);
  and (_10754_, _10699_, word_in[12]);
  or (_10755_, _10754_, _10753_);
  and (_10756_, _10755_, _10698_);
  and (_10757_, _10696_, _09518_);
  or (_10758_, _10757_, _10694_);
  or (_10759_, _10758_, _10756_);
  or (_10760_, _10695_, _09402_);
  and (_08504_, _10760_, _10759_);
  and (_10762_, _10696_, _09523_);
  not (_10763_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_10764_, _10701_, _10763_);
  and (_10765_, _10701_, word_in[5]);
  or (_10766_, _10765_, _10764_);
  and (_10767_, _10766_, _10700_);
  and (_10768_, _10699_, word_in[13]);
  or (_10769_, _10768_, _10767_);
  and (_10770_, _10769_, _10698_);
  or (_10771_, _10770_, _10762_);
  and (_10772_, _10771_, _10695_);
  and (_10773_, _10694_, _09414_);
  or (_08508_, _10773_, _10772_);
  and (_10774_, _10696_, _09548_);
  not (_10775_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_10776_, _10701_, _10775_);
  and (_10777_, _10701_, word_in[6]);
  or (_10778_, _10777_, _10776_);
  and (_10779_, _10778_, _10700_);
  and (_10780_, _10699_, word_in[14]);
  or (_10781_, _10780_, _10779_);
  and (_10782_, _10781_, _10698_);
  or (_10783_, _10782_, _10774_);
  and (_10784_, _10783_, _10695_);
  and (_10785_, _10694_, _09426_);
  or (_08510_, _10785_, _10784_);
  and (_10786_, _10696_, _08769_);
  nor (_10787_, _10701_, _08579_);
  and (_10788_, _10701_, word_in[7]);
  or (_10789_, _10788_, _10787_);
  and (_10790_, _10789_, _10700_);
  and (_10791_, _10699_, word_in[15]);
  or (_10792_, _10791_, _10790_);
  and (_10793_, _10792_, _10698_);
  or (_10794_, _10793_, _10786_);
  and (_10795_, _10794_, _10695_);
  and (_10796_, _10694_, _08774_);
  or (_08513_, _10796_, _10795_);
  nand (_10797_, _10587_, _06032_);
  or (_10798_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_10799_, _10798_, _04856_);
  and (_08582_, _10799_, _10797_);
  and (_10800_, _08745_, _08540_);
  not (_10801_, _10800_);
  and (_10802_, _08749_, _08514_);
  and (_10803_, _10802_, _09349_);
  not (_10804_, _10802_);
  and (_10805_, _09441_, _08573_);
  and (_10806_, _09445_, _08757_);
  and (_10807_, _10806_, word_in[0]);
  not (_10808_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_10809_, _10806_, _10808_);
  nor (_10810_, _10809_, _10807_);
  nor (_10811_, _10810_, _10805_);
  and (_10812_, _10805_, word_in[8]);
  or (_10813_, _10812_, _10811_);
  and (_10814_, _10813_, _10804_);
  or (_10815_, _10814_, _10803_);
  and (_10817_, _10815_, _10801_);
  and (_10818_, _10800_, _09801_);
  or (_13238_, _10818_, _10817_);
  not (_10819_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_10820_, _10806_, _10819_);
  and (_10821_, _10806_, _09466_);
  or (_10822_, _10821_, _10820_);
  or (_10823_, _10822_, _10805_);
  not (_10824_, _10805_);
  or (_10825_, _10824_, word_in[9]);
  and (_10826_, _10825_, _10823_);
  and (_10827_, _10826_, _10804_);
  and (_10828_, _10802_, _09464_);
  or (_10829_, _10828_, _10800_);
  or (_10830_, _10829_, _10827_);
  or (_10831_, _10801_, _09366_);
  and (_13239_, _10831_, _10830_);
  and (_10832_, _10806_, word_in[2]);
  not (_10833_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_10834_, _10806_, _10833_);
  nor (_10835_, _10834_, _10832_);
  nor (_10836_, _10835_, _10805_);
  and (_10837_, _10805_, word_in[10]);
  or (_10838_, _10837_, _10836_);
  and (_10839_, _10838_, _10804_);
  and (_10840_, _10802_, _09478_);
  or (_10841_, _10840_, _10800_);
  or (_10842_, _10841_, _10839_);
  or (_10843_, _10801_, _09368_);
  and (_13240_, _10843_, _10842_);
  not (_10844_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_10845_, _10806_, _10844_);
  and (_10846_, _10806_, _09495_);
  or (_10847_, _10846_, _10845_);
  or (_10848_, _10847_, _10805_);
  or (_10849_, _10824_, word_in[11]);
  and (_10851_, _10849_, _10848_);
  or (_10852_, _10851_, _10802_);
  or (_10853_, _10804_, _09493_);
  and (_10854_, _10853_, _10852_);
  or (_10855_, _10854_, _10800_);
  or (_10856_, _10801_, _09380_);
  and (_13241_, _10856_, _10855_);
  not (_10857_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_10858_, _10806_, _10857_);
  and (_10859_, _10806_, _09510_);
  or (_10860_, _10859_, _10858_);
  or (_10861_, _10860_, _10805_);
  or (_10862_, _10824_, word_in[12]);
  and (_10863_, _10862_, _10861_);
  or (_10864_, _10863_, _10802_);
  or (_10865_, _10804_, _09518_);
  and (_10867_, _10865_, _10864_);
  or (_10868_, _10867_, _10800_);
  or (_10870_, _10801_, _09402_);
  and (_13242_, _10870_, _10868_);
  not (_10871_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_10872_, _10806_, _10871_);
  and (_10873_, _10806_, _09525_);
  or (_10874_, _10873_, _10872_);
  or (_10875_, _10874_, _10805_);
  or (_10876_, _10824_, word_in[13]);
  and (_10877_, _10876_, _10875_);
  or (_10878_, _10877_, _10802_);
  or (_10879_, _10804_, _09523_);
  and (_10880_, _10879_, _10878_);
  or (_10881_, _10880_, _10800_);
  or (_10882_, _10801_, _09414_);
  and (_13243_, _10882_, _10881_);
  not (_10884_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_10885_, _10806_, _10884_);
  and (_10886_, _10806_, _09541_);
  or (_10887_, _10886_, _10885_);
  or (_10888_, _10887_, _10805_);
  or (_10890_, _10824_, word_in[14]);
  and (_10891_, _10890_, _10888_);
  or (_10892_, _10891_, _10802_);
  or (_10894_, _10804_, _09548_);
  and (_10895_, _10894_, _10892_);
  or (_10896_, _10895_, _10800_);
  or (_10897_, _10801_, _09426_);
  and (_13244_, _10897_, _10896_);
  nor (_10898_, _10806_, _08464_);
  and (_10899_, _10806_, _08760_);
  or (_10900_, _10899_, _10898_);
  or (_10901_, _10900_, _10805_);
  nand (_10903_, _10805_, _08764_);
  and (_10904_, _10903_, _10901_);
  or (_10905_, _10904_, _10802_);
  or (_10906_, _10804_, _08769_);
  and (_10907_, _10906_, _10905_);
  or (_10909_, _10907_, _10800_);
  or (_10910_, _10801_, _08774_);
  and (_13245_, _10910_, _10909_);
  and (_10912_, _08745_, _08514_);
  not (_10913_, _10912_);
  and (_10914_, _08749_, _08548_);
  and (_10915_, _10914_, _09349_);
  not (_10916_, _10914_);
  and (_10917_, _09569_, _08573_);
  and (_10918_, _09572_, _08741_);
  and (_10920_, _10918_, word_in[0]);
  not (_10921_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  nor (_10922_, _10918_, _10921_);
  nor (_10923_, _10922_, _10920_);
  nor (_10924_, _10923_, _10917_);
  and (_10925_, _10917_, word_in[8]);
  or (_10926_, _10925_, _10924_);
  and (_10927_, _10926_, _10916_);
  or (_10928_, _10927_, _10915_);
  and (_10929_, _10928_, _10913_);
  and (_10930_, _10912_, _09801_);
  or (_13246_, _10930_, _10929_);
  not (_10931_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_10932_, _10918_, _10931_);
  and (_10933_, _10918_, word_in[1]);
  nor (_10934_, _10933_, _10932_);
  nor (_10935_, _10934_, _10917_);
  and (_10936_, _10917_, word_in[9]);
  or (_10937_, _10936_, _10935_);
  and (_10938_, _10937_, _10916_);
  and (_10939_, _10914_, _09464_);
  or (_10940_, _10939_, _10912_);
  or (_10941_, _10940_, _10938_);
  or (_10942_, _10913_, _09366_);
  and (_08691_, _10942_, _10941_);
  not (_10943_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_10944_, _10918_, _10943_);
  and (_10945_, _10918_, word_in[2]);
  or (_10946_, _10945_, _10944_);
  or (_10947_, _10946_, _10917_);
  not (_10948_, _10917_);
  or (_10949_, _10948_, word_in[10]);
  and (_10950_, _10949_, _10947_);
  or (_10951_, _10950_, _10914_);
  or (_10952_, _10916_, _09478_);
  and (_10953_, _10952_, _10951_);
  or (_10954_, _10953_, _10912_);
  or (_10955_, _10913_, _09368_);
  and (_08694_, _10955_, _10954_);
  or (_10956_, _10948_, word_in[11]);
  not (_10957_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_10958_, _10918_, _10957_);
  and (_10959_, _10918_, word_in[3]);
  or (_10960_, _10959_, _10958_);
  or (_10961_, _10960_, _10917_);
  and (_10962_, _10961_, _10956_);
  or (_10963_, _10962_, _10914_);
  or (_10964_, _10916_, _09493_);
  and (_10965_, _10964_, _10963_);
  or (_10966_, _10965_, _10912_);
  or (_10967_, _10913_, _09380_);
  and (_08697_, _10967_, _10966_);
  not (_10968_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_10969_, _10918_, _10968_);
  and (_10970_, _10918_, word_in[4]);
  nor (_10971_, _10970_, _10969_);
  nor (_10972_, _10971_, _10917_);
  and (_10973_, _10917_, word_in[12]);
  or (_10974_, _10973_, _10972_);
  and (_10975_, _10974_, _10916_);
  and (_10976_, _10914_, _09518_);
  or (_10977_, _10976_, _10912_);
  or (_10978_, _10977_, _10975_);
  or (_10979_, _10913_, _09402_);
  and (_13247_, _10979_, _10978_);
  or (_10980_, _10916_, _09523_);
  not (_10981_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_10982_, _10918_, _10981_);
  and (_10983_, _10918_, word_in[5]);
  or (_10984_, _10983_, _10982_);
  or (_10985_, _10984_, _10917_);
  or (_10986_, _10948_, word_in[13]);
  and (_10987_, _10986_, _10985_);
  or (_10988_, _10987_, _10914_);
  and (_10989_, _10988_, _10980_);
  or (_10990_, _10989_, _10912_);
  or (_10991_, _10913_, _09414_);
  and (_08702_, _10991_, _10990_);
  and (_10993_, _10914_, _09548_);
  not (_10994_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_10995_, _10918_, _10994_);
  and (_10996_, _10918_, word_in[6]);
  nor (_10997_, _10996_, _10995_);
  nor (_10998_, _10997_, _10917_);
  and (_10999_, _10917_, word_in[14]);
  or (_11000_, _10999_, _10998_);
  and (_11001_, _11000_, _10916_);
  or (_11002_, _11001_, _10993_);
  and (_11003_, _11002_, _10913_);
  and (_11004_, _10912_, _09426_);
  or (_08705_, _11004_, _11003_);
  nand (_11005_, _10917_, _08764_);
  nor (_11006_, _10918_, _08574_);
  and (_11007_, _10918_, word_in[7]);
  or (_11008_, _11007_, _11006_);
  or (_11009_, _11008_, _10917_);
  and (_11010_, _11009_, _11005_);
  or (_11011_, _11010_, _10914_);
  or (_11012_, _10916_, _08769_);
  and (_11013_, _11012_, _11011_);
  or (_11014_, _11013_, _10912_);
  or (_11015_, _10913_, _08774_);
  and (_08709_, _11015_, _11014_);
  and (_11016_, _08758_, word_in[0]);
  not (_11017_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_11018_, _08758_, _11017_);
  nor (_11019_, _11018_, _11016_);
  nor (_11020_, _11019_, _08753_);
  and (_11021_, _08753_, word_in[8]);
  or (_11022_, _11021_, _11020_);
  and (_11023_, _11022_, _08768_);
  and (_11024_, _09349_, _08750_);
  or (_11025_, _11024_, _11023_);
  and (_11026_, _11025_, _08773_);
  and (_11027_, _09801_, _08746_);
  or (_13248_, _11027_, _11026_);
  not (_11028_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_11029_, _08758_, _11028_);
  and (_11030_, _09466_, _08758_);
  or (_11031_, _11030_, _11029_);
  or (_11032_, _11031_, _08753_);
  not (_11033_, _08753_);
  or (_11034_, _11033_, word_in[9]);
  and (_11035_, _11034_, _11032_);
  or (_11036_, _11035_, _08750_);
  or (_11037_, _09464_, _08768_);
  and (_11038_, _11037_, _11036_);
  or (_11039_, _11038_, _08746_);
  or (_11040_, _09366_, _08773_);
  and (_13249_, _11040_, _11039_);
  and (_11041_, _08758_, word_in[2]);
  not (_11043_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_11044_, _08758_, _11043_);
  nor (_11045_, _11044_, _11041_);
  nor (_11046_, _11045_, _08753_);
  and (_11047_, _08753_, word_in[10]);
  or (_11048_, _11047_, _11046_);
  and (_11049_, _11048_, _08768_);
  and (_11050_, _09478_, _08750_);
  or (_11051_, _11050_, _11049_);
  and (_11052_, _11051_, _08773_);
  and (_11053_, _09368_, _08746_);
  or (_13250_, _11053_, _11052_);
  and (_11054_, _08758_, word_in[3]);
  not (_11056_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_11057_, _08758_, _11056_);
  nor (_11059_, _11057_, _11054_);
  nor (_11060_, _11059_, _08753_);
  and (_11061_, _08753_, word_in[11]);
  or (_11062_, _11061_, _11060_);
  and (_11063_, _11062_, _08768_);
  and (_11064_, _09493_, _08750_);
  or (_11065_, _11064_, _11063_);
  and (_11066_, _11065_, _08773_);
  and (_11067_, _09380_, _08746_);
  or (_13251_, _11067_, _11066_);
  not (_11068_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_11069_, _08758_, _11068_);
  and (_11070_, _09510_, _08758_);
  or (_11071_, _11070_, _11069_);
  or (_11072_, _11071_, _08753_);
  or (_11073_, _11033_, word_in[12]);
  and (_11074_, _11073_, _11072_);
  or (_11075_, _11074_, _08750_);
  or (_11076_, _09518_, _08768_);
  and (_11077_, _11076_, _11075_);
  or (_11078_, _11077_, _08746_);
  or (_11079_, _09402_, _08773_);
  and (_13252_, _11079_, _11078_);
  not (_11080_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_11081_, _08758_, _11080_);
  and (_11082_, _09525_, _08758_);
  or (_11083_, _11082_, _11081_);
  or (_11084_, _11083_, _08753_);
  or (_11085_, _11033_, word_in[13]);
  and (_11086_, _11085_, _11084_);
  or (_11087_, _11086_, _08750_);
  or (_11088_, _09523_, _08768_);
  and (_11090_, _11088_, _11087_);
  or (_11091_, _11090_, _08746_);
  or (_11092_, _09414_, _08773_);
  and (_13253_, _11092_, _11091_);
  not (_11093_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_11094_, _08758_, _11093_);
  and (_11095_, _09541_, _08758_);
  or (_11096_, _11095_, _11094_);
  or (_11097_, _11096_, _08753_);
  or (_11098_, _11033_, word_in[14]);
  and (_11099_, _11098_, _11097_);
  or (_11100_, _11099_, _08750_);
  or (_11101_, _09548_, _08768_);
  and (_11102_, _11101_, _11100_);
  or (_11103_, _11102_, _08746_);
  or (_11104_, _09426_, _08773_);
  and (_13254_, _11104_, _11103_);
  and (_11105_, _06410_, _05671_);
  and (_11106_, _06696_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  or (_11107_, _11106_, _11105_);
  and (_08879_, _11107_, _04856_);
  nor (_08881_, _07651_, rst);
  and (_11108_, _08277_, _04986_);
  nand (_11109_, _11108_, _06088_);
  or (_11110_, _11108_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_11111_, _11110_, _06935_);
  and (_11112_, _11111_, _11109_);
  and (_11113_, _06934_, _06033_);
  or (_11114_, _11113_, _11112_);
  and (_09036_, _11114_, _04856_);
  and (_11115_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  and (_11116_, _06686_, _05718_);
  or (_11117_, _11116_, _11115_);
  and (_09073_, _11117_, _04856_);
  and (_11118_, _06705_, _05671_);
  and (_11119_, _06696_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or (_11120_, _11119_, _11118_);
  and (_09492_, _11120_, _04856_);
  or (_11121_, _05793_, _06812_);
  or (_11122_, _05729_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_11123_, _11122_, _04856_);
  and (_09513_, _11123_, _11121_);
  or (_11124_, _05818_, _06812_);
  or (_11125_, _05729_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_11126_, _11125_, _04856_);
  and (_09521_, _11126_, _11124_);
  or (_11127_, _05870_, _06812_);
  or (_11128_, _05729_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_11129_, _11128_, _04856_);
  and (_09529_, _11129_, _11127_);
  and (_11130_, _08451_, word_in[0]);
  nand (_11131_, _08361_, _10357_);
  or (_11132_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_11133_, _11132_, _11131_);
  and (_11134_, _11133_, _08416_);
  or (_11135_, _11134_, _08425_);
  nand (_11136_, _08361_, _10808_);
  or (_11137_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_11138_, _11137_, _11136_);
  and (_11139_, _11138_, _08393_);
  nand (_11140_, _08361_, _11017_);
  or (_11141_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_11142_, _11141_, _11140_);
  and (_11143_, _11142_, _08406_);
  nand (_11144_, _08361_, _10593_);
  or (_11145_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_11146_, _11145_, _11144_);
  and (_11147_, _11146_, _08397_);
  or (_11148_, _11147_, _11143_);
  or (_11149_, _11148_, _11139_);
  or (_11151_, _11149_, _11135_);
  nand (_11152_, _08361_, _09443_);
  or (_11153_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_11154_, _11153_, _11152_);
  and (_11155_, _11154_, _08416_);
  or (_11156_, _11155_, _08375_);
  nand (_11157_, _08361_, _09900_);
  or (_11158_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_11159_, _11158_, _11157_);
  and (_11160_, _11159_, _08393_);
  nand (_11161_, _08361_, _10123_);
  or (_11162_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_11163_, _11162_, _11161_);
  and (_11164_, _11163_, _08406_);
  nand (_11165_, _08361_, _09676_);
  or (_11166_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_11167_, _11166_, _11165_);
  and (_11168_, _11167_, _08397_);
  or (_11169_, _11168_, _11164_);
  or (_11170_, _11169_, _11160_);
  or (_11171_, _11170_, _11156_);
  and (_11172_, _11171_, _11151_);
  and (_11173_, _11172_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _11173_, _11130_);
  and (_11175_, _08451_, word_in[1]);
  nand (_11176_, _08361_, _10373_);
  or (_11177_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_11178_, _11177_, _11176_);
  and (_11179_, _11178_, _08416_);
  nand (_11180_, _08361_, _10612_);
  or (_11181_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_11182_, _11181_, _11180_);
  and (_11183_, _11182_, _08397_);
  nand (_11184_, _08361_, _10819_);
  or (_11185_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_11186_, _11185_, _11184_);
  and (_11187_, _11186_, _08393_);
  or (_11188_, _11187_, _11183_);
  or (_11189_, _11188_, _11179_);
  nand (_11190_, _08361_, _11028_);
  or (_11191_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_11192_, _11191_, _11190_);
  and (_11193_, _11192_, _08406_);
  or (_11194_, _11193_, _08425_);
  or (_11195_, _11194_, _11189_);
  nand (_11196_, _08361_, _09468_);
  or (_11197_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_11198_, _11197_, _11196_);
  and (_11199_, _11198_, _08416_);
  nand (_11200_, _08361_, _09691_);
  or (_11201_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_11202_, _11201_, _11200_);
  and (_11203_, _11202_, _08397_);
  nand (_11204_, _08361_, _09911_);
  or (_11205_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_11206_, _11205_, _11204_);
  and (_11207_, _11206_, _08393_);
  or (_11208_, _11207_, _11203_);
  or (_11209_, _11208_, _11199_);
  nand (_11210_, _08361_, _10134_);
  or (_11211_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_11212_, _11211_, _11210_);
  and (_11213_, _11212_, _08406_);
  or (_11214_, _11213_, _08375_);
  or (_11215_, _11214_, _11209_);
  and (_11216_, _11215_, _11195_);
  and (_11217_, _11216_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _11217_, _11175_);
  and (_11218_, _08451_, word_in[2]);
  nand (_11219_, _08361_, _10386_);
  or (_11220_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_11221_, _11220_, _11219_);
  and (_11222_, _11221_, _08416_);
  or (_11223_, _11222_, _08425_);
  nand (_11224_, _08361_, _10833_);
  or (_11225_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_11226_, _11225_, _11224_);
  and (_11227_, _11226_, _08393_);
  nand (_11228_, _08361_, _11043_);
  or (_11229_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_11230_, _11229_, _11228_);
  and (_11231_, _11230_, _08406_);
  nand (_11232_, _08361_, _10624_);
  or (_11233_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_11234_, _11233_, _11232_);
  and (_11235_, _11234_, _08397_);
  or (_11237_, _11235_, _11231_);
  or (_11238_, _11237_, _11227_);
  or (_11239_, _11238_, _11223_);
  nand (_11240_, _08361_, _09482_);
  or (_11241_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_11242_, _11241_, _11240_);
  and (_11243_, _11242_, _08416_);
  or (_11244_, _11243_, _08375_);
  nand (_11245_, _08361_, _09924_);
  or (_11246_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_11248_, _11246_, _11245_);
  and (_11249_, _11248_, _08393_);
  nand (_11250_, _08361_, _10149_);
  or (_11251_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_11252_, _11251_, _11250_);
  and (_11253_, _11252_, _08406_);
  nand (_11254_, _08361_, _09702_);
  or (_11255_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_11256_, _11255_, _11254_);
  and (_11257_, _11256_, _08397_);
  or (_11258_, _11257_, _11253_);
  or (_11259_, _11258_, _11249_);
  or (_11260_, _11259_, _11244_);
  and (_11261_, _11260_, _11239_);
  and (_11262_, _11261_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _11262_, _11218_);
  and (_11263_, _08451_, word_in[3]);
  nand (_11264_, _08361_, _10398_);
  or (_11265_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_11266_, _11265_, _11264_);
  and (_11267_, _11266_, _08416_);
  nand (_11268_, _08361_, _10636_);
  or (_11269_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_11270_, _11269_, _11268_);
  and (_11271_, _11270_, _08397_);
  nand (_11272_, _08361_, _10844_);
  or (_11273_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_11274_, _11273_, _11272_);
  and (_11275_, _11274_, _08393_);
  or (_11276_, _11275_, _11271_);
  or (_11277_, _11276_, _11267_);
  nand (_11278_, _08361_, _11056_);
  or (_11279_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_11280_, _11279_, _11278_);
  and (_11281_, _11280_, _08406_);
  or (_11282_, _11281_, _08425_);
  or (_11283_, _11282_, _11277_);
  nand (_11284_, _08361_, _09497_);
  or (_11285_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_11286_, _11285_, _11284_);
  and (_11287_, _11286_, _08416_);
  nand (_11288_, _08361_, _09715_);
  or (_11289_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_11290_, _11289_, _11288_);
  and (_11291_, _11290_, _08397_);
  nand (_11293_, _08361_, _09939_);
  or (_11294_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_11295_, _11294_, _11293_);
  and (_11296_, _11295_, _08393_);
  or (_11297_, _11296_, _11291_);
  or (_11298_, _11297_, _11287_);
  nand (_11299_, _08361_, _10160_);
  or (_11300_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_11301_, _11300_, _11299_);
  and (_11302_, _11301_, _08406_);
  or (_11303_, _11302_, _08375_);
  or (_11304_, _11303_, _11298_);
  and (_11305_, _11304_, _11283_);
  and (_11306_, _11305_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _11306_, _11263_);
  and (_11307_, _08451_, word_in[4]);
  nand (_11308_, _08361_, _10409_);
  or (_11309_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_11310_, _11309_, _11308_);
  and (_11311_, _11310_, _08416_);
  nand (_11313_, _08361_, _10646_);
  or (_11314_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_11315_, _11314_, _11313_);
  and (_11316_, _11315_, _08397_);
  nand (_11317_, _08361_, _10857_);
  or (_11318_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_11319_, _11318_, _11317_);
  and (_11320_, _11319_, _08393_);
  or (_11321_, _11320_, _11316_);
  or (_11322_, _11321_, _11311_);
  nand (_11323_, _08361_, _11068_);
  or (_11324_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_11325_, _11324_, _11323_);
  and (_11326_, _11325_, _08406_);
  or (_11328_, _11326_, _08425_);
  or (_11329_, _11328_, _11322_);
  nand (_11330_, _08361_, _09508_);
  or (_11331_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_11332_, _11331_, _11330_);
  and (_11333_, _11332_, _08416_);
  nand (_11334_, _08361_, _09728_);
  or (_11335_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_11336_, _11335_, _11334_);
  and (_11337_, _11336_, _08397_);
  nand (_11338_, _08361_, _09961_);
  or (_11339_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_11340_, _11339_, _11338_);
  and (_11341_, _11340_, _08393_);
  or (_11342_, _11341_, _11337_);
  or (_11344_, _11342_, _11333_);
  nand (_11345_, _08361_, _10175_);
  or (_11346_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_11348_, _11346_, _11345_);
  and (_11349_, _11348_, _08406_);
  or (_11351_, _11349_, _08375_);
  or (_11352_, _11351_, _11344_);
  and (_11353_, _11352_, _11329_);
  and (_11354_, _11353_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _11354_, _11307_);
  and (_11356_, _08451_, word_in[5]);
  nand (_11358_, _08361_, _10425_);
  or (_11359_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_11360_, _11359_, _11358_);
  and (_11361_, _11360_, _08416_);
  nand (_11362_, _08361_, _10660_);
  or (_11363_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_11364_, _11363_, _11362_);
  and (_11365_, _11364_, _08397_);
  nand (_11366_, _08361_, _10871_);
  or (_11367_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_11368_, _11367_, _11366_);
  and (_11369_, _11368_, _08393_);
  or (_11371_, _11369_, _11365_);
  or (_11372_, _11371_, _11361_);
  nand (_11373_, _08361_, _11080_);
  or (_11374_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_11375_, _11374_, _11373_);
  and (_11376_, _11375_, _08406_);
  or (_11377_, _11376_, _08425_);
  or (_11378_, _11377_, _11372_);
  nand (_11379_, _08361_, _09527_);
  or (_11380_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_11381_, _11380_, _11379_);
  and (_11382_, _11381_, _08416_);
  nand (_11383_, _08361_, _09740_);
  or (_11384_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_11385_, _11384_, _11383_);
  and (_11386_, _11385_, _08397_);
  nand (_11387_, _08361_, _09971_);
  or (_11388_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_11389_, _11388_, _11387_);
  and (_11390_, _11389_, _08393_);
  or (_11391_, _11390_, _11386_);
  or (_11392_, _11391_, _11382_);
  nand (_11393_, _08361_, _10187_);
  or (_11394_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_11395_, _11394_, _11393_);
  and (_11396_, _11395_, _08406_);
  or (_11397_, _11396_, _08375_);
  or (_11398_, _11397_, _11392_);
  and (_11399_, _11398_, _11378_);
  and (_11400_, _11399_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _11400_, _11356_);
  and (_11401_, _08451_, word_in[6]);
  nand (_11402_, _08361_, _10439_);
  or (_11403_, _08361_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_11404_, _11403_, _11402_);
  and (_11405_, _11404_, _08416_);
  nand (_11407_, _08361_, _10671_);
  or (_11408_, _08361_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_11409_, _11408_, _11407_);
  and (_11410_, _11409_, _08397_);
  nand (_11411_, _08361_, _10884_);
  or (_11413_, _08361_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_11414_, _11413_, _11411_);
  and (_11415_, _11414_, _08393_);
  or (_11416_, _11415_, _11410_);
  or (_11417_, _11416_, _11405_);
  nand (_11418_, _08361_, _11093_);
  or (_11419_, _08361_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_11420_, _11419_, _11418_);
  and (_11421_, _11420_, _08406_);
  or (_11422_, _11421_, _08425_);
  or (_11423_, _11422_, _11417_);
  nand (_11424_, _08361_, _09539_);
  or (_11425_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_11427_, _11425_, _11424_);
  and (_11429_, _11427_, _08416_);
  nand (_11430_, _08361_, _09752_);
  or (_11431_, _08361_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_11432_, _11431_, _11430_);
  and (_11433_, _11432_, _08397_);
  nand (_11434_, _08361_, _09983_);
  or (_11436_, _08361_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_11437_, _11436_, _11434_);
  and (_11438_, _11437_, _08393_);
  or (_11440_, _11438_, _11433_);
  or (_11441_, _11440_, _11429_);
  nand (_11442_, _08361_, _10203_);
  or (_11444_, _08361_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_11445_, _11444_, _11442_);
  and (_11446_, _11445_, _08406_);
  or (_11447_, _11446_, _08375_);
  or (_11448_, _11447_, _11441_);
  and (_11449_, _11448_, _11423_);
  and (_11450_, _11449_, _08450_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _11450_, _11401_);
  and (_11452_, _08557_, word_in[8]);
  nand (_11453_, _08361_, _10481_);
  or (_11454_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_11455_, _11454_, _11453_);
  and (_11456_, _11455_, _08559_);
  nand (_11457_, _08361_, _10246_);
  or (_11458_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_11459_, _11458_, _11457_);
  and (_11460_, _11459_, _08558_);
  or (_11461_, _11460_, _11456_);
  and (_11462_, _11461_, _08523_);
  nand (_11463_, _08361_, _09571_);
  or (_11465_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_11466_, _11465_, _11463_);
  and (_11468_, _11466_, _08559_);
  nand (_11469_, _08361_, _09332_);
  or (_11470_, _08361_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_11471_, _11470_, _11469_);
  and (_11472_, _11471_, _08558_);
  or (_11473_, _11472_, _11468_);
  and (_11474_, _11473_, _08525_);
  nand (_11475_, _08361_, _10016_);
  or (_11477_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_11478_, _11477_, _11475_);
  and (_11479_, _11478_, _08559_);
  nand (_11480_, _08361_, _09790_);
  or (_11481_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_11482_, _11481_, _11480_);
  and (_11483_, _11482_, _08558_);
  or (_11484_, _11483_, _11479_);
  and (_11485_, _11484_, _08600_);
  or (_11486_, _11485_, _11474_);
  nand (_11487_, _08361_, _10921_);
  or (_11488_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_11489_, _11488_, _11487_);
  and (_11490_, _11489_, _08559_);
  nand (_11491_, _08361_, _10703_);
  or (_11492_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_11493_, _11492_, _11491_);
  and (_11494_, _11493_, _08558_);
  or (_11495_, _11494_, _11490_);
  and (_11496_, _11495_, _08573_);
  or (_11497_, _11496_, _11486_);
  nor (_11498_, _11497_, _11462_);
  nor (_11499_, _11498_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _11499_, _11452_);
  and (_11500_, _08557_, word_in[9]);
  nand (_11501_, _08361_, _10495_);
  or (_11502_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_11503_, _11502_, _11501_);
  and (_11504_, _11503_, _08559_);
  nand (_11505_, _08361_, _10263_);
  or (_11506_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_11507_, _11506_, _11505_);
  and (_11508_, _11507_, _08558_);
  or (_11509_, _11508_, _11504_);
  and (_11510_, _11509_, _08523_);
  nand (_11511_, _08361_, _09586_);
  or (_11512_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_11513_, _11512_, _11511_);
  and (_11514_, _11513_, _08559_);
  and (_11515_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_11516_, _08361_, _09468_);
  or (_11517_, _11516_, _11515_);
  and (_11518_, _11517_, _08558_);
  or (_11519_, _11518_, _11514_);
  and (_11520_, _11519_, _08525_);
  nand (_11521_, _08361_, _10026_);
  or (_11523_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_11524_, _11523_, _11521_);
  and (_11525_, _11524_, _08559_);
  nand (_11526_, _08361_, _09804_);
  or (_11527_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_11528_, _11527_, _11526_);
  and (_11529_, _11528_, _08558_);
  or (_11530_, _11529_, _11525_);
  and (_11531_, _11530_, _08600_);
  or (_11532_, _11531_, _11520_);
  nand (_11533_, _08361_, _10931_);
  or (_11534_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_11535_, _11534_, _11533_);
  and (_11536_, _11535_, _08559_);
  nand (_11537_, _08361_, _10714_);
  or (_11538_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_11539_, _11538_, _11537_);
  and (_11540_, _11539_, _08558_);
  or (_11541_, _11540_, _11536_);
  and (_11542_, _11541_, _08573_);
  or (_11544_, _11542_, _11532_);
  nor (_11545_, _11544_, _11510_);
  nor (_11546_, _11545_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _11546_, _11500_);
  and (_11547_, _08557_, word_in[10]);
  nand (_11548_, _08361_, _10510_);
  or (_11549_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_11550_, _11549_, _11548_);
  and (_11551_, _11550_, _08559_);
  nand (_11552_, _08361_, _10276_);
  or (_11553_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_11554_, _11553_, _11552_);
  and (_11555_, _11554_, _08558_);
  or (_11556_, _11555_, _11551_);
  and (_11557_, _11556_, _08523_);
  nand (_11558_, _08361_, _09599_);
  or (_11559_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_11560_, _11559_, _11558_);
  and (_11561_, _11560_, _08559_);
  and (_11562_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_11563_, _08361_, _09482_);
  or (_11564_, _11563_, _11562_);
  and (_11566_, _11564_, _08558_);
  or (_11567_, _11566_, _11561_);
  and (_11568_, _11567_, _08525_);
  nand (_11569_, _08361_, _10040_);
  or (_11570_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_11571_, _11570_, _11569_);
  and (_11572_, _11571_, _08559_);
  nand (_11573_, _08361_, _09818_);
  or (_11574_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_11575_, _11574_, _11573_);
  and (_11576_, _11575_, _08558_);
  or (_11577_, _11576_, _11572_);
  and (_11578_, _11577_, _08600_);
  or (_11580_, _11578_, _11568_);
  nand (_11581_, _08361_, _10943_);
  or (_11582_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_11583_, _11582_, _11581_);
  and (_11584_, _11583_, _08559_);
  nand (_11585_, _08361_, _10726_);
  or (_11586_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_11587_, _11586_, _11585_);
  and (_11588_, _11587_, _08558_);
  or (_11589_, _11588_, _11584_);
  and (_11590_, _11589_, _08573_);
  or (_11591_, _11590_, _11580_);
  nor (_11592_, _11591_, _11557_);
  nor (_11593_, _11592_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _11593_, _11547_);
  and (_11594_, _08557_, word_in[11]);
  nand (_11596_, _08361_, _10522_);
  or (_11597_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_11599_, _11597_, _11596_);
  and (_11600_, _11599_, _08559_);
  nand (_11601_, _08361_, _10288_);
  or (_11603_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_11604_, _11603_, _11601_);
  and (_11606_, _11604_, _08558_);
  or (_11607_, _11606_, _11600_);
  and (_11608_, _11607_, _08523_);
  nand (_11609_, _08361_, _10957_);
  or (_11611_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_11612_, _11611_, _11609_);
  and (_11613_, _11612_, _08559_);
  nand (_11614_, _08361_, _10737_);
  or (_11615_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_11617_, _11615_, _11614_);
  and (_11619_, _11617_, _08558_);
  or (_11621_, _11619_, _11613_);
  and (_11622_, _11621_, _08573_);
  nand (_11623_, _08361_, _10053_);
  or (_11625_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_11626_, _11625_, _11623_);
  and (_11627_, _11626_, _08559_);
  nand (_11628_, _08361_, _09834_);
  or (_11629_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_11631_, _11629_, _11628_);
  and (_11632_, _11631_, _08558_);
  or (_11633_, _11632_, _11627_);
  and (_11634_, _11633_, _08600_);
  nand (_11635_, _08361_, _09610_);
  or (_11636_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_11637_, _11636_, _11635_);
  and (_11639_, _11637_, _08559_);
  and (_11640_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_11642_, _08361_, _09497_);
  or (_11643_, _11642_, _11640_);
  and (_11644_, _11643_, _08558_);
  or (_11645_, _11644_, _11639_);
  and (_11647_, _11645_, _08525_);
  or (_11648_, _11647_, _11634_);
  or (_11649_, _11648_, _11622_);
  nor (_11650_, _11649_, _11608_);
  nor (_11651_, _11650_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _11651_, _11594_);
  and (_11652_, _08557_, word_in[12]);
  nand (_11653_, _08361_, _10535_);
  or (_11654_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_11655_, _11654_, _11653_);
  and (_11656_, _11655_, _08559_);
  nand (_11657_, _08361_, _10302_);
  or (_11659_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_11660_, _11659_, _11657_);
  and (_11661_, _11660_, _08558_);
  or (_11662_, _11661_, _11656_);
  and (_11663_, _11662_, _08523_);
  nand (_11664_, _08361_, _09622_);
  or (_11665_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_11666_, _11665_, _11664_);
  and (_11667_, _11666_, _08559_);
  and (_11668_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_11669_, _08361_, _09508_);
  or (_11670_, _11669_, _11668_);
  and (_11671_, _11670_, _08558_);
  or (_11672_, _11671_, _11667_);
  and (_11673_, _11672_, _08525_);
  nand (_11674_, _08361_, _10066_);
  or (_11675_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_11676_, _11675_, _11674_);
  and (_11677_, _11676_, _08559_);
  nand (_11678_, _08361_, _09846_);
  or (_11679_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_11680_, _11679_, _11678_);
  and (_11681_, _11680_, _08558_);
  or (_11682_, _11681_, _11677_);
  and (_11683_, _11682_, _08600_);
  or (_11684_, _11683_, _11673_);
  nand (_11685_, _08361_, _10968_);
  or (_11686_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_11687_, _11686_, _11685_);
  and (_11688_, _11687_, _08559_);
  nand (_11689_, _08361_, _10749_);
  or (_11690_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_11691_, _11690_, _11689_);
  and (_11692_, _11691_, _08558_);
  or (_11693_, _11692_, _11688_);
  and (_11694_, _11693_, _08573_);
  or (_11695_, _11694_, _11684_);
  nor (_11696_, _11695_, _11663_);
  nor (_11697_, _11696_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _11697_, _11652_);
  and (_11699_, _08557_, word_in[13]);
  nand (_11700_, _08361_, _10548_);
  or (_11701_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_11702_, _11701_, _11700_);
  and (_11703_, _11702_, _08559_);
  nand (_11705_, _08361_, _10315_);
  or (_11706_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_11707_, _11706_, _11705_);
  and (_11708_, _11707_, _08558_);
  or (_11709_, _11708_, _11703_);
  and (_11711_, _11709_, _08523_);
  nand (_11712_, _08361_, _09635_);
  or (_11713_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_11714_, _11713_, _11712_);
  and (_11716_, _11714_, _08559_);
  and (_11717_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_11719_, _08361_, _09527_);
  or (_11721_, _11719_, _11717_);
  and (_11722_, _11721_, _08558_);
  or (_11724_, _11722_, _11716_);
  and (_11725_, _11724_, _08525_);
  nand (_11727_, _08361_, _10080_);
  or (_11728_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_11730_, _11728_, _11727_);
  and (_11731_, _11730_, _08559_);
  nand (_11732_, _08361_, _09858_);
  or (_11733_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_11734_, _11733_, _11732_);
  and (_11735_, _11734_, _08558_);
  or (_11737_, _11735_, _11731_);
  and (_11738_, _11737_, _08600_);
  or (_11739_, _11738_, _11725_);
  nand (_11740_, _08361_, _10981_);
  or (_11741_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_11742_, _11741_, _11740_);
  and (_11743_, _11742_, _08559_);
  nand (_11744_, _08361_, _10763_);
  or (_11745_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_11746_, _11745_, _11744_);
  and (_11747_, _11746_, _08558_);
  or (_11748_, _11747_, _11743_);
  and (_11749_, _11748_, _08573_);
  or (_11750_, _11749_, _11739_);
  nor (_11752_, _11750_, _11711_);
  nor (_11753_, _11752_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _11753_, _11699_);
  and (_11755_, _08557_, word_in[14]);
  nand (_11756_, _08361_, _10564_);
  or (_11757_, _08361_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_11758_, _11757_, _11756_);
  and (_11759_, _11758_, _08559_);
  nand (_11760_, _08361_, _10328_);
  or (_11761_, _08361_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_11762_, _11761_, _11760_);
  and (_11763_, _11762_, _08558_);
  or (_11764_, _11763_, _11759_);
  and (_11765_, _11764_, _08523_);
  nand (_11766_, _08361_, _10994_);
  or (_11767_, _08361_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_11768_, _11767_, _11766_);
  and (_11769_, _11768_, _08559_);
  nand (_11770_, _08361_, _10775_);
  or (_11771_, _08361_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_11772_, _11771_, _11770_);
  and (_11773_, _11772_, _08558_);
  or (_11774_, _11773_, _11769_);
  and (_11775_, _11774_, _08573_);
  nand (_11776_, _08361_, _10092_);
  or (_11777_, _08361_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_11778_, _11777_, _11776_);
  and (_11779_, _11778_, _08559_);
  nand (_11780_, _08361_, _09870_);
  or (_11781_, _08361_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_11782_, _11781_, _11780_);
  and (_11783_, _11782_, _08558_);
  or (_11784_, _11783_, _11779_);
  and (_11785_, _11784_, _08600_);
  nand (_11786_, _08361_, _09647_);
  or (_11787_, _08361_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_11788_, _11787_, _11786_);
  and (_11789_, _11788_, _08559_);
  and (_11790_, _08361_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_11791_, _08361_, _09539_);
  or (_11793_, _11791_, _11790_);
  and (_11794_, _11793_, _08558_);
  or (_11795_, _11794_, _11789_);
  and (_11796_, _11795_, _08525_);
  or (_11797_, _11796_, _11785_);
  or (_11798_, _11797_, _11775_);
  nor (_11799_, _11798_, _11765_);
  nor (_11800_, _11799_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _11800_, _11755_);
  and (_11802_, _08654_, word_in[16]);
  and (_11803_, _11154_, _08406_);
  and (_11804_, _11163_, _08393_);
  or (_11806_, _11804_, _11803_);
  and (_11807_, _11159_, _08397_);
  and (_11808_, _11167_, _08416_);
  or (_11809_, _11808_, _11807_);
  or (_11810_, _11809_, _11806_);
  or (_11811_, _11810_, _08619_);
  and (_11812_, _11138_, _08397_);
  and (_11813_, _11133_, _08406_);
  or (_11814_, _11813_, _11812_);
  and (_11815_, _11142_, _08393_);
  and (_11816_, _11146_, _08416_);
  or (_11817_, _11816_, _11815_);
  nor (_11818_, _11817_, _11814_);
  nand (_11819_, _11818_, _08619_);
  nand (_11820_, _11819_, _11811_);
  nor (_11821_, _11820_, _08654_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _11821_, _11802_);
  and (_11822_, _08654_, word_in[17]);
  and (_11823_, _11206_, _08397_);
  and (_11824_, _11198_, _08406_);
  or (_11826_, _11824_, _11823_);
  and (_11827_, _11212_, _08393_);
  and (_11828_, _11202_, _08416_);
  or (_11829_, _11828_, _11827_);
  or (_11831_, _11829_, _11826_);
  or (_11832_, _11831_, _08619_);
  and (_11833_, _11186_, _08397_);
  and (_11834_, _11178_, _08406_);
  or (_11835_, _11834_, _11833_);
  and (_11836_, _11192_, _08393_);
  and (_11837_, _11182_, _08416_);
  or (_11838_, _11837_, _11836_);
  nor (_11839_, _11838_, _11835_);
  nand (_11840_, _11839_, _08619_);
  nand (_11841_, _11840_, _11832_);
  nor (_11842_, _11841_, _08654_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _11842_, _11822_);
  and (_11843_, _08654_, word_in[18]);
  and (_11845_, _11248_, _08397_);
  and (_11846_, _11242_, _08406_);
  or (_11847_, _11846_, _11845_);
  and (_11849_, _11252_, _08393_);
  and (_11850_, _11256_, _08416_);
  or (_11851_, _11850_, _11849_);
  or (_11852_, _11851_, _11847_);
  or (_11853_, _11852_, _08619_);
  and (_11854_, _11226_, _08397_);
  and (_11855_, _11221_, _08406_);
  or (_11857_, _11855_, _11854_);
  and (_11858_, _11230_, _08393_);
  and (_11859_, _11234_, _08416_);
  or (_11860_, _11859_, _11858_);
  nor (_11861_, _11860_, _11857_);
  nand (_11862_, _11861_, _08619_);
  nand (_11863_, _11862_, _11853_);
  nor (_11864_, _11863_, _08654_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _11864_, _11843_);
  and (_11865_, _08654_, word_in[19]);
  and (_11866_, _11295_, _08397_);
  and (_11867_, _11286_, _08406_);
  or (_11868_, _11867_, _11866_);
  and (_11869_, _11301_, _08393_);
  and (_11870_, _11290_, _08416_);
  or (_11871_, _11870_, _11869_);
  or (_11872_, _11871_, _11868_);
  or (_11873_, _11872_, _08619_);
  and (_11874_, _11266_, _08406_);
  and (_11875_, _11280_, _08393_);
  or (_11876_, _11875_, _11874_);
  and (_11878_, _11274_, _08397_);
  and (_11879_, _11270_, _08416_);
  or (_11880_, _11879_, _11878_);
  nor (_11881_, _11880_, _11876_);
  nand (_11882_, _11881_, _08619_);
  nand (_11884_, _11882_, _11873_);
  nor (_11885_, _11884_, _08654_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _11885_, _11865_);
  and (_11886_, _08654_, word_in[20]);
  and (_11887_, _11332_, _08406_);
  and (_11889_, _11348_, _08393_);
  or (_11890_, _11889_, _11887_);
  and (_11892_, _11340_, _08397_);
  and (_11893_, _11336_, _08416_);
  or (_11894_, _11893_, _11892_);
  or (_11895_, _11894_, _11890_);
  or (_11896_, _11895_, _08619_);
  and (_11898_, _11319_, _08397_);
  and (_11899_, _11310_, _08406_);
  or (_11901_, _11899_, _11898_);
  and (_11902_, _11325_, _08393_);
  and (_11903_, _11315_, _08416_);
  or (_11905_, _11903_, _11902_);
  nor (_11906_, _11905_, _11901_);
  nand (_11908_, _11906_, _08619_);
  nand (_11909_, _11908_, _11896_);
  nor (_11911_, _11909_, _08654_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _11911_, _11886_);
  and (_11912_, _08654_, word_in[21]);
  and (_11913_, _11389_, _08397_);
  and (_11915_, _11381_, _08406_);
  or (_11916_, _11915_, _11913_);
  and (_11917_, _11395_, _08393_);
  and (_11918_, _11385_, _08416_);
  or (_11919_, _11918_, _11917_);
  or (_11920_, _11919_, _11916_);
  or (_11921_, _11920_, _08619_);
  and (_11922_, _11360_, _08406_);
  and (_11923_, _11375_, _08393_);
  or (_11925_, _11923_, _11922_);
  and (_11926_, _11368_, _08397_);
  and (_11928_, _11364_, _08416_);
  or (_11929_, _11928_, _11926_);
  nor (_11931_, _11929_, _11925_);
  nand (_11932_, _11931_, _08619_);
  nand (_11933_, _11932_, _11921_);
  nor (_11934_, _11933_, _08654_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _11934_, _11912_);
  and (_11935_, _08654_, word_in[22]);
  and (_11936_, _11427_, _08406_);
  and (_11937_, _11445_, _08393_);
  or (_11938_, _11937_, _11936_);
  and (_11939_, _11437_, _08397_);
  and (_11940_, _11432_, _08416_);
  or (_11941_, _11940_, _11939_);
  or (_11942_, _11941_, _11938_);
  or (_11943_, _11942_, _08619_);
  and (_11944_, _11404_, _08406_);
  and (_11946_, _11420_, _08393_);
  or (_11947_, _11946_, _11944_);
  and (_11948_, _11414_, _08397_);
  and (_11949_, _11409_, _08416_);
  or (_11950_, _11949_, _11948_);
  nor (_11951_, _11950_, _11947_);
  nand (_11952_, _11951_, _08619_);
  nand (_11953_, _11952_, _11943_);
  nor (_11954_, _11953_, _08654_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _11954_, _11935_);
  and (_11955_, _08717_, word_in[24]);
  and (_11956_, _11459_, _08559_);
  and (_11957_, _11455_, _08558_);
  or (_11958_, _11957_, _11956_);
  and (_11959_, _11958_, _08685_);
  and (_11960_, _11471_, _08559_);
  and (_11961_, _11466_, _08558_);
  or (_11962_, _11961_, _11960_);
  and (_11963_, _11962_, _08690_);
  and (_11964_, _11482_, _08559_);
  and (_11965_, _11478_, _08558_);
  or (_11966_, _11965_, _11964_);
  and (_11967_, _11966_, _08726_);
  and (_11968_, _11493_, _08559_);
  and (_11969_, _11489_, _08558_);
  or (_11970_, _11969_, _11968_);
  and (_11971_, _11970_, _08731_);
  or (_11972_, _11971_, _11967_);
  or (_11973_, _11972_, _11963_);
  nor (_11974_, _11973_, _11959_);
  nor (_11975_, _11974_, _08717_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _11975_, _11955_);
  and (_11976_, _08717_, word_in[25]);
  and (_11977_, _11507_, _08559_);
  and (_11978_, _11503_, _08558_);
  or (_11980_, _11978_, _11977_);
  and (_11981_, _11980_, _08685_);
  and (_11982_, _11517_, _08559_);
  and (_11983_, _11513_, _08558_);
  or (_11985_, _11983_, _11982_);
  and (_11986_, _11985_, _08690_);
  and (_11987_, _11528_, _08559_);
  and (_11988_, _11524_, _08558_);
  or (_11989_, _11988_, _11987_);
  and (_11990_, _11989_, _08726_);
  and (_11991_, _11539_, _08559_);
  and (_11992_, _11535_, _08558_);
  or (_11994_, _11992_, _11991_);
  and (_11996_, _11994_, _08731_);
  or (_11997_, _11996_, _11990_);
  or (_11998_, _11997_, _11986_);
  nor (_11999_, _11998_, _11981_);
  nor (_12000_, _11999_, _08717_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _12000_, _11976_);
  and (_12002_, _08717_, word_in[26]);
  and (_12003_, _11564_, _08559_);
  and (_12004_, _11560_, _08558_);
  or (_12005_, _12004_, _12003_);
  and (_12007_, _12005_, _08690_);
  and (_12008_, _11554_, _08559_);
  and (_12009_, _11550_, _08558_);
  or (_12010_, _12009_, _12008_);
  and (_12012_, _12010_, _08685_);
  and (_12013_, _11575_, _08559_);
  and (_12015_, _11571_, _08558_);
  or (_12016_, _12015_, _12013_);
  and (_12018_, _12016_, _08726_);
  and (_12019_, _11587_, _08559_);
  and (_12020_, _11583_, _08558_);
  or (_12021_, _12020_, _12019_);
  and (_12022_, _12021_, _08731_);
  or (_12023_, _12022_, _12018_);
  or (_12024_, _12023_, _12012_);
  nor (_12025_, _12024_, _12007_);
  nor (_12026_, _12025_, _08717_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _12026_, _12002_);
  and (_12027_, _08717_, word_in[27]);
  and (_12028_, _11643_, _08559_);
  and (_12029_, _11637_, _08558_);
  or (_12030_, _12029_, _12028_);
  and (_12031_, _12030_, _08690_);
  and (_12033_, _11604_, _08559_);
  and (_12034_, _11599_, _08558_);
  or (_12036_, _12034_, _12033_);
  and (_12037_, _12036_, _08685_);
  and (_12039_, _11631_, _08559_);
  and (_12041_, _11626_, _08558_);
  or (_12043_, _12041_, _12039_);
  and (_12044_, _12043_, _08726_);
  and (_12045_, _11617_, _08559_);
  and (_12046_, _11612_, _08558_);
  or (_12047_, _12046_, _12045_);
  and (_12048_, _12047_, _08731_);
  or (_12050_, _12048_, _12044_);
  or (_12051_, _12050_, _12037_);
  nor (_12052_, _12051_, _12031_);
  nor (_12053_, _12052_, _08717_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _12053_, _12027_);
  and (_12054_, _08717_, word_in[28]);
  and (_12055_, _11660_, _08559_);
  and (_12056_, _11655_, _08558_);
  or (_12057_, _12056_, _12055_);
  and (_12058_, _12057_, _08685_);
  and (_12059_, _11670_, _08559_);
  and (_12060_, _11666_, _08558_);
  or (_12061_, _12060_, _12059_);
  and (_12062_, _12061_, _08690_);
  and (_12063_, _11680_, _08559_);
  and (_12064_, _11676_, _08558_);
  or (_12065_, _12064_, _12063_);
  and (_12066_, _12065_, _08726_);
  and (_12067_, _11691_, _08559_);
  and (_12068_, _11687_, _08558_);
  or (_12069_, _12068_, _12067_);
  and (_12070_, _12069_, _08731_);
  or (_12071_, _12070_, _12066_);
  or (_12072_, _12071_, _12062_);
  nor (_12073_, _12072_, _12058_);
  nor (_12074_, _12073_, _08717_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _12074_, _12054_);
  and (_12075_, _08717_, word_in[29]);
  and (_12076_, _11707_, _08559_);
  and (_12078_, _11702_, _08558_);
  or (_12079_, _12078_, _12076_);
  and (_12080_, _12079_, _08685_);
  and (_12081_, _11721_, _08559_);
  and (_12083_, _11714_, _08558_);
  or (_12084_, _12083_, _12081_);
  and (_12085_, _12084_, _08690_);
  and (_12086_, _11734_, _08559_);
  and (_12087_, _11730_, _08558_);
  or (_12088_, _12087_, _12086_);
  and (_12089_, _12088_, _08726_);
  and (_12090_, _11746_, _08559_);
  and (_12091_, _11742_, _08558_);
  or (_12092_, _12091_, _12090_);
  and (_12094_, _12092_, _08731_);
  or (_12095_, _12094_, _12089_);
  or (_12096_, _12095_, _12085_);
  nor (_12097_, _12096_, _12080_);
  nor (_12098_, _12097_, _08717_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _12098_, _12075_);
  and (_12099_, _08717_, word_in[30]);
  and (_12100_, _11793_, _08559_);
  and (_12101_, _11788_, _08558_);
  or (_12102_, _12101_, _12100_);
  and (_12103_, _12102_, _08690_);
  and (_12104_, _11762_, _08559_);
  and (_12105_, _11758_, _08558_);
  or (_12106_, _12105_, _12104_);
  and (_12107_, _12106_, _08685_);
  and (_12108_, _11782_, _08559_);
  and (_12109_, _11778_, _08558_);
  or (_12110_, _12109_, _12108_);
  and (_12111_, _12110_, _08726_);
  and (_12112_, _11772_, _08559_);
  and (_12113_, _11768_, _08558_);
  or (_12114_, _12113_, _12112_);
  and (_12115_, _12114_, _08731_);
  or (_12116_, _12115_, _12111_);
  or (_12117_, _12116_, _12107_);
  nor (_12118_, _12117_, _12103_);
  nor (_12120_, _12118_, _08717_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _12120_, _12099_);
  or (_12121_, _05843_, _06812_);
  or (_12122_, _05729_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_12123_, _12122_, _04856_);
  and (_09782_, _12123_, _12121_);
  and (_09788_, _06849_, _04856_);
  or (_12124_, _05943_, _06812_);
  or (_12125_, _05729_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_12126_, _12125_, _04856_);
  and (_09791_, _12126_, _12124_);
  or (_12127_, _05983_, _05848_);
  and (_12129_, _12127_, _06777_);
  nor (_12131_, _06783_, _12129_);
  or (_09794_, _12131_, _06782_);
  or (_12132_, _05895_, _06812_);
  or (_12133_, _05729_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_12134_, _12133_, _04856_);
  and (_09806_, _12134_, _12132_);
  or (_12136_, _08164_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_12138_, _08168_, _08166_);
  or (_12139_, _12138_, _08159_);
  or (_12140_, _12139_, _12136_);
  and (_12142_, _12140_, _08181_);
  nor (_12143_, _08180_, _05957_);
  or (_12144_, _12143_, rst);
  or (_09810_, _12144_, _12142_);
  or (_12145_, _05767_, _06812_);
  or (_12146_, _05729_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_12148_, _12146_, _04856_);
  and (_09813_, _12148_, _12145_);
  and (_12149_, _05983_, _06772_);
  nor (_12150_, _06783_, _12149_);
  or (_09820_, _12150_, _06782_);
  and (_09822_, _06903_, _04856_);
  and (_12152_, _09950_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_12153_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_12155_, _12153_, _09954_);
  and (_12157_, _05718_, _05671_);
  or (_12158_, _12157_, _12155_);
  or (_12159_, _12158_, _12152_);
  and (_09831_, _12159_, _04856_);
  or (_12160_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand (_12161_, _08367_, _05906_);
  and (_12162_, _12161_, _04856_);
  and (_09984_, _12162_, _12160_);
  and (_12164_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  not (_12165_, _08367_);
  and (_12166_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or (_12167_, _12166_, _12164_);
  and (_09996_, _12167_, _04856_);
  and (_12168_, _06818_, _04856_);
  and (_10047_, _12168_, _06851_);
  nor (_12170_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_12171_, _12170_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_10060_, _12171_, _04856_);
  and (_02999_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _04856_);
  and (_12174_, _02999_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_10067_, _12174_, _10060_);
  nand (_12175_, _05726_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_10072_, _12175_, _04856_);
  and (_10114_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _04856_);
  nor (_12176_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_10135_, _12176_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_12177_, _08275_, _06142_);
  and (_12179_, _12177_, _04986_);
  or (_12180_, _12179_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_12182_, _06662_, _04993_);
  and (_12183_, _12182_, _06126_);
  not (_12185_, _12183_);
  and (_12186_, _12185_, _12180_);
  nand (_12187_, _12179_, _06088_);
  and (_12188_, _12187_, _12186_);
  nor (_12189_, _12185_, _06032_);
  or (_12190_, _12189_, _12188_);
  and (_10143_, _12190_, _04856_);
  and (_12191_, _12177_, _04990_);
  or (_12192_, _12191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_12193_, _12192_, _12185_);
  nand (_12194_, _12191_, _06088_);
  and (_12195_, _12194_, _12193_);
  and (_12196_, _12183_, _06997_);
  or (_12197_, _12196_, _12195_);
  and (_10146_, _12197_, _04856_);
  not (_12198_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  not (_12199_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_12200_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_12201_, _12200_, _12199_);
  nor (_12202_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  nor (_12203_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_12204_, _12203_, _12202_);
  and (_12205_, _12204_, _12201_);
  and (_12206_, _12205_, _12198_);
  and (_12207_, _12206_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_12208_, _12207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_10174_, _12208_, _04856_);
  and (_12209_, _05940_, _05839_);
  and (_12210_, _05815_, _05866_);
  and (_12212_, _12210_, _12209_);
  and (_12213_, _05731_, _04856_);
  and (_12214_, _12213_, _05915_);
  and (_12215_, _12214_, _05891_);
  and (_12216_, _05763_, _05789_);
  and (_12217_, _12216_, _12215_);
  and (_10190_, _12217_, _12212_);
  and (_12218_, _06134_, _04932_);
  and (_12219_, _12218_, _06662_);
  not (_12220_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_12221_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_12222_, _12221_, _12220_);
  or (_12223_, _12222_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_12224_, _12223_, _12219_);
  not (_12225_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_12226_, _06146_, _12225_);
  nand (_12227_, _12226_, _12177_);
  or (_12228_, _12227_, _06147_);
  and (_12230_, _12228_, _12224_);
  or (_12231_, _12230_, _12183_);
  nand (_12232_, _12183_, _05287_);
  and (_12233_, _12232_, _04856_);
  and (_10193_, _12233_, _12231_);
  and (_12235_, _12177_, _06091_);
  or (_12236_, _12235_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_12237_, _12236_, _12185_);
  nand (_12238_, _12235_, _06088_);
  and (_12240_, _12238_, _12237_);
  and (_12241_, _12183_, _05718_);
  or (_12242_, _12241_, _12240_);
  and (_10199_, _12242_, _04856_);
  and (_12243_, _12219_, _07857_);
  and (_12244_, _12219_, _04984_);
  not (_12245_, _12219_);
  nor (_12246_, _04989_, _04984_);
  or (_12247_, _12246_, _12245_);
  or (_12248_, _12247_, _12244_);
  and (_12249_, _12248_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_12250_, _12249_, _12183_);
  or (_12252_, _12250_, _12243_);
  or (_12253_, _12185_, _06410_);
  and (_12254_, _12253_, _04856_);
  and (_10202_, _12254_, _12252_);
  and (_12256_, _12219_, _07642_);
  or (_12257_, _05519_, _06090_);
  not (_12258_, _12257_);
  and (_12259_, _12219_, _12258_);
  not (_12260_, _12259_);
  nand (_12261_, _12260_, _12244_);
  and (_12262_, _12261_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  or (_12263_, _12262_, _12183_);
  or (_12264_, _12263_, _12256_);
  nand (_12265_, _12183_, _05669_);
  and (_12266_, _12265_, _04856_);
  and (_10208_, _12266_, _12264_);
  and (_12268_, _06705_, _05009_);
  nor (_12269_, _05009_, _07113_);
  or (_12270_, _12269_, _12268_);
  and (_10214_, _12270_, _04856_);
  nor (_12271_, _08367_, _08257_);
  and (_12272_, _08160_, _08154_);
  nor (_12273_, _12272_, _08095_);
  and (_12275_, _08103_, _08098_);
  nor (_12276_, _12275_, _08154_);
  nor (_12277_, _12276_, _12273_);
  not (_12278_, _12277_);
  and (_12279_, _08160_, _08146_);
  nor (_12281_, _12279_, _08116_);
  and (_12282_, _12281_, _08106_);
  and (_12283_, _08113_, _08102_);
  nor (_12284_, _12283_, _08138_);
  nor (_12285_, _12284_, _08152_);
  not (_12286_, _12285_);
  and (_12287_, _08109_, _08104_);
  not (_12288_, _08095_);
  and (_12289_, _08113_, _08098_);
  nor (_12290_, _12289_, _08110_);
  nor (_12291_, _12290_, _12288_);
  nor (_12292_, _12291_, _12287_);
  and (_12293_, _12292_, _12286_);
  and (_12294_, _12293_, _12282_);
  and (_12296_, _12294_, _12278_);
  not (_12297_, _12283_);
  nor (_12298_, _08136_, _08126_);
  and (_12299_, _12298_, _12297_);
  nor (_12301_, _12299_, _08092_);
  not (_12302_, _12301_);
  nor (_12304_, _08173_, _08122_);
  and (_12305_, _12304_, _12302_);
  and (_12306_, _08102_, _08097_);
  not (_12307_, _12306_);
  nor (_12308_, _08157_, _08109_);
  nor (_12309_, _12308_, _12307_);
  not (_12310_, _08120_);
  or (_12311_, _12306_, _12283_);
  not (_12312_, _12311_);
  and (_12313_, _08135_, _08098_);
  nor (_12314_, _12313_, _08104_);
  and (_12315_, _12314_, _12312_);
  nor (_12316_, _12315_, _12310_);
  nor (_12318_, _12316_, _12309_);
  and (_12319_, _12318_, _12305_);
  not (_12320_, _08147_);
  and (_12321_, _08125_, _05895_);
  and (_12322_, _08171_, _12321_);
  and (_12323_, _08158_, _05843_);
  and (_12324_, _12323_, _08093_);
  nor (_12325_, _12324_, _12322_);
  and (_12326_, _12325_, _12320_);
  and (_12327_, _12326_, _08142_);
  and (_12328_, _08146_, _08094_);
  nor (_12329_, _12328_, _08120_);
  not (_12330_, _08126_);
  nor (_12331_, _08146_, _08099_);
  and (_12332_, _12331_, _12330_);
  nor (_12333_, _12332_, _12329_);
  not (_12334_, _12333_);
  and (_12335_, _12334_, _08134_);
  and (_12336_, _12335_, _12327_);
  and (_12337_, _08136_, _08120_);
  and (_12339_, _08157_, _08153_);
  nor (_12340_, _12339_, _12337_);
  nor (_12341_, _08119_, _08094_);
  not (_12342_, _12341_);
  and (_12344_, _12342_, _08131_);
  not (_12345_, _08157_);
  nor (_12346_, _08126_, _08114_);
  nor (_12347_, _12346_, _12345_);
  nor (_12348_, _12347_, _12344_);
  and (_12349_, _12348_, _12340_);
  nor (_12350_, _12298_, _12288_);
  nor (_12351_, _12350_, _08156_);
  and (_12352_, _08154_, _08117_);
  and (_12353_, _12352_, _12342_);
  nor (_12354_, _12313_, _12306_);
  nor (_12355_, _12354_, _12288_);
  nor (_12356_, _12355_, _12353_);
  and (_12357_, _12356_, _12351_);
  and (_12358_, _12357_, _12349_);
  and (_12359_, _12358_, _12336_);
  and (_12360_, _12359_, _12319_);
  and (_12361_, _12360_, _12296_);
  or (_12362_, _12361_, _05737_);
  and (_12363_, _08125_, _08112_);
  and (_12364_, _12363_, _08160_);
  or (_12365_, _12306_, _08153_);
  and (_12366_, _12365_, _08109_);
  or (_12367_, _12366_, _12350_);
  nor (_12368_, _12367_, _12364_);
  and (_12369_, _12368_, _12304_);
  nand (_12370_, _12369_, _12282_);
  or (_12371_, _12370_, _12361_);
  and (_12373_, _12371_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_12374_, _12361_, _05737_);
  and (_12375_, _12374_, _12362_);
  nand (_12376_, _12375_, _12373_);
  nand (_12377_, _12376_, _12362_);
  and (_12378_, _12377_, _05730_);
  and (_12379_, _12378_, _05736_);
  nor (_12380_, _12378_, _05736_);
  nor (_12381_, _12380_, _12379_);
  nor (_12382_, _12381_, _12271_);
  and (_12383_, _05741_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_12384_, _12383_, _12271_);
  and (_12385_, _12384_, _12370_);
  or (_12386_, _12385_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_12387_, _12386_, _12382_);
  and (_10221_, _12387_, _04856_);
  and (_12388_, _06125_, _06091_);
  and (_12389_, _12388_, _12182_);
  not (_12390_, _12389_);
  nor (_12391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_12392_, _12391_, _12221_);
  and (_12393_, _12392_, _07391_);
  and (_12394_, _12393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  not (_12395_, _12393_);
  and (_12396_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not (_12397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_12398_, \oc8051_top_1.oc8051_sfr1.pres_ow , _12397_);
  nor (_12399_, _12398_, _12396_);
  not (_12400_, _12399_);
  and (_12401_, _12400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_12402_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_12403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_12404_, _12403_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_12405_, _12404_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_12406_, _12405_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_12407_, _12406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_12408_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_12409_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_12410_, _12409_, _12408_);
  and (_12411_, _12410_, _12407_);
  and (_12412_, _12411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_12413_, _12412_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_12414_, _12413_, _12402_);
  and (_12415_, _12414_, _12401_);
  nand (_12416_, _12415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_12417_, _12415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_12418_, _12417_, _12416_);
  and (_12419_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_12420_, _12419_, _12414_);
  and (_12421_, _12391_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not (_12422_, _12421_);
  and (_12423_, _12422_, _12401_);
  and (_12424_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_12425_, _12424_, _12420_);
  or (_12426_, _12425_, _12418_);
  and (_12427_, _12426_, _12395_);
  or (_12428_, _12427_, _12394_);
  and (_12429_, _07855_, _06125_);
  and (_12430_, _12429_, _12182_);
  not (_12431_, _12430_);
  and (_12432_, _12431_, _12428_);
  and (_12433_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_12434_, _12433_, _12432_);
  and (_12435_, _12434_, _12390_);
  nor (_12436_, _12390_, _05287_);
  or (_12437_, _12436_, _12435_);
  and (_10247_, _12437_, _04856_);
  and (_12438_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  not (_12439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_12440_, _12413_, _12401_);
  and (_12441_, _12440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_12442_, _12441_, _12439_);
  and (_12443_, _12441_, _12439_);
  or (_12444_, _12443_, _12442_);
  and (_12446_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_12447_, _12446_, _12420_);
  or (_12448_, _12447_, _12393_);
  or (_12449_, _12448_, _12444_);
  not (_12450_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  nand (_12451_, _12393_, _12450_);
  and (_12452_, _12451_, _12449_);
  nor (_12453_, _12430_, _12389_);
  and (_12454_, _12453_, _12452_);
  and (_12455_, _12389_, _05718_);
  or (_12456_, _12455_, _12454_);
  or (_12457_, _12456_, _12438_);
  and (_10250_, _12457_, _04856_);
  or (_12458_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  nor (_12459_, _12440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  nor (_12460_, _12459_, _12441_);
  or (_12461_, _12460_, _12393_);
  and (_12462_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_12463_, _12462_, _12420_);
  or (_12464_, _12463_, _12461_);
  and (_12465_, _12464_, _12458_);
  and (_12466_, _12465_, _12453_);
  and (_12467_, _12389_, _06410_);
  and (_12468_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_12469_, _12468_, _12467_);
  or (_12470_, _12469_, _12466_);
  and (_10257_, _12470_, _04856_);
  and (_10265_, _07384_, _04856_);
  and (_10297_, _07365_, _04856_);
  and (_10301_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _04856_);
  not (_12471_, _06809_);
  and (_12472_, _08217_, _06858_);
  and (_12473_, _12472_, _12471_);
  nor (_12474_, _12473_, _05994_);
  and (_12475_, _12474_, _06810_);
  nor (_12476_, _06268_, _06124_);
  and (_12477_, _12476_, _07996_);
  and (_12478_, _12477_, _12475_);
  not (_12479_, _12478_);
  nor (_12480_, _08206_, _05874_);
  not (_12481_, _12474_);
  not (_12483_, _07789_);
  and (_12484_, _07680_, _05617_);
  and (_12486_, _12484_, _05597_);
  and (_12487_, _12486_, _06508_);
  and (_12488_, _12487_, _06561_);
  and (_12490_, _12488_, _06810_);
  and (_12492_, _12490_, _12483_);
  and (_12494_, _12492_, _12481_);
  and (_12495_, _12494_, _07871_);
  and (_12497_, _12495_, _05634_);
  not (_12498_, _12497_);
  and (_12499_, _12475_, _06062_);
  nor (_12500_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_12501_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_12502_, _12501_, _12500_);
  nor (_12503_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_12504_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_12505_, _12504_, _12503_);
  and (_12506_, _12505_, _12502_);
  and (_12507_, _12506_, _06807_);
  and (_12508_, _06809_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_12509_, _12508_, _12507_);
  not (_12510_, _12509_);
  nor (_12511_, _12510_, _12499_);
  and (_12512_, _12511_, _12498_);
  or (_12513_, _12512_, _08218_);
  nor (_12514_, _12513_, _12480_);
  or (_12515_, _06635_, _06737_);
  and (_12516_, _12515_, _05983_);
  not (_12517_, _12516_);
  not (_12518_, _07511_);
  nor (_12519_, _09066_, _06610_);
  and (_12520_, _12519_, _12518_);
  and (_12521_, _06638_, _06612_);
  nor (_12522_, _12521_, _08214_);
  and (_12523_, _12522_, _12520_);
  and (_12524_, _12523_, _12517_);
  and (_12525_, _12524_, _12512_);
  nor (_12526_, _12525_, _12514_);
  nor (_12527_, _08213_, _09088_);
  and (_12528_, _12527_, _06824_);
  not (_12529_, _12528_);
  nor (_12530_, _12529_, _12526_);
  nor (_12531_, _12530_, _06647_);
  and (_12532_, _05949_, _05849_);
  nor (_12533_, _12532_, _05954_);
  nor (_12534_, _06799_, _12533_);
  nor (_12535_, _12534_, _06847_);
  not (_12536_, _12535_);
  nor (_12537_, _12536_, _12531_);
  not (_12538_, _06807_);
  nor (_12539_, _12538_, _06678_);
  nor (_12540_, _08277_, _07951_);
  and (_12541_, _12540_, _06935_);
  nor (_12542_, _12541_, _12471_);
  nor (_12543_, _12542_, _12539_);
  not (_12544_, _12543_);
  nor (_12545_, _12544_, _12537_);
  and (_12546_, _12545_, _07993_);
  and (_12547_, _12546_, _12479_);
  nand (_12548_, _12547_, _06901_);
  nor (_10310_, _12548_, rst);
  not (_12549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nand (_12550_, _12393_, _12549_);
  and (_12551_, _12407_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_12552_, _12551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_12553_, _12552_, _12401_);
  and (_12554_, _12553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nand (_12555_, _12554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_12556_, _12554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_12557_, _12556_, _12555_);
  or (_12558_, _12557_, _12393_);
  and (_12559_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_12560_, _12559_, _12420_);
  or (_12561_, _12560_, _12558_);
  and (_12562_, _12561_, _12550_);
  and (_12563_, _12562_, _12453_);
  nor (_12564_, _12390_, _06032_);
  and (_12565_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_12566_, _12565_, _12564_);
  or (_12567_, _12566_, _12563_);
  and (_10337_, _12567_, _04856_);
  or (_12568_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_12569_, _12553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor (_12570_, _12569_, _12554_);
  or (_12571_, _12570_, _12393_);
  and (_12572_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_12573_, _12572_, _12420_);
  or (_12574_, _12573_, _12571_);
  and (_12575_, _12574_, _12568_);
  and (_12576_, _12575_, _12453_);
  and (_12577_, _12389_, _06997_);
  and (_12578_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_12579_, _12578_, _12577_);
  or (_12581_, _12579_, _12576_);
  and (_10344_, _12581_, _04856_);
  or (_12582_, _12401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_12583_, _12401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_12584_, _12422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_12585_, _12584_, _12420_);
  nand (_12586_, _12585_, _12583_);
  and (_12587_, _12586_, _12582_);
  or (_12588_, _12587_, _12393_);
  nor (_12589_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nor (_12590_, _12589_, _12430_);
  and (_12591_, _12590_, _12588_);
  and (_12592_, _12430_, _06997_);
  or (_12593_, _12592_, _12389_);
  or (_12594_, _12593_, _12591_);
  or (_12595_, _12390_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_12596_, _12595_, _04856_);
  and (_10374_, _12596_, _12594_);
  nor (_12597_, _12431_, _05287_);
  or (_12598_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_12599_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_12600_, _12599_, _12420_);
  and (_12601_, _12407_, _12401_);
  and (_12602_, _12601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_12603_, _12601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_12604_, _12603_, _12602_);
  or (_12605_, _12604_, _12393_);
  or (_12606_, _12605_, _12600_);
  nand (_12607_, _12606_, _12598_);
  nor (_12608_, _12607_, _12430_);
  or (_12609_, _12608_, _12389_);
  or (_12610_, _12609_, _12597_);
  or (_12611_, _12390_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_12612_, _12611_, _04856_);
  and (_10416_, _12612_, _12610_);
  or (_12613_, _12431_, _05718_);
  and (_12614_, _12406_, _12401_);
  nor (_12615_, _12614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nor (_12616_, _12615_, _12601_);
  and (_12617_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_12618_, _12617_, _12420_);
  or (_12619_, _12618_, _12616_);
  and (_12620_, _12619_, _12395_);
  and (_12622_, _12393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_12623_, _12622_, _12620_);
  or (_12624_, _12623_, _12430_);
  and (_12625_, _12624_, _12613_);
  or (_12626_, _12625_, _12389_);
  not (_12627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand (_12628_, _12389_, _12627_);
  and (_12629_, _12628_, _04856_);
  and (_10419_, _12629_, _12626_);
  or (_12630_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_12631_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_12632_, _12631_, _12420_);
  not (_12633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand (_12634_, _12405_, _12401_);
  and (_12635_, _12634_, _12633_);
  nor (_12636_, _12635_, _12614_);
  or (_12637_, _12636_, _12393_);
  or (_12638_, _12637_, _12632_);
  and (_12639_, _12638_, _12630_);
  or (_12640_, _12639_, _12430_);
  or (_12641_, _12431_, _06410_);
  and (_12642_, _12641_, _12640_);
  or (_12643_, _12642_, _12389_);
  nand (_12644_, _12389_, _12633_);
  and (_12645_, _12644_, _04856_);
  and (_10424_, _12645_, _12643_);
  and (_12647_, _12404_, _12401_);
  or (_12648_, _12647_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_12649_, _12648_, _12634_);
  and (_12650_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_12651_, _12650_, _12420_);
  or (_12652_, _12651_, _12649_);
  and (_12653_, _12652_, _12395_);
  and (_12654_, _12393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_12655_, _12654_, _12653_);
  or (_12656_, _12655_, _12430_);
  nand (_12657_, _12430_, _05669_);
  and (_12658_, _12657_, _12656_);
  or (_12659_, _12658_, _12389_);
  nand (_12660_, _12389_, _08788_);
  and (_12661_, _12660_, _04856_);
  and (_10427_, _12661_, _12659_);
  and (_12662_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_12663_, _12662_, _12420_);
  nand (_12664_, _12403_, _12401_);
  and (_12665_, _12664_, _08898_);
  nor (_12666_, _12665_, _12647_);
  or (_12667_, _12666_, _12393_);
  or (_12668_, _12667_, _12663_);
  or (_12669_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  nand (_12671_, _12669_, _12668_);
  nor (_12672_, _12671_, _12430_);
  and (_12674_, _12430_, _06705_);
  or (_12675_, _12674_, _12389_);
  or (_12676_, _12675_, _12672_);
  nand (_12677_, _12389_, _08898_);
  and (_12678_, _12677_, _04856_);
  and (_10434_, _12678_, _12676_);
  and (_12680_, _06721_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_12681_, _08197_, _06878_);
  and (_12682_, _06594_, _05998_);
  or (_12683_, _12682_, _06726_);
  and (_12684_, _08198_, _05773_);
  or (_12685_, _06625_, _12684_);
  or (_12686_, _12685_, _12683_);
  or (_12687_, _12686_, _12681_);
  or (_12688_, _06865_, _06729_);
  and (_12689_, _06624_, _06731_);
  and (_12691_, _06745_, _06598_);
  or (_12692_, _12691_, _12689_);
  or (_12693_, _12692_, _12688_);
  and (_12695_, _06857_, _06598_);
  or (_12696_, _08193_, _12695_);
  and (_12697_, _06598_, _06612_);
  or (_12698_, _08246_, _06789_);
  or (_12699_, _12698_, _12697_);
  or (_12700_, _12699_, _12696_);
  and (_12701_, _06857_, _06638_);
  or (_12703_, _09075_, _06628_);
  or (_12704_, _12703_, _12701_);
  or (_12705_, _06835_, _06746_);
  or (_12707_, _12705_, _12704_);
  or (_12708_, _12707_, _12700_);
  or (_12709_, _12708_, _12693_);
  or (_12710_, _12709_, _12687_);
  and (_12711_, _12710_, _06770_);
  or (_10443_, _12711_, _12680_);
  and (_12713_, _06125_, _05520_);
  and (_12714_, _12713_, _12182_);
  not (_12715_, _12714_);
  and (_12716_, _12421_, _12221_);
  not (_12717_, _12716_);
  and (_12718_, _06494_, _06125_);
  and (_12719_, _12718_, _12182_);
  nor (_12720_, _12719_, _12717_);
  or (_12721_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nand (_12722_, _12720_, _08901_);
  and (_12723_, _12722_, _12721_);
  and (_12724_, _12723_, _12715_);
  and (_12725_, _12714_, _06705_);
  or (_12726_, _12725_, _12724_);
  and (_10471_, _12726_, _04856_);
  or (_12727_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  not (_12728_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nand (_12729_, _12720_, _12728_);
  and (_12730_, _12729_, _12727_);
  or (_12731_, _12730_, _12714_);
  nand (_12732_, _12714_, _06032_);
  and (_12733_, _12732_, _04856_);
  and (_10473_, _12733_, _12731_);
  or (_12734_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  not (_12735_, _12720_);
  or (_12737_, _12735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_12738_, _12737_, _12734_);
  or (_12739_, _12738_, _12714_);
  nand (_12740_, _12714_, _06369_);
  and (_12741_, _12740_, _04856_);
  and (_10478_, _12741_, _12739_);
  and (_12742_, _12735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_12743_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_12744_, _12743_, _12742_);
  and (_12745_, _12744_, _12715_);
  and (_12746_, _12714_, _06410_);
  or (_12747_, _12746_, _12745_);
  and (_10499_, _12747_, _04856_);
  nand (_12748_, _12714_, _05287_);
  and (_12749_, _12735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  and (_12751_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_12752_, _12751_, _12749_);
  or (_12753_, _12752_, _12714_);
  and (_12754_, _12753_, _04856_);
  and (_10507_, _12754_, _12748_);
  or (_12755_, _12715_, _05718_);
  nor (_12756_, _12720_, _12450_);
  and (_12757_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_12758_, _12757_, _12756_);
  or (_12759_, _12758_, _12714_);
  and (_12760_, _12759_, _04856_);
  and (_10514_, _12760_, _12755_);
  nor (_12761_, _10231_, _10232_);
  and (_12762_, _08067_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_12763_, _12762_, _10230_);
  or (_12764_, _12763_, _12761_);
  and (_12765_, _12764_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_12766_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _09249_);
  nand (_12767_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_12768_, _12767_, _08087_);
  or (_12769_, _12768_, _12766_);
  or (_12770_, _12769_, _12765_);
  and (_10531_, _12770_, _04856_);
  not (_12771_, _12719_);
  or (_12772_, _12771_, _06705_);
  and (_12773_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_12774_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  or (_12775_, _12774_, _12773_);
  or (_12776_, _12775_, _12719_);
  and (_12777_, _12776_, _12715_);
  and (_12778_, _12777_, _12772_);
  and (_12779_, _12714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_12780_, _12779_, _12778_);
  and (_10547_, _12780_, _04856_);
  nor (_12781_, _12771_, _05287_);
  and (_12782_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_12783_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_12784_, _12783_, _12782_);
  nor (_12785_, _12784_, _12719_);
  or (_12786_, _12785_, _12714_);
  or (_12787_, _12786_, _12781_);
  or (_12788_, _12715_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_12789_, _12788_, _04856_);
  and (_10549_, _12789_, _12787_);
  or (_12790_, _12771_, _05718_);
  not (_12791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  nor (_12792_, _12716_, _12791_);
  and (_12793_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_12794_, _12793_, _12792_);
  or (_12795_, _12794_, _12719_);
  and (_12796_, _12795_, _12715_);
  and (_12797_, _12796_, _12790_);
  and (_12798_, _12714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  or (_12799_, _12798_, _12797_);
  and (_10553_, _12799_, _04856_);
  or (_12800_, _12771_, _06410_);
  and (_12801_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_12802_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_12803_, _12802_, _12801_);
  or (_12804_, _12803_, _12719_);
  and (_12805_, _12804_, _12715_);
  and (_12806_, _12805_, _12800_);
  and (_12807_, _12714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_12808_, _12807_, _12806_);
  and (_10557_, _12808_, _04856_);
  nand (_12809_, _12719_, _05669_);
  and (_12810_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_12811_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_12812_, _12811_, _12810_);
  or (_12813_, _12812_, _12719_);
  and (_12814_, _12813_, _12715_);
  and (_12815_, _12814_, _12809_);
  and (_12816_, _12714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_12817_, _12816_, _12815_);
  and (_10566_, _12817_, _04856_);
  nor (_12818_, _12761_, _09249_);
  or (_12820_, _12818_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_12821_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _09249_);
  or (_12822_, _12821_, _08087_);
  and (_12823_, _12822_, _04856_);
  and (_10761_, _12823_, _12820_);
  and (_10850_, _05847_, _04856_);
  not (_12824_, _05823_);
  and (_12825_, _06612_, _12824_);
  nor (_12826_, _12825_, _06610_);
  nand (_12827_, _12826_, _12472_);
  nand (_12828_, _12827_, _05959_);
  and (_12829_, _05962_, _12532_);
  not (_12830_, _12829_);
  and (_12831_, _06822_, _05962_);
  and (_12832_, _12831_, _05983_);
  nor (_12833_, _12832_, _06847_);
  and (_12834_, _12833_, _12830_);
  nand (_12835_, _12834_, _12828_);
  or (_12836_, _12835_, _07261_);
  and (_12837_, _12834_, _12828_);
  nor (_12838_, _05730_, _05177_);
  and (_12839_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12840_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  and (_12841_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_12842_, _12841_, _12840_);
  and (_12843_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_12844_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_12845_, _12844_, _12843_);
  and (_12846_, _12845_, _12842_);
  and (_12847_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_12848_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_12849_, _12848_, _12847_);
  and (_12850_, _12849_, _12846_);
  nor (_12851_, _12850_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12852_, _12851_, _12839_);
  nor (_12853_, _12852_, _08257_);
  nor (_12854_, _12853_, _12838_);
  or (_12855_, _12854_, _12837_);
  and (_12856_, _12855_, _12836_);
  or (_12857_, _12856_, _05183_);
  nand (_12858_, _12856_, _05183_);
  and (_12859_, _12858_, _12857_);
  not (_12860_, _07191_);
  and (_12861_, _12837_, _12860_);
  nor (_12862_, _05730_, _05060_);
  and (_12863_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12864_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_12865_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_12866_, _12865_, _12864_);
  and (_12867_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_12868_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nor (_12869_, _12868_, _12867_);
  and (_12870_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  and (_12871_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  nor (_12872_, _12871_, _12870_);
  and (_12873_, _12872_, _12869_);
  and (_12874_, _12873_, _12866_);
  nor (_12875_, _12874_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12876_, _12875_, _12863_);
  nor (_12877_, _12876_, _08257_);
  nor (_12878_, _12877_, _12862_);
  not (_12879_, _12878_);
  and (_12880_, _12879_, _12835_);
  nor (_12881_, _12880_, _12861_);
  not (_12882_, _12881_);
  and (_12883_, _12882_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  not (_12884_, _12883_);
  not (_12885_, _07142_);
  and (_12886_, _12837_, _12885_);
  nor (_12887_, _05730_, _05082_);
  and (_12888_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12889_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  and (_12890_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_12891_, _12890_, _12889_);
  and (_12892_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_12893_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_12894_, _12893_, _12892_);
  and (_12895_, _12894_, _12891_);
  and (_12896_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_12897_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_12898_, _12897_, _12896_);
  and (_12899_, _12898_, _12895_);
  nor (_12900_, _12899_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12901_, _12900_, _12888_);
  nor (_12902_, _12901_, _08257_);
  nor (_12903_, _12902_, _12887_);
  not (_12904_, _12903_);
  and (_12905_, _12904_, _12835_);
  nor (_12906_, _12905_, _12886_);
  and (_12907_, _12906_, _05087_);
  nor (_12908_, _12906_, _05087_);
  or (_12909_, _12835_, _07089_);
  nor (_12910_, _05730_, _05154_);
  and (_12911_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12912_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_12913_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_12914_, _12913_, _12912_);
  and (_12915_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_12916_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_12917_, _12916_, _12915_);
  and (_12918_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_12919_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_12920_, _12919_, _12918_);
  and (_12921_, _12920_, _12917_);
  and (_12922_, _12921_, _12914_);
  nor (_12923_, _12922_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12924_, _12923_, _12911_);
  nor (_12925_, _12924_, _08257_);
  nor (_12926_, _12925_, _12910_);
  or (_12927_, _12926_, _12837_);
  and (_12928_, _12927_, _12909_);
  or (_12929_, _12928_, _05159_);
  not (_12930_, _12929_);
  not (_12931_, _07032_);
  or (_12932_, _12835_, _12931_);
  nor (_12933_, _05730_, _05135_);
  and (_12934_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12935_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  and (_12936_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_12937_, _12936_, _12935_);
  and (_12938_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_12939_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_12940_, _12939_, _12938_);
  and (_12941_, _12940_, _12937_);
  and (_12942_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_12943_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_12944_, _12943_, _12942_);
  and (_12945_, _12944_, _12941_);
  nor (_12946_, _12945_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12947_, _12946_, _12934_);
  nor (_12948_, _12947_, _08257_);
  nor (_12949_, _12948_, _12933_);
  nand (_12950_, _12949_, _12835_);
  and (_12952_, _12950_, _12932_);
  nand (_12953_, _12952_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_12954_, _06925_);
  and (_12955_, _12837_, _12954_);
  nor (_12956_, _05730_, _05106_);
  and (_12957_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12958_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_12959_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_12960_, _12959_, _12958_);
  and (_12961_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_12962_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_12963_, _12962_, _12961_);
  and (_12964_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_12965_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_12966_, _12965_, _12964_);
  and (_12967_, _12966_, _12963_);
  and (_12968_, _12967_, _12960_);
  nor (_12969_, _12968_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12970_, _12969_, _12957_);
  nor (_12971_, _12970_, _08257_);
  nor (_12972_, _12971_, _12956_);
  not (_12973_, _12972_);
  and (_12974_, _12973_, _12835_);
  or (_12975_, _12974_, _12955_);
  and (_12976_, _12975_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_12977_, _12952_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_12978_, _12977_, _12953_);
  and (_12979_, _12978_, _12976_);
  not (_12980_, _12979_);
  nand (_12981_, _12980_, _12953_);
  nand (_12982_, _12928_, _05159_);
  and (_12983_, _12982_, _12929_);
  and (_12984_, _12983_, _12981_);
  or (_12985_, _12984_, _12930_);
  nor (_12986_, _12985_, _12908_);
  nor (_12987_, _12986_, _12907_);
  nor (_12988_, _12882_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_12989_, _12988_, _12883_);
  nand (_12990_, _12989_, _12987_);
  nand (_12991_, _12990_, _12884_);
  and (_12992_, _12991_, _12859_);
  not (_12993_, _12992_);
  nand (_12994_, _12993_, _12857_);
  not (_12995_, _07294_);
  and (_12996_, _12837_, _12995_);
  nor (_12997_, _05730_, _05011_);
  and (_12998_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12999_, _05929_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_13000_, _05742_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_13001_, _13000_, _12999_);
  and (_13003_, _05933_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_13004_, _05935_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_13005_, _13004_, _13003_);
  and (_13006_, _13005_, _13001_);
  and (_13007_, _05927_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_13008_, _05758_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_13009_, _13008_, _13007_);
  and (_13010_, _13009_, _13006_);
  nor (_13011_, _13010_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_13012_, _13011_, _12998_);
  nor (_13013_, _13012_, _08257_);
  nor (_13014_, _13013_, _12997_);
  nor (_13015_, _13014_, _12837_);
  nor (_13016_, _13015_, _12996_);
  nor (_13017_, _13016_, _05026_);
  and (_13018_, _13016_, _05026_);
  nor (_13019_, _13018_, _13017_);
  nand (_13020_, _13019_, _12994_);
  or (_13021_, _13019_, _12994_);
  and (_13022_, _09088_, _05959_);
  nor (_13023_, _13022_, _12534_);
  or (_13024_, _13023_, _12835_);
  nor (_13025_, _12521_, _08207_);
  and (_13026_, _13025_, _12472_);
  and (_13027_, _12527_, _12520_);
  and (_13028_, _13027_, _13026_);
  nor (_13029_, _13028_, _06647_);
  or (_13030_, _13029_, _12832_);
  and (_13031_, _13030_, _13024_);
  and (_13032_, _13031_, _13021_);
  and (_13033_, _13032_, _13020_);
  not (_13034_, _06488_);
  nor (_13035_, _13030_, _12835_);
  and (_13036_, _13035_, _13023_);
  or (_13037_, _13036_, _13022_);
  and (_13038_, _13037_, _13034_);
  and (_13039_, _05983_, _05962_);
  and (_13040_, _13039_, _06822_);
  or (_13041_, _13029_, _13040_);
  nor (_13042_, _13041_, _13024_);
  and (_13043_, _13042_, _12995_);
  and (_13044_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_13045_, _13015_, _12534_);
  or (_13046_, _13045_, _13044_);
  or (_13047_, _13046_, _13043_);
  or (_13048_, _13047_, _13038_);
  or (_13049_, _13048_, _13033_);
  and (_13050_, _13049_, _12547_);
  and (_13051_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_13052_, _13051_, _08368_);
  and (_13053_, _13052_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_13055_, _13053_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_13056_, _13053_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_13057_, _13056_, _13055_);
  nor (_13058_, _13057_, _12547_);
  or (_13059_, _13058_, _13050_);
  and (_10866_, _13059_, _04856_);
  not (_13060_, _07897_);
  and (_13061_, _13037_, _13060_);
  nor (_13062_, _12854_, _12830_);
  not (_13063_, _07261_);
  and (_13065_, _13042_, _13063_);
  and (_13066_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_13067_, _13066_, _13065_);
  or (_13068_, _13067_, _13062_);
  or (_13069_, _13068_, _13061_);
  and (_13070_, _13041_, _13024_);
  nor (_13071_, _12991_, _12859_);
  nor (_13072_, _13071_, _12992_);
  and (_13073_, _13072_, _13070_);
  or (_13074_, _13073_, _13069_);
  and (_13075_, _13074_, _12547_);
  nor (_13076_, _13052_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_13077_, _13076_, _13053_);
  nor (_13078_, _13077_, _12547_);
  or (_13079_, _13078_, _13075_);
  and (_10869_, _13079_, _04856_);
  nor (_10883_, _13014_, rst);
  nor (_13080_, _07774_, _06901_);
  and (_13081_, _12829_, _12931_);
  or (_13082_, _13081_, _13080_);
  and (_13083_, _13042_, _05943_);
  and (_13084_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_13085_, _13084_, _13083_);
  or (_13086_, _13085_, _13082_);
  not (_13087_, _07380_);
  and (_13088_, _12837_, _13087_);
  not (_13089_, _08273_);
  and (_13090_, _12835_, _13089_);
  nor (_13091_, _13090_, _13088_);
  not (_13092_, _13091_);
  nor (_13093_, _13091_, _05327_);
  not (_13094_, _13017_);
  and (_13095_, _13091_, _05327_);
  nor (_13096_, _13095_, _13094_);
  nor (_13097_, _13096_, _13093_);
  nand (_13098_, _12883_, _12859_);
  nand (_13099_, _13098_, _12857_);
  nor (_13100_, _13095_, _13093_);
  and (_13101_, _13100_, _13019_);
  nand (_13102_, _13101_, _13099_);
  and (_13103_, _13102_, _13097_);
  and (_13104_, _12989_, _12859_);
  and (_13105_, _13101_, _13104_);
  nand (_13106_, _13105_, _12987_);
  and (_13107_, _13106_, _13103_);
  and (_13108_, _13107_, _05111_);
  and (_13109_, _13108_, _13092_);
  nor (_13110_, _13107_, _05111_);
  and (_13111_, _13110_, _13091_);
  nor (_13112_, _13111_, _13109_);
  nand (_13113_, _13112_, _05142_);
  or (_13114_, _13112_, _05142_);
  and (_13115_, _13114_, _13070_);
  and (_13116_, _13115_, _13113_);
  or (_13117_, _13116_, _13086_);
  nand (_13118_, _13022_, _07743_);
  nand (_13119_, _13118_, _12547_);
  or (_13120_, _13119_, _13117_);
  and (_13121_, _13055_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_13122_, _13121_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_13123_, _13122_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_13124_, _13122_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_13125_, _13124_, _13123_);
  or (_13126_, _13125_, _12547_);
  and (_13127_, _13126_, _04856_);
  and (_10889_, _13127_, _13120_);
  and (_13128_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_13129_, _06370_, _05679_);
  or (_13130_, _13129_, _13128_);
  and (_10893_, _13130_, _04856_);
  and (_13131_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_13132_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or (_13133_, _13132_, _13131_);
  and (_10902_, _13133_, _04856_);
  or (_13134_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  nand (_13135_, _08367_, _05861_);
  and (_13136_, _13135_, _04856_);
  and (_10908_, _13136_, _13134_);
  nor (_13137_, _13121_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_13138_, _13137_, _13122_);
  or (_13139_, _13138_, _12547_);
  and (_13140_, _13139_, _04856_);
  nor (_13141_, _13107_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_13142_, _13107_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_13143_, _13142_, _13141_);
  nor (_13144_, _13143_, _13092_);
  and (_13145_, _13143_, _13092_);
  or (_13146_, _13145_, _13144_);
  and (_13147_, _13146_, _13031_);
  and (_13148_, _13022_, _07676_);
  and (_13149_, _13042_, _05895_);
  and (_13150_, _12829_, _12954_);
  or (_13151_, _13150_, _13149_);
  and (_13152_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  not (_13153_, _07702_);
  and (_13154_, _13153_, _06847_);
  or (_13155_, _13154_, _13152_);
  or (_13156_, _13155_, _13151_);
  nor (_13157_, _13156_, _13148_);
  nand (_13159_, _13157_, _12547_);
  or (_13160_, _13159_, _13147_);
  and (_10911_, _13160_, _13140_);
  and (_13161_, _13020_, _13094_);
  nor (_13162_, _13161_, _13100_);
  and (_13163_, _13161_, _13100_);
  or (_13164_, _13163_, _13162_);
  and (_13166_, _13164_, _13031_);
  and (_13167_, _13037_, _05641_);
  and (_13169_, _12829_, _13089_);
  and (_13170_, _13088_, _12534_);
  and (_13171_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_13172_, _13171_, _13170_);
  or (_13173_, _13172_, _13169_);
  or (_13174_, _13173_, _13167_);
  or (_13175_, _13174_, _13166_);
  and (_13176_, _13175_, _12547_);
  nor (_13177_, _13055_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  or (_13178_, _13177_, _13121_);
  nor (_13179_, _13178_, _12547_);
  or (_13180_, _13179_, _13176_);
  and (_10919_, _13180_, _04856_);
  and (_13181_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _04856_);
  and (_13182_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _04856_);
  and (_13183_, _13182_, _12206_);
  or (_10992_, _13183_, _13181_);
  and (_11042_, _05772_, _04856_);
  and (_13184_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_13185_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or (_13186_, _13185_, _13184_);
  and (_11055_, _13186_, _04856_);
  and (_13187_, _12371_, _05730_);
  nand (_13189_, _13187_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_13190_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  or (_13191_, _13187_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_13192_, _13191_, _13190_);
  and (_11058_, _13192_, _13189_);
  or (_13193_, _12375_, _12373_);
  and (_13194_, _13193_, _12376_);
  or (_13195_, _13194_, _08257_);
  or (_13197_, _05730_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_13198_, _13197_, _13190_);
  and (_11089_, _13198_, _13195_);
  nor (_11150_, _07089_, rst);
  nor (_11174_, _07032_, rst);
  nand (_13199_, _12171_, _06586_);
  or (_13200_, _12171_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_13201_, _13200_, _04856_);
  and (_11236_, _13201_, _13199_);
  nand (_13202_, _12171_, _07702_);
  or (_13204_, _12171_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_13206_, _13204_, _04856_);
  and (_11247_, _13206_, _13202_);
  and (_13207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _04856_);
  and (_13208_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _04856_);
  and (_13209_, _13208_, _12206_);
  or (_11312_, _13209_, _13207_);
  and (_13210_, _12205_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_13211_, _13210_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_11327_, _13211_, _04856_);
  and (_13212_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_13214_, _12165_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_13215_, _13214_, _13212_);
  and (_11343_, _13215_, _04856_);
  or (_13216_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_13217_, _08367_, _05774_);
  and (_13218_, _13217_, _04856_);
  and (_11347_, _13218_, _13216_);
  and (_13219_, _08277_, _05520_);
  nand (_13220_, _13219_, _06088_);
  or (_13221_, _13219_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_13222_, _13221_, _06935_);
  and (_13223_, _13222_, _13220_);
  or (_13224_, _13223_, _06946_);
  and (_11350_, _13224_, _04856_);
  or (_13225_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand (_13226_, _08367_, _05911_);
  and (_13227_, _13226_, _04856_);
  and (_11355_, _13227_, _13225_);
  or (_13228_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nand (_13229_, _08367_, _05811_);
  and (_13230_, _13229_, _04856_);
  and (_11357_, _13230_, _13228_);
  or (_13231_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand (_13232_, _08367_, _05735_);
  and (_13233_, _13232_, _04856_);
  and (_11370_, _13233_, _13231_);
  and (_13234_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_13235_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  and (_13236_, _13235_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_13237_, _13235_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_00001_, _13237_, _13236_);
  or (_00002_, _00001_, _13234_);
  and (_11406_, _00002_, _04856_);
  and (_00003_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _08359_);
  and (_00004_, \oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00005_, _00004_, _00003_);
  and (_11412_, _00005_, _04856_);
  nor (_11426_, _12903_, rst);
  nor (_11428_, _12972_, rst);
  and (_00006_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_00007_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_00008_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_00009_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_00010_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_00011_, _00010_, _00008_);
  and (_00012_, _00011_, _00009_);
  nor (_00013_, _00012_, _00008_);
  not (_00014_, _00013_);
  nor (_00015_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_00016_, _00015_, _00007_);
  and (_00017_, _00016_, _00014_);
  nor (_00018_, _00017_, _00007_);
  nor (_00019_, _00018_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_00020_, _00018_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_00021_, _00020_, _00019_);
  not (_00022_, _12361_);
  nor (_00023_, _00011_, _00009_);
  nor (_00024_, _00023_, _00012_);
  nand (_00025_, _00024_, _00022_);
  nor (_00026_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_00027_, _00026_, _00009_);
  and (_00028_, _00027_, _12371_);
  or (_00029_, _00024_, _00022_);
  and (_00030_, _00029_, _00025_);
  nand (_00031_, _00030_, _00028_);
  nand (_00032_, _00031_, _00025_);
  nor (_00033_, _00016_, _00014_);
  nor (_00034_, _00033_, _00017_);
  and (_00035_, _00034_, _00032_);
  and (_00036_, _00035_, _00021_);
  nor (_00037_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00038_, _00037_, _13051_);
  nand (_00039_, _00038_, _00019_);
  or (_00040_, _00038_, _00019_);
  and (_00042_, _00040_, _00039_);
  not (_00043_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_00044_, _00037_, _00043_);
  and (_00045_, _00018_, _00044_);
  nand (_00046_, _00018_, _00037_);
  and (_00047_, _00046_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  or (_00048_, _00047_, _00045_);
  and (_00049_, _00048_, _00042_);
  and (_00050_, _00049_, _00036_);
  not (_00051_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_00052_, _00045_, _00051_);
  and (_00053_, _00045_, _00051_);
  or (_00054_, _00053_, _00052_);
  and (_00055_, _00054_, _00050_);
  nor (_00056_, _00054_, _00050_);
  nor (_00057_, _00056_, _00055_);
  or (_00058_, _00057_, _06911_);
  not (_00059_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00060_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_00061_, _00060_, _00059_);
  and (_00062_, _00061_, _00058_);
  or (_00063_, _00062_, _00006_);
  and (_11435_, _00063_, _04856_);
  and (_00064_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  nor (_00065_, _08367_, _05803_);
  or (_00066_, _00065_, _00064_);
  and (_11439_, _00066_, _04856_);
  and (_00067_, _00042_, _00036_);
  or (_00068_, _00048_, _00067_);
  nor (_00069_, _00050_, _06911_);
  and (_00070_, _00069_, _00068_);
  nor (_00071_, _06910_, _05183_);
  or (_00072_, _00071_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00073_, _00072_, _00070_);
  or (_00074_, _00059_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_00075_, _00074_, _04856_);
  and (_11443_, _00075_, _00073_);
  and (_00076_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_00077_, _08367_, _05754_);
  or (_00078_, _00077_, _00076_);
  and (_11451_, _00078_, _04856_);
  and (_00079_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_00080_, _08367_, _05850_);
  or (_00081_, _00080_, _00079_);
  and (_11464_, _00081_, _04856_);
  nor (_00082_, _00042_, _00036_);
  nor (_00083_, _00082_, _00067_);
  or (_00084_, _00083_, _06911_);
  or (_00085_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_00086_, _00085_, _00059_);
  and (_00087_, _00086_, _00084_);
  and (_00088_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00089_, _00088_, _00087_);
  and (_11467_, _00089_, _04856_);
  and (_00090_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  nor (_00091_, _08367_, _05824_);
  or (_00092_, _00091_, _00090_);
  and (_11476_, _00092_, _04856_);
  and (_00093_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_00094_, _00035_, _00021_);
  nor (_00095_, _00094_, _00036_);
  or (_00096_, _00095_, _06911_);
  or (_00097_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_00098_, _00097_, _00059_);
  and (_00099_, _00098_, _00096_);
  or (_00100_, _00099_, _00093_);
  and (_11522_, _00100_, _04856_);
  and (_00101_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_00102_, _00034_, _00032_);
  nor (_00103_, _00102_, _00035_);
  or (_00104_, _00103_, _06911_);
  or (_00105_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_00106_, _00105_, _00059_);
  and (_00107_, _00106_, _00104_);
  or (_00108_, _00107_, _00101_);
  and (_11543_, _00108_, _04856_);
  or (_00109_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  nand (_00110_, _08367_, _05855_);
  and (_00111_, _00110_, _04856_);
  and (_11565_, _00111_, _00109_);
  and (_00112_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _08359_);
  and (_00113_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00114_, _00113_, _00112_);
  and (_11579_, _00114_, _04856_);
  nor (_11595_, _12878_, rst);
  and (_00117_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_00118_, _08367_, _05861_);
  or (_00119_, _00118_, _00117_);
  and (_11598_, _00119_, _04856_);
  and (_00120_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nor (_00122_, _08367_, _05881_);
  or (_00123_, _00122_, _00120_);
  and (_11602_, _00123_, _04856_);
  and (_00125_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_00127_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_00128_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  not (_00129_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_00131_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_00132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_00134_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_00135_, _00044_, _00051_);
  and (_00136_, _00135_, _00134_);
  and (_00138_, _00136_, _00132_);
  and (_00139_, _00138_, _00131_);
  and (_00141_, _00139_, _00018_);
  and (_00142_, _00141_, _00129_);
  and (_00143_, _00142_, _00128_);
  nor (_00145_, _00143_, _00127_);
  and (_00146_, _00143_, _00127_);
  nor (_00147_, _00146_, _00145_);
  not (_00148_, _00147_);
  nor (_00149_, _00142_, _00128_);
  nor (_00151_, _00149_, _00143_);
  not (_00152_, _00151_);
  nor (_00153_, _00141_, _00129_);
  nor (_00154_, _00153_, _00142_);
  not (_00155_, _00154_);
  and (_00156_, _00138_, _00018_);
  nor (_00158_, _00156_, _00131_);
  nor (_00159_, _00158_, _00141_);
  not (_00160_, _00159_);
  not (_00161_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  not (_00162_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_00163_, _00136_, _00018_);
  and (_00164_, _00163_, _00162_);
  nor (_00166_, _00164_, _00161_);
  or (_00167_, _00166_, _00156_);
  nor (_00169_, _00163_, _00162_);
  nor (_00171_, _00169_, _00164_);
  nor (_00172_, _00053_, _00134_);
  nor (_00173_, _00172_, _00163_);
  not (_00174_, _00173_);
  and (_00175_, _00174_, _00055_);
  not (_00176_, _00175_);
  nor (_00178_, _00176_, _00171_);
  and (_00179_, _00178_, _00167_);
  and (_00180_, _00179_, _00160_);
  and (_00181_, _00180_, _00155_);
  and (_00182_, _00181_, _00152_);
  and (_00183_, _00182_, _00148_);
  nor (_00184_, _00182_, _00148_);
  nor (_00185_, _00184_, _00183_);
  or (_00186_, _00185_, _06911_);
  or (_00187_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_00188_, _00187_, _00059_);
  and (_00189_, _00188_, _00186_);
  or (_00190_, _00189_, _00125_);
  and (_11605_, _00190_, _04856_);
  and (_00191_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_00192_, _00181_, _00152_);
  nor (_00193_, _00192_, _00182_);
  or (_00194_, _00193_, _06911_);
  or (_00195_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_00197_, _00195_, _00059_);
  and (_00198_, _00197_, _00194_);
  or (_00199_, _00198_, _00191_);
  and (_11610_, _00199_, _04856_);
  nor (_00200_, _00180_, _00155_);
  nor (_00201_, _00200_, _00181_);
  or (_00202_, _00201_, _06911_);
  or (_00203_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_00204_, _00203_, _00059_);
  and (_00206_, _00204_, _00202_);
  and (_00207_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00208_, _00207_, _00206_);
  and (_11616_, _00208_, _04856_);
  nor (_00210_, _00179_, _00160_);
  nor (_00211_, _00210_, _00180_);
  or (_00212_, _00211_, _06911_);
  or (_00213_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_00214_, _00213_, _00059_);
  and (_00215_, _00214_, _00212_);
  and (_00216_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_00217_, _00216_, _00215_);
  and (_11618_, _00217_, _04856_);
  or (_00218_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand (_00219_, _08367_, _05808_);
  and (_00220_, _00219_, _04856_);
  and (_11620_, _00220_, _00218_);
  nor (_00221_, _00178_, _00167_);
  nor (_00222_, _00221_, _00179_);
  or (_00223_, _00222_, _06911_);
  or (_00224_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00225_, _00224_, _00059_);
  and (_00226_, _00225_, _00223_);
  and (_00227_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_00228_, _00227_, _00226_);
  and (_11624_, _00228_, _04856_);
  and (_00229_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _08359_);
  and (_00230_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00231_, _00230_, _00229_);
  and (_11630_, _00231_, _04856_);
  nor (_11638_, _12854_, rst);
  and (_00232_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_00233_, _08367_, _05884_);
  or (_00234_, _00233_, _00232_);
  and (_11641_, _00234_, _04856_);
  and (_00235_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_00236_, _00176_, _00171_);
  nor (_00237_, _00236_, _00178_);
  or (_00238_, _00237_, _06911_);
  or (_00239_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_00240_, _00239_, _00059_);
  and (_00241_, _00240_, _00238_);
  or (_00242_, _00241_, _00235_);
  and (_11646_, _00242_, _04856_);
  and (_00243_, \oc8051_top_1.oc8051_memory_interface1.cdata [5], _08359_);
  and (_00244_, \oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00245_, _00244_, _00243_);
  and (_11658_, _00245_, _04856_);
  not (_00246_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_00247_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _00246_);
  or (_00248_, _00247_, _08060_);
  nor (_00249_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  and (_00250_, _00249_, _00248_);
  or (_00251_, _00250_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_00252_, _00251_, _09259_);
  not (_00253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_00254_, _04990_, _00253_);
  nand (_00255_, _00254_, _09259_);
  or (_00256_, _00255_, _07708_);
  and (_00257_, _00256_, _00252_);
  or (_00258_, _00257_, _09263_);
  nand (_00259_, _09263_, _06369_);
  and (_00260_, _00259_, _04856_);
  and (_11698_, _00260_, _00258_);
  and (_00261_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  nor (_00262_, _08367_, _05749_);
  or (_00263_, _00262_, _00261_);
  and (_11704_, _00263_, _04856_);
  and (_00264_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_00265_, _08367_, _05805_);
  or (_00266_, _00265_, _00264_);
  and (_11710_, _00266_, _04856_);
  and (_00267_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  nor (_00268_, _08367_, _05782_);
  or (_00269_, _00268_, _00267_);
  and (_11715_, _00269_, _04856_);
  and (_00270_, _08277_, _07855_);
  nand (_00271_, _00270_, _06088_);
  or (_00272_, _00270_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_00273_, _00272_, _06935_);
  and (_00274_, _00273_, _00271_);
  or (_00275_, _00274_, _06937_);
  and (_11718_, _00275_, _04856_);
  and (_00276_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nor (_00277_, _08367_, _05909_);
  or (_00278_, _00277_, _00276_);
  and (_11720_, _00278_, _04856_);
  and (_00279_, _06163_, _05510_);
  or (_00280_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00281_, _00280_, _04856_);
  nand (_00282_, _00279_, _05287_);
  and (_11723_, _00282_, _00281_);
  and (_00283_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  and (_00284_, _12165_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_00285_, _00284_, _00283_);
  and (_11726_, _00285_, _04856_);
  or (_00286_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00287_, _00286_, _04856_);
  not (_00288_, _00279_);
  or (_00289_, _00288_, _05718_);
  and (_11729_, _00289_, _00287_);
  and (_00290_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_00291_, _08367_, _05778_);
  or (_00292_, _00291_, _00290_);
  and (_11736_, _00292_, _04856_);
  and (_00293_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_00294_, _08367_, _05834_);
  or (_00295_, _00294_, _00293_);
  and (_11751_, _00295_, _04856_);
  nor (_11754_, _07294_, rst);
  nor (_11792_, _12926_, rst);
  nor (_11801_, _12949_, rst);
  and (_00296_, _06721_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_00297_, _06834_, _06733_);
  or (_00298_, _12682_, _12695_);
  or (_00299_, _00298_, _06866_);
  or (_00300_, _00299_, _00297_);
  and (_00301_, _06598_, _05950_);
  or (_00302_, _09088_, _00301_);
  or (_00303_, _00302_, _05988_);
  or (_00304_, _06763_, _06799_);
  or (_00305_, _00304_, _09097_);
  or (_00306_, _00305_, _06756_);
  or (_00308_, _06786_, _06760_);
  or (_00309_, _00308_, _00306_);
  or (_00310_, _00309_, _00303_);
  or (_00311_, _09081_, _06740_);
  or (_00312_, _00311_, _00310_);
  or (_00313_, _00312_, _00300_);
  or (_00314_, _05999_, _05962_);
  nor (_00315_, rst, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_00316_, _00315_, _00314_);
  and (_00317_, _00316_, _00313_);
  or (_11805_, _00317_, _00296_);
  or (_00318_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_00319_, _00318_, _04856_);
  or (_00320_, _00288_, _06410_);
  and (_11825_, _00320_, _00319_);
  or (_00321_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_00322_, _00321_, _04856_);
  nand (_00323_, _00279_, _05669_);
  and (_11830_, _00323_, _00322_);
  and (_00324_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _08359_);
  and (_00325_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00326_, _00325_, _00324_);
  and (_11848_, _00326_, _04856_);
  and (_00327_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _08359_);
  and (_00328_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00329_, _00328_, _00327_);
  and (_11856_, _00329_, _04856_);
  and (_00330_, _12429_, _05517_);
  and (_00331_, _00330_, _05288_);
  and (_00332_, _12718_, _05517_);
  and (_00333_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_00334_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00335_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _00334_);
  and (_00336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00337_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00338_, _00337_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00339_, _00338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00340_, _00339_, _00336_);
  and (_00341_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_00342_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_00343_, _00342_, _00341_);
  and (_00344_, _00343_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  not (_00345_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_00346_, \oc8051_top_1.oc8051_sfr1.pres_ow , _00345_);
  not (_00347_, t0_i);
  and (_00348_, _00347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_00349_, _00348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff );
  or (_00350_, _00349_, _00346_);
  and (_00351_, _00350_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_00352_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00353_, _00352_, _00351_);
  and (_00354_, _00353_, _00344_);
  and (_00355_, _00354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_00356_, _00355_, _00340_);
  nor (_00357_, _00356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00358_, _00356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nor (_00359_, _00358_, _00357_);
  and (_00360_, _00359_, _00335_);
  nor (_00361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00362_, _00343_, _00351_);
  and (_00363_, _00362_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_00364_, _00363_, _00340_);
  nand (_00365_, _00364_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_00366_, _00364_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00367_, _00366_, _00365_);
  and (_00368_, _00367_, _00361_);
  and (_00369_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_00370_, _00369_, _00339_);
  and (_00371_, _00370_, _00336_);
  and (_00372_, _00371_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_00373_, _00372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_00374_, _00372_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00375_, _00374_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00376_, _00375_, _00373_);
  or (_00377_, _00376_, _00368_);
  or (_00378_, _00377_, _00360_);
  nor (_00379_, _00332_, _00330_);
  and (_00380_, _00379_, _00378_);
  or (_00381_, _00380_, _00333_);
  or (_00382_, _00381_, _00331_);
  and (_11877_, _00382_, _04856_);
  and (_00383_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _08359_);
  and (_00384_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00385_, _00384_, _00383_);
  and (_11883_, _00385_, _04856_);
  and (_00386_, _00330_, _06410_);
  and (_00387_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00388_, _00355_, _00339_);
  or (_00389_, _00388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00390_, _00388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_00391_, _00390_);
  and (_00392_, _00391_, _00335_);
  and (_00393_, _00392_, _00389_);
  and (_00394_, _00339_, _00344_);
  and (_00395_, _00394_, _00351_);
  nor (_00396_, _00395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00397_, _00395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_00398_, _00397_, _00396_);
  and (_00399_, _00398_, _00361_);
  not (_00400_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00401_, _00370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nor (_00402_, _00401_, _00400_);
  and (_00403_, _00401_, _00400_);
  or (_00404_, _00403_, _00402_);
  and (_00405_, _00404_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_00406_, _00405_, _00399_);
  or (_00407_, _00406_, _00393_);
  and (_00408_, _00407_, _00379_);
  or (_00409_, _00408_, _00387_);
  or (_00410_, _00409_, _00386_);
  and (_11888_, _00410_, _04856_);
  and (_00411_, _00330_, _05718_);
  and (_00412_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00413_, _07460_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_00414_, _00413_, _00335_);
  and (_00415_, _00390_, _00334_);
  or (_00416_, _00415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_00417_, _00415_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00418_, _00417_, _00416_);
  and (_00419_, _00418_, _00414_);
  and (_00420_, _00370_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_00421_, _00420_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not (_00422_, _00371_);
  and (_00423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00424_, _00423_, _00422_);
  and (_00425_, _00424_, _00421_);
  nand (_00426_, _00397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_00427_, _00397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00428_, _00427_, _00426_);
  and (_00429_, _00428_, _00361_);
  or (_00430_, _00429_, _00425_);
  or (_00431_, _00430_, _00419_);
  and (_00432_, _00431_, _00379_);
  or (_00433_, _00432_, _00412_);
  or (_00434_, _00433_, _00411_);
  and (_11891_, _00434_, _04856_);
  and (_00435_, _00330_, _06705_);
  and (_00436_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00437_, _00355_, _00338_);
  and (_00438_, _00352_, _00344_);
  and (_00439_, _00438_, _00351_);
  and (_00440_, _00439_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_00441_, _00440_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_00442_, _00441_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_00443_, _00442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_00444_, _00443_, _00335_);
  nor (_00445_, _00444_, _00437_);
  and (_00446_, _00363_, _00337_);
  or (_00447_, _00446_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  not (_00448_, _00361_);
  and (_00449_, _00363_, _00338_);
  nor (_00450_, _00449_, _00448_);
  and (_00451_, _00450_, _00447_);
  and (_00452_, _00369_, _00337_);
  and (_00453_, _00452_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_00454_, _00453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_00455_, _00453_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00456_, _00455_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00457_, _00456_, _00454_);
  or (_00458_, _00457_, _00451_);
  or (_00459_, _00458_, _00445_);
  and (_00460_, _00459_, _00379_);
  or (_00461_, _00460_, _00436_);
  or (_00462_, _00461_, _00435_);
  and (_11897_, _00462_, _04856_);
  and (_00463_, _00330_, _05670_);
  and (_00464_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_00465_, _00437_, _00334_);
  or (_00466_, _00465_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_00467_, _00388_);
  or (_00468_, _00467_, _00413_);
  and (_00469_, _00468_, _00414_);
  and (_00470_, _00469_, _00466_);
  and (_00471_, _00369_, _00338_);
  or (_00472_, _00471_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_00473_, _00370_);
  and (_00474_, _00423_, _00473_);
  and (_00475_, _00474_, _00472_);
  not (_00476_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_00477_, _00449_, _00476_);
  and (_00478_, _00449_, _00476_);
  or (_00479_, _00478_, _00477_);
  and (_00480_, _00479_, _00361_);
  or (_00481_, _00480_, _00475_);
  or (_00482_, _00481_, _00470_);
  and (_00483_, _00482_, _00379_);
  or (_00484_, _00483_, _00464_);
  or (_00485_, _00484_, _00463_);
  and (_11900_, _00485_, _04856_);
  not (_00486_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  nor (_00487_, _13234_, _00486_);
  nor (_00488_, _00487_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_00489_, _00487_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_00490_, _00489_, _00488_);
  nor (_11904_, _00490_, rst);
  not (_00491_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_00492_, _00355_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_00493_, _00492_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  nand (_00494_, _00493_, _00491_);
  not (_00495_, _00442_);
  or (_00496_, _00413_, _00495_);
  and (_00497_, _00496_, _00414_);
  and (_00499_, _00497_, _00494_);
  and (_00500_, _00369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_00501_, _00500_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_00502_, _00452_);
  and (_00503_, _00423_, _00502_);
  and (_00504_, _00503_, _00501_);
  and (_00505_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_00506_, _00505_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_00507_, _00446_, _00448_);
  and (_00508_, _00507_, _00506_);
  or (_00509_, _00508_, _00504_);
  or (_00510_, _00509_, _00499_);
  and (_00511_, _00510_, _00379_);
  and (_00512_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00513_, _00330_, _06033_);
  or (_00514_, _00513_, _00512_);
  or (_00515_, _00514_, _00511_);
  and (_11907_, _00515_, _04856_);
  not (_00516_, _00332_);
  or (_00517_, _00516_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_00518_, _00517_, _04856_);
  nand (_00519_, _00330_, _06369_);
  and (_00520_, _00440_, _00334_);
  or (_00521_, _00520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_00522_, _00521_, _00493_);
  and (_00523_, _00522_, _00414_);
  or (_00524_, _00369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_00525_, _00524_, _00423_);
  nor (_00526_, _00525_, _00500_);
  nor (_00527_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_00528_, _00527_, _00505_);
  and (_00529_, _00528_, _00361_);
  or (_00530_, _00529_, _00526_);
  or (_00531_, _00530_, _00523_);
  or (_00532_, _00531_, _00330_);
  and (_00533_, _00532_, _00519_);
  or (_00534_, _00533_, _00332_);
  and (_11910_, _00534_, _00518_);
  and (_00535_, _13234_, _00486_);
  nor (_00536_, _00535_, _00487_);
  and (_11914_, _00536_, _04856_);
  nand (_00537_, _00279_, _06032_);
  or (_00538_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00539_, _00538_, _04856_);
  and (_11924_, _00539_, _00537_);
  or (_00540_, _00288_, _06705_);
  or (_00541_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_00542_, _00541_, _04856_);
  and (_11927_, _00542_, _00540_);
  nor (_00543_, _00279_, _07460_);
  and (_00544_, _00279_, _06997_);
  or (_00545_, _00544_, _00543_);
  and (_11930_, _00545_, _04856_);
  and (_00546_, _06721_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  and (_00547_, _06612_, _05848_);
  or (_00548_, _00547_, _09068_);
  or (_00549_, _00548_, _09067_);
  or (_00550_, _05999_, _05988_);
  or (_00551_, _12689_, _06762_);
  or (_00552_, _00551_, _00550_);
  or (_00553_, _00552_, _06839_);
  or (_00554_, _00553_, _00549_);
  not (_00555_, _07509_);
  or (_00556_, _08051_, _00555_);
  or (_00557_, _12698_, _06760_);
  and (_00558_, _06822_, _06598_);
  and (_00559_, _06638_, _06635_);
  or (_00560_, _00559_, _00558_);
  or (_00561_, _00560_, _00557_);
  or (_00562_, _00561_, _06727_);
  or (_00563_, _00562_, _00556_);
  or (_00564_, _00563_, _00554_);
  and (_00565_, _00564_, _00316_);
  or (_11945_, _00565_, _00546_);
  and (_00566_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  nor (_00567_, _08367_, _05904_);
  or (_00568_, _00567_, _00566_);
  and (_11979_, _00568_, _04856_);
  and (_00569_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  and (_00570_, _12165_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  or (_00571_, _00570_, _00569_);
  and (_11984_, _00571_, _04856_);
  or (_00572_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nand (_00573_, _08367_, _05784_);
  and (_00575_, _00573_, _04856_);
  and (_11993_, _00575_, _00572_);
  or (_00576_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand (_00577_, _08367_, _05829_);
  and (_00578_, _00577_, _04856_);
  and (_11995_, _00578_, _00576_);
  and (_00579_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_00580_, _12165_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  or (_00581_, _00580_, _00579_);
  and (_12001_, _00581_, _04856_);
  or (_00582_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand (_00583_, _08367_, _05875_);
  and (_00584_, _00583_, _04856_);
  and (_12006_, _00584_, _00582_);
  or (_00585_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_00586_, _08367_, _05826_);
  and (_00587_, _00586_, _04856_);
  and (_12011_, _00587_, _00585_);
  not (_00588_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_00589_, t1_i);
  and (_00590_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _00589_);
  nor (_00591_, _00590_, _00588_);
  not (_00592_, _00591_);
  not (_00593_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_00594_, _00593_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_00595_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  not (_00596_, _00595_);
  and (_00597_, _00596_, _00594_);
  and (_00598_, _00597_, _00592_);
  and (_00599_, _00598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_00600_, _00599_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_00601_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_00602_, _00601_, _00598_);
  or (_00603_, _00602_, _00600_);
  and (_00604_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_00605_, _12388_, _05517_);
  nor (_00606_, _00605_, _00604_);
  nand (_00607_, _00606_, _00603_);
  or (_00608_, _00606_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_00609_, _00608_, _00607_);
  and (_00610_, _12713_, _05517_);
  not (_00611_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_00612_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _00611_);
  and (_00613_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_00614_, _00613_, _00601_);
  and (_00615_, _00614_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00616_, _00615_, _00598_);
  and (_00617_, _00616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_00618_, _00617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_00619_, _00618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_00620_, _00619_, _00612_);
  nand (_00621_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_00622_, _00621_, _00605_);
  or (_00623_, _00622_, _00610_);
  or (_00624_, _00623_, _00609_);
  nand (_00625_, _00610_, _06032_);
  and (_00626_, _00625_, _04856_);
  and (_12014_, _00626_, _00624_);
  and (_00627_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00628_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_00629_, _00628_, _00627_);
  and (_00630_, _00629_, _00615_);
  nand (_00631_, _00630_, _00612_);
  or (_00632_, _00631_, _00605_);
  nand (_00633_, _00632_, _00606_);
  and (_00634_, _00633_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_00635_, _00598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_00636_, _00635_, _00599_);
  and (_00637_, _00636_, _00606_);
  or (_00638_, _00637_, _00610_);
  or (_00639_, _00638_, _00634_);
  nand (_00640_, _00610_, _06369_);
  and (_00641_, _00640_, _04856_);
  and (_12017_, _00641_, _00639_);
  not (_00642_, _00606_);
  and (_00643_, _00642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_00644_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_00645_, _00602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_00646_, _00602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_00647_, _00646_, _00645_);
  nor (_00648_, _00647_, _00604_);
  nor (_00649_, _00648_, _00644_);
  nor (_00650_, _00649_, _00605_);
  or (_00651_, _00650_, _00610_);
  or (_00652_, _00651_, _00643_);
  not (_00653_, _00610_);
  or (_00654_, _00653_, _06705_);
  and (_00655_, _00654_, _04856_);
  and (_12032_, _00655_, _00652_);
  or (_00656_, _00653_, _06410_);
  and (_00657_, _00642_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00658_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00659_, _00613_, _00602_);
  or (_00660_, _00659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_00661_, _00616_, _00604_);
  and (_00662_, _00661_, _00660_);
  nor (_00663_, _00662_, _00658_);
  nor (_00664_, _00663_, _00605_);
  or (_00665_, _00664_, _00657_);
  or (_00666_, _00665_, _00610_);
  and (_00667_, _00666_, _04856_);
  and (_12035_, _00667_, _00656_);
  nor (_00668_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_00669_, _00668_, _00659_);
  and (_00671_, _00669_, _00606_);
  nor (_00672_, _00606_, _08808_);
  or (_00673_, _00672_, _00671_);
  nand (_00674_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_00675_, _00674_, _00605_);
  or (_00676_, _00675_, _00610_);
  or (_00677_, _00676_, _00673_);
  nand (_00678_, _00610_, _05669_);
  and (_00679_, _00678_, _04856_);
  and (_12038_, _00679_, _00677_);
  or (_00680_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand (_00681_, _08367_, _05745_);
  and (_00682_, _00681_, _04856_);
  and (_12040_, _00682_, _00680_);
  or (_00683_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_00684_, _08367_, _05879_);
  and (_00685_, _00684_, _04856_);
  and (_12042_, _00685_, _00683_);
  or (_00686_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nand (_00687_, _08367_, _05852_);
  and (_00688_, _00687_, _04856_);
  and (_12049_, _00688_, _00686_);
  nand (_00689_, _00610_, _05287_);
  not (_00690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00691_, _00690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  nor (_00692_, _00691_, _00612_);
  nor (_00693_, _00605_, _00692_);
  not (_00694_, _00693_);
  and (_00695_, _00694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_00696_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00697_, _00696_, _00605_);
  nor (_00698_, _00617_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_00699_, _00698_, _00618_);
  and (_00700_, _00699_, _00693_);
  or (_00701_, _00700_, _00697_);
  or (_00702_, _00701_, _00695_);
  or (_00703_, _00702_, _00610_);
  and (_00704_, _00703_, _04856_);
  and (_12077_, _00704_, _00689_);
  or (_00705_, _00653_, _05718_);
  not (_00706_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_00707_, _00693_, _00706_);
  and (_00708_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not (_00709_, _00692_);
  or (_00710_, _00616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nand (_00711_, _00710_, _00709_);
  nor (_00712_, _00711_, _00617_);
  nor (_00713_, _00712_, _00708_);
  nor (_00714_, _00713_, _00605_);
  or (_00715_, _00714_, _00707_);
  or (_00716_, _00715_, _00610_);
  and (_00717_, _00716_, _04856_);
  and (_12082_, _00717_, _00705_);
  and (_00718_, _12206_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_00719_, _00718_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_12093_, _00719_, _04856_);
  nand (_00720_, _00605_, _05287_);
  and (_00721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00722_, _00721_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_00723_, _00615_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00724_, _00723_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00725_, _00724_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00726_, _00725_, _00598_);
  and (_00727_, _00726_, _00722_);
  or (_00728_, _00727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00729_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  not (_00730_, _00729_);
  and (_00731_, _00727_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00732_, _00731_, _00730_);
  and (_00733_, _00732_, _00728_);
  and (_00734_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_00735_, _00598_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00736_, _00630_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00737_, _00736_, _00735_);
  and (_00738_, _00737_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00739_, _00738_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00740_, _00739_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_00741_, _00740_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_00742_, _00740_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nand (_00743_, _00742_, _00691_);
  nor (_00744_, _00743_, _00741_);
  or (_00745_, _00744_, _00734_);
  or (_00746_, _00745_, _00733_);
  or (_00747_, _00746_, _00605_);
  and (_00748_, _00747_, _00720_);
  or (_00749_, _00748_, _00610_);
  or (_00750_, _00653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_00751_, _00750_, _04856_);
  and (_12119_, _00751_, _00749_);
  nand (_00752_, _00723_, _00598_);
  nor (_00753_, _00752_, _00730_);
  and (_00754_, _00691_, _00598_);
  and (_00755_, _00754_, _00630_);
  or (_00756_, _00755_, _00753_);
  and (_00757_, _00756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_00758_, _00757_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_00759_, _00726_, _00730_);
  or (_00760_, _00759_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_00761_, _00737_, _00611_);
  nand (_00762_, _00761_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_00763_, _00762_, _00760_);
  and (_00764_, _00763_, _00758_);
  or (_00765_, _00764_, _00605_);
  not (_00766_, _00605_);
  or (_00767_, _00766_, _06705_);
  and (_00768_, _00767_, _00765_);
  or (_00769_, _00768_, _00610_);
  or (_00770_, _00653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00771_, _00770_, _04856_);
  and (_12128_, _00771_, _00769_);
  nand (_00772_, _00605_, _05669_);
  or (_00773_, _00737_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  not (_00774_, _00691_);
  nor (_00775_, _00738_, _00774_);
  and (_00776_, _00775_, _00773_);
  and (_00777_, _00726_, _00729_);
  or (_00778_, _00777_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_00779_, _00760_, _08812_);
  and (_00780_, _00779_, _00778_);
  or (_00781_, _00780_, _00776_);
  or (_00782_, _00781_, _00605_);
  and (_00783_, _00782_, _00772_);
  or (_00784_, _00783_, _00610_);
  nand (_00785_, _00610_, _08812_);
  and (_00786_, _00785_, _04856_);
  and (_12130_, _00786_, _00784_);
  or (_00787_, _00766_, _06410_);
  or (_00788_, _00738_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_00789_, _00739_, _00774_);
  and (_00790_, _00789_, _00788_);
  and (_00791_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00792_, _00726_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_00793_, _00792_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00794_, _00792_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nor (_00795_, _00794_, _00730_);
  and (_00796_, _00795_, _00793_);
  or (_00797_, _00796_, _00791_);
  or (_00798_, _00797_, _00790_);
  or (_00799_, _00798_, _00605_);
  and (_00800_, _00799_, _00787_);
  or (_00801_, _00800_, _00610_);
  or (_00802_, _00653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00803_, _00802_, _04856_);
  and (_12135_, _00803_, _00801_);
  or (_00804_, _00766_, _05718_);
  not (_00805_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_00806_, _00739_, _00611_);
  not (_00807_, _00806_);
  nor (_00808_, _00795_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00809_, _00808_, _00807_);
  and (_00810_, _00809_, _00805_);
  nor (_00811_, _00809_, _00805_);
  or (_00812_, _00811_, _00810_);
  or (_00813_, _00812_, _00605_);
  and (_00814_, _00813_, _00804_);
  or (_00815_, _00814_, _00610_);
  nand (_00816_, _00610_, _00805_);
  and (_00817_, _00816_, _04856_);
  and (_12137_, _00817_, _00815_);
  or (_00818_, _12818_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  or (_00819_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _09249_);
  or (_00820_, _00819_, _08087_);
  and (_00821_, _00820_, _04856_);
  and (_12141_, _00821_, _00818_);
  nor (_00822_, _05669_, _06046_);
  and (_00823_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_00824_, _00823_, _05673_);
  or (_00825_, _00824_, _00822_);
  or (_00826_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_00827_, _00826_, _04856_);
  and (_12147_, _00827_, _00825_);
  nor (_00828_, _00756_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_00829_, _00828_, _00757_);
  or (_00830_, _00829_, _00605_);
  nand (_00831_, _00605_, _06032_);
  and (_00832_, _00831_, _00830_);
  or (_00833_, _00832_, _00610_);
  not (_00834_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nand (_00835_, _00610_, _00834_);
  and (_00836_, _00835_, _04856_);
  and (_12151_, _00836_, _00833_);
  or (_00837_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  not (_00838_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nand (_00839_, _06238_, _00838_);
  and (_00840_, _00839_, _04856_);
  and (_12154_, _00840_, _00837_);
  nand (_00841_, _00605_, _06369_);
  nand (_00842_, _00629_, _00616_);
  and (_00843_, _00842_, _00691_);
  or (_00844_, _00619_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00845_, _00844_, _00843_);
  and (_00846_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or (_00847_, _00616_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00848_, _00752_, _00729_);
  and (_00849_, _00848_, _00847_);
  or (_00850_, _00849_, _00846_);
  or (_00851_, _00850_, _00845_);
  or (_00852_, _00851_, _00605_);
  and (_00853_, _00852_, _00841_);
  or (_00854_, _00853_, _00610_);
  or (_00855_, _00653_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00856_, _00855_, _04856_);
  and (_12156_, _00856_, _00854_);
  and (_00857_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_00858_, _00332_, _06997_);
  and (_00859_, _00351_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_00860_, _00351_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_00861_, _00860_, _00859_);
  and (_00862_, _00413_, _00441_);
  or (_00863_, _00862_, _00861_);
  and (_00864_, _00863_, _00379_);
  or (_00866_, _00864_, _00858_);
  or (_00867_, _00866_, _00857_);
  and (_12163_, _00867_, _04856_);
  or (_00868_, _00516_, _06705_);
  and (_00869_, _00868_, _04856_);
  nor (_00870_, _04984_, _04947_);
  and (_00871_, _00870_, _04989_);
  and (_00872_, _00871_, _05517_);
  and (_00873_, _00872_, _05510_);
  and (_00874_, _00341_, _00351_);
  nor (_00875_, _00874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_00876_, _00874_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_00877_, _00876_, _00875_);
  and (_00878_, _00413_, _00440_);
  and (_00879_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_00880_, _00879_, _00877_);
  nor (_00881_, _00880_, _00873_);
  and (_00882_, _00873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_00883_, _00882_, _00881_);
  or (_00884_, _00883_, _00332_);
  and (_12169_, _00884_, _00869_);
  and (_00885_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_00886_, _00876_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_00887_, _00886_, _00362_);
  and (_00888_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_00889_, _00888_, _00887_);
  and (_00890_, _00889_, _00379_);
  or (_00891_, _00890_, _00885_);
  nor (_00892_, _00516_, _05669_);
  or (_00893_, _00892_, _00891_);
  and (_12172_, _00893_, _04856_);
  and (_00894_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_00895_, _00516_, _06032_);
  nor (_00896_, _00859_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_00897_, _00896_, _00874_);
  and (_00898_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_00899_, _00898_, _00897_);
  and (_00900_, _00899_, _00379_);
  or (_00901_, _00900_, _00895_);
  or (_00902_, _00901_, _00894_);
  and (_12173_, _00902_, _04856_);
  and (_00903_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_00904_, _00363_, _00448_);
  and (_00905_, _00904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor (_00906_, _00904_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nor (_00907_, _00906_, _00905_);
  and (_00908_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_00909_, _00908_, _00907_);
  and (_00910_, _00909_, _00379_);
  or (_00911_, _00910_, _00903_);
  and (_00912_, _00332_, _05718_);
  or (_00913_, _00912_, _00911_);
  and (_12178_, _00913_, _04856_);
  and (_00914_, _00330_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00915_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_00916_, _00448_, _00439_);
  or (_00917_, _00905_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00918_, _00917_, _00916_);
  or (_00919_, _00918_, _00915_);
  and (_00920_, _00919_, _00379_);
  or (_00921_, _00920_, _00914_);
  nor (_00922_, _00516_, _05287_);
  or (_00923_, _00922_, _00921_);
  and (_12181_, _00923_, _04856_);
  nor (_00924_, _00362_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_00925_, _00924_, _00363_);
  and (_00926_, _00413_, _00355_);
  and (_00927_, _00926_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_00928_, _00927_, _00925_);
  nor (_00929_, _00928_, _00873_);
  and (_00930_, _00873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_00931_, _00930_, _00929_);
  and (_00932_, _00931_, _00516_);
  and (_00933_, _00332_, _06410_);
  or (_00934_, _00933_, _00932_);
  and (_12184_, _00934_, _04856_);
  and (_12211_, _05963_, _04856_);
  or (_00935_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand (_00936_, _08367_, _05803_);
  and (_00937_, _00936_, _04856_);
  and (_12229_, _00937_, _00935_);
  or (_00938_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  nand (_00939_, _08367_, _05850_);
  and (_00940_, _00939_, _04856_);
  and (_12234_, _00940_, _00938_);
  and (_00941_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_00942_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  or (_00943_, _00942_, _00941_);
  and (_12239_, _00943_, _04856_);
  and (_00944_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_00945_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or (_00946_, _00945_, _00944_);
  and (_12251_, _00946_, _04856_);
  nand (_00947_, _12719_, _06369_);
  or (_00948_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_00949_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_00950_, _00949_, _00948_);
  or (_00951_, _00950_, _12719_);
  and (_00952_, _00951_, _00947_);
  or (_00953_, _00952_, _12714_);
  or (_00954_, _12715_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_00955_, _00954_, _04856_);
  and (_12255_, _00955_, _00953_);
  and (_00956_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_00957_, _06238_);
  and (_00958_, _00957_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  or (_00959_, _00958_, _00956_);
  and (_12267_, _00959_, _04856_);
  or (_00960_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nand (_00961_, _06238_, _05295_);
  and (_00962_, _00961_, _04856_);
  and (_12274_, _00962_, _00960_);
  nand (_00963_, _12171_, _06552_);
  or (_00964_, _12171_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_00965_, _00964_, _04856_);
  and (_12280_, _00965_, _00963_);
  nand (_00966_, _12171_, _07774_);
  or (_00967_, _12171_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_00968_, _00967_, _04856_);
  and (_12300_, _00968_, _00966_);
  and (_12303_, _07212_, _04856_);
  nor (_12317_, _06925_, rst);
  not (_00969_, _07815_);
  and (_00970_, _13037_, _00969_);
  and (_00971_, _12879_, _12829_);
  and (_00972_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_00973_, _12861_, _12534_);
  or (_00974_, _00973_, _00972_);
  or (_00975_, _00974_, _00971_);
  or (_00976_, _00975_, _00970_);
  or (_00977_, _12989_, _12987_);
  and (_00978_, _00977_, _12990_);
  and (_00979_, _00978_, _13070_);
  or (_00980_, _00979_, _00976_);
  and (_00981_, _00980_, _12547_);
  nor (_00982_, _08369_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_00983_, _00982_, _13052_);
  nor (_00984_, _00983_, _12547_);
  or (_00985_, _00984_, _00981_);
  and (_12338_, _00985_, _04856_);
  nand (_00986_, _13108_, _05142_);
  or (_00987_, _00986_, _13091_);
  nand (_00988_, _13111_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_00989_, _00988_, _00987_);
  nand (_00990_, _00989_, _05157_);
  or (_00991_, _00989_, _05157_);
  and (_00992_, _00991_, _13031_);
  and (_00993_, _00992_, _00990_);
  and (_00994_, _13022_, _07598_);
  and (_00995_, _13042_, _05919_);
  not (_00996_, _07089_);
  and (_00997_, _12829_, _00996_);
  or (_00998_, _00997_, _00995_);
  and (_00999_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01000_, _06901_, _06552_);
  or (_01001_, _01000_, _00999_);
  or (_01002_, _01001_, _00998_);
  nor (_01003_, _01002_, _00994_);
  nand (_01004_, _01003_, _12547_);
  or (_01005_, _01004_, _00993_);
  and (_01006_, _13124_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01007_, _13124_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_01008_, _01007_, _01006_);
  or (_01009_, _01008_, _12547_);
  and (_01010_, _01009_, _04856_);
  and (_12343_, _01010_, _01005_);
  or (_01011_, _12688_, _12683_);
  or (_01012_, _05988_, _05949_);
  or (_01013_, _06598_, _05965_);
  and (_01014_, _01013_, _01012_);
  or (_01015_, _01014_, _00548_);
  or (_01016_, _01015_, _01011_);
  and (_01017_, _06635_, _06730_);
  or (_01018_, _08194_, _07508_);
  or (_01019_, _01018_, _01017_);
  or (_01021_, _06747_, _06724_);
  or (_01022_, _01021_, _01019_);
  or (_01024_, _01022_, _01016_);
  and (_01025_, _01024_, _05730_);
  and (_01026_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_01027_, _06002_, _04859_);
  or (_01028_, _01027_, _01026_);
  or (_01029_, _01028_, _01025_);
  and (_12372_, _01029_, _04856_);
  and (_01030_, _05718_, _05675_);
  and (_01032_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_01033_, _01032_, _05673_);
  or (_01034_, _01033_, _01030_);
  or (_01035_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_01036_, _01035_, _04856_);
  and (_12445_, _01036_, _01034_);
  or (_12482_, _07102_, rst);
  and (_12485_, _07310_, _04856_);
  nor (_12489_, _07274_, rst);
  and (_12491_, _07223_, _04856_);
  nor (_12493_, _07154_, rst);
  nand (_12496_, _07067_, _04856_);
  nor (_12621_, _07191_, rst);
  nor (_12646_, _07142_, rst);
  and (_01038_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01039_, _00030_, _00028_);
  and (_01041_, _01039_, _00031_);
  or (_01042_, _01041_, _06911_);
  or (_01043_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01045_, _01043_, _00059_);
  and (_01046_, _01045_, _01042_);
  or (_01047_, _01046_, _01038_);
  and (_12670_, _01047_, _04856_);
  not (_01048_, _10587_);
  or (_01049_, _01048_, _06410_);
  or (_01050_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_01052_, _01050_, _04856_);
  and (_12673_, _01052_, _01049_);
  and (_01053_, _12206_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_01054_, _01053_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_12679_, _01054_, _04856_);
  nor (_01055_, _05287_, _06046_);
  and (_01056_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_01057_, _01056_, _05673_);
  or (_01058_, _01057_, _01055_);
  or (_01059_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_01060_, _01059_, _04856_);
  and (_12690_, _01060_, _01058_);
  and (_01061_, _12206_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_01062_, _01061_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_12694_, _01062_, _04856_);
  or (_01063_, _00027_, _12371_);
  nor (_01064_, _00028_, _06911_);
  and (_01065_, _01064_, _01063_);
  nor (_01067_, _06910_, _05109_);
  or (_01068_, _01067_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_01069_, _01068_, _01065_);
  or (_01070_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _00059_);
  and (_01071_, _01070_, _04856_);
  and (_12702_, _01071_, _01069_);
  and (_01072_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  not (_01073_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_01074_, _00146_, _01073_);
  and (_01075_, _00146_, _01073_);
  or (_01076_, _01075_, _01074_);
  nand (_01077_, _01076_, _00183_);
  or (_01078_, _01076_, _00183_);
  and (_01079_, _01078_, _01077_);
  or (_01080_, _01079_, _06911_);
  or (_01081_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01082_, _01081_, _00059_);
  and (_01083_, _01082_, _01080_);
  or (_01084_, _01083_, _01072_);
  and (_12706_, _01084_, _04856_);
  and (_01085_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7], \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nor (_01086_, _00174_, _00055_);
  nor (_01087_, _01086_, _00175_);
  or (_01088_, _01087_, _06911_);
  or (_01089_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_01090_, _01089_, _00059_);
  and (_01091_, _01090_, _01088_);
  or (_01092_, _01091_, _01085_);
  and (_12712_, _01092_, _04856_);
  nor (_12736_, _07261_, rst);
  and (_01093_, _12206_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_01094_, _01093_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_12750_, _01094_, _04856_);
  and (_12819_, _10047_, _06994_);
  nand (_01095_, _07774_, _06498_);
  not (_01096_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  nand (_01097_, _06497_, _01096_);
  and (_01098_, _01097_, _04856_);
  and (_12951_, _01098_, _01095_);
  nor (_01099_, _12257_, _08816_);
  or (_01100_, _01099_, _07642_);
  and (_01101_, _01100_, _09259_);
  and (_01102_, _09259_, _04984_);
  nor (_01103_, _01102_, _08816_);
  or (_01104_, _01103_, _09263_);
  or (_01105_, _01104_, _01101_);
  nand (_01106_, _09263_, _05669_);
  and (_01107_, _01106_, _04856_);
  and (_13002_, _01107_, _01105_);
  nor (_01108_, _07702_, _06497_);
  and (_01109_, _06497_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  or (_01111_, _01109_, _01108_);
  and (_13064_, _01111_, _04856_);
  not (_01113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_01114_, _08060_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_01116_, _01114_, _01113_);
  nor (_01117_, _01116_, _08922_);
  and (_01118_, _01116_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_01119_, _01118_, _01117_);
  or (_01120_, _01119_, _09259_);
  or (_01121_, _06494_, _08922_);
  nand (_01122_, _01121_, _09259_);
  or (_01123_, _01122_, _07602_);
  and (_01124_, _01123_, _01120_);
  or (_01125_, _01124_, _09263_);
  or (_01126_, _09264_, _06705_);
  and (_01127_, _01126_, _04856_);
  and (_13158_, _01127_, _01125_);
  nor (_01128_, _01006_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  and (_01129_, _01006_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_01130_, _01129_, _01128_);
  or (_01131_, _01130_, _12547_);
  and (_01132_, _01131_, _04856_);
  and (_01133_, _13022_, _07640_);
  and (_01134_, _12829_, _12885_);
  nor (_01135_, _06901_, _06586_);
  or (_01136_, _01135_, _01134_);
  and (_01137_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_01138_, _01137_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01139_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_01140_, _01139_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_01141_, \oc8051_top_1.oc8051_memory_interface1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_01142_, \oc8051_top_1.oc8051_memory_interface1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_01143_, _01142_, _01141_);
  and (_01144_, _01143_, _01140_);
  and (_01145_, _01144_, _01138_);
  and (_01146_, _01145_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_01148_, _01145_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_01149_, _01148_, _01146_);
  and (_01150_, _01149_, _13042_);
  and (_01151_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_01152_, _01151_, _01150_);
  or (_01153_, _01152_, _01136_);
  nor (_01155_, _01153_, _01133_);
  nand (_01156_, _01155_, _12547_);
  not (_01157_, _01138_);
  nor (_01159_, _01157_, _13107_);
  and (_01160_, _01159_, _13091_);
  nor (_01161_, _00986_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01162_, _01161_, _13092_);
  nor (_01163_, _01162_, _01160_);
  nand (_01165_, _01163_, _05089_);
  or (_01166_, _01163_, _05089_);
  and (_01167_, _01166_, _01165_);
  and (_01168_, _01167_, _13070_);
  or (_01169_, _01168_, _01156_);
  and (_13165_, _01169_, _01132_);
  and (_01170_, _09259_, _06091_);
  and (_01171_, _01170_, _06144_);
  nor (_01172_, _01170_, _00246_);
  or (_01173_, _01172_, _09263_);
  or (_01174_, _01173_, _01171_);
  or (_01175_, _09264_, _05718_);
  and (_01176_, _01175_, _04856_);
  and (_13168_, _01176_, _01174_);
  nand (_01177_, _01161_, _05089_);
  or (_01178_, _01177_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_01179_, _01178_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_01180_, _01179_, _13091_);
  and (_01181_, _01159_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01182_, _01181_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_01183_, _01182_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nand (_01184_, _01183_, _13091_);
  and (_01185_, _01184_, _01180_);
  nor (_01186_, _01185_, _05022_);
  and (_01187_, _01185_, _05022_);
  or (_01188_, _01187_, _01186_);
  and (_01189_, _01188_, _13031_);
  and (_01190_, _13022_, _06452_);
  nor (_01191_, _06901_, _06488_);
  and (_01192_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_01193_, _01146_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01194_, _01193_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_01195_, _01194_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01196_, _01194_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_01197_, _01196_, _01195_);
  and (_01198_, _01197_, _13042_);
  and (_01199_, _12829_, _12995_);
  or (_01200_, _01199_, _01198_);
  or (_01201_, _01200_, _01192_);
  or (_01202_, _01201_, _01191_);
  nor (_01203_, _01202_, _01190_);
  nand (_01204_, _01203_, _12547_);
  or (_01205_, _01204_, _01189_);
  and (_01206_, _01129_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_01207_, _01206_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01208_, _01207_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  and (_01209_, _01207_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_01210_, _01209_, _01208_);
  or (_01211_, _01210_, _12547_);
  and (_01212_, _01211_, _04856_);
  and (_13188_, _01212_, _01205_);
  and (_01213_, _01178_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  or (_01214_, _01213_, _01180_);
  or (_01215_, _01182_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01216_, _01215_, _01183_);
  or (_01217_, _01216_, _13092_);
  and (_01218_, _01217_, _13031_);
  and (_01219_, _01218_, _01214_);
  and (_01220_, _13022_, _07924_);
  nor (_01221_, _01193_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  nor (_01222_, _01221_, _01194_);
  and (_01223_, _01222_, _13042_);
  and (_01224_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_01225_, _01224_, _01223_);
  and (_01226_, _12829_, _13063_);
  nor (_01227_, _07897_, _06901_);
  or (_01228_, _01227_, _01226_);
  or (_01229_, _01228_, _01225_);
  nor (_01230_, _01229_, _01220_);
  nand (_01231_, _01230_, _12547_);
  or (_01232_, _01231_, _01219_);
  nor (_01233_, _01206_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_01234_, _01233_, _01207_);
  or (_01235_, _01234_, _12547_);
  and (_01236_, _01235_, _04856_);
  and (_13196_, _01236_, _01232_);
  nand (_01237_, _01177_, _13092_);
  or (_01238_, _01181_, _13092_);
  nand (_01239_, _01238_, _01237_);
  nand (_01240_, _01239_, _05067_);
  or (_01241_, _01239_, _05067_);
  and (_01242_, _01241_, _13031_);
  and (_01243_, _01242_, _01240_);
  and (_01244_, _13022_, _07853_);
  nor (_01245_, _07815_, _06901_);
  and (_01246_, _12829_, _12860_);
  or (_01247_, _01246_, _01245_);
  nor (_01248_, _01146_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_01249_, _01248_, _01193_);
  and (_01250_, _01249_, _13042_);
  and (_01251_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_01252_, _01251_, _01250_);
  or (_01253_, _01252_, _01247_);
  nor (_01254_, _01253_, _01244_);
  nand (_01255_, _01254_, _12547_);
  or (_01256_, _01255_, _01243_);
  nor (_01257_, _01129_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_01258_, _01257_, _01206_);
  or (_01259_, _01258_, _12547_);
  and (_01260_, _01259_, _04856_);
  and (_13203_, _01260_, _01256_);
  and (_01261_, _09259_, _07857_);
  not (_01262_, _09259_);
  or (_01263_, _12246_, _01262_);
  or (_01264_, _01263_, _01102_);
  and (_01265_, _01264_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_01266_, _01265_, _09263_);
  or (_01267_, _01266_, _01261_);
  or (_01268_, _09264_, _06410_);
  and (_01269_, _01268_, _04856_);
  and (_13205_, _01269_, _01267_);
  and (_01270_, _06370_, _05675_);
  nand (_01271_, _05675_, _04861_);
  and (_01272_, _01271_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  or (_01273_, _01272_, _01270_);
  and (_00041_, _01273_, _04856_);
  nand (_01274_, _00332_, _06284_);
  nand (_01275_, _00878_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01276_, _00916_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_01277_, _01276_, _01275_);
  nor (_01278_, _01277_, _00330_);
  or (_01279_, _00916_, _00330_);
  and (_01280_, _01279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_01281_, _01280_, _01278_);
  or (_01282_, _01281_, _00332_);
  and (_01283_, _01282_, _04856_);
  and (_00115_, _01283_, _01274_);
  nand (_01284_, _00330_, _06284_);
  and (_01285_, _00358_, _00334_);
  nand (_01286_, _01285_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01287_, _01285_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_01288_, _01287_, _01286_);
  and (_01289_, _01288_, _00414_);
  and (_01290_, _00369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_01291_, _01290_, _00340_);
  and (_01292_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01293_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_01294_, _01293_, _00423_);
  nor (_01295_, _01294_, _01292_);
  and (_01296_, _00344_, _00351_);
  and (_01297_, _00340_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_01298_, _01297_, _01296_);
  or (_01299_, _01298_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_01300_, _01297_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_01301_, _01300_, _01296_);
  and (_01302_, _01301_, _00361_);
  and (_01303_, _01302_, _01299_);
  or (_01304_, _01303_, _01295_);
  or (_01305_, _01304_, _00330_);
  or (_01306_, _01305_, _01289_);
  and (_01307_, _01306_, _00516_);
  and (_01308_, _01307_, _01284_);
  and (_01309_, _00332_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01310_, _01309_, _01308_);
  and (_00116_, _01310_, _04856_);
  and (_01311_, _00610_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_01312_, _00605_, _06284_);
  or (_01313_, _00741_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_01314_, _01313_, _00691_);
  and (_01315_, _00741_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_01316_, _01315_, _01314_);
  nand (_01318_, _00690_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_01319_, _01318_, _00732_);
  and (_01320_, _00731_, _00729_);
  or (_01321_, _01320_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_01322_, _01321_, _01319_);
  or (_01323_, _01322_, _01316_);
  or (_01324_, _01323_, _00605_);
  and (_01325_, _01324_, _00653_);
  and (_01326_, _01325_, _01312_);
  or (_01327_, _01326_, _01311_);
  and (_00121_, _01327_, _04856_);
  nor (_01328_, _00351_, _06099_);
  or (_01329_, _01300_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_01330_, _00361_, _00440_);
  nand (_01331_, _01330_, _01329_);
  nor (_01332_, _01331_, _01302_);
  or (_01333_, _01332_, _01328_);
  and (_01334_, _01333_, _04856_);
  and (_00124_, _01334_, _00379_);
  not (_01335_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_01336_, _00598_, _01335_);
  or (_01337_, _01336_, _01315_);
  and (_01338_, _01337_, _00691_);
  and (_01339_, _01320_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nand (_01340_, _00598_, _00611_);
  nor (_01341_, _00691_, _01335_);
  and (_01342_, _01341_, _01340_);
  or (_01343_, _01342_, _00620_);
  or (_01344_, _01343_, _01339_);
  or (_01345_, _01344_, _01338_);
  nor (_01346_, _00605_, rst);
  and (_01347_, _01346_, _00653_);
  and (_00126_, _01347_, _01345_);
  or (_01348_, _04989_, _06090_);
  not (_01349_, _01348_);
  or (_01350_, _01349_, _07855_);
  and (_01351_, _06668_, _06930_);
  and (_01352_, _01351_, _06670_);
  nand (_01353_, _01352_, _01350_);
  and (_01354_, _01353_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01355_, _01349_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  or (_01356_, _01355_, _07857_);
  and (_01357_, _01356_, _01352_);
  or (_01358_, _01357_, _01354_);
  and (_01359_, _01358_, _06093_);
  and (_01360_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01361_, _09122_, _06662_);
  nand (_01362_, _01361_, _07815_);
  or (_01363_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01364_, _01363_, _05510_);
  and (_01365_, _01364_, _01362_);
  or (_01366_, _01365_, _01360_);
  or (_01367_, _01366_, _01359_);
  and (_00130_, _01367_, _04856_);
  nand (_01368_, _00610_, _06284_);
  and (_01369_, _00694_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_01370_, _00620_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_01371_, _00618_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_01372_, _01371_, _00619_);
  and (_01373_, _01372_, _00709_);
  nor (_01374_, _01373_, _01370_);
  nor (_01375_, _01374_, _00605_);
  or (_01376_, _01375_, _01369_);
  or (_01377_, _01376_, _00610_);
  and (_01378_, _01377_, _04856_);
  and (_00133_, _01378_, _01368_);
  not (_01379_, _12547_);
  and (_01380_, _13037_, _13153_);
  and (_01381_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_01382_, _12973_, _12829_);
  and (_01383_, _12955_, _12534_);
  or (_01384_, _01383_, _01382_);
  or (_01385_, _01384_, _01381_);
  or (_01386_, _01385_, _01380_);
  nor (_01387_, _12975_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_01388_, _01387_, _12976_);
  and (_01389_, _01388_, _13070_);
  or (_01390_, _01389_, _01386_);
  or (_01391_, _01390_, _01379_);
  or (_01392_, _12547_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_01393_, _01392_, _04856_);
  and (_00137_, _01393_, _01391_);
  and (_00140_, t1_i, _04856_);
  and (_01394_, _01352_, _05520_);
  and (_01395_, _01394_, _06088_);
  nor (_01396_, _01394_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_01398_, _01396_, _06094_);
  nor (_01399_, _01398_, _01395_);
  and (_01400_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  not (_01401_, _01361_);
  and (_01402_, _01401_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nor (_01403_, _01401_, _06586_);
  or (_01404_, _01403_, _01402_);
  and (_01405_, _01404_, _05510_);
  or (_01407_, _01405_, _01400_);
  or (_01408_, _01407_, _01399_);
  and (_00144_, _01408_, _04856_);
  and (_00150_, t0_i, _04856_);
  not (_01409_, _06586_);
  and (_01410_, _13037_, _01409_);
  and (_01411_, _12904_, _12829_);
  and (_01413_, _12886_, _12534_);
  and (_01414_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_01416_, _01414_, _01413_);
  or (_01417_, _01416_, _01411_);
  or (_01418_, _01417_, _01410_);
  or (_01419_, _12907_, _12908_);
  and (_01420_, _01419_, _12985_);
  nor (_01421_, _01419_, _12985_);
  or (_01422_, _01421_, _01420_);
  and (_01423_, _01422_, _13070_);
  or (_01424_, _01423_, _01418_);
  or (_01425_, _01424_, _01379_);
  or (_01426_, _12547_, _08371_);
  and (_01428_, _01426_, _04856_);
  and (_00157_, _01428_, _01425_);
  or (_01429_, _00279_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_01430_, _01429_, _04856_);
  nand (_01431_, _00279_, _06284_);
  and (_00165_, _01431_, _01430_);
  and (_01433_, _01352_, _06146_);
  nand (_01434_, _01433_, _06088_);
  or (_01435_, _01433_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01436_, _01435_, _06093_);
  and (_01438_, _01436_, _01434_);
  and (_01439_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_01440_, _01361_, _06488_);
  or (_01441_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_01442_, _01441_, _05510_);
  and (_01443_, _01442_, _01440_);
  or (_01444_, _01443_, _01439_);
  or (_01445_, _01444_, _01438_);
  and (_00168_, _01445_, _04856_);
  not (_01446_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_01447_, _00369_, _01446_);
  or (_01448_, _01447_, _01292_);
  and (_01449_, _00423_, _04856_);
  and (_01450_, _01449_, _01448_);
  and (_00170_, _01450_, _00379_);
  and (_01451_, _06847_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  not (_01452_, _06552_);
  and (_01453_, _13037_, _01452_);
  nor (_01454_, _12926_, _12830_);
  and (_01455_, _13042_, _00996_);
  or (_01456_, _01455_, _01454_);
  or (_01457_, _01456_, _01453_);
  nor (_01458_, _12983_, _12981_);
  nor (_01459_, _01458_, _12984_);
  and (_01460_, _01459_, _13070_);
  or (_01461_, _01460_, _01457_);
  or (_01462_, _01461_, _01451_);
  and (_01463_, _01462_, _12547_);
  and (_01464_, _01379_, _08387_);
  or (_01465_, _01464_, _01463_);
  and (_00177_, _01465_, _04856_);
  and (_01466_, _12548_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_01467_, _12952_, _12534_);
  not (_01468_, _07774_);
  and (_01469_, _13037_, _01468_);
  or (_01470_, _01469_, _01467_);
  nor (_01471_, _12978_, _12976_);
  nor (_01472_, _01471_, _12979_);
  and (_01473_, _01472_, _13070_);
  or (_01474_, _01473_, _01470_);
  and (_01475_, _01474_, _12547_);
  or (_01476_, _01475_, _01466_);
  and (_00196_, _01476_, _04856_);
  and (_01477_, _01352_, _04986_);
  nand (_01478_, _01477_, _06088_);
  or (_01479_, _01477_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_01480_, _01479_, _06093_);
  and (_01481_, _01480_, _01478_);
  and (_01482_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_01483_, _01401_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nor (_01484_, _01401_, _07774_);
  or (_01485_, _01484_, _01483_);
  and (_01486_, _01485_, _05510_);
  or (_01487_, _01486_, _01482_);
  or (_01488_, _01487_, _01481_);
  and (_00205_, _01488_, _04856_);
  or (_01489_, _01401_, _06144_);
  or (_01490_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_01491_, _01490_, _06093_);
  and (_01492_, _01491_, _01489_);
  and (_01493_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_01495_, _01361_, _07702_);
  and (_01496_, _01495_, _05510_);
  and (_01497_, _01496_, _01490_);
  or (_01498_, _01497_, _01493_);
  or (_01499_, _01498_, _01492_);
  and (_00209_, _01499_, _04856_);
  nor (_01500_, _06346_, rst);
  or (_01501_, _06338_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand (_01502_, _06338_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_01503_, _01502_, _01501_);
  and (_00307_, _01503_, _01500_);
  and (_01504_, _06721_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_01505_, _12825_, _06872_);
  or (_01506_, _12697_, _08209_);
  or (_01507_, _01506_, _01505_);
  or (_01509_, _00298_, _06878_);
  or (_01510_, _01509_, _01507_);
  or (_01511_, _12693_, _08249_);
  or (_01512_, _01511_, _01510_);
  and (_01513_, _01512_, _06770_);
  or (_00498_, _01513_, _01504_);
  and (_01514_, _06410_, _05675_);
  and (_01515_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_01516_, _01515_, _05673_);
  or (_01518_, _01516_, _01514_);
  or (_01519_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_01520_, _01519_, _04856_);
  and (_00574_, _01520_, _01518_);
  and (_01521_, _07176_, _07228_);
  and (_01522_, _01521_, _07499_);
  and (_01523_, _01522_, _06661_);
  nor (_01524_, _01523_, _12477_);
  and (_01525_, _07445_, _06410_);
  and (_01526_, _07074_, _05288_);
  or (_01527_, _01526_, _01525_);
  and (_01528_, _01527_, _07406_);
  and (_01529_, _07406_, _05718_);
  and (_01530_, _07127_, _06033_);
  or (_01531_, _01530_, _01529_);
  and (_01532_, _01531_, _07461_);
  and (_01533_, _07127_, _05670_);
  and (_01534_, _07406_, _09282_);
  or (_01535_, _01534_, _01533_);
  and (_01536_, _01535_, _07452_);
  or (_01537_, _01536_, _01532_);
  and (_01538_, _07445_, _06997_);
  and (_01539_, _07074_, _06705_);
  or (_01540_, _01539_, _01538_);
  and (_01541_, _01540_, _07127_);
  or (_01542_, _01541_, _01537_);
  nor (_01543_, _01542_, _01528_);
  nor (_01544_, _01543_, _01524_);
  or (_01545_, _07394_, _07228_);
  or (_01546_, _01545_, _07402_);
  or (_01548_, _07939_, _07406_);
  or (_01549_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_01550_, _01549_, _07445_);
  and (_01551_, _01550_, _01548_);
  and (_01552_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_01553_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_01554_, _01553_, _01552_);
  and (_01555_, _01554_, _07074_);
  or (_01556_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_01558_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_01560_, _01558_, _07461_);
  and (_01561_, _01560_, _01556_);
  or (_01562_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_01564_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_01565_, _01564_, _07452_);
  and (_01566_, _01565_, _01562_);
  or (_01567_, _01566_, _01561_);
  or (_01568_, _01567_, _01555_);
  nor (_01569_, _01568_, _01551_);
  nor (_01571_, _01569_, _01546_);
  or (_01572_, _07399_, _07398_);
  or (_01573_, _07337_, _07176_);
  or (_01574_, _01573_, _07400_);
  or (_01575_, _01574_, _01572_);
  and (_01576_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_01577_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_01578_, _01577_, _01576_);
  and (_01579_, _01578_, _07452_);
  or (_01581_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_01582_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_01584_, _01582_, _07074_);
  and (_01585_, _01584_, _01581_);
  and (_01587_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_01588_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  or (_01589_, _01588_, _01587_);
  and (_01590_, _01589_, _07445_);
  or (_01591_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_01592_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_01594_, _01592_, _07461_);
  and (_01595_, _01594_, _01591_);
  or (_01596_, _01595_, _01590_);
  or (_01598_, _01596_, _01585_);
  nor (_01600_, _01598_, _01579_);
  nor (_01601_, _01600_, _01575_);
  nand (_01602_, _07482_, _07176_);
  and (_01603_, _08841_, _07127_);
  or (_01604_, _07531_, p1_in[7]);
  or (_01605_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_01606_, _01605_, _01604_);
  and (_01607_, _01606_, _07406_);
  or (_01608_, _01607_, _01603_);
  and (_01609_, _01608_, _07452_);
  or (_01610_, _08940_, _07406_);
  or (_01611_, _07531_, p1_in[6]);
  or (_01612_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_01613_, _01612_, _01611_);
  or (_01614_, _01613_, _07127_);
  and (_01615_, _01614_, _07074_);
  and (_01616_, _01615_, _01610_);
  or (_01617_, _07531_, p1_in[4]);
  or (_01618_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_01619_, _01618_, _01617_);
  and (_01620_, _01619_, _07406_);
  and (_01621_, _07555_, _07127_);
  or (_01622_, _01621_, _01620_);
  and (_01623_, _01622_, _07445_);
  nor (_01624_, _07531_, p1_in[1]);
  not (_01625_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_01626_, _07531_, _01625_);
  nor (_01627_, _01626_, _01624_);
  or (_01628_, _01627_, _07406_);
  nor (_01629_, _07531_, p1_in[5]);
  not (_01630_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_01631_, _07531_, _01630_);
  nor (_01632_, _01631_, _01629_);
  or (_01633_, _01632_, _07127_);
  and (_01634_, _01633_, _07461_);
  and (_01635_, _01634_, _01628_);
  or (_01636_, _01635_, _01623_);
  or (_01637_, _01636_, _01616_);
  nor (_01638_, _01637_, _01609_);
  nor (_01639_, _01638_, _01602_);
  and (_01640_, _07394_, _07398_);
  and (_01641_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_01642_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_01643_, _01642_, _01641_);
  and (_01645_, _01643_, _07461_);
  and (_01646_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_01647_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_01648_, _01647_, _01646_);
  and (_01649_, _01648_, _07452_);
  or (_01650_, _01649_, _01645_);
  and (_01651_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_01652_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_01653_, _01652_, _01651_);
  and (_01654_, _01653_, _07445_);
  and (_01655_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_01656_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_01657_, _01656_, _01655_);
  and (_01658_, _01657_, _07074_);
  or (_01659_, _01658_, _01654_);
  or (_01660_, _01659_, _01650_);
  and (_01661_, _01660_, _07447_);
  and (_01662_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and (_01663_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_01664_, _01663_, _01662_);
  and (_01665_, _01664_, _07461_);
  and (_01666_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_01667_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  or (_01668_, _01667_, _01666_);
  and (_01670_, _01668_, _07452_);
  or (_01671_, _01670_, _01665_);
  and (_01672_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_01673_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_01674_, _01673_, _01672_);
  and (_01675_, _01674_, _07445_);
  and (_01676_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_01677_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_01678_, _01677_, _01676_);
  and (_01679_, _01678_, _07074_);
  or (_01680_, _01679_, _01675_);
  or (_01681_, _01680_, _01671_);
  and (_01682_, _01681_, _07386_);
  or (_01683_, _01682_, _01661_);
  and (_01684_, _01683_, _01640_);
  or (_01685_, _01684_, _01639_);
  or (_01686_, _01685_, _01601_);
  or (_01687_, _07401_, _07279_);
  or (_01688_, _01545_, _01687_);
  and (_01689_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_01690_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_01691_, _01690_, _01689_);
  and (_01692_, _01691_, _07452_);
  or (_01693_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_01694_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_01695_, _01694_, _07074_);
  and (_01696_, _01695_, _01693_);
  and (_01697_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01698_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_01699_, _01698_, _01697_);
  and (_01700_, _01699_, _07445_);
  or (_01701_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_01702_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_01703_, _01702_, _07461_);
  and (_01704_, _01703_, _01701_);
  or (_01705_, _01704_, _01700_);
  or (_01706_, _01705_, _01696_);
  nor (_01707_, _01706_, _01692_);
  nor (_01708_, _01707_, _01688_);
  or (_01709_, _07991_, _04858_);
  and (_01711_, _01688_, _01602_);
  nand (_01712_, _07447_, _07176_);
  and (_01713_, _01712_, _01575_);
  and (_01714_, _01713_, _01711_);
  not (_01715_, _01546_);
  nor (_01716_, _01715_, _01522_);
  and (_01717_, _01521_, _07386_);
  nand (_01718_, _07385_, _07394_);
  nand (_01719_, _01718_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_01720_, _01719_, _01717_);
  and (_01721_, _01720_, _01716_);
  nand (_01722_, _01721_, _01714_);
  nand (_01723_, _01722_, _01709_);
  or (_01724_, _01723_, _01708_);
  and (_01725_, _08836_, _07452_);
  nor (_01726_, _07531_, p0_in[1]);
  not (_01727_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_01728_, _07531_, _01727_);
  nor (_01729_, _01728_, _01726_);
  and (_01730_, _01729_, _07461_);
  or (_01731_, _01730_, _07406_);
  or (_01732_, _01731_, _01725_);
  or (_01733_, _07531_, p0_in[7]);
  or (_01734_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_01735_, _01734_, _01733_);
  and (_01736_, _01735_, _07452_);
  nor (_01737_, _07531_, p0_in[5]);
  not (_01738_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01739_, _07531_, _01738_);
  nor (_01740_, _01739_, _01737_);
  and (_01741_, _01740_, _07461_);
  or (_01742_, _01741_, _07127_);
  or (_01743_, _01742_, _01736_);
  and (_01744_, _01743_, _01732_);
  or (_01745_, _07531_, p0_in[6]);
  or (_01746_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_01747_, _01746_, _01745_);
  and (_01748_, _01747_, _07406_);
  and (_01749_, _08944_, _07127_);
  or (_01750_, _01749_, _01748_);
  and (_01751_, _01750_, _07074_);
  or (_01752_, _07531_, p0_in[4]);
  or (_01753_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_01754_, _01753_, _01752_);
  and (_01755_, _01754_, _07406_);
  and (_01756_, _07550_, _07127_);
  or (_01757_, _01756_, _01755_);
  and (_01758_, _01757_, _07445_);
  or (_01759_, _01758_, _01751_);
  or (_01760_, _01759_, _01744_);
  and (_01761_, _01760_, _01717_);
  and (_01762_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_01763_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_01764_, _01763_, _01762_);
  and (_01765_, _01764_, _07452_);
  or (_01766_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_01767_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_01768_, _01767_, _07074_);
  and (_01769_, _01768_, _01766_);
  and (_01770_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_01771_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_01772_, _01771_, _01770_);
  and (_01773_, _01772_, _07445_);
  or (_01774_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_01775_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01777_, _01775_, _07461_);
  and (_01778_, _01777_, _01774_);
  or (_01779_, _01778_, _01773_);
  or (_01780_, _01779_, _01769_);
  or (_01781_, _01780_, _01765_);
  and (_01782_, _01781_, _01522_);
  or (_01783_, _01782_, _01761_);
  or (_01784_, _01783_, _01724_);
  or (_01786_, _01784_, _01686_);
  and (_01787_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_01788_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_01789_, _01788_, _01787_);
  and (_01790_, _01789_, _07445_);
  or (_01792_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_01793_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_01795_, _01793_, _07461_);
  and (_01797_, _01795_, _01792_);
  or (_01798_, _01797_, _01790_);
  and (_01800_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_01802_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_01804_, _01802_, _01800_);
  and (_01806_, _01804_, _07074_);
  or (_01807_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_01809_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_01810_, _01809_, _07452_);
  and (_01811_, _01810_, _01807_);
  or (_01813_, _01811_, _01806_);
  or (_01814_, _01813_, _01798_);
  and (_01815_, _01814_, _07387_);
  and (_01816_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_01818_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_01819_, _01818_, _01816_);
  and (_01820_, _01819_, _07445_);
  or (_01821_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_01822_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_01823_, _01822_, _07461_);
  and (_01825_, _01823_, _01821_);
  or (_01826_, _01825_, _01820_);
  and (_01827_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_01828_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  or (_01830_, _01828_, _01827_);
  and (_01831_, _01830_, _07074_);
  or (_01832_, _07127_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_01833_, _07406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_01834_, _01833_, _07452_);
  and (_01835_, _01834_, _01832_);
  or (_01836_, _01835_, _01831_);
  or (_01837_, _01836_, _01826_);
  and (_01838_, _01837_, _07448_);
  or (_01839_, _01838_, _01815_);
  and (_01840_, _01839_, _07394_);
  and (_01841_, _08953_, _07127_);
  or (_01842_, _07531_, p2_in[6]);
  or (_01843_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_01844_, _01843_, _01842_);
  and (_01845_, _01844_, _07406_);
  or (_01847_, _01845_, _01841_);
  and (_01848_, _01847_, _07074_);
  nor (_01850_, _07531_, p2_in[5]);
  not (_01852_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_01854_, _07531_, _01852_);
  nor (_01855_, _01854_, _01850_);
  or (_01857_, _01855_, _07127_);
  nor (_01858_, _07531_, p2_in[1]);
  not (_01860_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_01861_, _07531_, _01860_);
  nor (_01862_, _01861_, _01858_);
  or (_01863_, _01862_, _07406_);
  and (_01864_, _01863_, _07461_);
  and (_01865_, _01864_, _01857_);
  or (_01866_, _01865_, _01848_);
  or (_01867_, _07531_, p2_in[4]);
  or (_01868_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_01869_, _01868_, _01867_);
  and (_01870_, _01869_, _07406_);
  and (_01871_, _07536_, _07127_);
  or (_01872_, _01871_, _01870_);
  and (_01873_, _01872_, _07445_);
  or (_01874_, _08847_, _07406_);
  or (_01875_, _07531_, p2_in[7]);
  or (_01876_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_01877_, _01876_, _01875_);
  or (_01878_, _01877_, _07127_);
  and (_01879_, _01878_, _07452_);
  and (_01880_, _01879_, _01874_);
  or (_01881_, _01880_, _01873_);
  or (_01882_, _01881_, _01866_);
  and (_01883_, _01882_, _07228_);
  nor (_01885_, _07531_, p3_in[1]);
  not (_01886_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_01887_, _07531_, _01886_);
  nor (_01888_, _01887_, _01885_);
  and (_01889_, _01888_, _07127_);
  nor (_01890_, _07531_, p3_in[5]);
  not (_01891_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_01892_, _07531_, _01891_);
  nor (_01893_, _01892_, _01890_);
  and (_01894_, _01893_, _07406_);
  or (_01895_, _01894_, _01889_);
  and (_01896_, _01895_, _07461_);
  or (_01897_, _07531_, p3_in[4]);
  or (_01898_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_01899_, _01898_, _01897_);
  or (_01900_, _01899_, _07127_);
  or (_01901_, _07544_, _07406_);
  and (_01902_, _01901_, _07445_);
  and (_01904_, _01902_, _01900_);
  or (_01905_, _01904_, _01896_);
  or (_01906_, _07531_, p3_in[6]);
  or (_01907_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_01908_, _01907_, _01906_);
  and (_01909_, _01908_, _07406_);
  and (_01910_, _08949_, _07127_);
  or (_01911_, _01910_, _01909_);
  and (_01912_, _01911_, _07074_);
  or (_01913_, _08852_, _07406_);
  or (_01914_, _07531_, p3_in[7]);
  or (_01915_, _07533_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_01916_, _01915_, _01914_);
  or (_01917_, _01916_, _07127_);
  and (_01918_, _01917_, _07452_);
  and (_01919_, _01918_, _01913_);
  or (_01921_, _01919_, _01912_);
  or (_01922_, _01921_, _01905_);
  and (_01923_, _01922_, _07398_);
  nor (_01925_, _01923_, _01883_);
  nor (_01926_, _01925_, _01712_);
  or (_01927_, _01926_, _01840_);
  or (_01928_, _01927_, _01786_);
  or (_01929_, _01928_, _01571_);
  or (_01930_, _01709_, _06144_);
  and (_01932_, _01930_, _01524_);
  and (_01933_, _01932_, _01929_);
  or (_01934_, _01933_, _01544_);
  and (_00670_, _01934_, _04856_);
  and (_01935_, _09254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_01936_, _01935_, _08063_);
  and (_01937_, _09253_, _01936_);
  or (_01938_, _01937_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  not (_01939_, rxd_i);
  nand (_01940_, _01937_, _01939_);
  and (_01941_, _01940_, _04856_);
  and (_00865_, _01941_, _01938_);
  or (_01942_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  or (_01944_, _01942_, _12219_);
  not (_01945_, _06268_);
  nand (_01946_, _01945_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_01947_, _01946_, _12177_);
  or (_01948_, _01947_, _06657_);
  and (_01949_, _01948_, _01944_);
  or (_01950_, _01949_, _12183_);
  nand (_01951_, _12183_, _06284_);
  and (_01952_, _01951_, _04856_);
  and (_01020_, _01952_, _01950_);
  nor (_01954_, _12453_, _12220_);
  not (_01956_, _12391_);
  nor (_01957_, _12393_, _01956_);
  and (_01958_, _01957_, _12401_);
  and (_01959_, _01958_, _12420_);
  and (_01961_, _01959_, _12453_);
  or (_01963_, _01961_, _01954_);
  and (_01023_, _01963_, _04856_);
  and (_01965_, _12401_, _01956_);
  and (_01966_, _01965_, _12453_);
  not (_01967_, _01966_);
  or (_01968_, _01967_, _12420_);
  or (_01969_, _01966_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_01970_, _01969_, _04856_);
  and (_01031_, _01970_, _01968_);
  and (_01971_, _05674_, _04861_);
  and (_01972_, _01971_, _05718_);
  not (_01973_, _01971_);
  and (_01974_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_01975_, _01974_, _01972_);
  and (_01037_, _01975_, _04856_);
  nand (_01976_, _12389_, _06284_);
  and (_01977_, _12393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  not (_01978_, _01977_);
  and (_01979_, _01978_, _12416_);
  nor (_01980_, _01979_, _12430_);
  or (_01981_, _01980_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  nand (_01982_, _12422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_01983_, _01982_, _12401_);
  nand (_01984_, _01983_, _12420_);
  and (_01985_, _01984_, _12395_);
  or (_01986_, _01985_, _01977_);
  or (_01987_, _01986_, _12430_);
  and (_01988_, _01987_, _01981_);
  or (_01989_, _01988_, _12389_);
  and (_01990_, _01989_, _04856_);
  and (_01040_, _01990_, _01976_);
  nand (_01991_, _12430_, _06284_);
  and (_01992_, _12393_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  nor (_01993_, _12602_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nor (_01994_, _01993_, _12553_);
  and (_01995_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_01996_, _01995_, _12420_);
  or (_01997_, _01996_, _01994_);
  and (_01998_, _01997_, _12395_);
  nor (_01999_, _01998_, _01992_);
  nand (_02000_, _01999_, _12431_);
  and (_02001_, _02000_, _12390_);
  and (_02002_, _02001_, _01991_);
  and (_02003_, _12389_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_02004_, _02003_, _02002_);
  and (_01044_, _02004_, _04856_);
  or (_02005_, _09251_, _08065_);
  or (_02006_, _09253_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_02007_, _02006_, _04856_);
  and (_01051_, _02007_, _02005_);
  nand (_02008_, _12714_, _06284_);
  and (_02009_, _12735_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_02010_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_02011_, _02010_, _02009_);
  or (_02012_, _02011_, _12714_);
  and (_02013_, _02012_, _04856_);
  and (_01066_, _02013_, _02008_);
  nor (_01110_, _07927_, rst);
  and (_01112_, _07573_, _04856_);
  and (_01115_, _07862_, _04856_);
  nor (_01147_, _07712_, rst);
  and (_02014_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_02015_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_02017_, _06238_, _02015_);
  or (_02018_, _02017_, _02014_);
  and (_01154_, _02018_, _04856_);
  and (_02019_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  not (_02020_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_02021_, _06238_, _02020_);
  or (_02023_, _02021_, _02019_);
  and (_01158_, _02023_, _04856_);
  and (_01317_, _07780_, _04856_);
  nand (_02024_, _12719_, _06284_);
  and (_02025_, _12717_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_02026_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_02027_, _02026_, _02025_);
  or (_02028_, _02027_, _12719_);
  and (_02029_, _02028_, _12715_);
  and (_02030_, _02029_, _02024_);
  and (_02031_, _12714_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_02032_, _02031_, _02030_);
  and (_01397_, _02032_, _04856_);
  and (_01406_, t2ex_i, _04856_);
  nor (_02033_, t2ex_i, rst);
  and (_01412_, _02033_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r );
  nor (_02034_, t2_i, rst);
  and (_01415_, _02034_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  or (_02035_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_02037_, _06238_, _05089_);
  and (_02038_, _02037_, _04856_);
  and (_01427_, _02038_, _02035_);
  and (_02039_, _09282_, _05671_);
  and (_02040_, _06696_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  or (_02041_, _02040_, _02039_);
  and (_01437_, _02041_, _04856_);
  and (_01494_, t2_i, _04856_);
  and (_02043_, _09251_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not (_02044_, _08062_);
  nor (_02045_, _01935_, _02044_);
  or (_02046_, _02045_, _02043_);
  and (_02047_, _09254_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02048_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02050_, _02048_, _04856_);
  and (_01508_, _02050_, _02046_);
  and (_02051_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_02052_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_01557_, _02052_, _02051_);
  and (_02053_, _06297_, _07855_);
  nand (_02055_, _02053_, _06088_);
  or (_02056_, _02053_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_02057_, _02056_, _06305_);
  and (_02058_, _02057_, _02055_);
  and (_02059_, _06410_, _06304_);
  or (_02060_, _02059_, _02058_);
  and (_01559_, _02060_, _04856_);
  and (_02061_, _06297_, _04986_);
  nand (_02063_, _02061_, _06088_);
  or (_02064_, _02061_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_02065_, _02064_, _06305_);
  and (_02066_, _02065_, _02063_);
  nor (_02067_, _06305_, _06032_);
  or (_02068_, _02067_, _02066_);
  and (_01563_, _02068_, _04856_);
  and (_02069_, _06270_, _07855_);
  or (_02070_, _02069_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_02071_, _02070_, _06276_);
  nand (_02073_, _02069_, _06088_);
  and (_02074_, _02073_, _02071_);
  and (_02075_, _06410_, _06275_);
  or (_02076_, _02075_, _02074_);
  and (_01570_, _02076_, _04856_);
  and (_02077_, _06270_, _04986_);
  or (_02078_, _02077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_02079_, _02078_, _06276_);
  nand (_02080_, _02077_, _06088_);
  and (_02081_, _02080_, _02079_);
  nor (_02083_, _06276_, _06032_);
  or (_02084_, _02083_, _02081_);
  and (_01580_, _02084_, _04856_);
  and (_02085_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_01583_, _02085_, _08058_);
  or (_02086_, _12716_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  not (_02087_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nand (_02088_, _12716_, _02087_);
  and (_02089_, _02088_, _02086_);
  or (_02090_, _02089_, _12719_);
  nand (_02092_, _12719_, _06032_);
  and (_02093_, _02092_, _02090_);
  or (_02094_, _02093_, _12714_);
  not (_02095_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  nand (_02096_, _12714_, _02095_);
  and (_02097_, _02096_, _04856_);
  and (_01586_, _02097_, _02094_);
  not (_02098_, _06225_);
  nor (_02099_, _02098_, _06202_);
  nand (_02100_, _06249_, _02099_);
  and (_02101_, _06249_, _06202_);
  or (_02102_, _02101_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and (_02103_, _02102_, _04856_);
  and (_01593_, _02103_, _02100_);
  nand (_02104_, _06288_, _02099_);
  and (_02105_, _06288_, _06202_);
  or (_02106_, _02105_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and (_02107_, _02106_, _04856_);
  and (_01597_, _02107_, _02104_);
  or (_02108_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_02109_, _02108_, _06206_);
  not (_02110_, _06208_);
  or (_02111_, _02110_, _06105_);
  not (_02112_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_02113_, _06218_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_02114_, _02113_, _02112_);
  and (_02115_, _06216_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_02116_, _02115_, _06221_);
  nand (_02117_, _02116_, _02114_);
  not (_02118_, _06210_);
  or (_02119_, _06222_, _06105_);
  and (_02120_, _02119_, _02118_);
  and (_02121_, _02120_, _02117_);
  and (_02122_, _02108_, _06210_);
  or (_02123_, _02122_, _06208_);
  or (_02124_, _02123_, _02121_);
  and (_02125_, _02124_, _02111_);
  or (_02126_, _02125_, _06205_);
  nand (_02127_, _02126_, _02109_);
  nand (_02128_, _02127_, _02099_);
  and (_02129_, _06194_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_02130_, _02129_, _02112_);
  nor (_02131_, _06190_, _06104_);
  nor (_02132_, _02131_, _06198_);
  nand (_02133_, _02132_, _02130_);
  or (_02134_, _06199_, _06105_);
  and (_02135_, _02134_, _02133_);
  or (_02136_, _02135_, _06184_);
  not (_02138_, _06182_);
  not (_02139_, _06184_);
  or (_02140_, _02108_, _02139_);
  and (_02141_, _02140_, _02138_);
  and (_02142_, _02141_, _02136_);
  and (_02143_, _06182_, _06105_);
  or (_02144_, _02143_, _06179_);
  or (_02145_, _02144_, _02142_);
  or (_02146_, _02108_, _06180_);
  and (_02147_, _02146_, _02145_);
  or (_02148_, _02147_, _06228_);
  and (_02149_, _02148_, _02128_);
  or (_02150_, _02149_, _06172_);
  nor (_02151_, _06172_, _06226_);
  or (_02152_, _02151_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_02153_, _02152_, _04856_);
  and (_01599_, _02153_, _02150_);
  not (_02154_, _05994_);
  and (_02155_, _06859_, _02154_);
  or (_02156_, _06872_, _06856_);
  or (_02157_, _02156_, _06616_);
  or (_02158_, _12685_, _06878_);
  or (_02160_, _02158_, _12688_);
  or (_02161_, _02160_, _02157_);
  and (_02162_, _02161_, _05962_);
  or (_02163_, _02162_, _02155_);
  and (_01644_, _02163_, _04856_);
  and (_02164_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_02165_, _01971_, _06033_);
  or (_02166_, _02165_, _02164_);
  and (_01776_, _02166_, _04856_);
  and (_02167_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_02168_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_01785_, _02168_, _02167_);
  and (_02169_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_02170_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_01791_, _02170_, _02169_);
  and (_02171_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_02172_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  or (_01794_, _02172_, _02171_);
  nor (_02173_, _06218_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_02174_, _02173_, _06216_);
  or (_02175_, _02174_, _06221_);
  and (_02176_, _02175_, _02118_);
  or (_02177_, _02176_, _06208_);
  and (_02178_, _02099_, _06206_);
  and (_02179_, _02178_, _02177_);
  or (_02180_, _06194_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_02181_, _02180_, _06190_);
  or (_02182_, _02181_, _06198_);
  and (_02183_, _02182_, _02139_);
  or (_02184_, _02183_, _06182_);
  and (_02185_, _06202_, _06180_);
  and (_02186_, _02185_, _02184_);
  or (_02187_, _02186_, _06172_);
  or (_02188_, _02187_, _02179_);
  nand (_02189_, _06172_, _12199_);
  and (_02190_, _02189_, _04856_);
  and (_01796_, _02190_, _02188_);
  and (_02191_, _06297_, _06091_);
  and (_02192_, _02191_, _06088_);
  nor (_02193_, _02191_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_02194_, _02193_, _02192_);
  nand (_02195_, _02194_, _06305_);
  or (_02196_, _06305_, _05718_);
  and (_02197_, _02196_, _04856_);
  and (_01799_, _02197_, _02195_);
  and (_02199_, _06270_, _06091_);
  or (_02200_, _02199_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_02201_, _02200_, _06276_);
  nand (_02202_, _02199_, _06088_);
  and (_02203_, _02202_, _02201_);
  and (_02204_, _06275_, _05718_);
  or (_02205_, _02204_, _02203_);
  and (_01801_, _02205_, _04856_);
  and (_02206_, _06136_, _04990_);
  or (_02207_, _02206_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_02209_, _02207_, _06129_);
  nand (_02210_, _02206_, _06088_);
  and (_02211_, _02210_, _02209_);
  and (_02212_, _06997_, _06127_);
  or (_02213_, _02212_, _02211_);
  and (_01803_, _02213_, _04856_);
  nand (_02214_, _10587_, _05287_);
  or (_02215_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_02216_, _02215_, _04856_);
  and (_01805_, _02216_, _02214_);
  or (_02217_, _06235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_02218_, _02217_, _04856_);
  or (_02219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_02220_, _02219_, _06180_);
  or (_02221_, _02220_, _06186_);
  and (_02222_, _06198_, _06110_);
  or (_02223_, _02129_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nand (_02225_, _02223_, _02132_);
  nand (_02226_, _02225_, _06185_);
  or (_02227_, _02226_, _02222_);
  and (_02228_, _02227_, _02221_);
  and (_02229_, _06179_, _06110_);
  or (_02230_, _02229_, _02228_);
  and (_02231_, _02230_, _06202_);
  and (_02232_, _02098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_02233_, _06205_, _06110_);
  and (_02234_, _02219_, _06206_);
  or (_02236_, _02234_, _06212_);
  or (_02237_, _02113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_02238_, _02237_, _02116_);
  nand (_02240_, _06221_, _06110_);
  nand (_02241_, _02240_, _06211_);
  or (_02242_, _02241_, _02238_);
  and (_02243_, _02242_, _02236_);
  or (_02244_, _02243_, _02233_);
  and (_02245_, _02244_, _06225_);
  or (_02246_, _02245_, _02232_);
  and (_02247_, _02246_, _06228_);
  or (_02248_, _02247_, _02231_);
  or (_02249_, _02248_, _06172_);
  and (_01808_, _02249_, _02218_);
  and (_02250_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  not (_02251_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_02252_, _06238_, _02251_);
  or (_02253_, _02252_, _02250_);
  and (_01812_, _02253_, _04856_);
  or (_02254_, _06221_, _06210_);
  and (_02255_, _06219_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_02256_, _02255_, _02254_);
  and (_02257_, _02256_, _02110_);
  and (_02258_, _02257_, _02178_);
  or (_02259_, _06198_, _06184_);
  and (_02260_, _06196_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_02261_, _02260_, _02259_);
  and (_02262_, _02261_, _02138_);
  and (_02263_, _02262_, _02185_);
  or (_02264_, _02263_, _06172_);
  or (_02265_, _02264_, _02258_);
  or (_02266_, _06235_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_02267_, _02266_, _04856_);
  and (_01817_, _02267_, _02265_);
  and (_02268_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_02269_, _06370_, _05674_);
  or (_02270_, _02269_, _02268_);
  and (_01824_, _02270_, _04856_);
  and (_02271_, _08057_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_02272_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_01829_, _02272_, _02271_);
  and (_02273_, _06172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_02274_, _02273_, _02151_);
  and (_01846_, _02274_, _04856_);
  and (_01849_, _13181_, _06172_);
  and (_02275_, _06172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_02276_, _02275_, _02151_);
  and (_01851_, _02276_, _04856_);
  and (_01853_, _13207_, _06172_);
  and (_02277_, _06222_, _06212_);
  nand (_02278_, _02277_, _06203_);
  or (_02279_, _02278_, _06219_);
  nor (_02280_, _02279_, _06202_);
  and (_02281_, _06172_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  or (_02282_, _06172_, _06198_);
  nor (_02283_, _02282_, _06177_);
  not (_02284_, _06186_);
  nor (_02285_, _06196_, _02284_);
  and (_02286_, _02285_, _02283_);
  or (_02287_, _02286_, _02281_);
  or (_02288_, _02287_, _02280_);
  and (_01856_, _02288_, _04856_);
  nand (_02289_, _06288_, _06226_);
  nor (_02290_, _06172_, _06202_);
  or (_02291_, _02290_, _06104_);
  and (_02292_, _02291_, _04856_);
  and (_01859_, _02292_, _02289_);
  or (_02293_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_02294_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  and (_02295_, _02294_, _12420_);
  nand (_02296_, _12412_, _12401_);
  and (_02297_, _02296_, _08794_);
  nor (_02298_, _02297_, _12440_);
  or (_02299_, _02298_, _12393_);
  or (_02300_, _02299_, _02295_);
  nand (_02301_, _02300_, _02293_);
  nor (_02302_, _02301_, _12430_);
  and (_02303_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  or (_02304_, _02303_, _12389_);
  or (_02305_, _02304_, _02302_);
  nand (_02306_, _12389_, _05669_);
  and (_02307_, _02306_, _04856_);
  and (_01884_, _02307_, _02305_);
  and (_02308_, _09259_, _06268_);
  nand (_02309_, _02308_, _06088_);
  or (_02310_, _02308_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_02311_, _02310_, _09264_);
  and (_02312_, _02311_, _02309_);
  nor (_02313_, _09264_, _06284_);
  or (_02314_, _02313_, _02312_);
  and (_01903_, _02314_, _04856_);
  or (_02315_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_02316_, _02315_, _04856_);
  nand (_02317_, _09200_, _06284_);
  and (_01920_, _02317_, _02316_);
  and (_02318_, _04856_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_02319_, _02318_, _09206_);
  and (_02320_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  nor (_02321_, _09206_, rst);
  and (_02322_, _02321_, _02320_);
  or (_01924_, _02322_, _02319_);
  not (_02323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_02324_, _02323_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_02325_, _02324_, _06179_);
  nor (_02326_, _02325_, _06186_);
  nand (_02327_, _06198_, _06109_);
  nor (_02328_, _06190_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_02329_, _02328_, _06198_);
  nand (_02330_, _06194_, _06104_);
  and (_02331_, _02330_, _02323_);
  or (_02332_, _02331_, _02329_);
  and (_02333_, _02332_, _06185_);
  and (_02334_, _02333_, _02327_);
  or (_02335_, _02334_, _02326_);
  nand (_02336_, _06179_, _06109_);
  and (_02337_, _02336_, _02335_);
  nand (_02338_, _02337_, _06202_);
  nor (_02339_, _02324_, _06205_);
  or (_02341_, _02339_, _06212_);
  and (_02342_, _06218_, _06104_);
  or (_02343_, _02342_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_02344_, _06216_, _06104_);
  nor (_02345_, _02344_, _06221_);
  and (_02346_, _02345_, _02343_);
  nand (_02347_, _06221_, _06109_);
  nand (_02348_, _02347_, _06211_);
  or (_02349_, _02348_, _02346_);
  and (_02350_, _02349_, _02341_);
  and (_02351_, _06205_, _06109_);
  or (_02352_, _02351_, _06202_);
  or (_02353_, _02352_, _02098_);
  or (_02354_, _02353_, _02350_);
  and (_02355_, _02354_, _02338_);
  or (_02356_, _02355_, _06172_);
  or (_02357_, _02151_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_02358_, _02357_, _04856_);
  and (_01931_, _02358_, _02356_);
  not (_02359_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  nor (_02360_, _02151_, _02359_);
  or (_02361_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _06104_);
  or (_02362_, _02361_, _06180_);
  and (_02363_, _02362_, _06202_);
  and (_02364_, _02330_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_02365_, _02364_, _02329_);
  or (_02366_, _06199_, _06103_);
  and (_02367_, _02366_, _02365_);
  or (_02368_, _02367_, _06184_);
  or (_02369_, _02361_, _02139_);
  and (_02370_, _02369_, _02138_);
  and (_02371_, _02370_, _02368_);
  and (_02372_, _06182_, _06103_);
  or (_02373_, _02372_, _06179_);
  or (_02374_, _02373_, _02371_);
  and (_02375_, _02374_, _02363_);
  or (_02376_, _02342_, _02359_);
  nand (_02377_, _02376_, _02345_);
  or (_02379_, _06222_, _06103_);
  and (_02381_, _02379_, _02377_);
  or (_02382_, _02381_, _06210_);
  or (_02383_, _02361_, _02118_);
  and (_02384_, _02383_, _02110_);
  and (_02385_, _02384_, _02382_);
  and (_02386_, _06208_, _06103_);
  or (_02387_, _02386_, _06205_);
  or (_02388_, _02387_, _02385_);
  or (_02389_, _02361_, _06206_);
  and (_02390_, _02389_, _02099_);
  and (_02391_, _02390_, _02388_);
  or (_02392_, _02391_, _02375_);
  and (_02394_, _02392_, _06235_);
  or (_02395_, _02394_, _02360_);
  and (_01943_, _02395_, _04856_);
  and (_01953_, _07173_, _04856_);
  and (_01960_, _07124_, _04856_);
  and (_01962_, _07053_, _04856_);
  and (_01964_, _06991_, _04856_);
  and (_02396_, _07855_, _06143_);
  or (_02397_, _02396_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_02398_, _02397_, _06129_);
  nand (_02399_, _02396_, _06088_);
  and (_02400_, _02399_, _02398_);
  and (_02401_, _06410_, _06127_);
  or (_02402_, _02401_, _02400_);
  and (_02016_, _02402_, _04856_);
  and (_02403_, _06494_, _06143_);
  or (_02404_, _02403_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_02405_, _02404_, _06129_);
  nand (_02406_, _02403_, _06088_);
  and (_02407_, _02406_, _02405_);
  and (_02409_, _06705_, _06127_);
  or (_02410_, _02409_, _02407_);
  and (_02022_, _02410_, _04856_);
  and (_02411_, _06270_, _04990_);
  or (_02412_, _02411_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_02413_, _02412_, _06276_);
  nand (_02414_, _02411_, _06088_);
  and (_02415_, _02414_, _02413_);
  and (_02416_, _06997_, _06275_);
  or (_02417_, _02416_, _02415_);
  and (_02036_, _02417_, _04856_);
  and (_02418_, _06269_, _06135_);
  and (_02419_, _07642_, _02418_);
  nand (_02420_, _02418_, _04984_);
  and (_02421_, _02418_, _12258_);
  or (_02422_, _02421_, _02420_);
  and (_02423_, _02422_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  or (_02425_, _02423_, _06275_);
  or (_02426_, _02425_, _02419_);
  nand (_02427_, _06275_, _05669_);
  and (_02428_, _02427_, _04856_);
  and (_02042_, _02428_, _02426_);
  not (_02429_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  nor (_02430_, _02421_, _02429_);
  or (_02431_, _02430_, _06275_);
  and (_02432_, _04985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_02433_, _02432_, _07602_);
  and (_02434_, _02433_, _06270_);
  or (_02435_, _02434_, _02431_);
  or (_02436_, _06705_, _06276_);
  and (_02437_, _02436_, _04856_);
  and (_02049_, _02437_, _02435_);
  and (_02439_, _06270_, _06146_);
  or (_02440_, _02439_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_02441_, _02440_, _06276_);
  nand (_02442_, _02439_, _06088_);
  and (_02443_, _02442_, _02441_);
  nor (_02444_, _06276_, _05287_);
  or (_02445_, _02444_, _02443_);
  and (_02054_, _02445_, _04856_);
  and (_02446_, _06297_, _04990_);
  and (_02447_, _02446_, _06088_);
  nor (_02448_, _02446_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_02449_, _02448_, _02447_);
  nand (_02450_, _02449_, _06305_);
  nand (_02451_, _06369_, _06304_);
  and (_02453_, _02451_, _04856_);
  and (_02062_, _02453_, _02450_);
  and (_02455_, _06297_, _05520_);
  nand (_02456_, _02455_, _06088_);
  or (_02457_, _02455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_02458_, _02457_, _06305_);
  and (_02459_, _02458_, _02456_);
  nor (_02460_, _06305_, _05669_);
  or (_02462_, _02460_, _02459_);
  and (_02072_, _02462_, _04856_);
  and (_02463_, _04985_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_02464_, _02463_, _07602_);
  and (_02465_, _02464_, _06297_);
  nand (_02466_, _06297_, _12258_);
  and (_02467_, _02466_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_02468_, _02467_, _06304_);
  or (_02469_, _02468_, _02465_);
  or (_02470_, _06705_, _06305_);
  and (_02471_, _02470_, _04856_);
  and (_02082_, _02471_, _02469_);
  and (_02472_, _06297_, _06146_);
  nand (_02473_, _02472_, _06088_);
  or (_02474_, _02472_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  and (_02475_, _02474_, _06305_);
  and (_02476_, _02475_, _02473_);
  nor (_02477_, _06305_, _05287_);
  or (_02478_, _02477_, _02476_);
  and (_02091_, _02478_, _04856_);
  and (_02479_, _09212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_02480_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_02482_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  or (_02484_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  nand (_02485_, _02482_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_02487_, _02485_, _02484_);
  and (_02137_, _02487_, _02321_);
  not (_02488_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  and (_02489_, _09215_, _02488_);
  and (_02490_, _02489_, _09236_);
  nor (_02491_, _09215_, _01113_);
  or (_02492_, _02491_, _02490_);
  and (_02493_, _02492_, _09212_);
  nand (_02494_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nor (_02495_, _02494_, _09211_);
  nor (_02496_, _02495_, _02493_);
  nor (_02497_, _02496_, _09210_);
  or (_02498_, _02497_, _09237_);
  and (_02159_, _02498_, _02321_);
  nand (_02499_, _02490_, _09211_);
  nand (_02500_, _02499_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_02501_, _02500_, _09237_);
  or (_02502_, _02501_, _09206_);
  and (_02198_, _02502_, _04856_);
  or (_02504_, _12818_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_02505_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _09249_);
  or (_02506_, _02505_, _08087_);
  and (_02507_, _02506_, _04856_);
  and (_02208_, _02507_, _02504_);
  nor (_02508_, _02479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_02509_, _02508_, _02480_);
  and (_02224_, _02509_, _02321_);
  or (_02510_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nand (_02511_, _06238_, _02015_);
  and (_02513_, _02511_, _04856_);
  and (_02235_, _02513_, _02510_);
  nor (_02514_, _09212_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_02515_, _02514_, _02479_);
  and (_02239_, _02515_, _02321_);
  and (_02340_, _06347_, _04856_);
  and (_02516_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  not (_02517_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nor (_02518_, _06238_, _02517_);
  or (_02519_, _02518_, _02516_);
  and (_02378_, _02519_, _04856_);
  and (_02521_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  and (_02522_, _08790_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_02523_, _07411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_02524_, _02523_, _02522_);
  and (_02525_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_02526_, _07429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_02527_, _02526_, _02525_);
  or (_02528_, _02527_, _02524_);
  and (_02529_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_02530_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_02531_, _02530_, _02529_);
  and (_02532_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_02533_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_02534_, _02533_, _02532_);
  or (_02535_, _02534_, _02531_);
  or (_02536_, _02535_, _02528_);
  and (_02537_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_02538_, _07463_, _00593_);
  or (_02539_, _02538_, _02537_);
  and (_02540_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_02541_, _07473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_02542_, _02541_, _02540_);
  or (_02544_, _02542_, _02539_);
  not (_02546_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_02547_, _07486_, _02546_);
  and (_02549_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  or (_02551_, _02549_, _02547_);
  and (_02553_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_02554_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_02556_, _02554_, _02553_);
  or (_02557_, _02556_, _02551_);
  or (_02559_, _02557_, _02544_);
  or (_02561_, _02559_, _02536_);
  and (_02562_, _08028_, _07346_);
  and (_02563_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  or (_02564_, _02563_, _02562_);
  and (_02565_, _07389_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_02566_, _07494_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_02567_, _02566_, _02565_);
  or (_02568_, _02567_, _02564_);
  and (_02569_, _01877_, _07507_);
  and (_02570_, _01916_, _07539_);
  or (_02571_, _02570_, _02569_);
  and (_02572_, _01735_, _07547_);
  and (_02574_, _01606_, _07552_);
  or (_02576_, _02574_, _02572_);
  or (_02578_, _02576_, _02571_);
  or (_02579_, _02578_, _02568_);
  and (_02580_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_02581_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_02582_, _02581_, _02580_);
  or (_02583_, _02582_, _02579_);
  or (_02584_, _02583_, _02561_);
  and (_02585_, _02584_, _08004_);
  or (_02586_, _02585_, _07390_);
  or (_02587_, _02586_, _02521_);
  or (_02589_, _08786_, _05641_);
  and (_02591_, _02589_, _04856_);
  and (_02393_, _02591_, _02587_);
  nor (_02593_, _02480_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_02594_, _02593_, _02482_);
  and (_02408_, _02594_, _02321_);
  nor (_02595_, _07390_, rst);
  and (_02424_, _02595_, _08787_);
  and (_02596_, _09023_, _04987_);
  and (_02597_, _02596_, _05510_);
  and (_02598_, _02597_, _08070_);
  and (_02599_, _02598_, _06705_);
  and (_02600_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  and (_02601_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  nor (_02602_, _02601_, _02600_);
  nor (_02603_, _02602_, _09206_);
  and (_02604_, _02597_, _08060_);
  and (_02605_, _02604_, _05670_);
  or (_02606_, _02605_, _02603_);
  or (_02607_, _02606_, _02599_);
  and (_02438_, _02607_, _04856_);
  and (_02608_, _08067_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_02609_, _02608_, _10230_);
  or (_02610_, _02609_, _10232_);
  and (_02611_, _08085_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_02612_, _02611_, _02610_);
  nand (_02613_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _04856_);
  nor (_02614_, _02613_, _12818_);
  or (_02452_, _02614_, _02612_);
  and (_02615_, _02604_, _06705_);
  and (_02616_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_02617_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nor (_02618_, _02617_, _02616_);
  nor (_02619_, _02618_, _09206_);
  and (_02620_, _02598_, _06033_);
  or (_02621_, _02620_, _02619_);
  or (_02622_, _02621_, _02615_);
  and (_02454_, _02622_, _04856_);
  and (_02623_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  and (_02624_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nor (_02626_, _02624_, _02623_);
  nor (_02628_, _02626_, _09206_);
  and (_02629_, _09223_, _05718_);
  or (_02630_, _02629_, _02628_);
  and (_02631_, _09207_, _05288_);
  or (_02632_, _02631_, _02630_);
  and (_02461_, _02632_, _04856_);
  not (_02633_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_02634_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_02635_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_02636_, _06316_, _02635_);
  nor (_02638_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _02546_);
  or (_02639_, _02638_, _02636_);
  nor (_02640_, _02639_, _02634_);
  nand (_02641_, _02640_, _02633_);
  nor (_02642_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor (_02643_, _02642_, _02640_);
  nand (_02644_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_02645_, _02644_, _02643_);
  and (_02646_, _02645_, _04856_);
  and (_02481_, _02646_, _02641_);
  and (_02483_, _02643_, _04856_);
  not (_02647_, _08082_);
  or (_02648_, _08068_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or (_02649_, _02648_, _02044_);
  and (_02650_, _02649_, _02647_);
  or (_02651_, _02650_, rxd_i);
  and (_02652_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], rxd_i);
  nor (_02653_, _02652_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  and (_02654_, _02653_, _08067_);
  and (_02656_, _02654_, _08062_);
  nor (_02657_, _02656_, _10231_);
  and (_02658_, _02657_, _02651_);
  or (_02659_, _02658_, _09249_);
  not (_02660_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  or (_02661_, _08087_, _09249_);
  nand (_02663_, _02661_, _02660_);
  and (_02665_, _02663_, _04856_);
  and (_02486_, _02665_, _02659_);
  and (_02666_, _10232_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_02667_, _08077_, _08072_);
  or (_02669_, _02667_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_02671_, _08077_, _08069_);
  and (_02672_, _02671_, _02647_);
  and (_02674_, _02672_, _02669_);
  or (_02675_, _02674_, _02666_);
  and (_02676_, _02675_, _08085_);
  or (_02503_, _02676_, _02271_);
  not (_02677_, _12761_);
  or (_02678_, _02677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_02679_, _08087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_02680_, _02679_, _08085_);
  and (_02681_, _02680_, _02678_);
  or (_02520_, _02681_, _02167_);
  and (_02682_, _09017_, _06146_);
  nand (_02683_, _02682_, _06088_);
  or (_02684_, _02682_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_02685_, _02684_, _06093_);
  and (_02686_, _02685_, _02683_);
  nand (_02687_, _09024_, _05287_);
  or (_02689_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_02690_, _02689_, _05510_);
  and (_02692_, _02690_, _02687_);
  and (_02694_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_02695_, _02694_, rst);
  or (_02696_, _02695_, _02692_);
  or (_02543_, _02696_, _02686_);
  and (_02698_, _08988_, _07855_);
  nand (_02699_, _02698_, _06088_);
  or (_02700_, _02698_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02701_, _02700_, _06093_);
  and (_02702_, _02701_, _02699_);
  not (_02703_, _08994_);
  or (_02704_, _02703_, _06410_);
  or (_02705_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02706_, _02705_, _05510_);
  and (_02707_, _02706_, _02704_);
  and (_02709_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_02711_, _02709_, rst);
  or (_02713_, _02711_, _02707_);
  or (_02545_, _02713_, _02702_);
  not (_02714_, _05631_);
  or (_02715_, _06054_, _02714_);
  or (_02716_, _05631_, _06053_);
  and (_02717_, _02716_, _05583_);
  and (_02718_, _02717_, _02715_);
  and (_02719_, _05497_, ABINPUT000000[0]);
  and (_02721_, _05499_, ABINPUT000[0]);
  or (_02722_, _02721_, _02719_);
  nand (_02723_, _05431_, _05340_);
  and (_02725_, _05433_, _05455_);
  and (_02727_, _02725_, _02723_);
  or (_02729_, _02727_, _02722_);
  or (_02730_, _02729_, _02718_);
  and (_02731_, _02730_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_02732_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  and (_02733_, _02732_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_02734_, _02733_, _08277_);
  or (_02735_, _02734_, _02731_);
  not (_02736_, _06494_);
  nand (_02737_, _02736_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  nand (_02738_, _02737_, _08277_);
  or (_02739_, _02738_, _07602_);
  and (_02741_, _02739_, _06935_);
  and (_02742_, _02741_, _02735_);
  and (_02743_, _06934_, _06705_);
  or (_02744_, _02743_, _02742_);
  and (_02548_, _02744_, _04856_);
  and (_02745_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_02746_, _02745_, _12766_);
  and (_02550_, _02746_, _04856_);
  and (_02747_, _09132_, _07855_);
  nand (_02748_, _02747_, _06088_);
  or (_02750_, _02747_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_02752_, _02750_, _06093_);
  and (_02753_, _02752_, _02748_);
  and (_02754_, _09138_, _06410_);
  and (_02755_, _09139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_02757_, _02755_, _02754_);
  and (_02758_, _02757_, _05510_);
  and (_02759_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_02760_, _02759_, rst);
  or (_02761_, _02760_, _02758_);
  or (_02552_, _02761_, _02753_);
  and (_02762_, _09116_, _06494_);
  or (_02764_, _02762_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_02765_, _02764_, _06093_);
  nand (_02766_, _02762_, _06088_);
  and (_02767_, _02766_, _02765_);
  and (_02769_, _09123_, _06705_);
  and (_02770_, _09124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_02772_, _02770_, _02769_);
  and (_02773_, _02772_, _05510_);
  and (_02774_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_02775_, _02774_, rst);
  or (_02777_, _02775_, _02773_);
  or (_02555_, _02777_, _02767_);
  and (_02778_, _09116_, _06091_);
  or (_02779_, _02778_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_02780_, _02779_, _06093_);
  nand (_02781_, _02778_, _06088_);
  and (_02783_, _02781_, _02780_);
  and (_02784_, _09123_, _05718_);
  nor (_02785_, _09123_, _01891_);
  or (_02786_, _02785_, _02784_);
  and (_02788_, _02786_, _05510_);
  nor (_02789_, _06092_, _01891_);
  or (_02790_, _02789_, rst);
  or (_02791_, _02790_, _02788_);
  or (_02558_, _02791_, _02783_);
  or (_02793_, _02045_, _09251_);
  and (_02794_, _02793_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_02795_, _02794_, _01937_);
  and (_02560_, _02795_, _04856_);
  and (_02796_, _09017_, _05520_);
  nand (_02797_, _02796_, _06088_);
  or (_02799_, _02796_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02800_, _02799_, _06093_);
  and (_02801_, _02800_, _02797_);
  nand (_02802_, _09024_, _05669_);
  or (_02803_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02805_, _02803_, _05510_);
  and (_02807_, _02805_, _02802_);
  nor (_02808_, _06092_, _08839_);
  or (_02810_, _02808_, rst);
  or (_02811_, _02810_, _02807_);
  or (_02573_, _02811_, _02801_);
  and (_02812_, _08988_, _05520_);
  nand (_02814_, _02812_, _06088_);
  or (_02815_, _02812_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_02817_, _02815_, _06093_);
  and (_02818_, _02817_, _02814_);
  nand (_02819_, _08994_, _05669_);
  or (_02820_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_02821_, _02820_, _05510_);
  and (_02822_, _02821_, _02819_);
  nor (_02823_, _06092_, _08834_);
  or (_02824_, _02823_, rst);
  or (_02825_, _02824_, _02822_);
  or (_02575_, _02825_, _02818_);
  and (_02826_, _08988_, _06146_);
  nand (_02827_, _02826_, _06088_);
  or (_02828_, _02826_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02830_, _02828_, _06093_);
  and (_02831_, _02830_, _02827_);
  nand (_02832_, _08994_, _05287_);
  or (_02834_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02835_, _02834_, _05510_);
  and (_02837_, _02835_, _02832_);
  and (_02838_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_02840_, _02838_, rst);
  or (_02841_, _02840_, _02837_);
  or (_02577_, _02841_, _02831_);
  and (_02842_, _09132_, _06146_);
  nand (_02843_, _02842_, _06088_);
  or (_02844_, _02842_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_02845_, _02844_, _06093_);
  and (_02846_, _02845_, _02843_);
  nor (_02848_, _09139_, _05287_);
  and (_02849_, _09139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02850_, _02849_, _02848_);
  and (_02851_, _02850_, _05510_);
  and (_02852_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02853_, _02852_, rst);
  or (_02854_, _02853_, _02851_);
  or (_02588_, _02854_, _02846_);
  and (_02855_, _09116_, _04990_);
  or (_02856_, _02855_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_02857_, _02856_, _06093_);
  nand (_02858_, _02855_, _06088_);
  and (_02859_, _02858_, _02857_);
  and (_02861_, _09123_, _06997_);
  and (_02862_, _09124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_02863_, _02862_, _02861_);
  and (_02865_, _02863_, _05510_);
  and (_02866_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_02867_, _02866_, rst);
  or (_02868_, _02867_, _02865_);
  or (_02590_, _02868_, _02859_);
  and (_02870_, _09116_, _07855_);
  or (_02871_, _02870_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_02872_, _02871_, _06093_);
  nand (_02873_, _02870_, _06088_);
  and (_02874_, _02873_, _02872_);
  and (_02875_, _09123_, _06410_);
  and (_02876_, _09124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_02878_, _02876_, _02875_);
  and (_02879_, _02878_, _05510_);
  and (_02880_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_02881_, _02880_, rst);
  or (_02882_, _02881_, _02879_);
  or (_02592_, _02882_, _02874_);
  and (_02884_, _09132_, _05520_);
  nand (_02885_, _02884_, _06088_);
  or (_02886_, _02884_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_02888_, _02886_, _06093_);
  and (_02889_, _02888_, _02885_);
  nor (_02890_, _09139_, _05669_);
  nor (_02891_, _09138_, _08845_);
  or (_02892_, _02891_, _02890_);
  and (_02893_, _02892_, _05510_);
  nor (_02894_, _06092_, _08845_);
  or (_02895_, _02894_, rst);
  or (_02897_, _02895_, _02893_);
  or (_02625_, _02897_, _02889_);
  and (_02899_, _09132_, _06494_);
  nand (_02900_, _02899_, _06088_);
  or (_02901_, _02899_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_02902_, _02901_, _06093_);
  and (_02903_, _02902_, _02900_);
  and (_02904_, _09138_, _06705_);
  and (_02905_, _09139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02907_, _02905_, _02904_);
  and (_02908_, _02907_, _05510_);
  and (_02909_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02910_, _02909_, rst);
  or (_02912_, _02910_, _02908_);
  or (_02627_, _02912_, _02903_);
  nand (_02914_, _01352_, _12258_);
  and (_02915_, _02914_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_02916_, _04985_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_02917_, _02916_, _07602_);
  and (_02918_, _02917_, _01352_);
  or (_02919_, _02918_, _02915_);
  and (_02920_, _02919_, _06093_);
  and (_02921_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_02922_, _01361_, _06552_);
  or (_02924_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_02926_, _02924_, _05510_);
  and (_02927_, _02926_, _02922_);
  or (_02928_, _02927_, _02921_);
  or (_02929_, _02928_, _02920_);
  and (_02637_, _02929_, _04856_);
  and (_02930_, _01352_, _06091_);
  nand (_02931_, _02930_, _06088_);
  or (_02932_, _02930_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_02933_, _02932_, _06093_);
  and (_02935_, _02933_, _02931_);
  and (_02937_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_02938_, _01361_, _07897_);
  or (_02939_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_02940_, _02939_, _05510_);
  and (_02942_, _02940_, _02938_);
  or (_02943_, _02942_, _02937_);
  or (_02944_, _02943_, _02935_);
  and (_02655_, _02944_, _04856_);
  and (_02945_, _09132_, _04986_);
  nand (_02947_, _02945_, _06088_);
  or (_02948_, _02945_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_02949_, _02948_, _06093_);
  and (_02951_, _02949_, _02947_);
  nor (_02952_, _09139_, _06032_);
  nor (_02953_, _09138_, _01860_);
  or (_02955_, _02953_, _02952_);
  and (_02956_, _02955_, _05510_);
  nor (_02957_, _06092_, _01860_);
  or (_02958_, _02957_, rst);
  or (_02959_, _02958_, _02956_);
  or (_02662_, _02959_, _02951_);
  and (_02960_, _09132_, _04990_);
  nand (_02961_, _02960_, _06088_);
  or (_02963_, _02960_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_02965_, _02963_, _06093_);
  and (_02966_, _02965_, _02961_);
  and (_02967_, _09138_, _06997_);
  and (_02969_, _09139_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_02970_, _02969_, _02967_);
  and (_02971_, _02970_, _05510_);
  and (_02972_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_02973_, _02972_, rst);
  or (_02974_, _02973_, _02971_);
  or (_02664_, _02974_, _02966_);
  and (_02975_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  and (_02976_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  nor (_02977_, _02976_, _02975_);
  nor (_02978_, _02977_, _09206_);
  and (_02979_, _09223_, _06410_);
  or (_02980_, _02979_, _02978_);
  and (_02981_, _09207_, _05718_);
  or (_02982_, _02981_, _02980_);
  and (_02668_, _02982_, _04856_);
  nand (_02984_, _08988_, _12258_);
  and (_02985_, _02984_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02986_, _04985_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_02987_, _02986_, _07602_);
  and (_02989_, _02987_, _08988_);
  or (_02990_, _02989_, _02985_);
  and (_02991_, _02990_, _06093_);
  or (_02992_, _02703_, _06705_);
  or (_02993_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02994_, _02993_, _05510_);
  and (_02995_, _02994_, _02992_);
  and (_02996_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_02997_, _02996_, rst);
  or (_02998_, _02997_, _02995_);
  or (_02670_, _02998_, _02991_);
  and (_03000_, _05517_, _04999_);
  nand (_03002_, _03000_, _06088_);
  or (_03003_, _03000_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_03004_, _03003_, _06093_);
  and (_03005_, _03004_, _03002_);
  or (_03006_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  nand (_03007_, _08994_, _06032_);
  and (_03008_, _03007_, _05510_);
  and (_03009_, _03008_, _03006_);
  nor (_03010_, _06092_, _01727_);
  or (_03011_, _03010_, rst);
  or (_03012_, _03011_, _03009_);
  or (_02673_, _03012_, _03005_);
  nand (_03013_, _08988_, _04990_);
  or (_03014_, _03013_, _06144_);
  or (_03015_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_03016_, _03015_, _06093_);
  and (_03017_, _03016_, _03014_);
  nand (_03018_, _08994_, _06369_);
  and (_03019_, _03018_, _05510_);
  and (_03020_, _03019_, _03015_);
  and (_03021_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_03022_, _03021_, rst);
  or (_03023_, _03022_, _03020_);
  or (_02688_, _03023_, _03017_);
  and (_03024_, _09017_, _04986_);
  nand (_03025_, _03024_, _06088_);
  or (_03026_, _03024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_03027_, _03026_, _06093_);
  and (_03028_, _03027_, _03025_);
  or (_03029_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nand (_03030_, _09024_, _06032_);
  and (_03031_, _03030_, _05510_);
  and (_03032_, _03031_, _03029_);
  nor (_03033_, _06092_, _01625_);
  or (_03034_, _03033_, rst);
  or (_03035_, _03034_, _03032_);
  or (_02691_, _03035_, _03028_);
  nand (_03037_, _09017_, _04990_);
  or (_03038_, _03037_, _06144_);
  or (_03039_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_03040_, _03039_, _06093_);
  and (_03041_, _03040_, _03038_);
  nand (_03042_, _09024_, _06369_);
  and (_03043_, _03042_, _05510_);
  and (_03044_, _03043_, _03039_);
  and (_03045_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_03046_, _03045_, rst);
  or (_03047_, _03046_, _03044_);
  or (_02693_, _03047_, _03041_);
  and (_03048_, _09017_, _06091_);
  nand (_03049_, _03048_, _06088_);
  or (_03050_, _03048_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03051_, _03050_, _06093_);
  and (_03052_, _03051_, _03049_);
  not (_03053_, _09024_);
  or (_03054_, _03053_, _05718_);
  or (_03055_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_03056_, _03055_, _05510_);
  and (_03057_, _03056_, _03054_);
  nor (_03058_, _06092_, _01630_);
  or (_03059_, _03058_, rst);
  or (_03060_, _03059_, _03057_);
  or (_02697_, _03060_, _03052_);
  and (_03061_, _09116_, _06146_);
  or (_03063_, _03061_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_03064_, _03063_, _06093_);
  nand (_03065_, _03061_, _06088_);
  and (_03066_, _03065_, _03064_);
  nor (_03068_, _09124_, _05287_);
  and (_03069_, _09124_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_03070_, _03069_, _03068_);
  and (_03071_, _03070_, _05510_);
  and (_03072_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_03073_, _03072_, rst);
  or (_03075_, _03073_, _03071_);
  or (_02708_, _03075_, _03066_);
  and (_03076_, _09116_, _05520_);
  or (_03077_, _03076_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_03078_, _03077_, _06093_);
  nand (_03079_, _03076_, _06088_);
  and (_03080_, _03079_, _03078_);
  nor (_03081_, _09124_, _05669_);
  nor (_03082_, _09123_, _08850_);
  or (_03083_, _03082_, _03081_);
  and (_03084_, _03083_, _05510_);
  nor (_03085_, _06092_, _08850_);
  or (_03086_, _03085_, rst);
  or (_03087_, _03086_, _03084_);
  or (_02710_, _03087_, _03080_);
  nand (_03088_, _09115_, _04933_);
  or (_03089_, _03088_, _09132_);
  and (_03090_, _03089_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  nor (_03091_, _04986_, _01886_);
  or (_03092_, _03091_, _07713_);
  and (_03093_, _03092_, _09116_);
  or (_03094_, _03093_, _03090_);
  and (_03095_, _03094_, _06093_);
  nor (_03096_, _09124_, _06032_);
  nor (_03098_, _09123_, _01886_);
  or (_03099_, _03098_, _03096_);
  and (_03100_, _03099_, _05510_);
  nor (_03101_, _06092_, _01886_);
  or (_03103_, _03101_, rst);
  or (_03104_, _03103_, _03100_);
  or (_02712_, _03104_, _03095_);
  and (_03105_, _08988_, _06091_);
  nand (_03106_, _03105_, _06088_);
  or (_03107_, _03105_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03108_, _03107_, _06093_);
  and (_03109_, _03108_, _03106_);
  or (_03110_, _02703_, _05718_);
  or (_03111_, _08994_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_03112_, _03111_, _05510_);
  and (_03113_, _03112_, _03110_);
  nor (_03114_, _06092_, _01738_);
  or (_03115_, _03114_, rst);
  or (_03116_, _03115_, _03113_);
  or (_02720_, _03116_, _03109_);
  and (_03117_, _09017_, _07855_);
  nand (_03118_, _03117_, _06088_);
  or (_03119_, _03117_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03120_, _03119_, _06093_);
  and (_03121_, _03120_, _03118_);
  or (_03122_, _03053_, _06410_);
  or (_03123_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_03124_, _03123_, _05510_);
  and (_03125_, _03124_, _03122_);
  and (_03126_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_03127_, _03126_, rst);
  or (_03128_, _03127_, _03125_);
  or (_02724_, _03128_, _03121_);
  and (_03129_, _09017_, _06494_);
  nand (_03130_, _03129_, _06088_);
  or (_03131_, _03129_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03132_, _03131_, _06093_);
  and (_03133_, _03132_, _03130_);
  or (_03134_, _03053_, _06705_);
  or (_03135_, _09024_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_03136_, _03135_, _05510_);
  and (_03137_, _03136_, _03134_);
  and (_03138_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_03139_, _03138_, rst);
  or (_03140_, _03139_, _03137_);
  or (_02726_, _03140_, _03133_);
  and (_03141_, _09132_, _06091_);
  nand (_03142_, _03141_, _06088_);
  or (_03143_, _03141_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_03144_, _03143_, _06093_);
  and (_03145_, _03144_, _03142_);
  and (_03146_, _09138_, _05718_);
  nor (_03147_, _09138_, _01852_);
  or (_03148_, _03147_, _03146_);
  and (_03149_, _03148_, _05510_);
  nor (_03150_, _06092_, _01852_);
  or (_03151_, _03150_, rst);
  or (_03152_, _03151_, _03149_);
  or (_02728_, _03152_, _03145_);
  or (_03154_, _08087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  nand (_03155_, _01114_, _08073_);
  or (_03156_, _03155_, _08062_);
  nand (_03157_, _03156_, _03154_);
  nand (_02740_, _03157_, _08085_);
  and (_03158_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_03159_, _06238_, _00838_);
  or (_03160_, _03159_, _03158_);
  and (_02749_, _03160_, _04856_);
  and (_02751_, _07334_, _04856_);
  and (_03161_, _09255_, _08064_);
  and (_03162_, _09253_, _03161_);
  nand (_03163_, _03162_, _01939_);
  or (_03164_, _03162_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_03166_, _03164_, _04856_);
  and (_02756_, _03166_, _03163_);
  and (_02763_, _07346_, _04856_);
  and (_03167_, _09218_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_03168_, _09217_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_03169_, _03168_, _03167_);
  and (_03170_, _03169_, _02321_);
  or (_03171_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _02546_);
  and (_03172_, _03171_, _04856_);
  and (_03173_, _03172_, _09223_);
  or (_02768_, _03173_, _03170_);
  not (_03174_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor (_03175_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _08073_);
  not (_03176_, _03175_);
  nor (_03178_, _08060_, _09249_);
  and (_03179_, _03178_, _03176_);
  and (_03181_, _03179_, _02044_);
  nor (_03183_, _03181_, _03174_);
  and (_03184_, _03181_, rxd_i);
  or (_03185_, _03184_, rst);
  or (_02771_, _03185_, _03183_);
  and (_02776_, _07246_, _04856_);
  or (_03187_, _03174_, rxd_i);
  nand (_03188_, _03187_, _08071_);
  or (_03189_, _08072_, _08061_);
  and (_03191_, _03189_, _03188_);
  or (_03192_, _08081_, _08078_);
  or (_03193_, _03192_, _03191_);
  and (_02782_, _03193_, _08085_);
  not (_03194_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_03196_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_03197_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_03199_, _06316_, _03197_);
  or (_03201_, _03199_, _02638_);
  nor (_03203_, _03201_, _03196_);
  nand (_03205_, _03203_, _03194_);
  nor (_03206_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nor (_03207_, _03206_, _03203_);
  nand (_03208_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_03209_, _03208_, _03207_);
  and (_03210_, _03209_, _04856_);
  and (_02787_, _03210_, _03205_);
  and (_03212_, _06041_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_03213_, _09282_, _06043_);
  or (_03214_, _03213_, _03212_);
  and (_02792_, _03214_, _04856_);
  nand (_02798_, _07011_, _04856_);
  and (_03215_, _09282_, _05719_);
  and (_03216_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  or (_03217_, _03216_, _03215_);
  and (_02804_, _03217_, _04856_);
  and (_03218_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_03219_, _00957_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  or (_03220_, _03219_, _03218_);
  and (_02806_, _03220_, _04856_);
  or (_03222_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  not (_03223_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_03224_, _06238_, _03223_);
  and (_03225_, _03224_, _04856_);
  and (_02809_, _03225_, _03222_);
  or (_03226_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  not (_03227_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_03228_, _06238_, _03227_);
  and (_03229_, _03228_, _04856_);
  and (_02813_, _03229_, _03226_);
  and (_03230_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_03231_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_03232_, _06238_, _03231_);
  or (_03233_, _03232_, _03230_);
  and (_02816_, _03233_, _04856_);
  and (_03234_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_03235_, _06238_, _06342_);
  or (_03236_, _03235_, _03234_);
  and (_02829_, _03236_, _04856_);
  and (_03237_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  not (_03238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nor (_03239_, _06238_, _03238_);
  or (_03240_, _03239_, _03237_);
  and (_02833_, _03240_, _04856_);
  and (_03241_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_03242_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_03243_, _06238_, _03242_);
  or (_03244_, _03243_, _03241_);
  and (_02836_, _03244_, _04856_);
  nor (_03245_, _06284_, _06046_);
  and (_03246_, _06046_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_03247_, _03246_, _05673_);
  or (_03248_, _03247_, _03245_);
  or (_03250_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_03251_, _03250_, _04856_);
  and (_02839_, _03251_, _03248_);
  nand (_03252_, _10587_, _06284_);
  or (_03253_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_03254_, _03253_, _04856_);
  and (_02847_, _03254_, _03252_);
  nand (_03255_, _09200_, _06032_);
  or (_03256_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_03257_, _03256_, _04856_);
  and (_02860_, _03257_, _03255_);
  and (_03258_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  nor (_03259_, _01973_, _06284_);
  or (_03260_, _03259_, _03258_);
  and (_02864_, _03260_, _04856_);
  nor (_03261_, _01973_, _05287_);
  and (_03262_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  or (_03263_, _03262_, _03261_);
  and (_02869_, _03263_, _04856_);
  nor (_03264_, _06688_, _06284_);
  and (_03265_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_03266_, _03265_, _03264_);
  and (_02877_, _03266_, _04856_);
  nand (_03267_, _09200_, _06369_);
  or (_03268_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_03269_, _03268_, _04856_);
  and (_02883_, _03269_, _03267_);
  and (_03270_, _09282_, _05009_);
  and (_03271_, _05007_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_03272_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_03273_, _03272_, _05005_);
  or (_03274_, _03273_, _03271_);
  or (_03275_, _03274_, _03270_);
  and (_02887_, _03275_, _04856_);
  or (_03276_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  not (_03277_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_03278_, _06238_, _03277_);
  and (_03279_, _03278_, _04856_);
  and (_02896_, _03279_, _03276_);
  and (_03280_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_03281_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_03282_, _06238_, _03281_);
  or (_03283_, _03282_, _03280_);
  and (_02898_, _03283_, _04856_);
  and (_03284_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_03285_, _06238_, _03223_);
  or (_03286_, _03285_, _03284_);
  and (_02906_, _03286_, _04856_);
  or (_03287_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_03288_, _03287_, _04856_);
  or (_03289_, _09203_, _05718_);
  and (_02911_, _03289_, _03288_);
  and (_03290_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_03291_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_03292_, _06238_, _03291_);
  or (_03293_, _03292_, _03290_);
  and (_02913_, _03293_, _04856_);
  or (_03294_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_03295_, _03294_, _04856_);
  or (_03296_, _09203_, _06410_);
  and (_02923_, _03296_, _03295_);
  or (_03297_, _02677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_03298_, _08087_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_03299_, _03298_, _08085_);
  and (_03300_, _03299_, _03297_);
  or (_02925_, _03300_, _02169_);
  or (_03301_, _09200_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_03302_, _03301_, _04856_);
  nand (_03303_, _09200_, _05287_);
  and (_02934_, _03303_, _03302_);
  or (_03304_, _12818_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_03305_, _02661_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  and (_03306_, _03305_, _04856_);
  and (_02936_, _03306_, _03304_);
  nor (_02941_, _06314_, rst);
  or (_03307_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  not (_03308_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_03309_, _06238_, _03308_);
  and (_03310_, _03309_, _04856_);
  and (_02946_, _03310_, _03307_);
  and (_03311_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  nor (_03312_, _06238_, _03277_);
  or (_03313_, _03312_, _03311_);
  and (_02950_, _03313_, _04856_);
  or (_03314_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nand (_03315_, _06238_, _02517_);
  and (_03316_, _03315_, _04856_);
  and (_02962_, _03316_, _03314_);
  and (_03317_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_03318_, _06238_, _03308_);
  or (_03319_, _03318_, _03317_);
  and (_02964_, _03319_, _04856_);
  or (_03320_, _05678_, _05673_);
  and (_03321_, _03320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_03322_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_03323_, _03322_, _05677_);
  and (_03324_, _01971_, _06705_);
  or (_03325_, _03324_, _03323_);
  or (_03326_, _03325_, _03321_);
  and (_02968_, _03326_, _04856_);
  and (_03327_, _03320_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_03328_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  and (_03329_, _03328_, _05677_);
  nor (_03330_, _01973_, _05669_);
  or (_03331_, _03330_, _03329_);
  or (_03332_, _03331_, _03327_);
  and (_02983_, _03332_, _04856_);
  and (_02988_, _03207_, _04856_);
  and (_03333_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _04856_);
  and (_03334_, _03333_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_03335_, _01075_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_03336_, _01075_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_03337_, _03336_, _03335_);
  and (_03338_, _03337_, _01077_);
  nor (_03339_, _03337_, _01077_);
  or (_03340_, _03339_, _03338_);
  or (_03341_, _03340_, _06911_);
  or (_03342_, _06910_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_03343_, _03342_, _13190_);
  and (_03344_, _03343_, _03341_);
  or (_03001_, _03344_, _03334_);
  or (_03345_, _05919_, _06812_);
  or (_03346_, _05729_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_03347_, _03346_, _04856_);
  and (_03062_, _03347_, _03345_);
  not (_03348_, _00536_);
  and (_03349_, _03348_, _00490_);
  or (_03350_, _13236_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_03097_, _03350_, _04856_);
  and (_03351_, _03097_, _00002_);
  and (_03067_, _03351_, _03349_);
  and (_03352_, _01973_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_03353_, _01971_, _06410_);
  or (_03354_, _03353_, _03352_);
  and (_03074_, _03354_, _04856_);
  or (_03355_, _01048_, _05718_);
  or (_03356_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_03357_, _03356_, _04856_);
  and (_03102_, _03357_, _03355_);
  and (_03153_, _06816_, _04856_);
  and (_03358_, _06705_, _05679_);
  and (_03359_, _06688_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  or (_03360_, _03359_, _03358_);
  or (_03361_, _04861_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  and (_03362_, _03361_, _04856_);
  and (_03165_, _03362_, _03360_);
  and (_03363_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  and (_03364_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  or (_03365_, _03364_, _03363_);
  and (_03177_, _03365_, _04856_);
  and (_03366_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_03367_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  or (_03368_, _03367_, _03366_);
  and (_03180_, _03368_, _04856_);
  and (_03369_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  and (_03370_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  or (_03371_, _03370_, _03369_);
  and (_03182_, _03371_, _04856_);
  and (_03372_, _06598_, _06001_);
  or (_03373_, _03372_, _05956_);
  and (_03374_, _03373_, _05962_);
  not (_03375_, _12131_);
  and (_03376_, _03375_, _05995_);
  or (_03377_, _03376_, _05961_);
  or (_03378_, _03377_, _03374_);
  or (_03379_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _04859_);
  and (_03380_, _03379_, _04856_);
  and (_03186_, _03380_, _03378_);
  and (_03381_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_03382_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or (_03383_, _03382_, _03381_);
  and (_03195_, _03383_, _04856_);
  not (_03384_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_03385_, _01209_, _03384_);
  and (_03386_, _01209_, _03384_);
  or (_03388_, _03386_, _03385_);
  or (_03389_, _03388_, _12547_);
  and (_03390_, _03389_, _04856_);
  nor (_03391_, _13091_, _05022_);
  and (_03392_, _13091_, _05022_);
  nor (_03393_, _03392_, _03391_);
  and (_03394_, _03393_, _01185_);
  nand (_03395_, _03394_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  or (_03396_, _03394_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_03397_, _03396_, _13031_);
  and (_03398_, _03397_, _03395_);
  and (_03399_, _13022_, _05507_);
  and (_03400_, _06847_, _05641_);
  or (_03401_, _01196_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nand (_03402_, _01196_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_03403_, _03402_, _03401_);
  and (_03404_, _03403_, _13042_);
  and (_03405_, _13036_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_03406_, _12829_, _13087_);
  or (_03407_, _03406_, _03405_);
  or (_03408_, _03407_, _03404_);
  or (_03409_, _03408_, _03400_);
  nor (_03410_, _03409_, _03399_);
  nand (_03411_, _03410_, _12547_);
  or (_03412_, _03411_, _03398_);
  and (_03198_, _03412_, _03390_);
  nor (_03200_, _06938_, rst);
  and (_03413_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _08359_);
  and (_03414_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_03415_, _03414_, _03413_);
  and (_03202_, _03415_, _04856_);
  nand (_03416_, _05730_, _00059_);
  nand (_03417_, _03416_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_03418_, _03417_, _12206_);
  and (_03204_, _03418_, _04856_);
  and (_03419_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_03420_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  or (_03421_, _03420_, _03419_);
  and (_03211_, _03421_, _04856_);
  or (_03422_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nand (_03423_, _06238_, _03238_);
  and (_03424_, _03423_, _04856_);
  and (_03249_, _03424_, _03422_);
  and (_03425_, _06370_, _05000_);
  and (_03426_, _05723_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  or (_03427_, _03426_, _03425_);
  and (_03387_, _03427_, _04856_);
  and (_03428_, _01945_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_03429_, _03428_, _06657_);
  and (_03430_, _03429_, _08277_);
  or (_03431_, _07949_, _06144_);
  nor (_03432_, _07951_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_03433_, _03432_, _08277_);
  and (_03434_, _03433_, _03431_);
  or (_03435_, _03434_, _06934_);
  or (_03436_, _03435_, _03430_);
  nand (_03437_, _06934_, _06284_);
  and (_03438_, _03437_, _04856_);
  and (_03471_, _03438_, _03436_);
  and (_03439_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_03440_, _00957_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  or (_03441_, _03440_, _03439_);
  and (_03559_, _03441_, _04856_);
  or (_03442_, _06757_, _06752_);
  or (_03443_, _06787_, _06732_);
  or (_03444_, _06777_, _06620_);
  and (_03445_, _03444_, _06637_);
  or (_03446_, _03445_, _03443_);
  or (_03447_, _03446_, _03442_);
  and (_03448_, _06777_, _05965_);
  or (_03449_, _06835_, _03448_);
  or (_03450_, _07508_, _06871_);
  or (_03451_, _03450_, _03449_);
  and (_03452_, _05998_, _05969_);
  or (_03453_, _12689_, _08242_);
  or (_03454_, _03453_, _03452_);
  or (_03455_, _06786_, _06761_);
  or (_03456_, _03455_, _03454_);
  or (_03457_, _03456_, _03451_);
  or (_03458_, _09071_, _08208_);
  or (_03459_, _03458_, _09079_);
  or (_03460_, _03459_, _09099_);
  or (_03461_, _03460_, _03457_);
  or (_03462_, _03461_, _03447_);
  and (_03463_, _03462_, _05730_);
  and (_03464_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_03465_, _03464_, _03376_);
  or (_03466_, _03465_, _03463_);
  and (_03577_, _03466_, _04856_);
  nor (_03612_, _06947_, rst);
  or (_03467_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand (_03468_, _08367_, _05884_);
  and (_03469_, _03468_, _04856_);
  and (_03641_, _03469_, _03467_);
  and (_03470_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_03472_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or (_03473_, _03472_, _03470_);
  and (_03643_, _03473_, _04856_);
  or (_03474_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand (_03475_, _08367_, _05904_);
  and (_03476_, _03475_, _04856_);
  and (_03647_, _03476_, _03474_);
  and (_03477_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_03478_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  or (_03479_, _03478_, _03477_);
  and (_03653_, _03479_, _04856_);
  and (_03480_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_03481_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  or (_03482_, _03481_, _03480_);
  and (_03677_, _03482_, _04856_);
  and (_03483_, _06041_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  and (_03484_, _06043_, _05718_);
  or (_03485_, _03484_, _03483_);
  and (_03698_, _03485_, _04856_);
  and (_03486_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_03487_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or (_03488_, _03487_, _03486_);
  and (_03706_, _03488_, _04856_);
  and (_03489_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nor (_03490_, _07410_, _12633_);
  nor (_03491_, _07404_, _02635_);
  or (_03492_, _03491_, _03490_);
  and (_03493_, _07429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_03494_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_03495_, _03494_, _03493_);
  or (_03496_, _03495_, _03492_);
  and (_03497_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_03498_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_03499_, _03498_, _03497_);
  and (_03500_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_03501_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_03502_, _03501_, _03500_);
  or (_03503_, _03502_, _03499_);
  or (_03504_, _03503_, _03496_);
  and (_03505_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_03506_, _07463_, _00611_);
  or (_03507_, _03506_, _03505_);
  and (_03508_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_03509_, _07473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_03510_, _03509_, _03508_);
  or (_03511_, _03510_, _03507_);
  nor (_03512_, _07486_, _08073_);
  and (_03513_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_03514_, _03513_, _03512_);
  and (_03515_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_03516_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or (_03517_, _03516_, _03515_);
  or (_03518_, _03517_, _03514_);
  or (_03519_, _03518_, _03511_);
  or (_03520_, _03519_, _03504_);
  and (_03521_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_03522_, _08028_, _07223_);
  or (_03523_, _03522_, _03521_);
  and (_03524_, _07494_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  and (_03525_, _07389_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  or (_03526_, _03525_, _03524_);
  or (_03527_, _03526_, _03523_);
  and (_03528_, _01899_, _07539_);
  and (_03529_, _01869_, _07507_);
  or (_03530_, _03529_, _03528_);
  and (_03531_, _01754_, _07547_);
  and (_03532_, _01619_, _07552_);
  or (_03533_, _03532_, _03531_);
  or (_03534_, _03533_, _03530_);
  or (_03535_, _03534_, _03527_);
  and (_03536_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_03537_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  or (_03538_, _03537_, _03536_);
  or (_03539_, _03538_, _03535_);
  or (_03540_, _03539_, _03520_);
  and (_03541_, _03540_, _08004_);
  or (_03542_, _03541_, _07390_);
  or (_03543_, _03542_, _03489_);
  nand (_03544_, _07390_, _07815_);
  and (_03545_, _03544_, _04856_);
  and (_03708_, _03545_, _03543_);
  and (_03546_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nor (_03547_, _07991_, _04904_);
  nand (_03548_, _03547_, _04858_);
  nand (_03549_, _07943_, _06661_);
  and (_03550_, _07996_, _07997_);
  nand (_03551_, _03550_, _06141_);
  and (_03552_, _03551_, _03549_);
  and (_03553_, _03552_, _03548_);
  nand (_03554_, _03553_, _07958_);
  or (_03555_, _07404_, _12397_);
  or (_03556_, _07410_, _02087_);
  and (_03557_, _03556_, _03555_);
  or (_03558_, _07428_, _12728_);
  or (_03560_, _07420_, _02095_);
  and (_03561_, _03560_, _03558_);
  and (_03562_, _03561_, _03557_);
  nand (_03563_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_03564_, _07441_, _12549_);
  and (_03565_, _03564_, _03563_);
  nand (_03566_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  nand (_03567_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_03568_, _03567_, _03566_);
  and (_03569_, _03568_, _03565_);
  and (_03570_, _03569_, _03562_);
  or (_03571_, _07463_, _00334_);
  nand (_03572_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_03573_, _03572_, _03571_);
  or (_03574_, _07472_, _00834_);
  nand (_03575_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_03576_, _03575_, _03574_);
  and (_03578_, _03576_, _03573_);
  or (_03579_, _07486_, _09271_);
  nand (_03580_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  and (_03581_, _03580_, _03579_);
  nand (_03582_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nand (_03583_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_03584_, _03583_, _03582_);
  and (_03585_, _03584_, _03581_);
  and (_03586_, _03585_, _03578_);
  and (_03587_, _03586_, _03570_);
  nand (_03588_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  or (_03589_, _07503_, _07067_);
  and (_03590_, _03589_, _03588_);
  or (_03591_, _07953_, _08340_);
  or (_03592_, _08025_, _01096_);
  and (_03593_, _03592_, _03591_);
  and (_03595_, _03593_, _03590_);
  nand (_03596_, _01862_, _07507_);
  nand (_03597_, _01888_, _07539_);
  and (_03598_, _03597_, _03596_);
  nand (_03599_, _01627_, _07552_);
  nand (_03600_, _01729_, _07547_);
  and (_03601_, _03600_, _03599_);
  and (_03602_, _03601_, _03598_);
  and (_03603_, _03602_, _03595_);
  nand (_03604_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  nand (_03605_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_03606_, _03605_, _03604_);
  and (_03607_, _03606_, _03603_);
  and (_03608_, _03607_, _03587_);
  or (_03609_, _03608_, _03554_);
  nand (_03610_, _03609_, _08786_);
  or (_03611_, _03610_, _03546_);
  nand (_03613_, _07390_, _07774_);
  and (_03614_, _03613_, _04856_);
  and (_03712_, _03614_, _03611_);
  and (_03615_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_03616_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or (_03617_, _03616_, _03615_);
  and (_03719_, _03617_, _04856_);
  and (_03618_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_03619_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  or (_03620_, _03619_, _03618_);
  and (_03721_, _03620_, _04856_);
  and (_03621_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_03622_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  or (_03623_, _03622_, _03621_);
  and (_03724_, _03623_, _04856_);
  or (_03624_, _12720_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nand (_03625_, _12720_, _08794_);
  and (_03626_, _03625_, _03624_);
  and (_03627_, _03626_, _12715_);
  nor (_03628_, _12715_, _05669_);
  or (_03629_, _03628_, _03627_);
  and (_03726_, _03629_, _04856_);
  or (_03630_, _01048_, _06705_);
  or (_03631_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_03632_, _03631_, _04856_);
  and (_03728_, _03632_, _03630_);
  and (_03633_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  or (_03634_, _07404_, _03197_);
  or (_03635_, _07410_, _12627_);
  and (_03636_, _03635_, _03634_);
  or (_03637_, _07420_, _12791_);
  or (_03638_, _07428_, _12439_);
  and (_03639_, _03638_, _03637_);
  and (_03640_, _03639_, _03636_);
  nand (_03642_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_03644_, _07441_, _12450_);
  and (_03645_, _03644_, _03642_);
  nand (_03646_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nand (_03648_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_03649_, _03648_, _03646_);
  and (_03650_, _03649_, _03645_);
  and (_03651_, _03650_, _03640_);
  or (_03652_, _07463_, _00690_);
  or (_03654_, _07465_, _00706_);
  and (_03655_, _03654_, _03652_);
  or (_03656_, _07472_, _00805_);
  nand (_03657_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_03658_, _03657_, _03656_);
  and (_03659_, _03658_, _03655_);
  or (_03660_, _07486_, _00246_);
  nand (_03661_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  and (_03662_, _03661_, _03660_);
  nand (_03663_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nand (_03664_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_03665_, _03664_, _03663_);
  and (_03666_, _03665_, _03662_);
  and (_03667_, _03666_, _03659_);
  and (_03668_, _03667_, _03651_);
  nand (_03669_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  or (_03670_, _07503_, _07274_);
  and (_03671_, _03670_, _03669_);
  or (_03672_, _08025_, _08313_);
  or (_03673_, _07953_, _08327_);
  and (_03674_, _03673_, _03672_);
  and (_03675_, _03674_, _03671_);
  nand (_03676_, _01893_, _07539_);
  nand (_03678_, _01855_, _07507_);
  and (_03679_, _03678_, _03676_);
  nand (_03680_, _01740_, _07547_);
  nand (_03681_, _01632_, _07552_);
  and (_03682_, _03681_, _03680_);
  and (_03683_, _03682_, _03679_);
  and (_03684_, _03683_, _03675_);
  nand (_03685_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  nand (_03686_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_03687_, _03686_, _03685_);
  and (_03688_, _03687_, _03684_);
  and (_03689_, _03688_, _03668_);
  or (_03690_, _03689_, _03554_);
  nand (_03691_, _03690_, _08786_);
  or (_03692_, _03691_, _03633_);
  nand (_03693_, _07390_, _07897_);
  and (_03694_, _03693_, _04856_);
  and (_03746_, _03694_, _03692_);
  nand (_03695_, _10587_, _05669_);
  or (_03696_, _10587_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_03697_, _03696_, _04856_);
  and (_03751_, _03697_, _03695_);
  or (_03699_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  nand (_03700_, _08367_, _05805_);
  and (_03701_, _03700_, _04856_);
  and (_03754_, _03701_, _03699_);
  or (_03702_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand (_03703_, _08367_, _05782_);
  and (_03704_, _03703_, _04856_);
  and (_03756_, _03704_, _03702_);
  or (_03705_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand (_03707_, _08367_, _05824_);
  and (_03709_, _03707_, _04856_);
  and (_03760_, _03709_, _03705_);
  or (_03710_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand (_03711_, _08367_, _05749_);
  and (_03713_, _03711_, _04856_);
  and (_03763_, _03713_, _03710_);
  and (_03714_, _08037_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_03715_, _07411_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_03716_, _07404_, _12225_);
  or (_03717_, _03716_, _03715_);
  and (_03718_, _07422_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_03720_, _07429_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_03722_, _03720_, _03718_);
  or (_03723_, _03722_, _03717_);
  and (_03725_, _07437_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03727_, _07442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_03729_, _03727_, _03725_);
  and (_03730_, _07449_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03731_, _07455_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_03732_, _03731_, _03730_);
  or (_03733_, _03732_, _03729_);
  or (_03734_, _03733_, _03723_);
  nor (_03735_, _07463_, _00588_);
  and (_03736_, _07466_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  or (_03737_, _03736_, _03735_);
  and (_03738_, _07470_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_03739_, _07473_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_03740_, _03739_, _03738_);
  or (_03741_, _03740_, _03737_);
  and (_03742_, _07487_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_03743_, _07484_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or (_03744_, _03743_, _03742_);
  and (_03745_, _07477_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_03747_, _07479_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_03748_, _03747_, _03745_);
  or (_03749_, _03748_, _03744_);
  or (_03750_, _03749_, _03741_);
  or (_03752_, _03750_, _03734_);
  and (_03753_, _08028_, _07310_);
  and (_03755_, _07500_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_03757_, _03755_, _03753_);
  and (_03758_, _07494_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  and (_03759_, _07389_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  or (_03761_, _03759_, _03758_);
  or (_03762_, _03761_, _03757_);
  and (_03764_, _01747_, _07547_);
  and (_03766_, _01613_, _07552_);
  or (_03767_, _03766_, _03764_);
  and (_03768_, _01844_, _07507_);
  and (_03769_, _01908_, _07539_);
  or (_03770_, _03769_, _03768_);
  or (_03771_, _03770_, _03767_);
  or (_03772_, _03771_, _03762_);
  and (_03773_, _07561_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_03774_, _07943_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_03775_, _03774_, _03773_);
  or (_03776_, _03775_, _03772_);
  or (_03777_, _03776_, _03752_);
  and (_03778_, _03777_, _08004_);
  or (_03780_, _03778_, _07390_);
  or (_03781_, _03780_, _03714_);
  nand (_03782_, _07390_, _06488_);
  and (_03783_, _03782_, _04856_);
  and (_03765_, _03783_, _03781_);
  nand (_03784_, _12393_, _02095_);
  or (_03785_, _12583_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_03786_, _03785_, _12664_);
  or (_03787_, _03786_, _12393_);
  and (_03788_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_03790_, _03788_, _12420_);
  or (_03792_, _03790_, _03787_);
  and (_03793_, _03792_, _03784_);
  or (_03794_, _03793_, _12430_);
  nand (_03795_, _12430_, _06032_);
  and (_03796_, _03795_, _03794_);
  or (_03797_, _03796_, _12389_);
  nand (_03799_, _12389_, _02087_);
  and (_03800_, _03799_, _04856_);
  and (_03779_, _03800_, _03797_);
  or (_03802_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand (_03804_, _08367_, _05881_);
  and (_03806_, _03804_, _04856_);
  and (_03789_, _03806_, _03802_);
  or (_03807_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand (_03808_, _08367_, _05778_);
  and (_03809_, _03808_, _04856_);
  and (_03791_, _03809_, _03807_);
  or (_03810_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand (_03811_, _08367_, _05834_);
  and (_03812_, _03811_, _04856_);
  and (_03798_, _03812_, _03810_);
  or (_03813_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  nand (_03814_, _08367_, _05754_);
  and (_03815_, _03814_, _04856_);
  and (_03801_, _03815_, _03813_);
  or (_03816_, _08367_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand (_03817_, _08367_, _05909_);
  and (_03818_, _03817_, _04856_);
  and (_03803_, _03818_, _03816_);
  and (_03819_, _08367_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_03820_, _12165_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  or (_03821_, _03820_, _03819_);
  and (_03805_, _03821_, _04856_);
  and (_03823_, _12423_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_03824_, _03823_, _12420_);
  and (_03825_, _12411_, _12401_);
  or (_03826_, _03825_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_03827_, _03826_, _02296_);
  or (_03828_, _03827_, _12393_);
  or (_03829_, _03828_, _03824_);
  or (_03830_, _12395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nand (_03831_, _03830_, _03829_);
  nor (_03832_, _03831_, _12430_);
  and (_03833_, _12430_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_03834_, _03833_, _12389_);
  or (_03835_, _03834_, _03832_);
  or (_03836_, _12390_, _06705_);
  and (_03837_, _03836_, _04856_);
  and (_03822_, _03837_, _03835_);
  and (_03838_, _06721_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_03839_, _08242_, _06736_);
  and (_03840_, _06597_, _05848_);
  or (_03841_, _07508_, _03840_);
  or (_03842_, _03841_, _03839_);
  and (_03843_, _03842_, _05773_);
  or (_03844_, _12521_, _06763_);
  or (_03845_, _03844_, _06750_);
  or (_03846_, _03845_, _06889_);
  or (_03847_, _03443_, _08212_);
  or (_03848_, _03847_, _03846_);
  or (_03849_, _06624_, _06612_);
  and (_03850_, _03849_, _05998_);
  or (_03851_, _08208_, _03850_);
  or (_03852_, _03851_, _09083_);
  or (_03853_, _03852_, _06758_);
  or (_03854_, _03853_, _03848_);
  or (_03855_, _03854_, _03843_);
  and (_03856_, _03855_, _06770_);
  or (_03857_, _03856_, _03838_);
  and (_03858_, _12260_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_03859_, _03858_, _12183_);
  and (_03860_, _04985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_03862_, _03860_, _07602_);
  and (_03863_, _03862_, _12177_);
  or (_03864_, _03863_, _03859_);
  or (_03866_, _12185_, _06705_);
  and (_03867_, _03866_, _04856_);
  and (_03861_, _03867_, _03864_);
  and (_03868_, _06238_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_03869_, _06238_, _03227_);
  or (_03870_, _03869_, _03868_);
  and (_03865_, _03870_, _04856_);
  or (_03871_, _01401_, _05641_);
  or (_03872_, _01361_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03873_, _03872_, _05510_);
  and (_03874_, _03873_, _03871_);
  and (_03875_, _08999_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03876_, _01352_, _06268_);
  nand (_03877_, _03876_, _06088_);
  or (_03878_, _03876_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03879_, _03878_, _06093_);
  and (_03880_, _03879_, _03877_);
  or (_03881_, _03880_, _03875_);
  or (_03882_, _03881_, _03874_);
  and (_03916_, _03882_, _04856_);
  and (_03883_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_03884_, _03883_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_03885_, _03231_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_03886_, _03885_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_03887_, _03886_, _03884_);
  nor (_03888_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_03889_, _03888_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_03890_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _03281_);
  and (_03891_, _03890_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_03892_, _03891_, _03889_);
  and (_03893_, _03892_, _03887_);
  and (_03894_, _03893_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_03895_, _03888_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_03896_, _03890_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_03897_, _03896_, _03895_);
  and (_03898_, _03883_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_03899_, _03885_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_03900_, _03899_, _03898_);
  and (_03901_, _03900_, _03897_);
  and (_03902_, _03901_, _06261_);
  nor (_03903_, _03902_, _03894_);
  nor (_03904_, _03903_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_03905_, _03904_);
  and (_03906_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08439_);
  nor (_03907_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_03908_, _03907_, _03906_);
  nor (_03909_, _03908_, _06261_);
  nor (_03910_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_03911_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _09148_);
  nor (_03912_, _03911_, _03910_);
  nor (_03913_, _03912_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_03914_, _03913_, _03909_);
  and (_03915_, _03914_, _03885_);
  nor (_03917_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_03918_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08363_);
  nor (_03919_, _03918_, _03917_);
  nor (_03920_, _03919_, _06261_);
  and (_03921_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_03922_, _06241_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_03923_, _03922_, _03921_);
  and (_03924_, _03923_, _06261_);
  nor (_03925_, _03924_, _03920_);
  and (_03926_, _03925_, _03890_);
  nor (_03927_, _03926_, _03915_);
  nor (_03928_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_03929_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08408_);
  nor (_03930_, _03929_, _03928_);
  nor (_03931_, _03930_, _06261_);
  nor (_03932_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_03933_, _06241_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_03934_, _03933_, _03932_);
  nor (_03935_, _03934_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_03936_, _03935_, _03931_);
  and (_03937_, _03936_, _03883_);
  and (_03938_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _09193_);
  nor (_03939_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_03940_, _03939_, _03938_);
  nor (_03941_, _03940_, _06261_);
  and (_03942_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_03943_, _06241_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_03944_, _03943_, _03942_);
  and (_03945_, _03944_, _06261_);
  nor (_03946_, _03945_, _03941_);
  and (_03947_, _03946_, _03888_);
  nor (_03948_, _03947_, _03937_);
  and (_03949_, _03948_, _03927_);
  and (_03950_, _03885_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_03951_, _03883_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_03952_, _03951_, _03950_);
  and (_03953_, _03888_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_03954_, _03890_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_03955_, _03954_, _03953_);
  and (_03956_, _03955_, _03952_);
  and (_03957_, _03956_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_03958_, _03888_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_03959_, _03890_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_03960_, _03959_, _03958_);
  and (_03961_, _03883_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_03962_, _03885_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_03963_, _03962_, _03961_);
  and (_03964_, _03963_, _03960_);
  and (_03965_, _03964_, _06261_);
  nor (_03966_, _03965_, _03957_);
  nor (_03967_, _03966_, _06241_);
  nor (_03968_, _03967_, _03949_);
  and (_03969_, _03968_, _03905_);
  nor (_03970_, _03969_, _03308_);
  and (_03971_, _03969_, _03308_);
  or (_03972_, _03971_, _03970_);
  and (_03973_, _03883_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_03974_, _03885_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_03975_, _03974_, _03973_);
  and (_03976_, _03888_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_03977_, _03890_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_03978_, _03977_, _03976_);
  and (_03979_, _03978_, _03975_);
  and (_03980_, _03979_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_03981_, _03888_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_03982_, _03890_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_03983_, _03982_, _03981_);
  and (_03984_, _03883_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_03985_, _03885_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_03986_, _03985_, _03984_);
  and (_03987_, _03986_, _03983_);
  and (_03988_, _03987_, _06261_);
  nor (_03989_, _03988_, _03980_);
  nor (_03990_, _03989_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_03991_, _03990_);
  and (_03992_, _03885_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_03993_, _03883_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_03994_, _03993_, _03992_);
  and (_03995_, _03888_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_03996_, _03890_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_03997_, _03996_, _03995_);
  and (_03998_, _03997_, _03994_);
  and (_03999_, _03998_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04000_, _03888_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_04001_, _03890_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_04002_, _04001_, _04000_);
  and (_04003_, _03883_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_04004_, _03885_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_04005_, _04004_, _04003_);
  and (_04006_, _04005_, _04002_);
  and (_04007_, _04006_, _06261_);
  nor (_04008_, _04007_, _03999_);
  nor (_04009_, _04008_, _06241_);
  nor (_04010_, _04009_, _03949_);
  and (_04011_, _04010_, _03991_);
  and (_04012_, _04011_, _03277_);
  nor (_04013_, _04011_, _03277_);
  or (_04015_, _04013_, _04012_);
  or (_04016_, _04015_, _03972_);
  and (_04017_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_04018_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  and (_04019_, _04018_, _04017_);
  and (_04020_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_04021_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04022_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_04023_, _04022_, _04021_);
  and (_04024_, _04023_, _04020_);
  and (_04025_, _04024_, _04019_);
  and (_04026_, _04025_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_04027_, _04025_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_04028_, _04027_, _04026_);
  nand (_04029_, _04028_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or (_04030_, _04028_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_04031_, _04030_, _04029_);
  and (_04032_, _03890_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_04033_, _04032_, _06261_);
  and (_04034_, _03885_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_04035_, _03883_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_04036_, _03888_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  or (_04037_, _04036_, _04035_);
  nor (_04038_, _04037_, _04034_);
  and (_04039_, _04038_, _04033_);
  and (_04040_, _03883_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_04041_, _03885_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nor (_04042_, _04041_, _04040_);
  and (_04043_, _03888_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_04044_, _03890_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_04045_, _04044_, _04043_);
  and (_04046_, _04045_, _04042_);
  and (_04047_, _04046_, _06261_);
  nor (_04048_, _04047_, _04039_);
  nor (_04049_, _04048_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  not (_04050_, _04049_);
  and (_04051_, _03885_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_04052_, _03883_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nor (_04053_, _04052_, _04051_);
  and (_04054_, _03888_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_04055_, _03890_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_04056_, _04055_, _04054_);
  and (_04057_, _04056_, _04053_);
  and (_04058_, _04057_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04059_, _03888_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_04060_, _03890_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nor (_04061_, _04060_, _04059_);
  and (_04062_, _03883_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_04063_, _03885_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nor (_04064_, _04063_, _04062_);
  and (_04066_, _04064_, _04061_);
  and (_04067_, _04066_, _06261_);
  nor (_04068_, _04067_, _04058_);
  nor (_04069_, _04068_, _06241_);
  nor (_04070_, _04069_, _03949_);
  and (_04071_, _04070_, _04050_);
  and (_04072_, _04071_, _02517_);
  nor (_04073_, _04071_, _02517_);
  or (_04074_, _04073_, _04072_);
  or (_04075_, _04074_, _04031_);
  or (_04076_, _04075_, _04016_);
  and (_04077_, _04026_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_04078_, _04077_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_04079_, _04077_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_04080_, _04079_, _04078_);
  nand (_04081_, _04080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  or (_04082_, _04080_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_04083_, _04082_, _04081_);
  nor (_04084_, _04026_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_04085_, _04084_, _04077_);
  and (_04086_, _04085_, _06342_);
  nor (_04087_, _04085_, _06342_);
  or (_04088_, _04087_, _04086_);
  or (_04089_, _04088_, _04083_);
  nor (_04090_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_04091_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_04092_, _04091_, _04090_);
  and (_04093_, _04079_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  or (_04094_, _04093_, _04092_);
  nand (_04095_, _04093_, _04092_);
  and (_04096_, _04095_, _04094_);
  nor (_04097_, _04079_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04098_, _04097_, _04093_);
  and (_04099_, _04098_, _00838_);
  nor (_04100_, _04098_, _00838_);
  or (_04101_, _04100_, _04099_);
  or (_04102_, _04101_, _04096_);
  or (_04103_, _04102_, _04089_);
  or (_04104_, _04103_, _04076_);
  not (_04105_, _03888_);
  and (_04106_, _03883_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04107_, _04106_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04108_, _04106_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_04109_, _04108_, _04107_);
  and (_04110_, _04109_, _08363_);
  not (_04111_, _03917_);
  nor (_04112_, _03883_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04113_, _04112_, _04106_);
  and (_04114_, _04113_, _04111_);
  not (_04115_, _04114_);
  nor (_04116_, _04115_, _04110_);
  not (_04117_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_04118_, _04109_, _04117_);
  and (_04119_, _04109_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_04120_, _04119_, _04118_);
  nor (_04121_, _04120_, _04113_);
  nor (_04122_, _04121_, _04116_);
  nor (_04123_, _04122_, _04105_);
  not (_04124_, _04123_);
  not (_04125_, _04113_);
  nor (_04126_, _04109_, \oc8051_symbolic_cxrom1.regvalid [6]);
  not (_04127_, _03890_);
  or (_04128_, _03906_, _04127_);
  or (_04129_, _04128_, _04126_);
  nor (_04130_, _04109_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not (_04131_, _03883_);
  or (_04132_, _03938_, _04131_);
  or (_04133_, _04132_, _04130_);
  and (_04134_, _04133_, _04129_);
  or (_04135_, _04134_, _04125_);
  not (_04136_, _04106_);
  not (_04137_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_04138_, _04109_, _04137_);
  and (_04139_, _04109_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_04140_, _04139_, _04138_);
  or (_04141_, _04140_, _04136_);
  not (_04142_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_04143_, _04109_, _04142_);
  and (_04144_, _04109_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_04145_, _04144_, _04143_);
  nand (_04146_, _04125_, _03890_);
  or (_04147_, _04146_, _04145_);
  and (_04148_, _04147_, _04141_);
  and (_04149_, _04148_, _04135_);
  not (_04150_, _03885_);
  and (_04151_, _04109_, _08408_);
  not (_04152_, _04151_);
  nor (_04153_, _03928_, _04125_);
  and (_04154_, _04153_, _04152_);
  nor (_04155_, _04109_, _08399_);
  and (_04156_, _04109_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_04157_, _04156_, _04155_);
  nor (_04158_, _04157_, _04113_);
  nor (_04159_, _04158_, _04154_);
  nor (_04160_, _04159_, _04150_);
  not (_04161_, _04160_);
  and (_04162_, _04161_, _04149_);
  and (_04163_, _04162_, _04124_);
  and (_04164_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_04165_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_04166_, _04165_, _04164_);
  and (_04167_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_04168_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_04169_, _04168_, _04167_);
  and (_04170_, _04169_, _04166_);
  and (_04171_, _04170_, _04125_);
  not (_04172_, _04109_);
  and (_04173_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_04174_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_04175_, _04174_, _04173_);
  and (_04176_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_04177_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_04178_, _04177_, _04176_);
  and (_04179_, _04178_, _04175_);
  and (_04180_, _04179_, _04113_);
  or (_04181_, _04180_, _04172_);
  nor (_04182_, _04181_, _04171_);
  and (_04183_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_04184_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_04185_, _04184_, _04183_);
  and (_04186_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_04187_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_04188_, _04187_, _04186_);
  and (_04189_, _04188_, _04185_);
  nor (_04190_, _04189_, _04113_);
  and (_04191_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_04192_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_04193_, _04192_, _04191_);
  and (_04194_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_04195_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_04196_, _04195_, _04194_);
  and (_04197_, _04196_, _04193_);
  nor (_04198_, _04197_, _04125_);
  or (_04199_, _04198_, _04190_);
  and (_04200_, _04199_, _04172_);
  nor (_04201_, _04200_, _04182_);
  nor (_04202_, _04201_, _04163_);
  nand (_04203_, _04202_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_04204_, _04202_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04205_, _04204_, _04203_);
  and (_04206_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_04207_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_04208_, _04207_, _04206_);
  and (_04209_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_04210_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_04211_, _04210_, _04209_);
  and (_04212_, _04211_, _04208_);
  and (_04213_, _04212_, _04125_);
  and (_04214_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_04215_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_04216_, _04215_, _04214_);
  and (_04217_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_04218_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_04219_, _04218_, _04217_);
  and (_04220_, _04219_, _04216_);
  and (_04221_, _04220_, _04113_);
  or (_04222_, _04221_, _04109_);
  nor (_04223_, _04222_, _04213_);
  and (_04224_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_04225_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_04226_, _04225_, _04224_);
  and (_04227_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_04228_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_04229_, _04228_, _04227_);
  and (_04230_, _04229_, _04226_);
  nor (_04231_, _04230_, _04113_);
  and (_04232_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_04233_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_04234_, _04233_, _04232_);
  and (_04235_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_04236_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_04237_, _04236_, _04235_);
  and (_04238_, _04237_, _04234_);
  nor (_04239_, _04238_, _04125_);
  or (_04240_, _04239_, _04231_);
  and (_04241_, _04240_, _04109_);
  nor (_04242_, _04241_, _04223_);
  nor (_04243_, _04242_, _04163_);
  and (_04244_, _04243_, _03291_);
  nor (_04245_, _04243_, _03291_);
  or (_04246_, _04245_, _04244_);
  or (_04247_, _04246_, _04205_);
  and (_04248_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_04249_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_04250_, _04249_, _04248_);
  and (_04251_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_04252_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_04253_, _04252_, _04251_);
  and (_04254_, _04253_, _04250_);
  and (_04255_, _04254_, _04125_);
  and (_04256_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_04257_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_04258_, _04257_, _04256_);
  and (_04259_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_04260_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_04261_, _04260_, _04259_);
  and (_04262_, _04261_, _04258_);
  and (_04263_, _04262_, _04113_);
  or (_04264_, _04263_, _04109_);
  nor (_04265_, _04264_, _04255_);
  and (_04266_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_04267_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_04268_, _04267_, _04266_);
  and (_04269_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_04270_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_04271_, _04270_, _04269_);
  and (_04272_, _04271_, _04268_);
  and (_04273_, _04272_, _04125_);
  and (_04274_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_04275_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_04276_, _04275_, _04274_);
  and (_04277_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_04278_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_04279_, _04278_, _04277_);
  and (_04280_, _04279_, _04276_);
  and (_04281_, _04280_, _04113_);
  or (_04282_, _04281_, _04172_);
  nor (_04283_, _04282_, _04273_);
  nor (_04284_, _04283_, _04265_);
  nor (_04285_, _04284_, _04163_);
  nand (_04286_, _04285_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_04287_, _04285_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04288_, _04287_, _04286_);
  and (_04289_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_04290_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_04291_, _04290_, _04289_);
  and (_04292_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_04293_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_04294_, _04293_, _04292_);
  and (_04295_, _04294_, _04291_);
  and (_04296_, _04295_, _04125_);
  and (_04297_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_04298_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_04299_, _04298_, _04297_);
  and (_04300_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_04301_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_04302_, _04301_, _04300_);
  and (_04303_, _04302_, _04299_);
  and (_04304_, _04303_, _04113_);
  nor (_04305_, _04304_, _04296_);
  nor (_04306_, _04305_, _04172_);
  and (_04307_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_04308_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_04309_, _04308_, _04307_);
  and (_04310_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_04311_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_04312_, _04311_, _04310_);
  and (_04313_, _04312_, _04309_);
  and (_04314_, _04313_, _04125_);
  and (_04315_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_04316_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_04317_, _04316_, _04315_);
  and (_04318_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_04319_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_04320_, _04319_, _04318_);
  and (_04321_, _04320_, _04317_);
  and (_04322_, _04321_, _04113_);
  nor (_04323_, _04322_, _04314_);
  nor (_04324_, _04323_, _04109_);
  nor (_04325_, _04324_, _04306_);
  not (_04326_, _04325_);
  nor (_04327_, _04326_, _04163_);
  nor (_04328_, _04327_, _02251_);
  and (_04329_, _04327_, _02251_);
  or (_04330_, _04329_, _04328_);
  or (_04331_, _04330_, _04288_);
  or (_04332_, _04331_, _04247_);
  and (_04333_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_04334_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_04335_, _04334_, _04333_);
  and (_04336_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  and (_04337_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_04338_, _04337_, _04336_);
  and (_04339_, _04338_, _04335_);
  and (_04340_, _04339_, _04125_);
  and (_04341_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_04342_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_04343_, _04342_, _04341_);
  and (_04344_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_04345_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_04346_, _04345_, _04344_);
  and (_04347_, _04346_, _04343_);
  and (_04348_, _04347_, _04113_);
  or (_04349_, _04348_, _04109_);
  nor (_04350_, _04349_, _04340_);
  and (_04351_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_04352_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_04353_, _04352_, _04351_);
  and (_04354_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_04355_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_04356_, _04355_, _04354_);
  and (_04357_, _04356_, _04353_);
  and (_04358_, _04357_, _04125_);
  and (_04359_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_04360_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_04361_, _04360_, _04359_);
  and (_04362_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_04363_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_04364_, _04363_, _04362_);
  and (_04365_, _04364_, _04361_);
  and (_04366_, _04365_, _04113_);
  or (_04367_, _04366_, _04172_);
  nor (_04368_, _04367_, _04358_);
  nor (_04369_, _04368_, _04350_);
  nor (_04370_, _04369_, _04163_);
  and (_04371_, _04370_, _03227_);
  nor (_04372_, _04370_, _03227_);
  or (_04373_, _04372_, _04371_);
  and (_04374_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_04375_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_04376_, _04375_, _04374_);
  and (_04377_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_04378_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_04379_, _04378_, _04377_);
  and (_04380_, _04379_, _04376_);
  and (_04381_, _04380_, _04125_);
  and (_04382_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_04383_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_04384_, _04383_, _04382_);
  and (_04385_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_04386_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_04387_, _04386_, _04385_);
  and (_04388_, _04387_, _04384_);
  and (_04389_, _04388_, _04113_);
  or (_04390_, _04389_, _04172_);
  nor (_04391_, _04390_, _04381_);
  and (_04392_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_04393_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_04394_, _04393_, _04392_);
  and (_04395_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_04396_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_04397_, _04396_, _04395_);
  and (_04398_, _04397_, _04394_);
  nor (_04399_, _04398_, _04113_);
  and (_04400_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_04401_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_04402_, _04401_, _04400_);
  and (_04403_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_04404_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_04405_, _04404_, _04403_);
  and (_04406_, _04405_, _04402_);
  nor (_04407_, _04406_, _04125_);
  or (_04408_, _04407_, _04399_);
  and (_04409_, _04408_, _04172_);
  nor (_04410_, _04409_, _04391_);
  nor (_04411_, _04410_, _04163_);
  and (_04412_, _04411_, _02015_);
  nor (_04413_, _04411_, _02015_);
  or (_04414_, _04413_, _04412_);
  or (_04415_, _04414_, _04373_);
  and (_04416_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_04417_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_04418_, _04417_, _04416_);
  and (_04419_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_04420_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_04421_, _04420_, _04419_);
  and (_04422_, _04421_, _04418_);
  and (_04423_, _04422_, _04125_);
  and (_04424_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_04425_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_04426_, _04425_, _04424_);
  and (_04427_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_04428_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_04429_, _04428_, _04427_);
  and (_04430_, _04429_, _04426_);
  and (_04431_, _04430_, _04113_);
  or (_04432_, _04431_, _04109_);
  nor (_04433_, _04432_, _04423_);
  and (_04434_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_04435_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor (_04436_, _04435_, _04434_);
  and (_04437_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_04438_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_04439_, _04438_, _04437_);
  and (_04440_, _04439_, _04436_);
  and (_04441_, _04440_, _04125_);
  and (_04442_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_04443_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_04444_, _04443_, _04442_);
  and (_04445_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_04446_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_04447_, _04446_, _04445_);
  and (_04448_, _04447_, _04444_);
  and (_04449_, _04448_, _04113_);
  or (_04450_, _04449_, _04172_);
  nor (_04451_, _04450_, _04441_);
  nor (_04452_, _04451_, _04433_);
  nor (_04453_, _04452_, _04163_);
  and (_04454_, _04453_, _03223_);
  nor (_04455_, _04453_, _03223_);
  or (_04456_, _04455_, _04454_);
  and (_04457_, _03890_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_04458_, _03885_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_04459_, _04458_, _04457_);
  and (_04460_, _03888_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_04461_, _03883_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_04462_, _04461_, _04460_);
  and (_04463_, _04462_, _04459_);
  and (_04464_, _04463_, _04125_);
  and (_04465_, _03885_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_04466_, _03888_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_04467_, _04466_, _04465_);
  and (_04468_, _03890_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_04469_, _03883_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_04470_, _04469_, _04468_);
  and (_04471_, _04470_, _04467_);
  and (_04472_, _04471_, _04113_);
  or (_04473_, _04472_, _04109_);
  nor (_04474_, _04473_, _04464_);
  and (_04475_, _03890_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_04476_, _03885_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_04477_, _04476_, _04475_);
  and (_04478_, _03888_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_04479_, _03883_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_04480_, _04479_, _04478_);
  and (_04481_, _04480_, _04477_);
  and (_04482_, _04481_, _04125_);
  and (_04483_, _03885_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_04484_, _03883_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_04485_, _04484_, _04483_);
  and (_04486_, _03890_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_04487_, _03888_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_04488_, _04487_, _04486_);
  and (_04489_, _04488_, _04485_);
  and (_04490_, _04489_, _04113_);
  or (_04491_, _04490_, _04172_);
  nor (_04492_, _04491_, _04482_);
  nor (_04493_, _04492_, _04474_);
  nor (_04494_, _04493_, _04163_);
  nor (_04495_, _04494_, _03238_);
  and (_04496_, _04494_, _03238_);
  or (_04497_, _04496_, _04495_);
  or (_04498_, _04497_, _04456_);
  or (_04499_, _04498_, _04415_);
  or (_04500_, _04499_, _04332_);
  or (_04501_, _04500_, _04104_);
  nor (_04502_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_04503_, _04502_, _02251_);
  not (_04504_, _04503_);
  and (_04505_, _04502_, _02251_);
  nor (_04506_, _04505_, _04504_);
  nor (_04507_, _04503_, _03242_);
  and (_04508_, _04503_, _03242_);
  nor (_04509_, _04508_, _04507_);
  and (_04510_, _04509_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_04511_, _03242_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_04512_, _04511_, _04510_);
  and (_04513_, _04512_, _04506_);
  not (_04514_, _04506_);
  nor (_04515_, _04509_, _04142_);
  and (_04516_, _04509_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_04517_, _04516_, _04515_);
  and (_04518_, _04517_, _04514_);
  or (_04519_, _04518_, _04513_);
  and (_04520_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04521_, _04520_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_04522_, _04521_);
  and (_04523_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_04524_, _04523_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04525_, _04524_, _04522_);
  not (_04526_, _04525_);
  nor (_04527_, _04521_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04528_, _04521_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_04529_, _04528_, _04527_);
  nor (_04530_, _04529_, _04137_);
  and (_04531_, _04529_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_04532_, _04531_, _04530_);
  and (_04533_, _04532_, _04526_);
  or (_04534_, _04529_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_04535_, _03242_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_04536_, _04535_, _04525_);
  and (_04537_, _04536_, _04534_);
  or (_04538_, _04537_, _04533_);
  and (_04539_, _04509_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_04540_, _03242_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_04541_, _04540_, _04514_);
  or (_04542_, _04541_, _04539_);
  nand (_04543_, _04509_, _08414_);
  or (_04544_, _04509_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_04545_, _04544_, _04543_);
  or (_04546_, _04545_, _04506_);
  and (_04547_, _04546_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04548_, _04547_, _04542_);
  or (_04549_, _03242_, \oc8051_symbolic_cxrom1.regvalid [15]);
  or (_04550_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_04551_, _04550_, _04549_);
  or (_04552_, _04551_, _02251_);
  or (_04553_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_04554_, _03242_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_04555_, _04554_, _04553_);
  or (_04556_, _04555_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04557_, _04556_, _04552_);
  and (_04558_, _04557_, _04548_);
  and (_04559_, _04558_, _04538_);
  and (_04560_, _04559_, _04519_);
  or (_04561_, _04560_, _02020_);
  or (_04562_, _04529_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_04563_, _03242_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_04564_, _04563_, _04525_);
  and (_04565_, _04564_, _04562_);
  or (_04566_, _04529_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_04567_, _04529_, _09148_);
  and (_04568_, _04567_, _04526_);
  and (_04569_, _04568_, _04566_);
  or (_04570_, _04569_, _04565_);
  or (_04571_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_04572_, _03242_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_04573_, _04572_, _04571_);
  or (_04574_, _04573_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04575_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [13]);
  or (_04576_, _04575_, _04540_);
  or (_04577_, _04576_, _02251_);
  and (_04578_, _04577_, _04574_);
  and (_04579_, _03242_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_04580_, _04509_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_04581_, _04580_, _04579_);
  and (_04582_, _04581_, _04506_);
  nor (_04583_, _04509_, _04137_);
  and (_04584_, _04509_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_04585_, _04584_, _04583_);
  and (_04586_, _04585_, _04514_);
  or (_04587_, _04586_, _04582_);
  and (_04588_, _04587_, _04578_);
  and (_04589_, _04588_, _04570_);
  or (_04590_, _04589_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_04591_, _04557_, _04548_);
  and (_04592_, _04591_, _04590_);
  and (_04593_, _04592_, _04561_);
  or (_04594_, _04593_, _03291_);
  and (_04595_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_04596_, _04511_, _02251_);
  or (_04597_, _04596_, _04595_);
  or (_04598_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_04599_, _03242_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_04600_, _04599_, _04598_);
  or (_04601_, _04600_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04602_, _04601_, _04597_);
  and (_04603_, _04602_, _02020_);
  or (_04604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_04605_, _03242_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_04606_, _04605_, _04520_);
  and (_04607_, _04606_, _04604_);
  and (_04608_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _02251_);
  and (_04609_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_04610_, _04609_, _04579_);
  and (_04611_, _04610_, _04608_);
  or (_04612_, _04611_, _04607_);
  or (_04613_, _04612_, _04603_);
  or (_04614_, _03242_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or (_04615_, _04529_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_04616_, _04615_, _04614_);
  or (_04617_, _04616_, _04526_);
  nand (_04618_, _04529_, _08414_);
  or (_04619_, _04529_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_04620_, _04619_, _04618_);
  or (_04621_, _04620_, _04525_);
  and (_04622_, _04621_, _04617_);
  nor (_04623_, _04509_, _08399_);
  and (_04624_, _04509_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_04625_, _04624_, _04623_);
  or (_04626_, _04625_, _04506_);
  and (_04627_, _04509_, \oc8051_symbolic_cxrom1.regvalid [15]);
  nand (_04628_, _03242_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand (_04629_, _04628_, _04506_);
  or (_04630_, _04629_, _04627_);
  or (_04631_, _04610_, _02251_);
  or (_04632_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_04633_, _03242_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_04634_, _04633_, _04632_);
  or (_04635_, _04634_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04636_, _04635_, _02020_);
  and (_04637_, _04636_, _04631_);
  and (_04638_, _04637_, _04630_);
  and (_04639_, _04638_, _04626_);
  and (_04640_, _04639_, _04622_);
  nor (_04641_, _04529_, _08399_);
  and (_04642_, _04529_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_04643_, _04642_, _04641_);
  or (_04644_, _04643_, _04525_);
  or (_04645_, _04529_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_04646_, _04645_, _04549_);
  or (_04647_, _04646_, _04526_);
  and (_04648_, _04647_, _04644_);
  and (_04649_, _04602_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04650_, _04649_, _04542_);
  and (_04651_, _04650_, _04546_);
  and (_04652_, _04651_, _04648_);
  or (_04653_, _04652_, _04640_);
  and (_04654_, _04653_, _04613_);
  or (_04655_, _04654_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_04656_, _03888_, _06261_);
  nor (_04657_, _04656_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04658_, _04656_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_04659_, _04658_, _04657_);
  or (_04660_, _04659_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nand (_04661_, _03888_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04662_, _04661_, _03929_);
  and (_04663_, _04662_, _04660_);
  or (_04664_, _04659_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_04665_, _03888_, _06261_);
  not (_04666_, _04659_);
  or (_04667_, _04666_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_04668_, _04667_, _04665_);
  and (_04669_, _04668_, _04664_);
  or (_04670_, _04669_, _04663_);
  nand (_04671_, _04659_, _08363_);
  nor (_04672_, _04665_, _04656_);
  and (_04673_, _04672_, _04111_);
  and (_04674_, _04673_, _04671_);
  not (_04675_, _04672_);
  nor (_04676_, _04659_, _04117_);
  and (_04677_, _04659_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_04678_, _04677_, _04676_);
  and (_04679_, _04678_, _04675_);
  or (_04680_, _04679_, _04674_);
  and (_04681_, _04680_, _03885_);
  or (_04682_, _04681_, _04670_);
  or (_04683_, _04659_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_04684_, _04675_, _03906_);
  and (_04685_, _04684_, _04683_);
  and (_04686_, _04659_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_04687_, _04659_, _04142_);
  or (_04688_, _04687_, _04686_);
  and (_04689_, _04688_, _04675_);
  or (_04690_, _04689_, _04685_);
  and (_04691_, _04690_, _03883_);
  or (_04692_, _04666_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_04693_, _04659_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_04694_, _04693_, _04675_);
  and (_04695_, _04694_, _04692_);
  or (_04696_, _04659_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_04697_, _04675_, _03938_);
  and (_04698_, _04697_, _04696_);
  or (_04699_, _04698_, _04695_);
  and (_04700_, _04699_, _03890_);
  or (_04701_, _04700_, _04691_);
  or (_04702_, _04701_, _04682_);
  and (_04703_, _03885_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_04704_, _03890_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  or (_04705_, _04704_, _04703_);
  and (_04706_, _03883_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_04707_, _03888_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  or (_04708_, _04707_, _04706_);
  or (_04709_, _04708_, _04705_);
  nand (_04710_, _03888_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  or (_04711_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nand (_04712_, _04711_, _03885_);
  and (_04713_, _04712_, _04710_);
  nand (_04714_, _03885_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nand (_04715_, _03890_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_04716_, _04715_, _04714_);
  and (_04717_, _04716_, _04713_);
  nand (_04718_, _03883_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  or (_04719_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nand (_04720_, _04719_, _03888_);
  and (_04721_, _04720_, _04718_);
  or (_04722_, \oc8051_symbolic_cxrom1.regarray[3] [3], \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nand (_04723_, _04722_, _03883_);
  or (_04724_, \oc8051_symbolic_cxrom1.regarray[1] [3], \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nand (_04725_, _04724_, _03890_);
  and (_04726_, _04725_, _04723_);
  and (_04727_, _04726_, _04721_);
  and (_04728_, _04727_, _04717_);
  and (_04729_, _04728_, _04709_);
  or (_04730_, _04729_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04731_, _03883_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_04732_, _03888_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  or (_04733_, _04732_, _04731_);
  and (_04734_, _03885_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_04735_, _03890_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  or (_04736_, _04735_, _04734_);
  or (_04737_, _04736_, _04733_);
  nand (_04738_, _03888_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  or (_04739_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nand (_04740_, _04739_, _03885_);
  and (_04741_, _04740_, _04738_);
  nand (_04742_, _03885_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nand (_04743_, _03890_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_04744_, _04743_, _04742_);
  and (_04745_, _04744_, _04741_);
  nand (_04746_, _03883_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  or (_04747_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nand (_04748_, _04747_, _03888_);
  and (_04749_, _04748_, _04746_);
  or (_04750_, \oc8051_symbolic_cxrom1.regarray[11] [3], \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nand (_04751_, _04750_, _03883_);
  or (_04752_, \oc8051_symbolic_cxrom1.regarray[9] [3], \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nand (_04753_, _04752_, _03890_);
  and (_04754_, _04753_, _04751_);
  and (_04755_, _04754_, _04749_);
  and (_04756_, _04755_, _04745_);
  and (_04757_, _04756_, _04737_);
  or (_04758_, _04757_, _06241_);
  and (_04759_, _04758_, _06261_);
  and (_04760_, _04759_, _04730_);
  and (_04761_, _03885_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_04762_, _03890_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  or (_04763_, _04762_, _04761_);
  and (_04764_, _03883_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_04765_, _03888_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  or (_04766_, _04765_, _04764_);
  or (_04767_, _04766_, _04763_);
  nand (_04768_, _03888_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  or (_04769_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nand (_04770_, _04769_, _03885_);
  and (_04771_, _04770_, _04768_);
  nand (_04772_, _03885_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nand (_04773_, _03890_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_04774_, _04773_, _04772_);
  and (_04775_, _04774_, _04771_);
  nand (_04776_, _03883_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  or (_04777_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nand (_04778_, _04777_, _03888_);
  and (_04779_, _04778_, _04776_);
  or (_04780_, \oc8051_symbolic_cxrom1.regarray[7] [3], \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nand (_04781_, _04780_, _03883_);
  or (_04782_, \oc8051_symbolic_cxrom1.regarray[5] [3], \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nand (_04783_, _04782_, _03890_);
  and (_04784_, _04783_, _04781_);
  and (_04785_, _04784_, _04779_);
  and (_04786_, _04785_, _04775_);
  and (_04787_, _04786_, _04767_);
  or (_04788_, _04787_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04789_, _03883_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_04790_, _03888_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  or (_04791_, _04790_, _04789_);
  and (_04792_, _03885_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_04793_, _03890_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  or (_04794_, _04793_, _04792_);
  or (_04795_, _04794_, _04791_);
  nand (_04796_, _03888_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  or (_04797_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nand (_04798_, _04797_, _03885_);
  and (_04799_, _04798_, _04796_);
  nand (_04800_, _03885_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nand (_04801_, _03890_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_04802_, _04801_, _04800_);
  and (_04803_, _04802_, _04799_);
  nand (_04804_, _03883_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  or (_04805_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nand (_04806_, _04805_, _03888_);
  and (_04807_, _04806_, _04804_);
  or (_04808_, \oc8051_symbolic_cxrom1.regarray[15] [3], \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nand (_04809_, _04808_, _03883_);
  or (_04810_, \oc8051_symbolic_cxrom1.regarray[13] [3], \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nand (_04811_, _04810_, _03890_);
  and (_04812_, _04811_, _04809_);
  and (_04813_, _04812_, _04807_);
  and (_04814_, _04813_, _04803_);
  and (_04815_, _04814_, _04795_);
  or (_04816_, _04815_, _06241_);
  and (_04817_, _04816_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04818_, _04817_, _04788_);
  or (_04819_, _04818_, _04760_);
  and (_04820_, _03936_, _03890_);
  and (_04821_, _03940_, _06261_);
  or (_04822_, _06241_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_04823_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_04824_, _04823_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04825_, _04824_, _04822_);
  or (_04826_, _04825_, _04821_);
  and (_04827_, _04826_, _03885_);
  or (_04828_, _04827_, _04820_);
  and (_04829_, _03914_, _03888_);
  and (_04830_, _03919_, _06261_);
  or (_04831_, _06241_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_04832_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_04833_, _04832_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04834_, _04833_, _04831_);
  or (_04835_, _04834_, _04830_);
  and (_04836_, _04835_, _03883_);
  or (_04837_, _04836_, _04829_);
  or (_04838_, _04837_, _04828_);
  nor (_04839_, _00957_, first_instr);
  nand (_04840_, _04839_, _04838_);
  nor (_04841_, _04840_, _03949_);
  nand (_04842_, _04841_, _04819_);
  nor (_04843_, _04842_, _04163_);
  and (_04844_, _04843_, _04702_);
  and (_04845_, _04844_, _04655_);
  and (_04846_, _04845_, _04594_);
  and (property_invalid_ajmp, _04846_, _04501_);
  and (_04847_, _00957_, first_instr);
  or (_00000_, _04847_, rst);
  dff (first_instr, _00000_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _13248_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _13249_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _13250_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _13251_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _13252_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _13253_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _13254_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _13255_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _13246_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _08691_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _08694_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _08697_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _13247_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _08702_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _08705_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _08709_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _13238_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _13239_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _13240_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _13241_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _13242_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _13243_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _13244_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _13245_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _08492_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _08497_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _08499_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _08501_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _08504_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _08508_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _08510_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _08513_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _08374_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _08379_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _08384_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _08388_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _08391_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _08395_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _08400_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _08402_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _08293_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _08297_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _08299_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _08300_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _08301_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _08302_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _08303_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _08307_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _13261_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _13262_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _13263_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _13264_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _13265_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _08227_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _08230_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _08234_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _08129_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _13256_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _13257_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _08141_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _13258_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _13259_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _08148_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _13260_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _08020_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _08023_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _08026_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _08030_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _08035_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _08039_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _08042_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _08045_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _07923_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _07926_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _07930_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _07934_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _07938_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _07941_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _07946_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _07950_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _07827_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _07830_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _07834_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _07839_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _07844_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _07849_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _07852_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _07856_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _07413_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _07416_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _07419_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _07421_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _07423_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _07427_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _07431_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _07434_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _07298_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _07302_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _07307_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _07313_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _07318_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _07324_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _07329_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _07332_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _07608_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _07611_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _07615_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _07618_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _07623_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _07627_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _07630_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _07635_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _07517_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _07520_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _07524_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _07529_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _07534_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _07537_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _07540_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _07543_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _07728_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _07731_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _07734_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _07738_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _07742_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _07745_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _07747_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _07750_);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _05859_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _05887_);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _05931_);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _05981_);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _06031_);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _06085_);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _06158_);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _06239_);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _06315_);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _06394_);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _06484_);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _06577_);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _06683_);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _06785_);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _06896_);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _05809_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _05508_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _05511_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _05514_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _05516_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _05518_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _05521_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _05523_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _05358_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], _12317_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], _11174_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _11150_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], _12621_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], _12736_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], _11754_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _05361_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _11428_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], _11426_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], _11595_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], _11638_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _10883_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _05364_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _09788_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _09822_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _03153_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _09794_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _09820_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _05116_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _09810_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _05182_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _09813_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _09782_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _09513_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _09521_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _09529_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _09806_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _09791_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _03062_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _05222_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _03577_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _05127_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _03857_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _05136_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _03594_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _04891_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _05200_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _06447_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _07107_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _03186_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _10443_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _05219_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _11805_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _11945_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _12372_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _05113_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _00498_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _05311_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _05302_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _08362_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _08582_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _03728_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _03751_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _12673_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _03102_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _01805_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _02847_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _00041_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _06640_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _04854_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _12147_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _00574_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _12445_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _12690_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _02839_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _01824_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _01776_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _02968_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _02983_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _03074_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _01037_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _02869_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _02864_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _10893_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _08283_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _03165_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _07837_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _05251_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _09073_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _04065_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _02877_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _07842_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _04849_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _09492_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _04850_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _08879_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _09831_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _03190_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _01437_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _03387_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _04970_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _04855_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _01669_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _05203_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _04852_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _06909_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _02804_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _01432_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _05235_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _04853_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _01710_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _01517_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _03698_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _01955_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _02792_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _13213_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _04983_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _10214_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _08279_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _01547_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _01164_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _13054_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _02887_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _11042_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _10850_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _12211_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _03612_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _03200_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _02913_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _01158_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _01812_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _02836_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _03865_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _01154_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _02833_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _02906_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _02950_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _02964_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _02378_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _01427_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _02829_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _04851_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _02749_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _12274_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _02816_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _02898_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _09528_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _09192_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _02813_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _02235_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _03249_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _02809_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _02896_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _02946_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _02962_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _03559_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _12295_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _02806_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _12154_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _12267_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _03763_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _03760_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _03756_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _03754_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _12234_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _03789_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _03805_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _03803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _03801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _03798_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _03791_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _12229_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _10908_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _03641_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _03653_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _03647_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _03643_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _12251_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _03677_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _03724_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _03721_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _03719_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _03706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _12239_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _10902_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _11055_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _03211_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _03195_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _03182_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _03180_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _03177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _09996_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _10265_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _01964_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _01962_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _01960_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _01953_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _12303_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _02776_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _02751_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _10297_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _12646_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _10310_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _10301_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _00137_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _00196_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _00177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _00157_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _12338_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _10869_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _10866_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _10919_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _10911_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _10889_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _12343_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _13165_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _13203_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _13196_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _13188_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _03198_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _12702_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _12670_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _11543_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _11522_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _11467_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _11443_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _11435_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _12712_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _11646_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _11624_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _11618_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _11616_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _11610_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _11605_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _12706_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03001_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _10135_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _03204_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _10114_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _12694_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _12679_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _10992_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _12093_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _12750_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _11327_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _11312_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _10174_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _11058_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _11089_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _10221_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], _11801_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], _11792_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _10190_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _11856_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _11848_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _11412_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _11579_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _11630_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _11658_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _11883_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03202_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _02999_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _03067_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _11914_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _11904_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _11406_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _03097_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _11704_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _11476_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _11715_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _11710_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _11464_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _11602_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _11726_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _11720_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _11451_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _11751_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _11736_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _11439_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _11598_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _11641_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _11984_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _11979_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _11370_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _11995_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _11993_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _11357_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11565_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _12006_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _12001_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _11355_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _12040_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _12011_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _11347_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _11620_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _12049_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _12042_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _11343_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _09984_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _10072_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _10067_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _10060_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _11247_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _12300_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _12280_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _11236_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _10047_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _02340_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _11844_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _11292_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _12580_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _00307_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _00670_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _02424_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _05133_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _03712_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _06111_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _05975_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _03708_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _03746_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _03765_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _02393_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _01644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _01147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _01317_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _06465_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _08881_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _01115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _01110_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _01112_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _04014_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _00209_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _00205_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _02637_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _00144_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _00130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _02655_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _00168_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _03916_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _05691_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _05706_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _05712_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _05709_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _05697_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _05695_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _02380_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _03221_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _13064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _12951_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _02954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _03036_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _05575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _05566_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _02512_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _04848_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _10675_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _01846_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _01851_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _01849_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _01796_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _01817_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _01856_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _01853_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _10459_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _01859_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _09163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _10162_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _01943_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _01931_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _10318_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _01599_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _01808_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _09318_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _01597_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _01593_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _10816_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _08683_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _08562_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _10480_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _01803_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _02022_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _02016_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _08584_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _02036_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _01580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _02049_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _02042_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _01570_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _01801_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _02054_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _10217_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _02062_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _01563_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _02082_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _02072_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _01559_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _01799_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _02091_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _10339_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _02688_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _02673_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _02670_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _02575_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _02545_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _02720_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _02577_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _06167_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _02693_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _02691_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _02726_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _02573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _02724_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _02697_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _02543_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _06247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _02664_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _02662_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _02627_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _02625_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _02552_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _02728_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _02588_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _06472_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _02590_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _02712_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _02555_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _02710_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _02592_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _02558_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _02708_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _06467_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _09036_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _02548_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _11350_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _11718_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _05539_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _05505_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _03471_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _02798_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _12496_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _12482_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _12493_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _12491_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _12489_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _12485_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _02763_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _12819_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _00150_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _00140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _12017_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _12014_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _12032_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _12038_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _12035_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _12082_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _12077_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _00133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _12156_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _12151_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _12128_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _12130_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _12135_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _12137_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _12119_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _00121_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _00126_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _00124_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _12163_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _12173_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _12169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _12172_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _12184_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _12178_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _12181_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _00115_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _11910_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _11907_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _11897_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _11900_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _11888_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _11891_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _11877_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _00116_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _00170_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _11930_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _11924_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _11927_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _11830_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _11825_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _11729_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _11723_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _00165_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _01494_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _01415_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _01412_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _01406_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _12255_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _01586_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _10547_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _10566_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _10557_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _10553_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _10549_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _01397_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _10478_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _10473_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _10471_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _03726_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _10499_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _10514_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _10507_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _01066_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _01031_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _10374_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _03779_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _10434_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _10427_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _10424_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _10419_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _10416_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _01044_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _10344_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _10337_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _03822_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _01884_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _10257_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _10250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _10247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _01040_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _01023_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _10146_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _10143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _03861_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _10208_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _10202_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _10199_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _10193_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _01020_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _02936_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _02208_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _10761_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _08118_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _05143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _12141_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _02925_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _02520_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _02503_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _02452_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _10531_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _02486_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _02941_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _02988_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _02787_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _02782_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _02740_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _02771_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _00865_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _02756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _01051_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _06914_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _01508_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _02560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _06954_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _01583_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _01557_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _01791_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _01785_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _01829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _01794_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _02550_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _02483_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _02481_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _02198_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _02159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _02239_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _02224_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _02408_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _02137_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _06884_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _06945_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _02454_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _02438_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _06881_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _02668_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _02461_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _06942_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _06975_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _02768_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _01924_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _02883_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _02860_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _06874_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _06939_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _02923_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _02911_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _02934_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _01920_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _11698_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _06933_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _13158_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _13002_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _13205_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _13168_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _06927_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _01903_);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [1], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [4], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [5], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], \oc8051_top_1.oc8051_memory_interface1.op3_buff [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], \oc8051_top_1.oc8051_memory_interface1.op3_buff [2]);
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [0], ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [1], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [2], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [3], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [4], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [5], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [6], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [7], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [8], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [9], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [10], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [11], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [12], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [13], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [14], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [15], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT [16], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [0], ABINPUT000[1]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [1], ABINPUT000[2]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [2], ABINPUT000[3]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [3], ABINPUT000[4]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [4], ABINPUT000[5]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [5], ABINPUT000[6]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [6], ABINPUT000[7]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc1 [7], ABINPUT000[8]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [0], ABINPUT000[9]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [1], ABINPUT000[10]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [2], ABINPUT000[11]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [3], ABINPUT000[12]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [4], ABINPUT000[13]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [5], ABINPUT000[14]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [6], ABINPUT000[15]);
  buf(\oc8051_top_1.oc8051_alu1.mulsrc2 [7], ABINPUT000[16]);
  buf(\oc8051_top_1.oc8051_alu1.mulOv , ABINPUT000[0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [0], ABINPUT000000[1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [1], ABINPUT000000[2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [2], ABINPUT000000[3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [3], ABINPUT000000[4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [4], ABINPUT000000[5]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [5], ABINPUT000000[6]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [6], ABINPUT000000[7]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc1 [7], ABINPUT000000[8]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [0], ABINPUT000000[9]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [1], ABINPUT000000[10]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], ABINPUT000000[11]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], ABINPUT000000[12]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], ABINPUT000000[13]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], ABINPUT000000[14]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], ABINPUT000000[15]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], ABINPUT000000[16]);
  buf(\oc8051_top_1.oc8051_alu1.divOv , ABINPUT000000[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [0], ABINPUT000000[0]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [1], ABINPUT000000[1]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [2], ABINPUT000000[2]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [3], ABINPUT000000[3]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [4], ABINPUT000000[4]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [5], ABINPUT000000[5]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [6], ABINPUT000000[6]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [7], ABINPUT000000[7]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [8], ABINPUT000000[8]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [9], ABINPUT000000[9]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [10], ABINPUT000000[10]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [11], ABINPUT000000[11]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [12], ABINPUT000000[12]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [13], ABINPUT000000[13]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [14], ABINPUT000000[14]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [15], ABINPUT000000[15]);
  buf(\oc8051_top_1.oc8051_alu1.ABINPUT000 [16], ABINPUT000000[16]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(\oc8051_top_1.ABINPUT000 [0], ABINPUT000[0]);
  buf(\oc8051_top_1.ABINPUT000 [1], ABINPUT000[1]);
  buf(\oc8051_top_1.ABINPUT000 [2], ABINPUT000[2]);
  buf(\oc8051_top_1.ABINPUT000 [3], ABINPUT000[3]);
  buf(\oc8051_top_1.ABINPUT000 [4], ABINPUT000[4]);
  buf(\oc8051_top_1.ABINPUT000 [5], ABINPUT000[5]);
  buf(\oc8051_top_1.ABINPUT000 [6], ABINPUT000[6]);
  buf(\oc8051_top_1.ABINPUT000 [7], ABINPUT000[7]);
  buf(\oc8051_top_1.ABINPUT000 [8], ABINPUT000[8]);
  buf(\oc8051_top_1.ABINPUT000 [9], ABINPUT000[9]);
  buf(\oc8051_top_1.ABINPUT000 [10], ABINPUT000[10]);
  buf(\oc8051_top_1.ABINPUT000 [11], ABINPUT000[11]);
  buf(\oc8051_top_1.ABINPUT000 [12], ABINPUT000[12]);
  buf(\oc8051_top_1.ABINPUT000 [13], ABINPUT000[13]);
  buf(\oc8051_top_1.ABINPUT000 [14], ABINPUT000[14]);
  buf(\oc8051_top_1.ABINPUT000 [15], ABINPUT000[15]);
  buf(\oc8051_top_1.ABINPUT000 [16], ABINPUT000[16]);
  buf(\oc8051_top_1.ABINPUT000000 [0], ABINPUT000000[0]);
  buf(\oc8051_top_1.ABINPUT000000 [1], ABINPUT000000[1]);
  buf(\oc8051_top_1.ABINPUT000000 [2], ABINPUT000000[2]);
  buf(\oc8051_top_1.ABINPUT000000 [3], ABINPUT000000[3]);
  buf(\oc8051_top_1.ABINPUT000000 [4], ABINPUT000000[4]);
  buf(\oc8051_top_1.ABINPUT000000 [5], ABINPUT000000[5]);
  buf(\oc8051_top_1.ABINPUT000000 [6], ABINPUT000000[6]);
  buf(\oc8051_top_1.ABINPUT000000 [7], ABINPUT000000[7]);
  buf(\oc8051_top_1.ABINPUT000000 [8], ABINPUT000000[8]);
  buf(\oc8051_top_1.ABINPUT000000 [9], ABINPUT000000[9]);
  buf(\oc8051_top_1.ABINPUT000000 [10], ABINPUT000000[10]);
  buf(\oc8051_top_1.ABINPUT000000 [11], ABINPUT000000[11]);
  buf(\oc8051_top_1.ABINPUT000000 [12], ABINPUT000000[12]);
  buf(\oc8051_top_1.ABINPUT000000 [13], ABINPUT000000[13]);
  buf(\oc8051_top_1.ABINPUT000000 [14], ABINPUT000000[14]);
  buf(\oc8051_top_1.ABINPUT000000 [15], ABINPUT000000[15]);
  buf(\oc8051_top_1.ABINPUT000000 [16], ABINPUT000000[16]);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(cy, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
