
module oc8051_fv_top(clk, rst, word_in, p0_in, p1_in, p2_in, p3_in, rxd_i, t0_i, t1_i, t2_i, t2ex_i, property_invalid, ABINPUT);
  wire _00000_;
  wire _00001_;
  wire _00002_;
  wire _00003_;
  wire _00004_;
  wire _00005_;
  wire _00006_;
  wire _00007_;
  wire _00008_;
  wire _00009_;
  wire _00010_;
  wire _00011_;
  wire _00012_;
  wire _00013_;
  wire _00014_;
  wire _00015_;
  wire _00016_;
  wire _00017_;
  wire _00018_;
  wire _00019_;
  wire _00020_;
  wire _00021_;
  wire _00022_;
  wire _00023_;
  wire _00024_;
  wire _00025_;
  wire _00026_;
  wire _00027_;
  wire _00028_;
  wire _00029_;
  wire _00030_;
  wire _00031_;
  wire _00032_;
  wire _00033_;
  wire _00034_;
  wire _00035_;
  wire _00036_;
  wire _00037_;
  wire _00038_;
  wire _00039_;
  wire _00040_;
  wire _00041_;
  wire _00042_;
  wire _00043_;
  wire _00044_;
  wire _00045_;
  wire _00046_;
  wire _00047_;
  wire _00048_;
  wire _00049_;
  wire _00050_;
  wire _00051_;
  wire _00052_;
  wire _00053_;
  wire _00054_;
  wire _00055_;
  wire _00056_;
  wire _00057_;
  wire _00058_;
  wire _00059_;
  wire _00060_;
  wire _00061_;
  wire _00062_;
  wire _00063_;
  wire _00064_;
  wire _00065_;
  wire _00066_;
  wire _00067_;
  wire _00068_;
  wire _00069_;
  wire _00070_;
  wire _00071_;
  wire _00072_;
  wire _00073_;
  wire _00074_;
  wire _00075_;
  wire _00076_;
  wire _00077_;
  wire _00078_;
  wire _00079_;
  wire _00080_;
  wire _00081_;
  wire _00082_;
  wire _00083_;
  wire _00084_;
  wire _00085_;
  wire _00086_;
  wire _00087_;
  wire _00088_;
  wire _00089_;
  wire _00090_;
  wire _00091_;
  wire _00092_;
  wire _00093_;
  wire _00094_;
  wire _00095_;
  wire _00096_;
  wire _00097_;
  wire _00098_;
  wire _00099_;
  wire _00100_;
  wire _00101_;
  wire _00102_;
  wire _00103_;
  wire _00104_;
  wire _00105_;
  wire _00106_;
  wire _00107_;
  wire _00108_;
  wire _00109_;
  wire _00110_;
  wire _00111_;
  wire _00112_;
  wire _00113_;
  wire _00114_;
  wire _00115_;
  wire _00116_;
  wire _00117_;
  wire _00118_;
  wire _00119_;
  wire _00120_;
  wire _00121_;
  wire _00122_;
  wire _00123_;
  wire _00124_;
  wire _00125_;
  wire _00126_;
  wire _00127_;
  wire _00128_;
  wire _00129_;
  wire _00130_;
  wire _00131_;
  wire _00132_;
  wire _00133_;
  wire _00134_;
  wire _00135_;
  wire _00136_;
  wire _00137_;
  wire _00138_;
  wire _00139_;
  wire _00140_;
  wire _00141_;
  wire _00142_;
  wire _00143_;
  wire _00144_;
  wire _00145_;
  wire _00146_;
  wire _00147_;
  wire _00148_;
  wire _00149_;
  wire _00150_;
  wire _00151_;
  wire _00152_;
  wire _00153_;
  wire _00154_;
  wire _00155_;
  wire _00156_;
  wire _00157_;
  wire _00158_;
  wire _00159_;
  wire _00160_;
  wire _00161_;
  wire _00162_;
  wire _00163_;
  wire _00164_;
  wire _00165_;
  wire _00166_;
  wire _00167_;
  wire _00168_;
  wire _00169_;
  wire _00170_;
  wire _00171_;
  wire _00172_;
  wire _00173_;
  wire _00174_;
  wire _00175_;
  wire _00176_;
  wire _00177_;
  wire _00178_;
  wire _00179_;
  wire _00180_;
  wire _00181_;
  wire _00182_;
  wire _00183_;
  wire _00184_;
  wire _00185_;
  wire _00186_;
  wire _00187_;
  wire _00188_;
  wire _00189_;
  wire _00190_;
  wire _00191_;
  wire _00192_;
  wire _00193_;
  wire _00194_;
  wire _00195_;
  wire _00196_;
  wire _00197_;
  wire _00198_;
  wire _00199_;
  wire _00200_;
  wire _00201_;
  wire _00202_;
  wire _00203_;
  wire _00204_;
  wire _00205_;
  wire _00206_;
  wire _00207_;
  wire _00208_;
  wire _00209_;
  wire _00210_;
  wire _00211_;
  wire _00212_;
  wire _00213_;
  wire _00214_;
  wire _00215_;
  wire _00216_;
  wire _00217_;
  wire _00218_;
  wire _00219_;
  wire _00220_;
  wire _00221_;
  wire _00222_;
  wire _00223_;
  wire _00224_;
  wire _00225_;
  wire _00226_;
  wire _00227_;
  wire _00228_;
  wire _00229_;
  wire _00230_;
  wire _00231_;
  wire _00232_;
  wire _00233_;
  wire _00234_;
  wire _00235_;
  wire _00236_;
  wire _00237_;
  wire _00238_;
  wire _00239_;
  wire _00240_;
  wire _00241_;
  wire _00242_;
  wire _00243_;
  wire _00244_;
  wire _00245_;
  wire _00246_;
  wire _00247_;
  wire _00248_;
  wire _00249_;
  wire _00250_;
  wire _00251_;
  wire _00252_;
  wire _00253_;
  wire _00254_;
  wire _00255_;
  wire _00256_;
  wire _00257_;
  wire _00258_;
  wire _00259_;
  wire _00260_;
  wire _00261_;
  wire _00262_;
  wire _00263_;
  wire _00264_;
  wire _00265_;
  wire _00266_;
  wire _00267_;
  wire _00268_;
  wire _00269_;
  wire _00270_;
  wire _00271_;
  wire _00272_;
  wire _00273_;
  wire _00274_;
  wire _00275_;
  wire _00276_;
  wire _00277_;
  wire _00278_;
  wire _00279_;
  wire _00280_;
  wire _00281_;
  wire _00282_;
  wire _00283_;
  wire _00284_;
  wire _00285_;
  wire _00286_;
  wire _00287_;
  wire _00288_;
  wire _00289_;
  wire _00290_;
  wire _00291_;
  wire _00292_;
  wire _00293_;
  wire _00294_;
  wire _00295_;
  wire _00296_;
  wire _00297_;
  wire _00298_;
  wire _00299_;
  wire _00300_;
  wire _00301_;
  wire _00302_;
  wire _00303_;
  wire _00304_;
  wire _00305_;
  wire _00306_;
  wire _00307_;
  wire _00308_;
  wire _00309_;
  wire _00310_;
  wire _00311_;
  wire _00312_;
  wire _00313_;
  wire _00314_;
  wire _00315_;
  wire _00316_;
  wire _00317_;
  wire _00318_;
  wire _00319_;
  wire _00320_;
  wire _00321_;
  wire _00322_;
  wire _00323_;
  wire _00324_;
  wire _00325_;
  wire _00326_;
  wire _00327_;
  wire _00328_;
  wire _00329_;
  wire _00330_;
  wire _00331_;
  wire _00332_;
  wire _00333_;
  wire _00334_;
  wire _00335_;
  wire _00336_;
  wire _00337_;
  wire _00338_;
  wire _00339_;
  wire _00340_;
  wire _00341_;
  wire _00342_;
  wire _00343_;
  wire _00344_;
  wire _00345_;
  wire _00346_;
  wire _00347_;
  wire _00348_;
  wire _00349_;
  wire _00350_;
  wire _00351_;
  wire _00352_;
  wire _00353_;
  wire _00354_;
  wire _00355_;
  wire _00356_;
  wire _00357_;
  wire _00358_;
  wire _00359_;
  wire _00360_;
  wire _00361_;
  wire _00362_;
  wire _00363_;
  wire _00364_;
  wire _00365_;
  wire _00366_;
  wire _00367_;
  wire _00368_;
  wire _00369_;
  wire _00370_;
  wire _00371_;
  wire _00372_;
  wire _00373_;
  wire _00374_;
  wire _00375_;
  wire _00376_;
  wire _00377_;
  wire _00378_;
  wire _00379_;
  wire _00380_;
  wire _00381_;
  wire _00382_;
  wire _00383_;
  wire _00384_;
  wire _00385_;
  wire _00386_;
  wire _00387_;
  wire _00388_;
  wire _00389_;
  wire _00390_;
  wire _00391_;
  wire _00392_;
  wire _00393_;
  wire _00394_;
  wire _00395_;
  wire _00396_;
  wire _00397_;
  wire _00398_;
  wire _00399_;
  wire _00400_;
  wire _00401_;
  wire _00402_;
  wire _00403_;
  wire _00404_;
  wire _00405_;
  wire _00406_;
  wire _00407_;
  wire _00408_;
  wire _00409_;
  wire _00410_;
  wire _00411_;
  wire _00412_;
  wire _00413_;
  wire _00414_;
  wire _00415_;
  wire _00416_;
  wire _00417_;
  wire _00418_;
  wire _00419_;
  wire _00420_;
  wire _00421_;
  wire _00422_;
  wire _00423_;
  wire _00424_;
  wire _00425_;
  wire _00426_;
  wire _00427_;
  wire _00428_;
  wire _00429_;
  wire _00430_;
  wire _00431_;
  wire _00432_;
  wire _00433_;
  wire _00434_;
  wire _00435_;
  wire _00436_;
  wire _00437_;
  wire _00438_;
  wire _00439_;
  wire _00440_;
  wire _00441_;
  wire _00442_;
  wire _00443_;
  wire _00444_;
  wire _00445_;
  wire _00446_;
  wire _00447_;
  wire _00448_;
  wire _00449_;
  wire _00450_;
  wire _00451_;
  wire _00452_;
  wire _00453_;
  wire _00454_;
  wire _00455_;
  wire _00456_;
  wire _00457_;
  wire _00458_;
  wire _00459_;
  wire _00460_;
  wire _00461_;
  wire _00462_;
  wire _00463_;
  wire _00464_;
  wire _00465_;
  wire _00466_;
  wire _00467_;
  wire _00468_;
  wire _00469_;
  wire _00470_;
  wire _00471_;
  wire _00472_;
  wire _00473_;
  wire _00474_;
  wire _00475_;
  wire _00476_;
  wire _00477_;
  wire _00478_;
  wire _00479_;
  wire _00480_;
  wire _00481_;
  wire _00482_;
  wire _00483_;
  wire _00484_;
  wire _00485_;
  wire _00486_;
  wire _00487_;
  wire _00488_;
  wire _00489_;
  wire _00490_;
  wire _00491_;
  wire _00492_;
  wire _00493_;
  wire _00494_;
  wire _00495_;
  wire _00496_;
  wire _00497_;
  wire _00498_;
  wire _00499_;
  wire _00500_;
  wire _00501_;
  wire _00502_;
  wire _00503_;
  wire _00504_;
  wire _00505_;
  wire _00506_;
  wire _00507_;
  wire _00508_;
  wire _00509_;
  wire _00510_;
  wire _00511_;
  wire _00512_;
  wire _00513_;
  wire _00514_;
  wire _00515_;
  wire _00516_;
  wire _00517_;
  wire _00518_;
  wire _00519_;
  wire _00520_;
  wire _00521_;
  wire _00522_;
  wire _00523_;
  wire _00524_;
  wire _00525_;
  wire _00526_;
  wire _00527_;
  wire _00528_;
  wire _00529_;
  wire _00530_;
  wire _00531_;
  wire _00532_;
  wire _00533_;
  wire _00534_;
  wire _00535_;
  wire _00536_;
  wire _00537_;
  wire _00538_;
  wire _00539_;
  wire _00540_;
  wire _00541_;
  wire _00542_;
  wire _00543_;
  wire _00544_;
  wire _00545_;
  wire _00546_;
  wire _00547_;
  wire _00548_;
  wire _00549_;
  wire _00550_;
  wire _00551_;
  wire _00552_;
  wire _00553_;
  wire _00554_;
  wire _00555_;
  wire _00556_;
  wire _00557_;
  wire _00558_;
  wire _00559_;
  wire _00560_;
  wire _00561_;
  wire _00562_;
  wire _00563_;
  wire _00564_;
  wire _00565_;
  wire _00566_;
  wire _00567_;
  wire _00568_;
  wire _00569_;
  wire _00570_;
  wire _00571_;
  wire _00572_;
  wire _00573_;
  wire _00574_;
  wire _00575_;
  wire _00576_;
  wire _00577_;
  wire _00578_;
  wire _00579_;
  wire _00580_;
  wire _00581_;
  wire _00582_;
  wire _00583_;
  wire _00584_;
  wire _00585_;
  wire _00586_;
  wire _00587_;
  wire _00588_;
  wire _00589_;
  wire _00590_;
  wire _00591_;
  wire _00592_;
  wire _00593_;
  wire _00594_;
  wire _00595_;
  wire _00596_;
  wire _00597_;
  wire _00598_;
  wire _00599_;
  wire _00600_;
  wire _00601_;
  wire _00602_;
  wire _00603_;
  wire _00604_;
  wire _00605_;
  wire _00606_;
  wire _00607_;
  wire _00608_;
  wire _00609_;
  wire _00610_;
  wire _00611_;
  wire _00612_;
  wire _00613_;
  wire _00614_;
  wire _00615_;
  wire _00616_;
  wire _00617_;
  wire _00618_;
  wire _00619_;
  wire _00620_;
  wire _00621_;
  wire _00622_;
  wire _00623_;
  wire _00624_;
  wire _00625_;
  wire _00626_;
  wire _00627_;
  wire _00628_;
  wire _00629_;
  wire _00630_;
  wire _00631_;
  wire _00632_;
  wire _00633_;
  wire _00634_;
  wire _00635_;
  wire _00636_;
  wire _00637_;
  wire _00638_;
  wire _00639_;
  wire _00640_;
  wire _00641_;
  wire _00642_;
  wire _00643_;
  wire _00644_;
  wire _00645_;
  wire _00646_;
  wire _00647_;
  wire _00648_;
  wire _00649_;
  wire _00650_;
  wire _00651_;
  wire _00652_;
  wire _00653_;
  wire _00654_;
  wire _00655_;
  wire _00656_;
  wire _00657_;
  wire _00658_;
  wire _00659_;
  wire _00660_;
  wire _00661_;
  wire _00662_;
  wire _00663_;
  wire _00664_;
  wire _00665_;
  wire _00666_;
  wire _00667_;
  wire _00668_;
  wire _00669_;
  wire _00670_;
  wire _00671_;
  wire _00672_;
  wire _00673_;
  wire _00674_;
  wire _00675_;
  wire _00676_;
  wire _00677_;
  wire _00678_;
  wire _00679_;
  wire _00680_;
  wire _00681_;
  wire _00682_;
  wire _00683_;
  wire _00684_;
  wire _00685_;
  wire _00686_;
  wire _00687_;
  wire _00688_;
  wire _00689_;
  wire _00690_;
  wire _00691_;
  wire _00692_;
  wire _00693_;
  wire _00694_;
  wire _00695_;
  wire _00696_;
  wire _00697_;
  wire _00698_;
  wire _00699_;
  wire _00700_;
  wire _00701_;
  wire _00702_;
  wire _00703_;
  wire _00704_;
  wire _00705_;
  wire _00706_;
  wire _00707_;
  wire _00708_;
  wire _00709_;
  wire _00710_;
  wire _00711_;
  wire _00712_;
  wire _00713_;
  wire _00714_;
  wire _00715_;
  wire _00716_;
  wire _00717_;
  wire _00718_;
  wire _00719_;
  wire _00720_;
  wire _00721_;
  wire _00722_;
  wire _00723_;
  wire _00724_;
  wire _00725_;
  wire _00726_;
  wire _00727_;
  wire _00728_;
  wire _00729_;
  wire _00730_;
  wire _00731_;
  wire _00732_;
  wire _00733_;
  wire _00734_;
  wire _00735_;
  wire _00736_;
  wire _00737_;
  wire _00738_;
  wire _00739_;
  wire _00740_;
  wire _00741_;
  wire _00742_;
  wire _00743_;
  wire _00744_;
  wire _00745_;
  wire _00746_;
  wire _00747_;
  wire _00748_;
  wire _00749_;
  wire _00750_;
  wire _00751_;
  wire _00752_;
  wire _00753_;
  wire _00754_;
  wire _00755_;
  wire _00756_;
  wire _00757_;
  wire _00758_;
  wire _00759_;
  wire _00760_;
  wire _00761_;
  wire _00762_;
  wire _00763_;
  wire _00764_;
  wire _00765_;
  wire _00766_;
  wire _00767_;
  wire _00768_;
  wire _00769_;
  wire _00770_;
  wire _00771_;
  wire _00772_;
  wire _00773_;
  wire _00774_;
  wire _00775_;
  wire _00776_;
  wire _00777_;
  wire _00778_;
  wire _00779_;
  wire _00780_;
  wire _00781_;
  wire _00782_;
  wire _00783_;
  wire _00784_;
  wire _00785_;
  wire _00786_;
  wire _00787_;
  wire _00788_;
  wire _00789_;
  wire _00790_;
  wire _00791_;
  wire _00792_;
  wire _00793_;
  wire _00794_;
  wire _00795_;
  wire _00796_;
  wire _00797_;
  wire _00798_;
  wire _00799_;
  wire _00800_;
  wire _00801_;
  wire _00802_;
  wire _00803_;
  wire _00804_;
  wire _00805_;
  wire _00806_;
  wire _00807_;
  wire _00808_;
  wire _00809_;
  wire _00810_;
  wire _00811_;
  wire _00812_;
  wire _00813_;
  wire _00814_;
  wire _00815_;
  wire _00816_;
  wire _00817_;
  wire _00818_;
  wire _00819_;
  wire _00820_;
  wire _00821_;
  wire _00822_;
  wire _00823_;
  wire _00824_;
  wire _00825_;
  wire _00826_;
  wire _00827_;
  wire _00828_;
  wire _00829_;
  wire _00830_;
  wire _00831_;
  wire _00832_;
  wire _00833_;
  wire _00834_;
  wire _00835_;
  wire _00836_;
  wire _00837_;
  wire _00838_;
  wire _00839_;
  wire _00840_;
  wire _00841_;
  wire _00842_;
  wire _00843_;
  wire _00844_;
  wire _00845_;
  wire _00846_;
  wire _00847_;
  wire _00848_;
  wire _00849_;
  wire _00850_;
  wire _00851_;
  wire _00852_;
  wire _00853_;
  wire _00854_;
  wire _00855_;
  wire _00856_;
  wire _00857_;
  wire _00858_;
  wire _00859_;
  wire _00860_;
  wire _00861_;
  wire _00862_;
  wire _00863_;
  wire _00864_;
  wire _00865_;
  wire _00866_;
  wire _00867_;
  wire _00868_;
  wire _00869_;
  wire _00870_;
  wire _00871_;
  wire _00872_;
  wire _00873_;
  wire _00874_;
  wire _00875_;
  wire _00876_;
  wire _00877_;
  wire _00878_;
  wire _00879_;
  wire _00880_;
  wire _00881_;
  wire _00882_;
  wire _00883_;
  wire _00884_;
  wire _00885_;
  wire _00886_;
  wire _00887_;
  wire _00888_;
  wire _00889_;
  wire _00890_;
  wire _00891_;
  wire _00892_;
  wire _00893_;
  wire _00894_;
  wire _00895_;
  wire _00896_;
  wire _00897_;
  wire _00898_;
  wire _00899_;
  wire _00900_;
  wire _00901_;
  wire _00902_;
  wire _00903_;
  wire _00904_;
  wire _00905_;
  wire _00906_;
  wire _00907_;
  wire _00908_;
  wire _00909_;
  wire _00910_;
  wire _00911_;
  wire _00912_;
  wire _00913_;
  wire _00914_;
  wire _00915_;
  wire _00916_;
  wire _00917_;
  wire _00918_;
  wire _00919_;
  wire _00920_;
  wire _00921_;
  wire _00922_;
  wire _00923_;
  wire _00924_;
  wire _00925_;
  wire _00926_;
  wire _00927_;
  wire _00928_;
  wire _00929_;
  wire _00930_;
  wire _00931_;
  wire _00932_;
  wire _00933_;
  wire _00934_;
  wire _00935_;
  wire _00936_;
  wire _00937_;
  wire _00938_;
  wire _00939_;
  wire _00940_;
  wire _00941_;
  wire _00942_;
  wire _00943_;
  wire _00944_;
  wire _00945_;
  wire _00946_;
  wire _00947_;
  wire _00948_;
  wire _00949_;
  wire _00950_;
  wire _00951_;
  wire _00952_;
  wire _00953_;
  wire _00954_;
  wire _00955_;
  wire _00956_;
  wire _00957_;
  wire _00958_;
  wire _00959_;
  wire _00960_;
  wire _00961_;
  wire _00962_;
  wire _00963_;
  wire _00964_;
  wire _00965_;
  wire _00966_;
  wire _00967_;
  wire _00968_;
  wire _00969_;
  wire _00970_;
  wire _00971_;
  wire _00972_;
  wire _00973_;
  wire _00974_;
  wire _00975_;
  wire _00976_;
  wire _00977_;
  wire _00978_;
  wire _00979_;
  wire _00980_;
  wire _00981_;
  wire _00982_;
  wire _00983_;
  wire _00984_;
  wire _00985_;
  wire _00986_;
  wire _00987_;
  wire _00988_;
  wire _00989_;
  wire _00990_;
  wire _00991_;
  wire _00992_;
  wire _00993_;
  wire _00994_;
  wire _00995_;
  wire _00996_;
  wire _00997_;
  wire _00998_;
  wire _00999_;
  wire _01000_;
  wire _01001_;
  wire _01002_;
  wire _01003_;
  wire _01004_;
  wire _01005_;
  wire _01006_;
  wire _01007_;
  wire _01008_;
  wire _01009_;
  wire _01010_;
  wire _01011_;
  wire _01012_;
  wire _01013_;
  wire _01014_;
  wire _01015_;
  wire _01016_;
  wire _01017_;
  wire _01018_;
  wire _01019_;
  wire _01020_;
  wire _01021_;
  wire _01022_;
  wire _01023_;
  wire _01024_;
  wire _01025_;
  wire _01026_;
  wire _01027_;
  wire _01028_;
  wire _01029_;
  wire _01030_;
  wire _01031_;
  wire _01032_;
  wire _01033_;
  wire _01034_;
  wire _01035_;
  wire _01036_;
  wire _01037_;
  wire _01038_;
  wire _01039_;
  wire _01040_;
  wire _01041_;
  wire _01042_;
  wire _01043_;
  wire _01044_;
  wire _01045_;
  wire _01046_;
  wire _01047_;
  wire _01048_;
  wire _01049_;
  wire _01050_;
  wire _01051_;
  wire _01052_;
  wire _01053_;
  wire _01054_;
  wire _01055_;
  wire _01056_;
  wire _01057_;
  wire _01058_;
  wire _01059_;
  wire _01060_;
  wire _01061_;
  wire _01062_;
  wire _01063_;
  wire _01064_;
  wire _01065_;
  wire _01066_;
  wire _01067_;
  wire _01068_;
  wire _01069_;
  wire _01070_;
  wire _01071_;
  wire _01072_;
  wire _01073_;
  wire _01074_;
  wire _01075_;
  wire _01076_;
  wire _01077_;
  wire _01078_;
  wire _01079_;
  wire _01080_;
  wire _01081_;
  wire _01082_;
  wire _01083_;
  wire _01084_;
  wire _01085_;
  wire _01086_;
  wire _01087_;
  wire _01088_;
  wire _01089_;
  wire _01090_;
  wire _01091_;
  wire _01092_;
  wire _01093_;
  wire _01094_;
  wire _01095_;
  wire _01096_;
  wire _01097_;
  wire _01098_;
  wire _01099_;
  wire _01100_;
  wire _01101_;
  wire _01102_;
  wire _01103_;
  wire _01104_;
  wire _01105_;
  wire _01106_;
  wire _01107_;
  wire _01108_;
  wire _01109_;
  wire _01110_;
  wire _01111_;
  wire _01112_;
  wire _01113_;
  wire _01114_;
  wire _01115_;
  wire _01116_;
  wire _01117_;
  wire _01118_;
  wire _01119_;
  wire _01120_;
  wire _01121_;
  wire _01122_;
  wire _01123_;
  wire _01124_;
  wire _01125_;
  wire _01126_;
  wire _01127_;
  wire _01128_;
  wire _01129_;
  wire _01130_;
  wire _01131_;
  wire _01132_;
  wire _01133_;
  wire _01134_;
  wire _01135_;
  wire _01136_;
  wire _01137_;
  wire _01138_;
  wire _01139_;
  wire _01140_;
  wire _01141_;
  wire _01142_;
  wire _01143_;
  wire _01144_;
  wire _01145_;
  wire _01146_;
  wire _01147_;
  wire _01148_;
  wire _01149_;
  wire _01150_;
  wire _01151_;
  wire _01152_;
  wire _01153_;
  wire _01154_;
  wire _01155_;
  wire _01156_;
  wire _01157_;
  wire _01158_;
  wire _01159_;
  wire _01160_;
  wire _01161_;
  wire _01162_;
  wire _01163_;
  wire _01164_;
  wire _01165_;
  wire _01166_;
  wire _01167_;
  wire _01168_;
  wire _01169_;
  wire _01170_;
  wire _01171_;
  wire _01172_;
  wire _01173_;
  wire _01174_;
  wire _01175_;
  wire _01176_;
  wire _01177_;
  wire _01178_;
  wire _01179_;
  wire _01180_;
  wire _01181_;
  wire _01182_;
  wire _01183_;
  wire _01184_;
  wire _01185_;
  wire _01186_;
  wire _01187_;
  wire _01188_;
  wire _01189_;
  wire _01190_;
  wire _01191_;
  wire _01192_;
  wire _01193_;
  wire _01194_;
  wire _01195_;
  wire _01196_;
  wire _01197_;
  wire _01198_;
  wire _01199_;
  wire _01200_;
  wire _01201_;
  wire _01202_;
  wire _01203_;
  wire _01204_;
  wire _01205_;
  wire _01206_;
  wire _01207_;
  wire _01208_;
  wire _01209_;
  wire _01210_;
  wire _01211_;
  wire _01212_;
  wire _01213_;
  wire _01214_;
  wire _01215_;
  wire _01216_;
  wire _01217_;
  wire _01218_;
  wire _01219_;
  wire _01220_;
  wire _01221_;
  wire _01222_;
  wire _01223_;
  wire _01224_;
  wire _01225_;
  wire _01226_;
  wire _01227_;
  wire _01228_;
  wire _01229_;
  wire _01230_;
  wire _01231_;
  wire _01232_;
  wire _01233_;
  wire _01234_;
  wire _01235_;
  wire _01236_;
  wire _01237_;
  wire _01238_;
  wire _01239_;
  wire _01240_;
  wire _01241_;
  wire _01242_;
  wire _01243_;
  wire _01244_;
  wire _01245_;
  wire _01246_;
  wire _01247_;
  wire _01248_;
  wire _01249_;
  wire _01250_;
  wire _01251_;
  wire _01252_;
  wire _01253_;
  wire _01254_;
  wire _01255_;
  wire _01256_;
  wire _01257_;
  wire _01258_;
  wire _01259_;
  wire _01260_;
  wire _01261_;
  wire _01262_;
  wire _01263_;
  wire _01264_;
  wire _01265_;
  wire _01266_;
  wire _01267_;
  wire _01268_;
  wire _01269_;
  wire _01270_;
  wire _01271_;
  wire _01272_;
  wire _01273_;
  wire _01274_;
  wire _01275_;
  wire _01276_;
  wire _01277_;
  wire _01278_;
  wire _01279_;
  wire _01280_;
  wire _01281_;
  wire _01282_;
  wire _01283_;
  wire _01284_;
  wire _01285_;
  wire _01286_;
  wire _01287_;
  wire _01288_;
  wire _01289_;
  wire _01290_;
  wire _01291_;
  wire _01292_;
  wire _01293_;
  wire _01294_;
  wire _01295_;
  wire _01296_;
  wire _01297_;
  wire _01298_;
  wire _01299_;
  wire _01300_;
  wire _01301_;
  wire _01302_;
  wire _01303_;
  wire _01304_;
  wire _01305_;
  wire _01306_;
  wire _01307_;
  wire _01308_;
  wire _01309_;
  wire _01310_;
  wire _01311_;
  wire _01312_;
  wire _01313_;
  wire _01314_;
  wire _01315_;
  wire _01316_;
  wire _01317_;
  wire _01318_;
  wire _01319_;
  wire _01320_;
  wire _01321_;
  wire _01322_;
  wire _01323_;
  wire _01324_;
  wire _01325_;
  wire _01326_;
  wire _01327_;
  wire _01328_;
  wire _01329_;
  wire _01330_;
  wire _01331_;
  wire _01332_;
  wire _01333_;
  wire _01334_;
  wire _01335_;
  wire _01336_;
  wire _01337_;
  wire _01338_;
  wire _01339_;
  wire _01340_;
  wire _01341_;
  wire _01342_;
  wire _01343_;
  wire _01344_;
  wire _01345_;
  wire _01346_;
  wire _01347_;
  wire _01348_;
  wire _01349_;
  wire _01350_;
  wire _01351_;
  wire _01352_;
  wire _01353_;
  wire _01354_;
  wire _01355_;
  wire _01356_;
  wire _01357_;
  wire _01358_;
  wire _01359_;
  wire _01360_;
  wire _01361_;
  wire _01362_;
  wire _01363_;
  wire _01364_;
  wire _01365_;
  wire _01366_;
  wire _01367_;
  wire _01368_;
  wire _01369_;
  wire _01370_;
  wire _01371_;
  wire _01372_;
  wire _01373_;
  wire _01374_;
  wire _01375_;
  wire _01376_;
  wire _01377_;
  wire _01378_;
  wire _01379_;
  wire _01380_;
  wire _01381_;
  wire _01382_;
  wire _01383_;
  wire _01384_;
  wire _01385_;
  wire _01386_;
  wire _01387_;
  wire _01388_;
  wire _01389_;
  wire _01390_;
  wire _01391_;
  wire _01392_;
  wire _01393_;
  wire _01394_;
  wire _01395_;
  wire _01396_;
  wire _01397_;
  wire _01398_;
  wire _01399_;
  wire _01400_;
  wire _01401_;
  wire _01402_;
  wire _01403_;
  wire _01404_;
  wire _01405_;
  wire _01406_;
  wire _01407_;
  wire _01408_;
  wire _01409_;
  wire _01410_;
  wire _01411_;
  wire _01412_;
  wire _01413_;
  wire _01414_;
  wire _01415_;
  wire _01416_;
  wire _01417_;
  wire _01418_;
  wire _01419_;
  wire _01420_;
  wire _01421_;
  wire _01422_;
  wire _01423_;
  wire _01424_;
  wire _01425_;
  wire _01426_;
  wire _01427_;
  wire _01428_;
  wire _01429_;
  wire _01430_;
  wire _01431_;
  wire _01432_;
  wire _01433_;
  wire _01434_;
  wire _01435_;
  wire _01436_;
  wire _01437_;
  wire _01438_;
  wire _01439_;
  wire _01440_;
  wire _01441_;
  wire _01442_;
  wire _01443_;
  wire _01444_;
  wire _01445_;
  wire _01446_;
  wire _01447_;
  wire _01448_;
  wire _01449_;
  wire _01450_;
  wire _01451_;
  wire _01452_;
  wire _01453_;
  wire _01454_;
  wire _01455_;
  wire _01456_;
  wire _01457_;
  wire _01458_;
  wire _01459_;
  wire _01460_;
  wire _01461_;
  wire _01462_;
  wire _01463_;
  wire _01464_;
  wire _01465_;
  wire _01466_;
  wire _01467_;
  wire _01468_;
  wire _01469_;
  wire _01470_;
  wire _01471_;
  wire _01472_;
  wire _01473_;
  wire _01474_;
  wire _01475_;
  wire _01476_;
  wire _01477_;
  wire _01478_;
  wire _01479_;
  wire _01480_;
  wire _01481_;
  wire _01482_;
  wire _01483_;
  wire _01484_;
  wire _01485_;
  wire _01486_;
  wire _01487_;
  wire _01488_;
  wire _01489_;
  wire _01490_;
  wire _01491_;
  wire _01492_;
  wire _01493_;
  wire _01494_;
  wire _01495_;
  wire _01496_;
  wire _01497_;
  wire _01498_;
  wire _01499_;
  wire _01500_;
  wire _01501_;
  wire _01502_;
  wire _01503_;
  wire _01504_;
  wire _01505_;
  wire _01506_;
  wire _01507_;
  wire _01508_;
  wire _01509_;
  wire _01510_;
  wire _01511_;
  wire _01512_;
  wire _01513_;
  wire _01514_;
  wire _01515_;
  wire _01516_;
  wire _01517_;
  wire _01518_;
  wire _01519_;
  wire _01520_;
  wire _01521_;
  wire _01522_;
  wire _01523_;
  wire _01524_;
  wire _01525_;
  wire _01526_;
  wire _01527_;
  wire _01528_;
  wire _01529_;
  wire _01530_;
  wire _01531_;
  wire _01532_;
  wire _01533_;
  wire _01534_;
  wire _01535_;
  wire _01536_;
  wire _01537_;
  wire _01538_;
  wire _01539_;
  wire _01540_;
  wire _01541_;
  wire _01542_;
  wire _01543_;
  wire _01544_;
  wire _01545_;
  wire _01546_;
  wire _01547_;
  wire _01548_;
  wire _01549_;
  wire _01550_;
  wire _01551_;
  wire _01552_;
  wire _01553_;
  wire _01554_;
  wire _01555_;
  wire _01556_;
  wire _01557_;
  wire _01558_;
  wire _01559_;
  wire _01560_;
  wire _01561_;
  wire _01562_;
  wire _01563_;
  wire _01564_;
  wire _01565_;
  wire _01566_;
  wire _01567_;
  wire _01568_;
  wire _01569_;
  wire _01570_;
  wire _01571_;
  wire _01572_;
  wire _01573_;
  wire _01574_;
  wire _01575_;
  wire _01576_;
  wire _01577_;
  wire _01578_;
  wire _01579_;
  wire _01580_;
  wire _01581_;
  wire _01582_;
  wire _01583_;
  wire _01584_;
  wire _01585_;
  wire _01586_;
  wire _01587_;
  wire _01588_;
  wire _01589_;
  wire _01590_;
  wire _01591_;
  wire _01592_;
  wire _01593_;
  wire _01594_;
  wire _01595_;
  wire _01596_;
  wire _01597_;
  wire _01598_;
  wire _01599_;
  wire _01600_;
  wire _01601_;
  wire _01602_;
  wire _01603_;
  wire _01604_;
  wire _01605_;
  wire _01606_;
  wire _01607_;
  wire _01608_;
  wire _01609_;
  wire _01610_;
  wire _01611_;
  wire _01612_;
  wire _01613_;
  wire _01614_;
  wire _01615_;
  wire _01616_;
  wire _01617_;
  wire _01618_;
  wire _01619_;
  wire _01620_;
  wire _01621_;
  wire _01622_;
  wire _01623_;
  wire _01624_;
  wire _01625_;
  wire _01626_;
  wire _01627_;
  wire _01628_;
  wire _01629_;
  wire _01630_;
  wire _01631_;
  wire _01632_;
  wire _01633_;
  wire _01634_;
  wire _01635_;
  wire _01636_;
  wire _01637_;
  wire _01638_;
  wire _01639_;
  wire _01640_;
  wire _01641_;
  wire _01642_;
  wire _01643_;
  wire _01644_;
  wire _01645_;
  wire _01646_;
  wire _01647_;
  wire _01648_;
  wire _01649_;
  wire _01650_;
  wire _01651_;
  wire _01652_;
  wire _01653_;
  wire _01654_;
  wire _01655_;
  wire _01656_;
  wire _01657_;
  wire _01658_;
  wire _01659_;
  wire _01660_;
  wire _01661_;
  wire _01662_;
  wire _01663_;
  wire _01664_;
  wire _01665_;
  wire _01666_;
  wire _01667_;
  wire _01668_;
  wire _01669_;
  wire _01670_;
  wire _01671_;
  wire _01672_;
  wire _01673_;
  wire _01674_;
  wire _01675_;
  wire _01676_;
  wire _01677_;
  wire _01678_;
  wire _01679_;
  wire _01680_;
  wire _01681_;
  wire _01682_;
  wire _01683_;
  wire _01684_;
  wire _01685_;
  wire _01686_;
  wire _01687_;
  wire _01688_;
  wire _01689_;
  wire _01690_;
  wire _01691_;
  wire _01692_;
  wire _01693_;
  wire _01694_;
  wire _01695_;
  wire _01696_;
  wire _01697_;
  wire _01698_;
  wire _01699_;
  wire _01700_;
  wire _01701_;
  wire _01702_;
  wire _01703_;
  wire _01704_;
  wire _01705_;
  wire _01706_;
  wire _01707_;
  wire _01708_;
  wire _01709_;
  wire _01710_;
  wire _01711_;
  wire _01712_;
  wire _01713_;
  wire _01714_;
  wire _01715_;
  wire _01716_;
  wire _01717_;
  wire _01718_;
  wire _01719_;
  wire _01720_;
  wire _01721_;
  wire _01722_;
  wire _01723_;
  wire _01724_;
  wire _01725_;
  wire _01726_;
  wire _01727_;
  wire _01728_;
  wire _01729_;
  wire _01730_;
  wire _01731_;
  wire _01732_;
  wire _01733_;
  wire _01734_;
  wire _01735_;
  wire _01736_;
  wire _01737_;
  wire _01738_;
  wire _01739_;
  wire _01740_;
  wire _01741_;
  wire _01742_;
  wire _01743_;
  wire _01744_;
  wire _01745_;
  wire _01746_;
  wire _01747_;
  wire _01748_;
  wire _01749_;
  wire _01750_;
  wire _01751_;
  wire _01752_;
  wire _01753_;
  wire _01754_;
  wire _01755_;
  wire _01756_;
  wire _01757_;
  wire _01758_;
  wire _01759_;
  wire _01760_;
  wire _01761_;
  wire _01762_;
  wire _01763_;
  wire _01764_;
  wire _01765_;
  wire _01766_;
  wire _01767_;
  wire _01768_;
  wire _01769_;
  wire _01770_;
  wire _01771_;
  wire _01772_;
  wire _01773_;
  wire _01774_;
  wire _01775_;
  wire _01776_;
  wire _01777_;
  wire _01778_;
  wire _01779_;
  wire _01780_;
  wire _01781_;
  wire _01782_;
  wire _01783_;
  wire _01784_;
  wire _01785_;
  wire _01786_;
  wire _01787_;
  wire _01788_;
  wire _01789_;
  wire _01790_;
  wire _01791_;
  wire _01792_;
  wire _01793_;
  wire _01794_;
  wire _01795_;
  wire _01796_;
  wire _01797_;
  wire _01798_;
  wire _01799_;
  wire _01800_;
  wire _01801_;
  wire _01802_;
  wire _01803_;
  wire _01804_;
  wire _01805_;
  wire _01806_;
  wire _01807_;
  wire _01808_;
  wire _01809_;
  wire _01810_;
  wire _01811_;
  wire _01812_;
  wire _01813_;
  wire _01814_;
  wire _01815_;
  wire _01816_;
  wire _01817_;
  wire _01818_;
  wire _01819_;
  wire _01820_;
  wire _01821_;
  wire _01822_;
  wire _01823_;
  wire _01824_;
  wire _01825_;
  wire _01826_;
  wire _01827_;
  wire _01828_;
  wire _01829_;
  wire _01830_;
  wire _01831_;
  wire _01832_;
  wire _01833_;
  wire _01834_;
  wire _01835_;
  wire _01836_;
  wire _01837_;
  wire _01838_;
  wire _01839_;
  wire _01840_;
  wire _01841_;
  wire _01842_;
  wire _01843_;
  wire _01844_;
  wire _01845_;
  wire _01846_;
  wire _01847_;
  wire _01848_;
  wire _01849_;
  wire _01850_;
  wire _01851_;
  wire _01852_;
  wire _01853_;
  wire _01854_;
  wire _01855_;
  wire _01856_;
  wire _01857_;
  wire _01858_;
  wire _01859_;
  wire _01860_;
  wire _01861_;
  wire _01862_;
  wire _01863_;
  wire _01864_;
  wire _01865_;
  wire _01866_;
  wire _01867_;
  wire _01868_;
  wire _01869_;
  wire _01870_;
  wire _01871_;
  wire _01872_;
  wire _01873_;
  wire _01874_;
  wire _01875_;
  wire _01876_;
  wire _01877_;
  wire _01878_;
  wire _01879_;
  wire _01880_;
  wire _01881_;
  wire _01882_;
  wire _01883_;
  wire _01884_;
  wire _01885_;
  wire _01886_;
  wire _01887_;
  wire _01888_;
  wire _01889_;
  wire _01890_;
  wire _01891_;
  wire _01892_;
  wire _01893_;
  wire _01894_;
  wire _01895_;
  wire _01896_;
  wire _01897_;
  wire _01898_;
  wire _01899_;
  wire _01900_;
  wire _01901_;
  wire _01902_;
  wire _01903_;
  wire _01904_;
  wire _01905_;
  wire _01906_;
  wire _01907_;
  wire _01908_;
  wire _01909_;
  wire _01910_;
  wire _01911_;
  wire _01912_;
  wire _01913_;
  wire _01914_;
  wire _01915_;
  wire _01916_;
  wire _01917_;
  wire _01918_;
  wire _01919_;
  wire _01920_;
  wire _01921_;
  wire _01922_;
  wire _01923_;
  wire _01924_;
  wire _01925_;
  wire _01926_;
  wire _01927_;
  wire _01928_;
  wire _01929_;
  wire _01930_;
  wire _01931_;
  wire _01932_;
  wire _01933_;
  wire _01934_;
  wire _01935_;
  wire _01936_;
  wire _01937_;
  wire _01938_;
  wire _01939_;
  wire _01940_;
  wire _01941_;
  wire _01942_;
  wire _01943_;
  wire _01944_;
  wire _01945_;
  wire _01946_;
  wire _01947_;
  wire _01948_;
  wire _01949_;
  wire _01950_;
  wire _01951_;
  wire _01952_;
  wire _01953_;
  wire _01954_;
  wire _01955_;
  wire _01956_;
  wire _01957_;
  wire _01958_;
  wire _01959_;
  wire _01960_;
  wire _01961_;
  wire _01962_;
  wire _01963_;
  wire _01964_;
  wire _01965_;
  wire _01966_;
  wire _01967_;
  wire _01968_;
  wire _01969_;
  wire _01970_;
  wire _01971_;
  wire _01972_;
  wire _01973_;
  wire _01974_;
  wire _01975_;
  wire _01976_;
  wire _01977_;
  wire _01978_;
  wire _01979_;
  wire _01980_;
  wire _01981_;
  wire _01982_;
  wire _01983_;
  wire _01984_;
  wire _01985_;
  wire _01986_;
  wire _01987_;
  wire _01988_;
  wire _01989_;
  wire _01990_;
  wire _01991_;
  wire _01992_;
  wire _01993_;
  wire _01994_;
  wire _01995_;
  wire _01996_;
  wire _01997_;
  wire _01998_;
  wire _01999_;
  wire _02000_;
  wire _02001_;
  wire _02002_;
  wire _02003_;
  wire _02004_;
  wire _02005_;
  wire _02006_;
  wire _02007_;
  wire _02008_;
  wire _02009_;
  wire _02010_;
  wire _02011_;
  wire _02012_;
  wire _02013_;
  wire _02014_;
  wire _02015_;
  wire _02016_;
  wire _02017_;
  wire _02018_;
  wire _02019_;
  wire _02020_;
  wire _02021_;
  wire _02022_;
  wire _02023_;
  wire _02024_;
  wire _02025_;
  wire _02026_;
  wire _02027_;
  wire _02028_;
  wire _02029_;
  wire _02030_;
  wire _02031_;
  wire _02032_;
  wire _02033_;
  wire _02034_;
  wire _02035_;
  wire _02036_;
  wire _02037_;
  wire _02038_;
  wire _02039_;
  wire _02040_;
  wire _02041_;
  wire _02042_;
  wire _02043_;
  wire _02044_;
  wire _02045_;
  wire _02046_;
  wire _02047_;
  wire _02048_;
  wire _02049_;
  wire _02050_;
  wire _02051_;
  wire _02052_;
  wire _02053_;
  wire _02054_;
  wire _02055_;
  wire _02056_;
  wire _02057_;
  wire _02058_;
  wire _02059_;
  wire _02060_;
  wire _02061_;
  wire _02062_;
  wire _02063_;
  wire _02064_;
  wire _02065_;
  wire _02066_;
  wire _02067_;
  wire _02068_;
  wire _02069_;
  wire _02070_;
  wire _02071_;
  wire _02072_;
  wire _02073_;
  wire _02074_;
  wire _02075_;
  wire _02076_;
  wire _02077_;
  wire _02078_;
  wire _02079_;
  wire _02080_;
  wire _02081_;
  wire _02082_;
  wire _02083_;
  wire _02084_;
  wire _02085_;
  wire _02086_;
  wire _02087_;
  wire _02088_;
  wire _02089_;
  wire _02090_;
  wire _02091_;
  wire _02092_;
  wire _02093_;
  wire _02094_;
  wire _02095_;
  wire _02096_;
  wire _02097_;
  wire _02098_;
  wire _02099_;
  wire _02100_;
  wire _02101_;
  wire _02102_;
  wire _02103_;
  wire _02104_;
  wire _02105_;
  wire _02106_;
  wire _02107_;
  wire _02108_;
  wire _02109_;
  wire _02110_;
  wire _02111_;
  wire _02112_;
  wire _02113_;
  wire _02114_;
  wire _02115_;
  wire _02116_;
  wire _02117_;
  wire _02118_;
  wire _02119_;
  wire _02120_;
  wire _02121_;
  wire _02122_;
  wire _02123_;
  wire _02124_;
  wire _02125_;
  wire _02126_;
  wire _02127_;
  wire _02128_;
  wire _02129_;
  wire _02130_;
  wire _02131_;
  wire _02132_;
  wire _02133_;
  wire _02134_;
  wire _02135_;
  wire _02136_;
  wire _02137_;
  wire _02138_;
  wire _02139_;
  wire _02140_;
  wire _02141_;
  wire _02142_;
  wire _02143_;
  wire _02144_;
  wire _02145_;
  wire _02146_;
  wire _02147_;
  wire _02148_;
  wire _02149_;
  wire _02150_;
  wire _02151_;
  wire _02152_;
  wire _02153_;
  wire _02154_;
  wire _02155_;
  wire _02156_;
  wire _02157_;
  wire _02158_;
  wire _02159_;
  wire _02160_;
  wire _02161_;
  wire _02162_;
  wire _02163_;
  wire _02164_;
  wire _02165_;
  wire _02166_;
  wire _02167_;
  wire _02168_;
  wire _02169_;
  wire _02170_;
  wire _02171_;
  wire _02172_;
  wire _02173_;
  wire _02174_;
  wire _02175_;
  wire _02176_;
  wire _02177_;
  wire _02178_;
  wire _02179_;
  wire _02180_;
  wire _02181_;
  wire _02182_;
  wire _02183_;
  wire _02184_;
  wire _02185_;
  wire _02186_;
  wire _02187_;
  wire _02188_;
  wire _02189_;
  wire _02190_;
  wire _02191_;
  wire _02192_;
  wire _02193_;
  wire _02194_;
  wire _02195_;
  wire _02196_;
  wire _02197_;
  wire _02198_;
  wire _02199_;
  wire _02200_;
  wire _02201_;
  wire _02202_;
  wire _02203_;
  wire _02204_;
  wire _02205_;
  wire _02206_;
  wire _02207_;
  wire _02208_;
  wire _02209_;
  wire _02210_;
  wire _02211_;
  wire _02212_;
  wire _02213_;
  wire _02214_;
  wire _02215_;
  wire _02216_;
  wire _02217_;
  wire _02218_;
  wire _02219_;
  wire _02220_;
  wire _02221_;
  wire _02222_;
  wire _02223_;
  wire _02224_;
  wire _02225_;
  wire _02226_;
  wire _02227_;
  wire _02228_;
  wire _02229_;
  wire _02230_;
  wire _02231_;
  wire _02232_;
  wire _02233_;
  wire _02234_;
  wire _02235_;
  wire _02236_;
  wire _02237_;
  wire _02238_;
  wire _02239_;
  wire _02240_;
  wire _02241_;
  wire _02242_;
  wire _02243_;
  wire _02244_;
  wire _02245_;
  wire _02246_;
  wire _02247_;
  wire _02248_;
  wire _02249_;
  wire _02250_;
  wire _02251_;
  wire _02252_;
  wire _02253_;
  wire _02254_;
  wire _02255_;
  wire _02256_;
  wire _02257_;
  wire _02258_;
  wire _02259_;
  wire _02260_;
  wire _02261_;
  wire _02262_;
  wire _02263_;
  wire _02264_;
  wire _02265_;
  wire _02266_;
  wire _02267_;
  wire _02268_;
  wire _02269_;
  wire _02270_;
  wire _02271_;
  wire _02272_;
  wire _02273_;
  wire _02274_;
  wire _02275_;
  wire _02276_;
  wire _02277_;
  wire _02278_;
  wire _02279_;
  wire _02280_;
  wire _02281_;
  wire _02282_;
  wire _02283_;
  wire _02284_;
  wire _02285_;
  wire _02286_;
  wire _02287_;
  wire _02288_;
  wire _02289_;
  wire _02290_;
  wire _02291_;
  wire _02292_;
  wire _02293_;
  wire _02294_;
  wire _02295_;
  wire _02296_;
  wire _02297_;
  wire _02298_;
  wire _02299_;
  wire _02300_;
  wire _02301_;
  wire _02302_;
  wire _02303_;
  wire _02304_;
  wire _02305_;
  wire _02306_;
  wire _02307_;
  wire _02308_;
  wire _02309_;
  wire _02310_;
  wire _02311_;
  wire _02312_;
  wire _02313_;
  wire _02314_;
  wire _02315_;
  wire _02316_;
  wire _02317_;
  wire _02318_;
  wire _02319_;
  wire _02320_;
  wire _02321_;
  wire _02322_;
  wire _02323_;
  wire _02324_;
  wire _02325_;
  wire _02326_;
  wire _02327_;
  wire _02328_;
  wire _02329_;
  wire _02330_;
  wire _02331_;
  wire _02332_;
  wire _02333_;
  wire _02334_;
  wire _02335_;
  wire _02336_;
  wire _02337_;
  wire _02338_;
  wire _02339_;
  wire _02340_;
  wire _02341_;
  wire _02342_;
  wire _02343_;
  wire _02344_;
  wire _02345_;
  wire _02346_;
  wire _02347_;
  wire _02348_;
  wire _02349_;
  wire _02350_;
  wire _02351_;
  wire _02352_;
  wire _02353_;
  wire _02354_;
  wire _02355_;
  wire _02356_;
  wire _02357_;
  wire _02358_;
  wire _02359_;
  wire _02360_;
  wire _02361_;
  wire _02362_;
  wire _02363_;
  wire _02364_;
  wire _02365_;
  wire _02366_;
  wire _02367_;
  wire _02368_;
  wire _02369_;
  wire _02370_;
  wire _02371_;
  wire _02372_;
  wire _02373_;
  wire _02374_;
  wire _02375_;
  wire _02376_;
  wire _02377_;
  wire _02378_;
  wire _02379_;
  wire _02380_;
  wire _02381_;
  wire _02382_;
  wire _02383_;
  wire _02384_;
  wire _02385_;
  wire _02386_;
  wire _02387_;
  wire _02388_;
  wire _02389_;
  wire _02390_;
  wire _02391_;
  wire _02392_;
  wire _02393_;
  wire _02394_;
  wire _02395_;
  wire _02396_;
  wire _02397_;
  wire _02398_;
  wire _02399_;
  wire _02400_;
  wire _02401_;
  wire _02402_;
  wire _02403_;
  wire _02404_;
  wire _02405_;
  wire _02406_;
  wire _02407_;
  wire _02408_;
  wire _02409_;
  wire _02410_;
  wire _02411_;
  wire _02412_;
  wire _02413_;
  wire _02414_;
  wire _02415_;
  wire _02416_;
  wire _02417_;
  wire _02418_;
  wire _02419_;
  wire _02420_;
  wire _02421_;
  wire _02422_;
  wire _02423_;
  wire _02424_;
  wire _02425_;
  wire _02426_;
  wire _02427_;
  wire _02428_;
  wire _02429_;
  wire _02430_;
  wire _02431_;
  wire _02432_;
  wire _02433_;
  wire _02434_;
  wire _02435_;
  wire _02436_;
  wire _02437_;
  wire _02438_;
  wire _02439_;
  wire _02440_;
  wire _02441_;
  wire _02442_;
  wire _02443_;
  wire _02444_;
  wire _02445_;
  wire _02446_;
  wire _02447_;
  wire _02448_;
  wire _02449_;
  wire _02450_;
  wire _02451_;
  wire _02452_;
  wire _02453_;
  wire _02454_;
  wire _02455_;
  wire _02456_;
  wire _02457_;
  wire _02458_;
  wire _02459_;
  wire _02460_;
  wire _02461_;
  wire _02462_;
  wire _02463_;
  wire _02464_;
  wire _02465_;
  wire _02466_;
  wire _02467_;
  wire _02468_;
  wire _02469_;
  wire _02470_;
  wire _02471_;
  wire _02472_;
  wire _02473_;
  wire _02474_;
  wire _02475_;
  wire _02476_;
  wire _02477_;
  wire _02478_;
  wire _02479_;
  wire _02480_;
  wire _02481_;
  wire _02482_;
  wire _02483_;
  wire _02484_;
  wire _02485_;
  wire _02486_;
  wire _02487_;
  wire _02488_;
  wire _02489_;
  wire _02490_;
  wire _02491_;
  wire _02492_;
  wire _02493_;
  wire _02494_;
  wire _02495_;
  wire _02496_;
  wire _02497_;
  wire _02498_;
  wire _02499_;
  wire _02500_;
  wire _02501_;
  wire _02502_;
  wire _02503_;
  wire _02504_;
  wire _02505_;
  wire _02506_;
  wire _02507_;
  wire _02508_;
  wire _02509_;
  wire _02510_;
  wire _02511_;
  wire _02512_;
  wire _02513_;
  wire _02514_;
  wire _02515_;
  wire _02516_;
  wire _02517_;
  wire _02518_;
  wire _02519_;
  wire _02520_;
  wire _02521_;
  wire _02522_;
  wire _02523_;
  wire _02524_;
  wire _02525_;
  wire _02526_;
  wire _02527_;
  wire _02528_;
  wire _02529_;
  wire _02530_;
  wire _02531_;
  wire _02532_;
  wire _02533_;
  wire _02534_;
  wire _02535_;
  wire _02536_;
  wire _02537_;
  wire _02538_;
  wire _02539_;
  wire _02540_;
  wire _02541_;
  wire _02542_;
  wire _02543_;
  wire _02544_;
  wire _02545_;
  wire _02546_;
  wire _02547_;
  wire _02548_;
  wire _02549_;
  wire _02550_;
  wire _02551_;
  wire _02552_;
  wire _02553_;
  wire _02554_;
  wire _02555_;
  wire _02556_;
  wire _02557_;
  wire _02558_;
  wire _02559_;
  wire _02560_;
  wire _02561_;
  wire _02562_;
  wire _02563_;
  wire _02564_;
  wire _02565_;
  wire _02566_;
  wire _02567_;
  wire _02568_;
  wire _02569_;
  wire _02570_;
  wire _02571_;
  wire _02572_;
  wire _02573_;
  wire _02574_;
  wire _02575_;
  wire _02576_;
  wire _02577_;
  wire _02578_;
  wire _02579_;
  wire _02580_;
  wire _02581_;
  wire _02582_;
  wire _02583_;
  wire _02584_;
  wire _02585_;
  wire _02586_;
  wire _02587_;
  wire _02588_;
  wire _02589_;
  wire _02590_;
  wire _02591_;
  wire _02592_;
  wire _02593_;
  wire _02594_;
  wire _02595_;
  wire _02596_;
  wire _02597_;
  wire _02598_;
  wire _02599_;
  wire _02600_;
  wire _02601_;
  wire _02602_;
  wire _02603_;
  wire _02604_;
  wire _02605_;
  wire _02606_;
  wire _02607_;
  wire _02608_;
  wire _02609_;
  wire _02610_;
  wire _02611_;
  wire _02612_;
  wire _02613_;
  wire _02614_;
  wire _02615_;
  wire _02616_;
  wire _02617_;
  wire _02618_;
  wire _02619_;
  wire _02620_;
  wire _02621_;
  wire _02622_;
  wire _02623_;
  wire _02624_;
  wire _02625_;
  wire _02626_;
  wire _02627_;
  wire _02628_;
  wire _02629_;
  wire _02630_;
  wire _02631_;
  wire _02632_;
  wire _02633_;
  wire _02634_;
  wire _02635_;
  wire _02636_;
  wire _02637_;
  wire _02638_;
  wire _02639_;
  wire _02640_;
  wire _02641_;
  wire _02642_;
  wire _02643_;
  wire _02644_;
  wire _02645_;
  wire _02646_;
  wire _02647_;
  wire _02648_;
  wire _02649_;
  wire _02650_;
  wire _02651_;
  wire _02652_;
  wire _02653_;
  wire _02654_;
  wire _02655_;
  wire _02656_;
  wire _02657_;
  wire _02658_;
  wire _02659_;
  wire _02660_;
  wire _02661_;
  wire _02662_;
  wire _02663_;
  wire _02664_;
  wire _02665_;
  wire _02666_;
  wire _02667_;
  wire _02668_;
  wire _02669_;
  wire _02670_;
  wire _02671_;
  wire _02672_;
  wire _02673_;
  wire _02674_;
  wire _02675_;
  wire _02676_;
  wire _02677_;
  wire _02678_;
  wire _02679_;
  wire _02680_;
  wire _02681_;
  wire _02682_;
  wire _02683_;
  wire _02684_;
  wire _02685_;
  wire _02686_;
  wire _02687_;
  wire _02688_;
  wire _02689_;
  wire _02690_;
  wire _02691_;
  wire _02692_;
  wire _02693_;
  wire _02694_;
  wire _02695_;
  wire _02696_;
  wire _02697_;
  wire _02698_;
  wire _02699_;
  wire _02700_;
  wire _02701_;
  wire _02702_;
  wire _02703_;
  wire _02704_;
  wire _02705_;
  wire _02706_;
  wire _02707_;
  wire _02708_;
  wire _02709_;
  wire _02710_;
  wire _02711_;
  wire _02712_;
  wire _02713_;
  wire _02714_;
  wire _02715_;
  wire _02716_;
  wire _02717_;
  wire _02718_;
  wire _02719_;
  wire _02720_;
  wire _02721_;
  wire _02722_;
  wire _02723_;
  wire _02724_;
  wire _02725_;
  wire _02726_;
  wire _02727_;
  wire _02728_;
  wire _02729_;
  wire _02730_;
  wire _02731_;
  wire _02732_;
  wire _02733_;
  wire _02734_;
  wire _02735_;
  wire _02736_;
  wire _02737_;
  wire _02738_;
  wire _02739_;
  wire _02740_;
  wire _02741_;
  wire _02742_;
  wire _02743_;
  wire _02744_;
  wire _02745_;
  wire _02746_;
  wire _02747_;
  wire _02748_;
  wire _02749_;
  wire _02750_;
  wire _02751_;
  wire _02752_;
  wire _02753_;
  wire _02754_;
  wire _02755_;
  wire _02756_;
  wire _02757_;
  wire _02758_;
  wire _02759_;
  wire _02760_;
  wire _02761_;
  wire _02762_;
  wire _02763_;
  wire _02764_;
  wire _02765_;
  wire _02766_;
  wire _02767_;
  wire _02768_;
  wire _02769_;
  wire _02770_;
  wire _02771_;
  wire _02772_;
  wire _02773_;
  wire _02774_;
  wire _02775_;
  wire _02776_;
  wire _02777_;
  wire _02778_;
  wire _02779_;
  wire _02780_;
  wire _02781_;
  wire _02782_;
  wire _02783_;
  wire _02784_;
  wire _02785_;
  wire _02786_;
  wire _02787_;
  wire _02788_;
  wire _02789_;
  wire _02790_;
  wire _02791_;
  wire _02792_;
  wire _02793_;
  wire _02794_;
  wire _02795_;
  wire _02796_;
  wire _02797_;
  wire _02798_;
  wire _02799_;
  wire _02800_;
  wire _02801_;
  wire _02802_;
  wire _02803_;
  wire _02804_;
  wire _02805_;
  wire _02806_;
  wire _02807_;
  wire _02808_;
  wire _02809_;
  wire _02810_;
  wire _02811_;
  wire _02812_;
  wire _02813_;
  wire _02814_;
  wire _02815_;
  wire _02816_;
  wire _02817_;
  wire _02818_;
  wire _02819_;
  wire _02820_;
  wire _02821_;
  wire _02822_;
  wire _02823_;
  wire _02824_;
  wire _02825_;
  wire _02826_;
  wire _02827_;
  wire _02828_;
  wire _02829_;
  wire _02830_;
  wire _02831_;
  wire _02832_;
  wire _02833_;
  wire _02834_;
  wire _02835_;
  wire _02836_;
  wire _02837_;
  wire _02838_;
  wire _02839_;
  wire _02840_;
  wire _02841_;
  wire _02842_;
  wire _02843_;
  wire _02844_;
  wire _02845_;
  wire _02846_;
  wire _02847_;
  wire _02848_;
  wire _02849_;
  wire _02850_;
  wire _02851_;
  wire _02852_;
  wire _02853_;
  wire _02854_;
  wire _02855_;
  wire _02856_;
  wire _02857_;
  wire _02858_;
  wire _02859_;
  wire _02860_;
  wire _02861_;
  wire _02862_;
  wire _02863_;
  wire _02864_;
  wire _02865_;
  wire _02866_;
  wire _02867_;
  wire _02868_;
  wire _02869_;
  wire _02870_;
  wire _02871_;
  wire _02872_;
  wire _02873_;
  wire _02874_;
  wire _02875_;
  wire _02876_;
  wire _02877_;
  wire _02878_;
  wire _02879_;
  wire _02880_;
  wire _02881_;
  wire _02882_;
  wire _02883_;
  wire _02884_;
  wire _02885_;
  wire _02886_;
  wire _02887_;
  wire _02888_;
  wire _02889_;
  wire _02890_;
  wire _02891_;
  wire _02892_;
  wire _02893_;
  wire _02894_;
  wire _02895_;
  wire _02896_;
  wire _02897_;
  wire _02898_;
  wire _02899_;
  wire _02900_;
  wire _02901_;
  wire _02902_;
  wire _02903_;
  wire _02904_;
  wire _02905_;
  wire _02906_;
  wire _02907_;
  wire _02908_;
  wire _02909_;
  wire _02910_;
  wire _02911_;
  wire _02912_;
  wire _02913_;
  wire _02914_;
  wire _02915_;
  wire _02916_;
  wire _02917_;
  wire _02918_;
  wire _02919_;
  wire _02920_;
  wire _02921_;
  wire _02922_;
  wire _02923_;
  wire _02924_;
  wire _02925_;
  wire _02926_;
  wire _02927_;
  wire _02928_;
  wire _02929_;
  wire _02930_;
  wire _02931_;
  wire _02932_;
  wire _02933_;
  wire _02934_;
  wire _02935_;
  wire _02936_;
  wire _02937_;
  wire _02938_;
  wire _02939_;
  wire _02940_;
  wire _02941_;
  wire _02942_;
  wire _02943_;
  wire _02944_;
  wire _02945_;
  wire _02946_;
  wire _02947_;
  wire _02948_;
  wire _02949_;
  wire _02950_;
  wire _02951_;
  wire _02952_;
  wire _02953_;
  wire _02954_;
  wire _02955_;
  wire _02956_;
  wire _02957_;
  wire _02958_;
  wire _02959_;
  wire _02960_;
  wire _02961_;
  wire _02962_;
  wire _02963_;
  wire _02964_;
  wire _02965_;
  wire _02966_;
  wire _02967_;
  wire _02968_;
  wire _02969_;
  wire _02970_;
  wire _02971_;
  wire _02972_;
  wire _02973_;
  wire _02974_;
  wire _02975_;
  wire _02976_;
  wire _02977_;
  wire _02978_;
  wire _02979_;
  wire _02980_;
  wire _02981_;
  wire _02982_;
  wire _02983_;
  wire _02984_;
  wire _02985_;
  wire _02986_;
  wire _02987_;
  wire _02988_;
  wire _02989_;
  wire _02990_;
  wire _02991_;
  wire _02992_;
  wire _02993_;
  wire _02994_;
  wire _02995_;
  wire _02996_;
  wire _02997_;
  wire _02998_;
  wire _02999_;
  wire _03000_;
  wire _03001_;
  wire _03002_;
  wire _03003_;
  wire _03004_;
  wire _03005_;
  wire _03006_;
  wire _03007_;
  wire _03008_;
  wire _03009_;
  wire _03010_;
  wire _03011_;
  wire _03012_;
  wire _03013_;
  wire _03014_;
  wire _03015_;
  wire _03016_;
  wire _03017_;
  wire _03018_;
  wire _03019_;
  wire _03020_;
  wire _03021_;
  wire _03022_;
  wire _03023_;
  wire _03024_;
  wire _03025_;
  wire _03026_;
  wire _03027_;
  wire _03028_;
  wire _03029_;
  wire _03030_;
  wire _03031_;
  wire _03032_;
  wire _03033_;
  wire _03034_;
  wire _03035_;
  wire _03036_;
  wire _03037_;
  wire _03038_;
  wire _03039_;
  wire _03040_;
  wire _03041_;
  wire _03042_;
  wire _03043_;
  wire _03044_;
  wire _03045_;
  wire _03046_;
  wire _03047_;
  wire _03048_;
  wire _03049_;
  wire _03050_;
  wire _03051_;
  wire _03052_;
  wire _03053_;
  wire _03054_;
  wire _03055_;
  wire _03056_;
  wire _03057_;
  wire _03058_;
  wire _03059_;
  wire _03060_;
  wire _03061_;
  wire _03062_;
  wire _03063_;
  wire _03064_;
  wire _03065_;
  wire _03066_;
  wire _03067_;
  wire _03068_;
  wire _03069_;
  wire _03070_;
  wire _03071_;
  wire _03072_;
  wire _03073_;
  wire _03074_;
  wire _03075_;
  wire _03076_;
  wire _03077_;
  wire _03078_;
  wire _03079_;
  wire _03080_;
  wire _03081_;
  wire _03082_;
  wire _03083_;
  wire _03084_;
  wire _03085_;
  wire _03086_;
  wire _03087_;
  wire _03088_;
  wire _03089_;
  wire _03090_;
  wire _03091_;
  wire _03092_;
  wire _03093_;
  wire _03094_;
  wire _03095_;
  wire _03096_;
  wire _03097_;
  wire _03098_;
  wire _03099_;
  wire _03100_;
  wire _03101_;
  wire _03102_;
  wire _03103_;
  wire _03104_;
  wire _03105_;
  wire _03106_;
  wire _03107_;
  wire _03108_;
  wire _03109_;
  wire _03110_;
  wire _03111_;
  wire _03112_;
  wire _03113_;
  wire _03114_;
  wire _03115_;
  wire _03116_;
  wire _03117_;
  wire _03118_;
  wire _03119_;
  wire _03120_;
  wire _03121_;
  wire _03122_;
  wire _03123_;
  wire _03124_;
  wire _03125_;
  wire _03126_;
  wire _03127_;
  wire _03128_;
  wire _03129_;
  wire _03130_;
  wire _03131_;
  wire _03132_;
  wire _03133_;
  wire _03134_;
  wire _03135_;
  wire _03136_;
  wire _03137_;
  wire _03138_;
  wire _03139_;
  wire _03140_;
  wire _03141_;
  wire _03142_;
  wire _03143_;
  wire _03144_;
  wire _03145_;
  wire _03146_;
  wire _03147_;
  wire _03148_;
  wire _03149_;
  wire _03150_;
  wire _03151_;
  wire _03152_;
  wire _03153_;
  wire _03154_;
  wire _03155_;
  wire _03156_;
  wire _03157_;
  wire _03158_;
  wire _03159_;
  wire _03160_;
  wire _03161_;
  wire _03162_;
  wire _03163_;
  wire _03164_;
  wire _03165_;
  wire _03166_;
  wire _03167_;
  wire _03168_;
  wire _03169_;
  wire _03170_;
  wire _03171_;
  wire _03172_;
  wire _03173_;
  wire _03174_;
  wire _03175_;
  wire _03176_;
  wire _03177_;
  wire _03178_;
  wire _03179_;
  wire _03180_;
  wire _03181_;
  wire _03182_;
  wire _03183_;
  wire _03184_;
  wire _03185_;
  wire _03186_;
  wire _03187_;
  wire _03188_;
  wire _03189_;
  wire _03190_;
  wire _03191_;
  wire _03192_;
  wire _03193_;
  wire _03194_;
  wire _03195_;
  wire _03196_;
  wire _03197_;
  wire _03198_;
  wire _03199_;
  wire _03200_;
  wire _03201_;
  wire _03202_;
  wire _03203_;
  wire _03204_;
  wire _03205_;
  wire _03206_;
  wire _03207_;
  wire _03208_;
  wire _03209_;
  wire _03210_;
  wire _03211_;
  wire _03212_;
  wire _03213_;
  wire _03214_;
  wire _03215_;
  wire _03216_;
  wire _03217_;
  wire _03218_;
  wire _03219_;
  wire _03220_;
  wire _03221_;
  wire _03222_;
  wire _03223_;
  wire _03224_;
  wire _03225_;
  wire _03226_;
  wire _03227_;
  wire _03228_;
  wire _03229_;
  wire _03230_;
  wire _03231_;
  wire _03232_;
  wire _03233_;
  wire _03234_;
  wire _03235_;
  wire _03236_;
  wire _03237_;
  wire _03238_;
  wire _03239_;
  wire _03240_;
  wire _03241_;
  wire _03242_;
  wire _03243_;
  wire _03244_;
  wire _03245_;
  wire _03246_;
  wire _03247_;
  wire _03248_;
  wire _03249_;
  wire _03250_;
  wire _03251_;
  wire _03252_;
  wire _03253_;
  wire _03254_;
  wire _03255_;
  wire _03256_;
  wire _03257_;
  wire _03258_;
  wire _03259_;
  wire _03260_;
  wire _03261_;
  wire _03262_;
  wire _03263_;
  wire _03264_;
  wire _03265_;
  wire _03266_;
  wire _03267_;
  wire _03268_;
  wire _03269_;
  wire _03270_;
  wire _03271_;
  wire _03272_;
  wire _03273_;
  wire _03274_;
  wire _03275_;
  wire _03276_;
  wire _03277_;
  wire _03278_;
  wire _03279_;
  wire _03280_;
  wire _03281_;
  wire _03282_;
  wire _03283_;
  wire _03284_;
  wire _03285_;
  wire _03286_;
  wire _03287_;
  wire _03288_;
  wire _03289_;
  wire _03290_;
  wire _03291_;
  wire _03292_;
  wire _03293_;
  wire _03294_;
  wire _03295_;
  wire _03296_;
  wire _03297_;
  wire _03298_;
  wire _03299_;
  wire _03300_;
  wire _03301_;
  wire _03302_;
  wire _03303_;
  wire _03304_;
  wire _03305_;
  wire _03306_;
  wire _03307_;
  wire _03308_;
  wire _03309_;
  wire _03310_;
  wire _03311_;
  wire _03312_;
  wire _03313_;
  wire _03314_;
  wire _03315_;
  wire _03316_;
  wire _03317_;
  wire _03318_;
  wire _03319_;
  wire _03320_;
  wire _03321_;
  wire _03322_;
  wire _03323_;
  wire _03324_;
  wire _03325_;
  wire _03326_;
  wire _03327_;
  wire _03328_;
  wire _03329_;
  wire _03330_;
  wire _03331_;
  wire _03332_;
  wire _03333_;
  wire _03334_;
  wire _03335_;
  wire _03336_;
  wire _03337_;
  wire _03338_;
  wire _03339_;
  wire _03340_;
  wire _03341_;
  wire _03342_;
  wire _03343_;
  wire _03344_;
  wire _03345_;
  wire _03346_;
  wire _03347_;
  wire _03348_;
  wire _03349_;
  wire _03350_;
  wire _03351_;
  wire _03352_;
  wire _03353_;
  wire _03354_;
  wire _03355_;
  wire _03356_;
  wire _03357_;
  wire _03358_;
  wire _03359_;
  wire _03360_;
  wire _03361_;
  wire _03362_;
  wire _03363_;
  wire _03364_;
  wire _03365_;
  wire _03366_;
  wire _03367_;
  wire _03368_;
  wire _03369_;
  wire _03370_;
  wire _03371_;
  wire _03372_;
  wire _03373_;
  wire _03374_;
  wire _03375_;
  wire _03376_;
  wire _03377_;
  wire _03378_;
  wire _03379_;
  wire _03380_;
  wire _03381_;
  wire _03382_;
  wire _03383_;
  wire _03384_;
  wire _03385_;
  wire _03386_;
  wire _03387_;
  wire _03388_;
  wire _03389_;
  wire _03390_;
  wire _03391_;
  wire _03392_;
  wire _03393_;
  wire _03394_;
  wire _03395_;
  wire _03396_;
  wire _03397_;
  wire _03398_;
  wire _03399_;
  wire _03400_;
  wire _03401_;
  wire _03402_;
  wire _03403_;
  wire _03404_;
  wire _03405_;
  wire _03406_;
  wire _03407_;
  wire _03408_;
  wire _03409_;
  wire _03410_;
  wire _03411_;
  wire _03412_;
  wire _03413_;
  wire _03414_;
  wire _03415_;
  wire _03416_;
  wire _03417_;
  wire _03418_;
  wire _03419_;
  wire _03420_;
  wire _03421_;
  wire _03422_;
  wire _03423_;
  wire _03424_;
  wire _03425_;
  wire _03426_;
  wire _03427_;
  wire _03428_;
  wire _03429_;
  wire _03430_;
  wire _03431_;
  wire _03432_;
  wire _03433_;
  wire _03434_;
  wire _03435_;
  wire _03436_;
  wire _03437_;
  wire _03438_;
  wire _03439_;
  wire _03440_;
  wire _03441_;
  wire _03442_;
  wire _03443_;
  wire _03444_;
  wire _03445_;
  wire _03446_;
  wire _03447_;
  wire _03448_;
  wire _03449_;
  wire _03450_;
  wire _03451_;
  wire _03452_;
  wire _03453_;
  wire _03454_;
  wire _03455_;
  wire _03456_;
  wire _03457_;
  wire _03458_;
  wire _03459_;
  wire _03460_;
  wire _03461_;
  wire _03462_;
  wire _03463_;
  wire _03464_;
  wire _03465_;
  wire _03466_;
  wire _03467_;
  wire _03468_;
  wire _03469_;
  wire _03470_;
  wire _03471_;
  wire _03472_;
  wire _03473_;
  wire _03474_;
  wire _03475_;
  wire _03476_;
  wire _03477_;
  wire _03478_;
  wire _03479_;
  wire _03480_;
  wire _03481_;
  wire _03482_;
  wire _03483_;
  wire _03484_;
  wire _03485_;
  wire _03486_;
  wire _03487_;
  wire _03488_;
  wire _03489_;
  wire _03490_;
  wire _03491_;
  wire _03492_;
  wire _03493_;
  wire _03494_;
  wire _03495_;
  wire _03496_;
  wire _03497_;
  wire _03498_;
  wire _03499_;
  wire _03500_;
  wire _03501_;
  wire _03502_;
  wire _03503_;
  wire _03504_;
  wire _03505_;
  wire _03506_;
  wire _03507_;
  wire _03508_;
  wire _03509_;
  wire _03510_;
  wire _03511_;
  wire _03512_;
  wire _03513_;
  wire _03514_;
  wire _03515_;
  wire _03516_;
  wire _03517_;
  wire _03518_;
  wire _03519_;
  wire _03520_;
  wire _03521_;
  wire _03522_;
  wire _03523_;
  wire _03524_;
  wire _03525_;
  wire _03526_;
  wire _03527_;
  wire _03528_;
  wire _03529_;
  wire _03530_;
  wire _03531_;
  wire _03532_;
  wire _03533_;
  wire _03534_;
  wire _03535_;
  wire _03536_;
  wire _03537_;
  wire _03538_;
  wire _03539_;
  wire _03540_;
  wire _03541_;
  wire _03542_;
  wire _03543_;
  wire _03544_;
  wire _03545_;
  wire _03546_;
  wire _03547_;
  wire _03548_;
  wire _03549_;
  wire _03550_;
  wire _03551_;
  wire _03552_;
  wire _03553_;
  wire _03554_;
  wire _03555_;
  wire _03556_;
  wire _03557_;
  wire _03558_;
  wire _03559_;
  wire _03560_;
  wire _03561_;
  wire _03562_;
  wire _03563_;
  wire _03564_;
  wire _03565_;
  wire _03566_;
  wire _03567_;
  wire _03568_;
  wire _03569_;
  wire _03570_;
  wire _03571_;
  wire _03572_;
  wire _03573_;
  wire _03574_;
  wire _03575_;
  wire _03576_;
  wire _03577_;
  wire _03578_;
  wire _03579_;
  wire _03580_;
  wire _03581_;
  wire _03582_;
  wire _03583_;
  wire _03584_;
  wire _03585_;
  wire _03586_;
  wire _03587_;
  wire _03588_;
  wire _03589_;
  wire _03590_;
  wire _03591_;
  wire _03592_;
  wire _03593_;
  wire _03594_;
  wire _03595_;
  wire _03596_;
  wire _03597_;
  wire _03598_;
  wire _03599_;
  wire _03600_;
  wire _03601_;
  wire _03602_;
  wire _03603_;
  wire _03604_;
  wire _03605_;
  wire _03606_;
  wire _03607_;
  wire _03608_;
  wire _03609_;
  wire _03610_;
  wire _03611_;
  wire _03612_;
  wire _03613_;
  wire _03614_;
  wire _03615_;
  wire _03616_;
  wire _03617_;
  wire _03618_;
  wire _03619_;
  wire _03620_;
  wire _03621_;
  wire _03622_;
  wire _03623_;
  wire _03624_;
  wire _03625_;
  wire _03626_;
  wire _03627_;
  wire _03628_;
  wire _03629_;
  wire _03630_;
  wire _03631_;
  wire _03632_;
  wire _03633_;
  wire _03634_;
  wire _03635_;
  wire _03636_;
  wire _03637_;
  wire _03638_;
  wire _03639_;
  wire _03640_;
  wire _03641_;
  wire _03642_;
  wire _03643_;
  wire _03644_;
  wire _03645_;
  wire _03646_;
  wire _03647_;
  wire _03648_;
  wire _03649_;
  wire _03650_;
  wire _03651_;
  wire _03652_;
  wire _03653_;
  wire _03654_;
  wire _03655_;
  wire _03656_;
  wire _03657_;
  wire _03658_;
  wire _03659_;
  wire _03660_;
  wire _03661_;
  wire _03662_;
  wire _03663_;
  wire _03664_;
  wire _03665_;
  wire _03666_;
  wire _03667_;
  wire _03668_;
  wire _03669_;
  wire _03670_;
  wire _03671_;
  wire _03672_;
  wire _03673_;
  wire _03674_;
  wire _03675_;
  wire _03676_;
  wire _03677_;
  wire _03678_;
  wire _03679_;
  wire _03680_;
  wire _03681_;
  wire _03682_;
  wire _03683_;
  wire _03684_;
  wire _03685_;
  wire _03686_;
  wire _03687_;
  wire _03688_;
  wire _03689_;
  wire _03690_;
  wire _03691_;
  wire _03692_;
  wire _03693_;
  wire _03694_;
  wire _03695_;
  wire _03696_;
  wire _03697_;
  wire _03698_;
  wire _03699_;
  wire _03700_;
  wire _03701_;
  wire _03702_;
  wire _03703_;
  wire _03704_;
  wire _03705_;
  wire _03706_;
  wire _03707_;
  wire _03708_;
  wire _03709_;
  wire _03710_;
  wire _03711_;
  wire _03712_;
  wire _03713_;
  wire _03714_;
  wire _03715_;
  wire _03716_;
  wire _03717_;
  wire _03718_;
  wire _03719_;
  wire _03720_;
  wire _03721_;
  wire _03722_;
  wire _03723_;
  wire _03724_;
  wire _03725_;
  wire _03726_;
  wire _03727_;
  wire _03728_;
  wire _03729_;
  wire _03730_;
  wire _03731_;
  wire _03732_;
  wire _03733_;
  wire _03734_;
  wire _03735_;
  wire _03736_;
  wire _03737_;
  wire _03738_;
  wire _03739_;
  wire _03740_;
  wire _03741_;
  wire _03742_;
  wire _03743_;
  wire _03744_;
  wire _03745_;
  wire _03746_;
  wire _03747_;
  wire _03748_;
  wire _03749_;
  wire _03750_;
  wire _03751_;
  wire _03752_;
  wire _03753_;
  wire _03754_;
  wire _03755_;
  wire _03756_;
  wire _03757_;
  wire _03758_;
  wire _03759_;
  wire _03760_;
  wire _03761_;
  wire _03762_;
  wire _03763_;
  wire _03764_;
  wire _03765_;
  wire _03766_;
  wire _03767_;
  wire _03768_;
  wire _03769_;
  wire _03770_;
  wire _03771_;
  wire _03772_;
  wire _03773_;
  wire _03774_;
  wire _03775_;
  wire _03776_;
  wire _03777_;
  wire _03778_;
  wire _03779_;
  wire _03780_;
  wire _03781_;
  wire _03782_;
  wire _03783_;
  wire _03784_;
  wire _03785_;
  wire _03786_;
  wire _03787_;
  wire _03788_;
  wire _03789_;
  wire _03790_;
  wire _03791_;
  wire _03792_;
  wire _03793_;
  wire _03794_;
  wire _03795_;
  wire _03796_;
  wire _03797_;
  wire _03798_;
  wire _03799_;
  wire _03800_;
  wire _03801_;
  wire _03802_;
  wire _03803_;
  wire _03804_;
  wire _03805_;
  wire _03806_;
  wire _03807_;
  wire _03808_;
  wire _03809_;
  wire _03810_;
  wire _03811_;
  wire _03812_;
  wire _03813_;
  wire _03814_;
  wire _03815_;
  wire _03816_;
  wire _03817_;
  wire _03818_;
  wire _03819_;
  wire _03820_;
  wire _03821_;
  wire _03822_;
  wire _03823_;
  wire _03824_;
  wire _03825_;
  wire _03826_;
  wire _03827_;
  wire _03828_;
  wire _03829_;
  wire _03830_;
  wire _03831_;
  wire _03832_;
  wire _03833_;
  wire _03834_;
  wire _03835_;
  wire _03836_;
  wire _03837_;
  wire _03838_;
  wire _03839_;
  wire _03840_;
  wire _03841_;
  wire _03842_;
  wire _03843_;
  wire _03844_;
  wire _03845_;
  wire _03846_;
  wire _03847_;
  wire _03848_;
  wire _03849_;
  wire _03850_;
  wire _03851_;
  wire _03852_;
  wire _03853_;
  wire _03854_;
  wire _03855_;
  wire _03856_;
  wire _03857_;
  wire _03858_;
  wire _03859_;
  wire _03860_;
  wire _03861_;
  wire _03862_;
  wire _03863_;
  wire _03864_;
  wire _03865_;
  wire _03866_;
  wire _03867_;
  wire _03868_;
  wire _03869_;
  wire _03870_;
  wire _03871_;
  wire _03872_;
  wire _03873_;
  wire _03874_;
  wire _03875_;
  wire _03876_;
  wire _03877_;
  wire _03878_;
  wire _03879_;
  wire _03880_;
  wire _03881_;
  wire _03882_;
  wire _03883_;
  wire _03884_;
  wire _03885_;
  wire _03886_;
  wire _03887_;
  wire _03888_;
  wire _03889_;
  wire _03890_;
  wire _03891_;
  wire _03892_;
  wire _03893_;
  wire _03894_;
  wire _03895_;
  wire _03896_;
  wire _03897_;
  wire _03898_;
  wire _03899_;
  wire _03900_;
  wire _03901_;
  wire _03902_;
  wire _03903_;
  wire _03904_;
  wire _03905_;
  wire _03906_;
  wire _03907_;
  wire _03908_;
  wire _03909_;
  wire _03910_;
  wire _03911_;
  wire _03912_;
  wire _03913_;
  wire _03914_;
  wire _03915_;
  wire _03916_;
  wire _03917_;
  wire _03918_;
  wire _03919_;
  wire _03920_;
  wire _03921_;
  wire _03922_;
  wire _03923_;
  wire _03924_;
  wire _03925_;
  wire _03926_;
  wire _03927_;
  wire _03928_;
  wire _03929_;
  wire _03930_;
  wire _03931_;
  wire _03932_;
  wire _03933_;
  wire _03934_;
  wire _03935_;
  wire _03936_;
  wire _03937_;
  wire _03938_;
  wire _03939_;
  wire _03940_;
  wire _03941_;
  wire _03942_;
  wire _03943_;
  wire _03944_;
  wire _03945_;
  wire _03946_;
  wire _03947_;
  wire _03948_;
  wire _03949_;
  wire _03950_;
  wire _03951_;
  wire _03952_;
  wire _03953_;
  wire _03954_;
  wire _03955_;
  wire _03956_;
  wire _03957_;
  wire _03958_;
  wire _03959_;
  wire _03960_;
  wire _03961_;
  wire _03962_;
  wire _03963_;
  wire _03964_;
  wire _03965_;
  wire _03966_;
  wire _03967_;
  wire _03968_;
  wire _03969_;
  wire _03970_;
  wire _03971_;
  wire _03972_;
  wire _03973_;
  wire _03974_;
  wire _03975_;
  wire _03976_;
  wire _03977_;
  wire _03978_;
  wire _03979_;
  wire _03980_;
  wire _03981_;
  wire _03982_;
  wire _03983_;
  wire _03984_;
  wire _03985_;
  wire _03986_;
  wire _03987_;
  wire _03988_;
  wire _03989_;
  wire _03990_;
  wire _03991_;
  wire _03992_;
  wire _03993_;
  wire _03994_;
  wire _03995_;
  wire _03996_;
  wire _03997_;
  wire _03998_;
  wire _03999_;
  wire _04000_;
  wire _04001_;
  wire _04002_;
  wire _04003_;
  wire _04004_;
  wire _04005_;
  wire _04006_;
  wire _04007_;
  wire _04008_;
  wire _04009_;
  wire _04010_;
  wire _04011_;
  wire _04012_;
  wire _04013_;
  wire _04014_;
  wire _04015_;
  wire _04016_;
  wire _04017_;
  wire _04018_;
  wire _04019_;
  wire _04020_;
  wire _04021_;
  wire _04022_;
  wire _04023_;
  wire _04024_;
  wire _04025_;
  wire _04026_;
  wire _04027_;
  wire _04028_;
  wire _04029_;
  wire _04030_;
  wire _04031_;
  wire _04032_;
  wire _04033_;
  wire _04034_;
  wire _04035_;
  wire _04036_;
  wire _04037_;
  wire _04038_;
  wire _04039_;
  wire _04040_;
  wire _04041_;
  wire _04042_;
  wire _04043_;
  wire _04044_;
  wire _04045_;
  wire _04046_;
  wire _04047_;
  wire _04048_;
  wire _04049_;
  wire _04050_;
  wire _04051_;
  wire _04052_;
  wire _04053_;
  wire _04054_;
  wire _04055_;
  wire _04056_;
  wire _04057_;
  wire _04058_;
  wire _04059_;
  wire _04060_;
  wire _04061_;
  wire _04062_;
  wire _04063_;
  wire _04064_;
  wire _04065_;
  wire _04066_;
  wire _04067_;
  wire _04068_;
  wire _04069_;
  wire _04070_;
  wire _04071_;
  wire _04072_;
  wire _04073_;
  wire _04074_;
  wire _04075_;
  wire _04076_;
  wire _04077_;
  wire _04078_;
  wire _04079_;
  wire _04080_;
  wire _04081_;
  wire _04082_;
  wire _04083_;
  wire _04084_;
  wire _04085_;
  wire _04086_;
  wire _04087_;
  wire _04088_;
  wire _04089_;
  wire _04090_;
  wire _04091_;
  wire _04092_;
  wire _04093_;
  wire _04094_;
  wire _04095_;
  wire _04096_;
  wire _04097_;
  wire _04098_;
  wire _04099_;
  wire _04100_;
  wire _04101_;
  wire _04102_;
  wire _04103_;
  wire _04104_;
  wire _04105_;
  wire _04106_;
  wire _04107_;
  wire _04108_;
  wire _04109_;
  wire _04110_;
  wire _04111_;
  wire _04112_;
  wire _04113_;
  wire _04114_;
  wire _04115_;
  wire _04116_;
  wire _04117_;
  wire _04118_;
  wire _04119_;
  wire _04120_;
  wire _04121_;
  wire _04122_;
  wire _04123_;
  wire _04124_;
  wire _04125_;
  wire _04126_;
  wire _04127_;
  wire _04128_;
  wire _04129_;
  wire _04130_;
  wire _04131_;
  wire _04132_;
  wire _04133_;
  wire _04134_;
  wire _04135_;
  wire _04136_;
  wire _04137_;
  wire _04138_;
  wire _04139_;
  wire _04140_;
  wire _04141_;
  wire _04142_;
  wire _04143_;
  wire _04144_;
  wire _04145_;
  wire _04146_;
  wire _04147_;
  wire _04148_;
  wire _04149_;
  wire _04150_;
  wire _04151_;
  wire _04152_;
  wire _04153_;
  wire _04154_;
  wire _04155_;
  wire _04156_;
  wire _04157_;
  wire _04158_;
  wire _04159_;
  wire _04160_;
  wire _04161_;
  wire _04162_;
  wire _04163_;
  wire _04164_;
  wire _04165_;
  wire _04166_;
  wire _04167_;
  wire _04168_;
  wire _04169_;
  wire _04170_;
  wire _04171_;
  wire _04172_;
  wire _04173_;
  wire _04174_;
  wire _04175_;
  wire _04176_;
  wire _04177_;
  wire _04178_;
  wire _04179_;
  wire _04180_;
  wire _04181_;
  wire _04182_;
  wire _04183_;
  wire _04184_;
  wire _04185_;
  wire _04186_;
  wire _04187_;
  wire _04188_;
  wire _04189_;
  wire _04190_;
  wire _04191_;
  wire _04192_;
  wire _04193_;
  wire _04194_;
  wire _04195_;
  wire _04196_;
  wire _04197_;
  wire _04198_;
  wire _04199_;
  wire _04200_;
  wire _04201_;
  wire _04202_;
  wire _04203_;
  wire _04204_;
  wire _04205_;
  wire _04206_;
  wire _04207_;
  wire _04208_;
  wire _04209_;
  wire _04210_;
  wire _04211_;
  wire _04212_;
  wire _04213_;
  wire _04214_;
  wire _04215_;
  wire _04216_;
  wire _04217_;
  wire _04218_;
  wire _04219_;
  wire _04220_;
  wire _04221_;
  wire _04222_;
  wire _04223_;
  wire _04224_;
  wire _04225_;
  wire _04226_;
  wire _04227_;
  wire _04228_;
  wire _04229_;
  wire _04230_;
  wire _04231_;
  wire _04232_;
  wire _04233_;
  wire _04234_;
  wire _04235_;
  wire _04236_;
  wire _04237_;
  wire _04238_;
  wire _04239_;
  wire _04240_;
  wire _04241_;
  wire _04242_;
  wire _04243_;
  wire _04244_;
  wire _04245_;
  wire _04246_;
  wire _04247_;
  wire _04248_;
  wire _04249_;
  wire _04250_;
  wire _04251_;
  wire _04252_;
  wire _04253_;
  wire _04254_;
  wire _04255_;
  wire _04256_;
  wire _04257_;
  wire _04258_;
  wire _04259_;
  wire _04260_;
  wire _04261_;
  wire _04262_;
  wire _04263_;
  wire _04264_;
  wire _04265_;
  wire _04266_;
  wire _04267_;
  wire _04268_;
  wire _04269_;
  wire _04270_;
  wire _04271_;
  wire _04272_;
  wire _04273_;
  wire _04274_;
  wire _04275_;
  wire _04276_;
  wire _04277_;
  wire _04278_;
  wire _04279_;
  wire _04280_;
  wire _04281_;
  wire _04282_;
  wire _04283_;
  wire _04284_;
  wire _04285_;
  wire _04286_;
  wire _04287_;
  wire _04288_;
  wire _04289_;
  wire _04290_;
  wire _04291_;
  wire _04292_;
  wire _04293_;
  wire _04294_;
  wire _04295_;
  wire _04296_;
  wire _04297_;
  wire _04298_;
  wire _04299_;
  wire _04300_;
  wire _04301_;
  wire _04302_;
  wire _04303_;
  wire _04304_;
  wire _04305_;
  wire _04306_;
  wire _04307_;
  wire _04308_;
  wire _04309_;
  wire _04310_;
  wire _04311_;
  wire _04312_;
  wire _04313_;
  wire _04314_;
  wire _04315_;
  wire _04316_;
  wire _04317_;
  wire _04318_;
  wire _04319_;
  wire _04320_;
  wire _04321_;
  wire _04322_;
  wire _04323_;
  wire _04324_;
  wire _04325_;
  wire _04326_;
  wire _04327_;
  wire _04328_;
  wire _04329_;
  wire _04330_;
  wire _04331_;
  wire _04332_;
  wire _04333_;
  wire _04334_;
  wire _04335_;
  wire _04336_;
  wire _04337_;
  wire _04338_;
  wire _04339_;
  wire _04340_;
  wire _04341_;
  wire _04342_;
  wire _04343_;
  wire _04344_;
  wire _04345_;
  wire _04346_;
  wire _04347_;
  wire _04348_;
  wire _04349_;
  wire _04350_;
  wire _04351_;
  wire _04352_;
  wire _04353_;
  wire _04354_;
  wire _04355_;
  wire _04356_;
  wire _04357_;
  wire _04358_;
  wire _04359_;
  wire _04360_;
  wire _04361_;
  wire _04362_;
  wire _04363_;
  wire _04364_;
  wire _04365_;
  wire _04366_;
  wire _04367_;
  wire _04368_;
  wire _04369_;
  wire _04370_;
  wire _04371_;
  wire _04372_;
  wire _04373_;
  wire _04374_;
  wire _04375_;
  wire _04376_;
  wire _04377_;
  wire _04378_;
  wire _04379_;
  wire _04380_;
  wire _04381_;
  wire _04382_;
  wire _04383_;
  wire _04384_;
  wire _04385_;
  wire _04386_;
  wire _04387_;
  wire _04388_;
  wire _04389_;
  wire _04390_;
  wire _04391_;
  wire _04392_;
  wire _04393_;
  wire _04394_;
  wire _04395_;
  wire _04396_;
  wire _04397_;
  wire _04398_;
  wire _04399_;
  wire _04400_;
  wire _04401_;
  wire _04402_;
  wire _04403_;
  wire _04404_;
  wire _04405_;
  wire _04406_;
  wire _04407_;
  wire _04408_;
  wire _04409_;
  wire _04410_;
  wire _04411_;
  wire _04412_;
  wire _04413_;
  wire _04414_;
  wire _04415_;
  wire _04416_;
  wire _04417_;
  wire _04418_;
  wire _04419_;
  wire _04420_;
  wire _04421_;
  wire _04422_;
  wire _04423_;
  wire _04424_;
  wire _04425_;
  wire _04426_;
  wire _04427_;
  wire _04428_;
  wire _04429_;
  wire _04430_;
  wire _04431_;
  wire _04432_;
  wire _04433_;
  wire _04434_;
  wire _04435_;
  wire _04436_;
  wire _04437_;
  wire _04438_;
  wire _04439_;
  wire _04440_;
  wire _04441_;
  wire _04442_;
  wire _04443_;
  wire _04444_;
  wire _04445_;
  wire _04446_;
  wire _04447_;
  wire _04448_;
  wire _04449_;
  wire _04450_;
  wire _04451_;
  wire _04452_;
  wire _04453_;
  wire _04454_;
  wire _04455_;
  wire _04456_;
  wire _04457_;
  wire _04458_;
  wire _04459_;
  wire _04460_;
  wire _04461_;
  wire _04462_;
  wire _04463_;
  wire _04464_;
  wire _04465_;
  wire _04466_;
  wire _04467_;
  wire _04468_;
  wire _04469_;
  wire _04470_;
  wire _04471_;
  wire _04472_;
  wire _04473_;
  wire _04474_;
  wire _04475_;
  wire _04476_;
  wire _04477_;
  wire _04478_;
  wire _04479_;
  wire _04480_;
  wire _04481_;
  wire _04482_;
  wire _04483_;
  wire _04484_;
  wire _04485_;
  wire _04486_;
  wire _04487_;
  wire _04488_;
  wire _04489_;
  wire _04490_;
  wire _04491_;
  wire _04492_;
  wire _04493_;
  wire _04494_;
  wire _04495_;
  wire _04496_;
  wire _04497_;
  wire _04498_;
  wire _04499_;
  wire _04500_;
  wire _04501_;
  wire _04502_;
  wire _04503_;
  wire _04504_;
  wire _04505_;
  wire _04506_;
  wire _04507_;
  wire _04508_;
  wire _04509_;
  wire _04510_;
  wire _04511_;
  wire _04512_;
  wire _04513_;
  wire _04514_;
  wire _04515_;
  wire _04516_;
  wire _04517_;
  wire _04518_;
  wire _04519_;
  wire _04520_;
  wire _04521_;
  wire _04522_;
  wire _04523_;
  wire _04524_;
  wire _04525_;
  wire _04526_;
  wire _04527_;
  wire _04528_;
  wire _04529_;
  wire _04530_;
  wire _04531_;
  wire _04532_;
  wire _04533_;
  wire _04534_;
  wire _04535_;
  wire _04536_;
  wire _04537_;
  wire _04538_;
  wire _04539_;
  wire _04540_;
  wire _04541_;
  wire _04542_;
  wire _04543_;
  wire _04544_;
  wire _04545_;
  wire _04546_;
  wire _04547_;
  wire _04548_;
  wire _04549_;
  wire _04550_;
  wire _04551_;
  wire _04552_;
  wire _04553_;
  wire _04554_;
  wire _04555_;
  wire _04556_;
  wire _04557_;
  wire _04558_;
  wire _04559_;
  wire _04560_;
  wire _04561_;
  wire _04562_;
  wire _04563_;
  wire _04564_;
  wire _04565_;
  wire _04566_;
  wire _04567_;
  wire _04568_;
  wire _04569_;
  wire _04570_;
  wire _04571_;
  wire _04572_;
  wire _04573_;
  wire _04574_;
  wire _04575_;
  wire _04576_;
  wire _04577_;
  wire _04578_;
  wire _04579_;
  wire _04580_;
  wire _04581_;
  wire _04582_;
  wire _04583_;
  wire _04584_;
  wire _04585_;
  wire _04586_;
  wire _04587_;
  wire _04588_;
  wire _04589_;
  wire _04590_;
  wire _04591_;
  wire _04592_;
  wire _04593_;
  wire _04594_;
  wire _04595_;
  wire _04596_;
  wire _04597_;
  wire _04598_;
  wire _04599_;
  wire _04600_;
  wire _04601_;
  wire _04602_;
  wire _04603_;
  wire _04604_;
  wire _04605_;
  wire _04606_;
  wire _04607_;
  wire _04608_;
  wire _04609_;
  wire _04610_;
  wire _04611_;
  wire _04612_;
  wire _04613_;
  wire _04614_;
  wire _04615_;
  wire _04616_;
  wire _04617_;
  wire _04618_;
  wire _04619_;
  wire _04620_;
  wire _04621_;
  wire _04622_;
  wire _04623_;
  wire _04624_;
  wire _04625_;
  wire _04626_;
  wire _04627_;
  wire _04628_;
  wire _04629_;
  wire _04630_;
  wire _04631_;
  wire _04632_;
  wire _04633_;
  wire _04634_;
  wire _04635_;
  wire _04636_;
  wire _04637_;
  wire _04638_;
  wire _04639_;
  wire _04640_;
  wire _04641_;
  wire _04642_;
  wire _04643_;
  wire _04644_;
  wire _04645_;
  wire _04646_;
  wire _04647_;
  wire _04648_;
  wire _04649_;
  wire _04650_;
  wire _04651_;
  wire _04652_;
  wire _04653_;
  wire _04654_;
  wire _04655_;
  wire _04656_;
  wire _04657_;
  wire _04658_;
  wire _04659_;
  wire _04660_;
  wire _04661_;
  wire _04662_;
  wire _04663_;
  wire _04664_;
  wire _04665_;
  wire _04666_;
  wire _04667_;
  wire _04668_;
  wire _04669_;
  wire _04670_;
  wire _04671_;
  wire _04672_;
  wire _04673_;
  wire _04674_;
  wire _04675_;
  wire _04676_;
  wire _04677_;
  wire _04678_;
  wire _04679_;
  wire _04680_;
  wire _04681_;
  wire _04682_;
  wire _04683_;
  wire _04684_;
  wire _04685_;
  wire _04686_;
  wire _04687_;
  wire _04688_;
  wire _04689_;
  wire _04690_;
  wire _04691_;
  wire _04692_;
  wire _04693_;
  wire _04694_;
  wire _04695_;
  wire _04696_;
  wire _04697_;
  wire _04698_;
  wire _04699_;
  wire _04700_;
  wire _04701_;
  wire _04702_;
  wire _04703_;
  wire _04704_;
  wire _04705_;
  wire _04706_;
  wire _04707_;
  wire _04708_;
  wire _04709_;
  wire _04710_;
  wire _04711_;
  wire _04712_;
  wire _04713_;
  wire _04714_;
  wire _04715_;
  wire _04716_;
  wire _04717_;
  wire _04718_;
  wire _04719_;
  wire _04720_;
  wire _04721_;
  wire _04722_;
  wire _04723_;
  wire _04724_;
  wire _04725_;
  wire _04726_;
  wire _04727_;
  wire _04728_;
  wire _04729_;
  wire _04730_;
  wire _04731_;
  wire _04732_;
  wire _04733_;
  wire _04734_;
  wire _04735_;
  wire _04736_;
  wire _04737_;
  wire _04738_;
  wire _04739_;
  wire _04740_;
  wire _04741_;
  wire _04742_;
  wire _04743_;
  wire _04744_;
  wire _04745_;
  wire _04746_;
  wire _04747_;
  wire _04748_;
  wire _04749_;
  wire _04750_;
  wire _04751_;
  wire _04752_;
  wire _04753_;
  wire _04754_;
  wire _04755_;
  wire _04756_;
  wire _04757_;
  wire _04758_;
  wire _04759_;
  wire _04760_;
  wire _04761_;
  wire _04762_;
  wire _04763_;
  wire _04764_;
  wire _04765_;
  wire _04766_;
  wire _04767_;
  wire _04768_;
  wire _04769_;
  wire _04770_;
  wire _04771_;
  wire _04772_;
  wire _04773_;
  wire _04774_;
  wire _04775_;
  wire _04776_;
  wire _04777_;
  wire _04778_;
  wire _04779_;
  wire _04780_;
  wire _04781_;
  wire _04782_;
  wire _04783_;
  wire _04784_;
  wire _04785_;
  wire _04786_;
  wire _04787_;
  wire _04788_;
  wire _04789_;
  wire _04790_;
  wire _04791_;
  wire _04792_;
  wire _04793_;
  wire _04794_;
  wire _04795_;
  wire _04796_;
  wire _04797_;
  wire _04798_;
  wire _04799_;
  wire _04800_;
  wire _04801_;
  wire _04802_;
  wire _04803_;
  wire _04804_;
  wire _04805_;
  wire _04806_;
  wire _04807_;
  wire _04808_;
  wire _04809_;
  wire _04810_;
  wire _04811_;
  wire _04812_;
  wire _04813_;
  wire _04814_;
  wire _04815_;
  wire _04816_;
  wire _04817_;
  wire _04818_;
  wire _04819_;
  wire _04820_;
  wire _04821_;
  wire _04822_;
  wire _04823_;
  wire _04824_;
  wire _04825_;
  wire _04826_;
  wire _04827_;
  wire _04828_;
  wire _04829_;
  wire _04830_;
  wire _04831_;
  wire _04832_;
  wire _04833_;
  wire _04834_;
  wire _04835_;
  wire _04836_;
  wire _04837_;
  wire _04838_;
  wire _04839_;
  wire _04840_;
  wire _04841_;
  wire _04842_;
  wire _04843_;
  wire _04844_;
  wire _04845_;
  wire _04846_;
  wire _04847_;
  wire _04848_;
  wire _04849_;
  wire _04850_;
  wire _04851_;
  wire _04852_;
  wire _04853_;
  wire _04854_;
  wire _04855_;
  wire _04856_;
  wire _04857_;
  wire _04858_;
  wire _04859_;
  wire _04860_;
  wire _04861_;
  wire _04862_;
  wire _04863_;
  wire _04864_;
  wire _04865_;
  wire _04866_;
  wire _04867_;
  wire _04868_;
  wire _04869_;
  wire _04870_;
  wire _04871_;
  wire _04872_;
  wire _04873_;
  wire _04874_;
  wire _04875_;
  wire _04876_;
  wire _04877_;
  wire _04878_;
  wire _04879_;
  wire _04880_;
  wire _04881_;
  wire _04882_;
  wire _04883_;
  wire _04884_;
  wire _04885_;
  wire _04886_;
  wire _04887_;
  wire _04888_;
  wire _04889_;
  wire _04890_;
  wire _04891_;
  wire _04892_;
  wire _04893_;
  wire _04894_;
  wire _04895_;
  wire _04896_;
  wire _04897_;
  wire _04898_;
  wire _04899_;
  wire _04900_;
  wire _04901_;
  wire _04902_;
  wire _04903_;
  wire _04904_;
  wire _04905_;
  wire _04906_;
  wire _04907_;
  wire _04908_;
  wire _04909_;
  wire _04910_;
  wire _04911_;
  wire _04912_;
  wire _04913_;
  wire _04914_;
  wire _04915_;
  wire _04916_;
  wire _04917_;
  wire _04918_;
  wire _04919_;
  wire _04920_;
  wire _04921_;
  wire _04922_;
  wire _04923_;
  wire _04924_;
  wire _04925_;
  wire _04926_;
  wire _04927_;
  wire _04928_;
  wire _04929_;
  wire _04930_;
  wire _04931_;
  wire _04932_;
  wire _04933_;
  wire _04934_;
  wire _04935_;
  wire _04936_;
  wire _04937_;
  wire _04938_;
  wire _04939_;
  wire _04940_;
  wire _04941_;
  wire _04942_;
  wire _04943_;
  wire _04944_;
  wire _04945_;
  wire _04946_;
  wire _04947_;
  wire _04948_;
  wire _04949_;
  wire _04950_;
  wire _04951_;
  wire _04952_;
  wire _04953_;
  wire _04954_;
  wire _04955_;
  wire _04956_;
  wire _04957_;
  wire _04958_;
  wire _04959_;
  wire _04960_;
  wire _04961_;
  wire _04962_;
  wire _04963_;
  wire _04964_;
  wire _04965_;
  wire _04966_;
  wire _04967_;
  wire _04968_;
  wire _04969_;
  wire _04970_;
  wire _04971_;
  wire _04972_;
  wire _04973_;
  wire _04974_;
  wire _04975_;
  wire _04976_;
  wire _04977_;
  wire _04978_;
  wire _04979_;
  wire _04980_;
  wire _04981_;
  wire _04982_;
  wire _04983_;
  wire _04984_;
  wire _04985_;
  wire _04986_;
  wire _04987_;
  wire _04988_;
  wire _04989_;
  wire _04990_;
  wire _04991_;
  wire _04992_;
  wire _04993_;
  wire _04994_;
  wire _04995_;
  wire _04996_;
  wire _04997_;
  wire _04998_;
  wire _04999_;
  wire _05000_;
  wire _05001_;
  wire _05002_;
  wire _05003_;
  wire _05004_;
  wire _05005_;
  wire _05006_;
  wire _05007_;
  wire _05008_;
  wire _05009_;
  wire _05010_;
  wire _05011_;
  wire _05012_;
  wire _05013_;
  wire _05014_;
  wire _05015_;
  wire _05016_;
  wire _05017_;
  wire _05018_;
  wire _05019_;
  wire _05020_;
  wire _05021_;
  wire _05022_;
  wire _05023_;
  wire _05024_;
  wire _05025_;
  wire _05026_;
  wire _05027_;
  wire _05028_;
  wire _05029_;
  wire _05030_;
  wire _05031_;
  wire _05032_;
  wire _05033_;
  wire _05034_;
  wire _05035_;
  wire _05036_;
  wire _05037_;
  wire _05038_;
  wire _05039_;
  wire _05040_;
  wire _05041_;
  wire _05042_;
  wire _05043_;
  wire _05044_;
  wire _05045_;
  wire _05046_;
  wire _05047_;
  wire _05048_;
  wire _05049_;
  wire _05050_;
  wire _05051_;
  wire _05052_;
  wire _05053_;
  wire _05054_;
  wire _05055_;
  wire _05056_;
  wire _05057_;
  wire _05058_;
  wire _05059_;
  wire _05060_;
  wire _05061_;
  wire _05062_;
  wire _05063_;
  wire _05064_;
  wire _05065_;
  wire _05066_;
  wire _05067_;
  wire _05068_;
  wire _05069_;
  wire _05070_;
  wire _05071_;
  wire _05072_;
  wire _05073_;
  wire _05074_;
  wire _05075_;
  wire _05076_;
  wire _05077_;
  wire _05078_;
  wire _05079_;
  wire _05080_;
  wire _05081_;
  wire _05082_;
  wire _05083_;
  wire _05084_;
  wire _05085_;
  wire _05086_;
  wire _05087_;
  wire _05088_;
  wire _05089_;
  wire _05090_;
  wire _05091_;
  wire _05092_;
  wire _05093_;
  wire _05094_;
  wire _05095_;
  wire _05096_;
  wire _05097_;
  wire _05098_;
  wire _05099_;
  wire _05100_;
  wire _05101_;
  wire _05102_;
  wire _05103_;
  wire _05104_;
  wire _05105_;
  wire _05106_;
  wire _05107_;
  wire _05108_;
  wire _05109_;
  wire _05110_;
  wire _05111_;
  wire _05112_;
  wire _05113_;
  wire _05114_;
  wire _05115_;
  wire _05116_;
  wire _05117_;
  wire _05118_;
  wire _05119_;
  wire _05120_;
  wire _05121_;
  wire _05122_;
  wire _05123_;
  wire _05124_;
  wire _05125_;
  wire _05126_;
  wire _05127_;
  wire _05128_;
  wire _05129_;
  wire _05130_;
  wire _05131_;
  wire _05132_;
  wire _05133_;
  wire _05134_;
  wire _05135_;
  wire _05136_;
  wire _05137_;
  wire _05138_;
  wire _05139_;
  wire _05140_;
  wire _05141_;
  wire _05142_;
  wire _05143_;
  wire _05144_;
  wire _05145_;
  wire _05146_;
  wire _05147_;
  wire _05148_;
  wire _05149_;
  wire _05150_;
  wire _05151_;
  wire _05152_;
  wire _05153_;
  wire _05154_;
  wire _05155_;
  wire _05156_;
  wire _05157_;
  wire _05158_;
  wire _05159_;
  wire _05160_;
  wire _05161_;
  wire _05162_;
  wire _05163_;
  wire _05164_;
  wire _05165_;
  wire _05166_;
  wire _05167_;
  wire _05168_;
  wire _05169_;
  wire _05170_;
  wire _05171_;
  wire _05172_;
  wire _05173_;
  wire _05174_;
  wire _05175_;
  wire _05176_;
  wire _05177_;
  wire _05178_;
  wire _05179_;
  wire _05180_;
  wire _05181_;
  wire _05182_;
  wire _05183_;
  wire _05184_;
  wire _05185_;
  wire _05186_;
  wire _05187_;
  wire _05188_;
  wire _05189_;
  wire _05190_;
  wire _05191_;
  wire _05192_;
  wire _05193_;
  wire _05194_;
  wire _05195_;
  wire _05196_;
  wire _05197_;
  wire _05198_;
  wire _05199_;
  wire _05200_;
  wire _05201_;
  wire _05202_;
  wire _05203_;
  wire _05204_;
  wire _05205_;
  wire _05206_;
  wire _05207_;
  wire _05208_;
  wire _05209_;
  wire _05210_;
  wire _05211_;
  wire _05212_;
  wire _05213_;
  wire _05214_;
  wire _05215_;
  wire _05216_;
  wire _05217_;
  wire _05218_;
  wire _05219_;
  wire _05220_;
  wire _05221_;
  wire _05222_;
  wire _05223_;
  wire _05224_;
  wire _05225_;
  wire _05226_;
  wire _05227_;
  wire _05228_;
  wire _05229_;
  wire _05230_;
  wire _05231_;
  wire _05232_;
  wire _05233_;
  wire _05234_;
  wire _05235_;
  wire _05236_;
  wire _05237_;
  wire _05238_;
  wire _05239_;
  wire _05240_;
  wire _05241_;
  wire _05242_;
  wire _05243_;
  wire _05244_;
  wire _05245_;
  wire _05246_;
  wire _05247_;
  wire _05248_;
  wire _05249_;
  wire _05250_;
  wire _05251_;
  wire _05252_;
  wire _05253_;
  wire _05254_;
  wire _05255_;
  wire _05256_;
  wire _05257_;
  wire _05258_;
  wire _05259_;
  wire _05260_;
  wire _05261_;
  wire _05262_;
  wire _05263_;
  wire _05264_;
  wire _05265_;
  wire _05266_;
  wire _05267_;
  wire _05268_;
  wire _05269_;
  wire _05270_;
  wire _05271_;
  wire _05272_;
  wire _05273_;
  wire _05274_;
  wire _05275_;
  wire _05276_;
  wire _05277_;
  wire _05278_;
  wire _05279_;
  wire _05280_;
  wire _05281_;
  wire _05282_;
  wire _05283_;
  wire _05284_;
  wire _05285_;
  wire _05286_;
  wire _05287_;
  wire _05288_;
  wire _05289_;
  wire _05290_;
  wire _05291_;
  wire _05292_;
  wire _05293_;
  wire _05294_;
  wire _05295_;
  wire _05296_;
  wire _05297_;
  wire _05298_;
  wire _05299_;
  wire _05300_;
  wire _05301_;
  wire _05302_;
  wire _05303_;
  wire _05304_;
  wire _05305_;
  wire _05306_;
  wire _05307_;
  wire _05308_;
  wire _05309_;
  wire _05310_;
  wire _05311_;
  wire _05312_;
  wire _05313_;
  wire _05314_;
  wire _05315_;
  wire _05316_;
  wire _05317_;
  wire _05318_;
  wire _05319_;
  wire _05320_;
  wire _05321_;
  wire _05322_;
  wire _05323_;
  wire _05324_;
  wire _05325_;
  wire _05326_;
  wire _05327_;
  wire _05328_;
  wire _05329_;
  wire _05330_;
  wire _05331_;
  wire _05332_;
  wire _05333_;
  wire _05334_;
  wire _05335_;
  wire _05336_;
  wire _05337_;
  wire _05338_;
  wire _05339_;
  wire _05340_;
  wire _05341_;
  wire _05342_;
  wire _05343_;
  wire _05344_;
  wire _05345_;
  wire _05346_;
  wire _05347_;
  wire _05348_;
  wire _05349_;
  wire _05350_;
  wire _05351_;
  wire _05352_;
  wire _05353_;
  wire _05354_;
  wire _05355_;
  wire _05356_;
  wire _05357_;
  wire _05358_;
  wire _05359_;
  wire _05360_;
  wire _05361_;
  wire _05362_;
  wire _05363_;
  wire _05364_;
  wire _05365_;
  wire _05366_;
  wire _05367_;
  wire _05368_;
  wire _05369_;
  wire _05370_;
  wire _05371_;
  wire _05372_;
  wire _05373_;
  wire _05374_;
  wire _05375_;
  wire _05376_;
  wire _05377_;
  wire _05378_;
  wire _05379_;
  wire _05380_;
  wire _05381_;
  wire _05382_;
  wire _05383_;
  wire _05384_;
  wire _05385_;
  wire _05386_;
  wire _05387_;
  wire _05388_;
  wire _05389_;
  wire _05390_;
  wire _05391_;
  wire _05392_;
  wire _05393_;
  wire _05394_;
  wire _05395_;
  wire _05396_;
  wire _05397_;
  wire _05398_;
  wire _05399_;
  wire _05400_;
  wire _05401_;
  wire _05402_;
  wire _05403_;
  wire _05404_;
  wire _05405_;
  wire _05406_;
  wire _05407_;
  wire _05408_;
  wire _05409_;
  wire _05410_;
  wire _05411_;
  wire _05412_;
  wire _05413_;
  wire _05414_;
  wire _05415_;
  wire _05416_;
  wire _05417_;
  wire _05418_;
  wire _05419_;
  wire _05420_;
  wire _05421_;
  wire _05422_;
  wire _05423_;
  wire _05424_;
  wire _05425_;
  wire _05426_;
  wire _05427_;
  wire _05428_;
  wire _05429_;
  wire _05430_;
  wire _05431_;
  wire _05432_;
  wire _05433_;
  wire _05434_;
  wire _05435_;
  wire _05436_;
  wire _05437_;
  wire _05438_;
  wire _05439_;
  wire _05440_;
  wire _05441_;
  wire _05442_;
  wire _05443_;
  wire _05444_;
  wire _05445_;
  wire _05446_;
  wire _05447_;
  wire _05448_;
  wire _05449_;
  wire _05450_;
  wire _05451_;
  wire _05452_;
  wire _05453_;
  wire _05454_;
  wire _05455_;
  wire _05456_;
  wire _05457_;
  wire _05458_;
  wire _05459_;
  wire _05460_;
  wire _05461_;
  wire _05462_;
  wire _05463_;
  wire _05464_;
  wire _05465_;
  wire _05466_;
  wire _05467_;
  wire _05468_;
  wire _05469_;
  wire _05470_;
  wire _05471_;
  wire _05472_;
  wire _05473_;
  wire _05474_;
  wire _05475_;
  wire _05476_;
  wire _05477_;
  wire _05478_;
  wire _05479_;
  wire _05480_;
  wire _05481_;
  wire _05482_;
  wire _05483_;
  wire _05484_;
  wire _05485_;
  wire _05486_;
  wire _05487_;
  wire _05488_;
  wire _05489_;
  wire _05490_;
  wire _05491_;
  wire _05492_;
  wire _05493_;
  wire _05494_;
  wire _05495_;
  wire _05496_;
  wire _05497_;
  wire _05498_;
  wire _05499_;
  wire _05500_;
  wire _05501_;
  wire _05502_;
  wire _05503_;
  wire _05504_;
  wire _05505_;
  wire _05506_;
  wire _05507_;
  wire _05508_;
  wire _05509_;
  wire _05510_;
  wire _05511_;
  wire _05512_;
  wire _05513_;
  wire _05514_;
  wire _05515_;
  wire _05516_;
  wire _05517_;
  wire _05518_;
  wire _05519_;
  wire _05520_;
  wire _05521_;
  wire _05522_;
  wire _05523_;
  wire _05524_;
  wire _05525_;
  wire _05526_;
  wire _05527_;
  wire _05528_;
  wire _05529_;
  wire _05530_;
  wire _05531_;
  wire _05532_;
  wire _05533_;
  wire _05534_;
  wire _05535_;
  wire _05536_;
  wire _05537_;
  wire _05538_;
  wire _05539_;
  wire _05540_;
  wire _05541_;
  wire _05542_;
  wire _05543_;
  wire _05544_;
  wire _05545_;
  wire _05546_;
  wire _05547_;
  wire _05548_;
  wire _05549_;
  wire _05550_;
  wire _05551_;
  wire _05552_;
  wire _05553_;
  wire _05554_;
  wire _05555_;
  wire _05556_;
  wire _05557_;
  wire _05558_;
  wire _05559_;
  wire _05560_;
  wire _05561_;
  wire _05562_;
  wire _05563_;
  wire _05564_;
  wire _05565_;
  wire _05566_;
  wire _05567_;
  wire _05568_;
  wire _05569_;
  wire _05570_;
  wire _05571_;
  wire _05572_;
  wire _05573_;
  wire _05574_;
  wire _05575_;
  wire _05576_;
  wire _05577_;
  wire _05578_;
  wire _05579_;
  wire _05580_;
  wire _05581_;
  wire _05582_;
  wire _05583_;
  wire _05584_;
  wire _05585_;
  wire _05586_;
  wire _05587_;
  wire _05588_;
  wire _05589_;
  wire _05590_;
  wire _05591_;
  wire _05592_;
  wire _05593_;
  wire _05594_;
  wire _05595_;
  wire _05596_;
  wire _05597_;
  wire _05598_;
  wire _05599_;
  wire _05600_;
  wire _05601_;
  wire _05602_;
  wire _05603_;
  wire _05604_;
  wire _05605_;
  wire _05606_;
  wire _05607_;
  wire _05608_;
  wire _05609_;
  wire _05610_;
  wire _05611_;
  wire _05612_;
  wire _05613_;
  wire _05614_;
  wire _05615_;
  wire _05616_;
  wire _05617_;
  wire _05618_;
  wire _05619_;
  wire _05620_;
  wire _05621_;
  wire _05622_;
  wire _05623_;
  wire _05624_;
  wire _05625_;
  wire _05626_;
  wire _05627_;
  wire _05628_;
  wire _05629_;
  wire _05630_;
  wire _05631_;
  wire _05632_;
  wire _05633_;
  wire _05634_;
  wire _05635_;
  wire _05636_;
  wire _05637_;
  wire _05638_;
  wire _05639_;
  wire _05640_;
  wire _05641_;
  wire _05642_;
  wire _05643_;
  wire _05644_;
  wire _05645_;
  wire _05646_;
  wire _05647_;
  wire _05648_;
  wire _05649_;
  wire _05650_;
  wire _05651_;
  wire _05652_;
  wire _05653_;
  wire _05654_;
  wire _05655_;
  wire _05656_;
  wire _05657_;
  wire _05658_;
  wire _05659_;
  wire _05660_;
  wire _05661_;
  wire _05662_;
  wire _05663_;
  wire _05664_;
  wire _05665_;
  wire _05666_;
  wire _05667_;
  wire _05668_;
  wire _05669_;
  wire _05670_;
  wire _05671_;
  wire _05672_;
  wire _05673_;
  wire _05674_;
  wire _05675_;
  wire _05676_;
  wire _05677_;
  wire _05678_;
  wire _05679_;
  wire _05680_;
  wire _05681_;
  wire _05682_;
  wire _05683_;
  wire _05684_;
  wire _05685_;
  wire _05686_;
  wire _05687_;
  wire _05688_;
  wire _05689_;
  wire _05690_;
  wire _05691_;
  wire _05692_;
  wire _05693_;
  wire _05694_;
  wire _05695_;
  wire _05696_;
  wire _05697_;
  wire _05698_;
  wire _05699_;
  wire _05700_;
  wire _05701_;
  wire _05702_;
  wire _05703_;
  wire _05704_;
  wire _05705_;
  wire _05706_;
  wire _05707_;
  wire _05708_;
  wire _05709_;
  wire _05710_;
  wire _05711_;
  wire _05712_;
  wire _05713_;
  wire _05714_;
  wire _05715_;
  wire _05716_;
  wire _05717_;
  wire _05718_;
  wire _05719_;
  wire _05720_;
  wire _05721_;
  wire _05722_;
  wire _05723_;
  wire _05724_;
  wire _05725_;
  wire _05726_;
  wire _05727_;
  wire _05728_;
  wire _05729_;
  wire _05730_;
  wire _05731_;
  wire _05732_;
  wire _05733_;
  wire _05734_;
  wire _05735_;
  wire _05736_;
  wire _05737_;
  wire _05738_;
  wire _05739_;
  wire _05740_;
  wire _05741_;
  wire _05742_;
  wire _05743_;
  wire _05744_;
  wire _05745_;
  wire _05746_;
  wire _05747_;
  wire _05748_;
  wire _05749_;
  wire _05750_;
  wire _05751_;
  wire _05752_;
  wire _05753_;
  wire _05754_;
  wire _05755_;
  wire _05756_;
  wire _05757_;
  wire _05758_;
  wire _05759_;
  wire _05760_;
  wire _05761_;
  wire _05762_;
  wire _05763_;
  wire _05764_;
  wire _05765_;
  wire _05766_;
  wire _05767_;
  wire _05768_;
  wire _05769_;
  wire _05770_;
  wire _05771_;
  wire _05772_;
  wire _05773_;
  wire _05774_;
  wire _05775_;
  wire _05776_;
  wire _05777_;
  wire _05778_;
  wire _05779_;
  wire _05780_;
  wire _05781_;
  wire _05782_;
  wire _05783_;
  wire _05784_;
  wire _05785_;
  wire _05786_;
  wire _05787_;
  wire _05788_;
  wire _05789_;
  wire _05790_;
  wire _05791_;
  wire _05792_;
  wire _05793_;
  wire _05794_;
  wire _05795_;
  wire _05796_;
  wire _05797_;
  wire _05798_;
  wire _05799_;
  wire _05800_;
  wire _05801_;
  wire _05802_;
  wire _05803_;
  wire _05804_;
  wire _05805_;
  wire _05806_;
  wire _05807_;
  wire _05808_;
  wire _05809_;
  wire _05810_;
  wire _05811_;
  wire _05812_;
  wire _05813_;
  wire _05814_;
  wire _05815_;
  wire _05816_;
  wire _05817_;
  wire _05818_;
  wire _05819_;
  wire _05820_;
  wire _05821_;
  wire _05822_;
  wire _05823_;
  wire _05824_;
  wire _05825_;
  wire _05826_;
  wire _05827_;
  wire _05828_;
  wire _05829_;
  wire _05830_;
  wire _05831_;
  wire _05832_;
  wire _05833_;
  wire _05834_;
  wire _05835_;
  wire _05836_;
  wire _05837_;
  wire _05838_;
  wire _05839_;
  wire _05840_;
  wire _05841_;
  wire _05842_;
  wire _05843_;
  wire _05844_;
  wire _05845_;
  wire _05846_;
  wire _05847_;
  wire _05848_;
  wire _05849_;
  wire _05850_;
  wire _05851_;
  wire _05852_;
  wire _05853_;
  wire _05854_;
  wire _05855_;
  wire _05856_;
  wire _05857_;
  wire _05858_;
  wire _05859_;
  wire _05860_;
  wire _05861_;
  wire _05862_;
  wire _05863_;
  wire _05864_;
  wire _05865_;
  wire _05866_;
  wire _05867_;
  wire _05868_;
  wire _05869_;
  wire _05870_;
  wire _05871_;
  wire _05872_;
  wire _05873_;
  wire _05874_;
  wire _05875_;
  wire _05876_;
  wire _05877_;
  wire _05878_;
  wire _05879_;
  wire _05880_;
  wire _05881_;
  wire _05882_;
  wire _05883_;
  wire _05884_;
  wire _05885_;
  wire _05886_;
  wire _05887_;
  wire _05888_;
  wire _05889_;
  wire _05890_;
  wire _05891_;
  wire _05892_;
  wire _05893_;
  wire _05894_;
  wire _05895_;
  wire _05896_;
  wire _05897_;
  wire _05898_;
  wire _05899_;
  wire _05900_;
  wire _05901_;
  wire _05902_;
  wire _05903_;
  wire _05904_;
  wire _05905_;
  wire _05906_;
  wire _05907_;
  wire _05908_;
  wire _05909_;
  wire _05910_;
  wire _05911_;
  wire _05912_;
  wire _05913_;
  wire _05914_;
  wire _05915_;
  wire _05916_;
  wire _05917_;
  wire _05918_;
  wire _05919_;
  wire _05920_;
  wire _05921_;
  wire _05922_;
  wire _05923_;
  wire _05924_;
  wire _05925_;
  wire _05926_;
  wire _05927_;
  wire _05928_;
  wire _05929_;
  wire _05930_;
  wire _05931_;
  wire _05932_;
  wire _05933_;
  wire _05934_;
  wire _05935_;
  wire _05936_;
  wire _05937_;
  wire _05938_;
  wire _05939_;
  wire _05940_;
  wire _05941_;
  wire _05942_;
  wire _05943_;
  wire _05944_;
  wire _05945_;
  wire _05946_;
  wire _05947_;
  wire _05948_;
  wire _05949_;
  wire _05950_;
  wire _05951_;
  wire _05952_;
  wire _05953_;
  wire _05954_;
  wire _05955_;
  wire _05956_;
  wire _05957_;
  wire _05958_;
  wire _05959_;
  wire _05960_;
  wire _05961_;
  wire _05962_;
  wire _05963_;
  wire _05964_;
  wire _05965_;
  wire _05966_;
  wire _05967_;
  wire _05968_;
  wire _05969_;
  wire _05970_;
  wire _05971_;
  wire _05972_;
  wire _05973_;
  wire _05974_;
  wire _05975_;
  wire _05976_;
  wire _05977_;
  wire _05978_;
  wire _05979_;
  wire _05980_;
  wire _05981_;
  wire _05982_;
  wire _05983_;
  wire _05984_;
  wire _05985_;
  wire _05986_;
  wire _05987_;
  wire _05988_;
  wire _05989_;
  wire _05990_;
  wire _05991_;
  wire _05992_;
  wire _05993_;
  wire _05994_;
  wire _05995_;
  wire _05996_;
  wire _05997_;
  wire _05998_;
  wire _05999_;
  wire _06000_;
  wire _06001_;
  wire _06002_;
  wire _06003_;
  wire _06004_;
  wire _06005_;
  wire _06006_;
  wire _06007_;
  wire _06008_;
  wire _06009_;
  wire _06010_;
  wire _06011_;
  wire _06012_;
  wire _06013_;
  wire _06014_;
  wire _06015_;
  wire _06016_;
  wire _06017_;
  wire _06018_;
  wire _06019_;
  wire _06020_;
  wire _06021_;
  wire _06022_;
  wire _06023_;
  wire _06024_;
  wire _06025_;
  wire _06026_;
  wire _06027_;
  wire _06028_;
  wire _06029_;
  wire _06030_;
  wire _06031_;
  wire _06032_;
  wire _06033_;
  wire _06034_;
  wire _06035_;
  wire _06036_;
  wire _06037_;
  wire _06038_;
  wire _06039_;
  wire _06040_;
  wire _06041_;
  wire _06042_;
  wire _06043_;
  wire _06044_;
  wire _06045_;
  wire _06046_;
  wire _06047_;
  wire _06048_;
  wire _06049_;
  wire _06050_;
  wire _06051_;
  wire _06052_;
  wire _06053_;
  wire _06054_;
  wire _06055_;
  wire _06056_;
  wire _06057_;
  wire _06058_;
  wire _06059_;
  wire _06060_;
  wire _06061_;
  wire _06062_;
  wire _06063_;
  wire _06064_;
  wire _06065_;
  wire _06066_;
  wire _06067_;
  wire _06068_;
  wire _06069_;
  wire _06070_;
  wire _06071_;
  wire _06072_;
  wire _06073_;
  wire _06074_;
  wire _06075_;
  wire _06076_;
  wire _06077_;
  wire _06078_;
  wire _06079_;
  wire _06080_;
  wire _06081_;
  wire _06082_;
  wire _06083_;
  wire _06084_;
  wire _06085_;
  wire _06086_;
  wire _06087_;
  wire _06088_;
  wire _06089_;
  wire _06090_;
  wire _06091_;
  wire _06092_;
  wire _06093_;
  wire _06094_;
  wire _06095_;
  wire _06096_;
  wire _06097_;
  wire _06098_;
  wire _06099_;
  wire _06100_;
  wire _06101_;
  wire _06102_;
  wire _06103_;
  wire _06104_;
  wire _06105_;
  wire _06106_;
  wire _06107_;
  wire _06108_;
  wire _06109_;
  wire _06110_;
  wire _06111_;
  wire _06112_;
  wire _06113_;
  wire _06114_;
  wire _06115_;
  wire _06116_;
  wire _06117_;
  wire _06118_;
  wire _06119_;
  wire _06120_;
  wire _06121_;
  wire _06122_;
  wire _06123_;
  wire _06124_;
  wire _06125_;
  wire _06126_;
  wire _06127_;
  wire _06128_;
  wire _06129_;
  wire _06130_;
  wire _06131_;
  wire _06132_;
  wire _06133_;
  wire _06134_;
  wire _06135_;
  wire _06136_;
  wire _06137_;
  wire _06138_;
  wire _06139_;
  wire _06140_;
  wire _06141_;
  wire _06142_;
  wire _06143_;
  wire _06144_;
  wire _06145_;
  wire _06146_;
  wire _06147_;
  wire _06148_;
  wire _06149_;
  wire _06150_;
  wire _06151_;
  wire _06152_;
  wire _06153_;
  wire _06154_;
  wire _06155_;
  wire _06156_;
  wire _06157_;
  wire _06158_;
  wire _06159_;
  wire _06160_;
  wire _06161_;
  wire _06162_;
  wire _06163_;
  wire _06164_;
  wire _06165_;
  wire _06166_;
  wire _06167_;
  wire _06168_;
  wire _06169_;
  wire _06170_;
  wire _06171_;
  wire _06172_;
  wire _06173_;
  wire _06174_;
  wire _06175_;
  wire _06176_;
  wire _06177_;
  wire _06178_;
  wire _06179_;
  wire _06180_;
  wire _06181_;
  wire _06182_;
  wire _06183_;
  wire _06184_;
  wire _06185_;
  wire _06186_;
  wire _06187_;
  wire _06188_;
  wire _06189_;
  wire _06190_;
  wire _06191_;
  wire _06192_;
  wire _06193_;
  wire _06194_;
  wire _06195_;
  wire _06196_;
  wire _06197_;
  wire _06198_;
  wire _06199_;
  wire _06200_;
  wire _06201_;
  wire _06202_;
  wire _06203_;
  wire _06204_;
  wire _06205_;
  wire _06206_;
  wire _06207_;
  wire _06208_;
  wire _06209_;
  wire _06210_;
  wire _06211_;
  wire _06212_;
  wire _06213_;
  wire _06214_;
  wire _06215_;
  wire _06216_;
  wire _06217_;
  wire _06218_;
  wire _06219_;
  wire _06220_;
  wire _06221_;
  wire _06222_;
  wire _06223_;
  wire _06224_;
  wire _06225_;
  wire _06226_;
  wire _06227_;
  wire _06228_;
  wire _06229_;
  wire _06230_;
  wire _06231_;
  wire _06232_;
  wire _06233_;
  wire _06234_;
  wire _06235_;
  wire _06236_;
  wire _06237_;
  wire _06238_;
  wire _06239_;
  wire _06240_;
  wire _06241_;
  wire _06242_;
  wire _06243_;
  wire _06244_;
  wire _06245_;
  wire _06246_;
  wire _06247_;
  wire _06248_;
  wire _06249_;
  wire _06250_;
  wire _06251_;
  wire _06252_;
  wire _06253_;
  wire _06254_;
  wire _06255_;
  wire _06256_;
  wire _06257_;
  wire _06258_;
  wire _06259_;
  wire _06260_;
  wire _06261_;
  wire _06262_;
  wire _06263_;
  wire _06264_;
  wire _06265_;
  wire _06266_;
  wire _06267_;
  wire _06268_;
  wire _06269_;
  wire _06270_;
  wire _06271_;
  wire _06272_;
  wire _06273_;
  wire _06274_;
  wire _06275_;
  wire _06276_;
  wire _06277_;
  wire _06278_;
  wire _06279_;
  wire _06280_;
  wire _06281_;
  wire _06282_;
  wire _06283_;
  wire _06284_;
  wire _06285_;
  wire _06286_;
  wire _06287_;
  wire _06288_;
  wire _06289_;
  wire _06290_;
  wire _06291_;
  wire _06292_;
  wire _06293_;
  wire _06294_;
  wire _06295_;
  wire _06296_;
  wire _06297_;
  wire _06298_;
  wire _06299_;
  wire _06300_;
  wire _06301_;
  wire _06302_;
  wire _06303_;
  wire _06304_;
  wire _06305_;
  wire _06306_;
  wire _06307_;
  wire _06308_;
  wire _06309_;
  wire _06310_;
  wire _06311_;
  wire _06312_;
  wire _06313_;
  wire _06314_;
  wire _06315_;
  wire _06316_;
  wire _06317_;
  wire _06318_;
  wire _06319_;
  wire _06320_;
  wire _06321_;
  wire _06322_;
  wire _06323_;
  wire _06324_;
  wire _06325_;
  wire _06326_;
  wire _06327_;
  wire _06328_;
  wire _06329_;
  wire _06330_;
  wire _06331_;
  wire _06332_;
  wire _06333_;
  wire _06334_;
  wire _06335_;
  wire _06336_;
  wire _06337_;
  wire _06338_;
  wire _06339_;
  wire _06340_;
  wire _06341_;
  wire _06342_;
  wire _06343_;
  wire _06344_;
  wire _06345_;
  wire _06346_;
  wire _06347_;
  wire _06348_;
  wire _06349_;
  wire _06350_;
  wire _06351_;
  wire _06352_;
  wire _06353_;
  wire _06354_;
  wire _06355_;
  wire _06356_;
  wire _06357_;
  wire _06358_;
  wire _06359_;
  wire _06360_;
  wire _06361_;
  wire _06362_;
  wire _06363_;
  wire _06364_;
  wire _06365_;
  wire _06366_;
  wire _06367_;
  wire _06368_;
  wire _06369_;
  wire _06370_;
  wire _06371_;
  wire _06372_;
  wire _06373_;
  wire _06374_;
  wire _06375_;
  wire _06376_;
  wire _06377_;
  wire _06378_;
  wire _06379_;
  wire _06380_;
  wire _06381_;
  wire _06382_;
  wire _06383_;
  wire _06384_;
  wire _06385_;
  wire _06386_;
  wire _06387_;
  wire _06388_;
  wire _06389_;
  wire _06390_;
  wire _06391_;
  wire _06392_;
  wire _06393_;
  wire _06394_;
  wire _06395_;
  wire _06396_;
  wire _06397_;
  wire _06398_;
  wire _06399_;
  wire _06400_;
  wire _06401_;
  wire _06402_;
  wire _06403_;
  wire _06404_;
  wire _06405_;
  wire _06406_;
  wire _06407_;
  wire _06408_;
  wire _06409_;
  wire _06410_;
  wire _06411_;
  wire _06412_;
  wire _06413_;
  wire _06414_;
  wire _06415_;
  wire _06416_;
  wire _06417_;
  wire _06418_;
  wire _06419_;
  wire _06420_;
  wire _06421_;
  wire _06422_;
  wire _06423_;
  wire _06424_;
  wire _06425_;
  wire _06426_;
  wire _06427_;
  wire _06428_;
  wire _06429_;
  wire _06430_;
  wire _06431_;
  wire _06432_;
  wire _06433_;
  wire _06434_;
  wire _06435_;
  wire _06436_;
  wire _06437_;
  wire _06438_;
  wire _06439_;
  wire _06440_;
  wire _06441_;
  wire _06442_;
  wire _06443_;
  wire _06444_;
  wire _06445_;
  wire _06446_;
  wire _06447_;
  wire _06448_;
  wire _06449_;
  wire _06450_;
  wire _06451_;
  wire _06452_;
  wire _06453_;
  wire _06454_;
  wire _06455_;
  wire _06456_;
  wire _06457_;
  wire _06458_;
  wire _06459_;
  wire _06460_;
  wire _06461_;
  wire _06462_;
  wire _06463_;
  wire _06464_;
  wire _06465_;
  wire _06466_;
  wire _06467_;
  wire _06468_;
  wire _06469_;
  wire _06470_;
  wire _06471_;
  wire _06472_;
  wire _06473_;
  wire _06474_;
  wire _06475_;
  wire _06476_;
  wire _06477_;
  wire _06478_;
  wire _06479_;
  wire _06480_;
  wire _06481_;
  wire _06482_;
  wire _06483_;
  wire _06484_;
  wire _06485_;
  wire _06486_;
  wire _06487_;
  wire _06488_;
  wire _06489_;
  wire _06490_;
  wire _06491_;
  wire _06492_;
  wire _06493_;
  wire _06494_;
  wire _06495_;
  wire _06496_;
  wire _06497_;
  wire _06498_;
  wire _06499_;
  wire _06500_;
  wire _06501_;
  wire _06502_;
  wire _06503_;
  wire _06504_;
  wire _06505_;
  wire _06506_;
  wire _06507_;
  wire _06508_;
  wire _06509_;
  wire _06510_;
  wire _06511_;
  wire _06512_;
  wire _06513_;
  wire _06514_;
  wire _06515_;
  wire _06516_;
  wire _06517_;
  wire _06518_;
  wire _06519_;
  wire _06520_;
  wire _06521_;
  wire _06522_;
  wire _06523_;
  wire _06524_;
  wire _06525_;
  wire _06526_;
  wire _06527_;
  wire _06528_;
  wire _06529_;
  wire _06530_;
  wire _06531_;
  wire _06532_;
  wire _06533_;
  wire _06534_;
  wire _06535_;
  wire _06536_;
  wire _06537_;
  wire _06538_;
  wire _06539_;
  wire _06540_;
  wire _06541_;
  wire _06542_;
  wire _06543_;
  wire _06544_;
  wire _06545_;
  wire _06546_;
  wire _06547_;
  wire _06548_;
  wire _06549_;
  wire _06550_;
  wire _06551_;
  wire _06552_;
  wire _06553_;
  wire _06554_;
  wire _06555_;
  wire _06556_;
  wire _06557_;
  wire _06558_;
  wire _06559_;
  wire _06560_;
  wire _06561_;
  wire _06562_;
  wire _06563_;
  wire _06564_;
  wire _06565_;
  wire _06566_;
  wire _06567_;
  wire _06568_;
  wire _06569_;
  wire _06570_;
  wire _06571_;
  wire _06572_;
  wire _06573_;
  wire _06574_;
  wire _06575_;
  wire _06576_;
  wire _06577_;
  wire _06578_;
  wire _06579_;
  wire _06580_;
  wire _06581_;
  wire _06582_;
  wire _06583_;
  wire _06584_;
  wire _06585_;
  wire _06586_;
  wire _06587_;
  wire _06588_;
  wire _06589_;
  wire _06590_;
  wire _06591_;
  wire _06592_;
  wire _06593_;
  wire _06594_;
  wire _06595_;
  wire _06596_;
  wire _06597_;
  wire _06598_;
  wire _06599_;
  wire _06600_;
  wire _06601_;
  wire _06602_;
  wire _06603_;
  wire _06604_;
  wire _06605_;
  wire _06606_;
  wire _06607_;
  wire _06608_;
  wire _06609_;
  wire _06610_;
  wire _06611_;
  wire _06612_;
  wire _06613_;
  wire _06614_;
  wire _06615_;
  wire _06616_;
  wire _06617_;
  wire _06618_;
  wire _06619_;
  wire _06620_;
  wire _06621_;
  wire _06622_;
  wire _06623_;
  wire _06624_;
  wire _06625_;
  wire _06626_;
  wire _06627_;
  wire _06628_;
  wire _06629_;
  wire _06630_;
  wire _06631_;
  wire _06632_;
  wire _06633_;
  wire _06634_;
  wire _06635_;
  wire _06636_;
  wire _06637_;
  wire _06638_;
  wire _06639_;
  wire _06640_;
  wire _06641_;
  wire _06642_;
  wire _06643_;
  wire _06644_;
  wire _06645_;
  wire _06646_;
  wire _06647_;
  wire _06648_;
  wire _06649_;
  wire _06650_;
  wire _06651_;
  wire _06652_;
  wire _06653_;
  wire _06654_;
  wire _06655_;
  wire _06656_;
  wire _06657_;
  wire _06658_;
  wire _06659_;
  wire _06660_;
  wire _06661_;
  wire _06662_;
  wire _06663_;
  wire _06664_;
  wire _06665_;
  wire _06666_;
  wire _06667_;
  wire _06668_;
  wire _06669_;
  wire _06670_;
  wire _06671_;
  wire _06672_;
  wire _06673_;
  wire _06674_;
  wire _06675_;
  wire _06676_;
  wire _06677_;
  wire _06678_;
  wire _06679_;
  wire _06680_;
  wire _06681_;
  wire _06682_;
  wire _06683_;
  wire _06684_;
  wire _06685_;
  wire _06686_;
  wire _06687_;
  wire _06688_;
  wire _06689_;
  wire _06690_;
  wire _06691_;
  wire _06692_;
  wire _06693_;
  wire _06694_;
  wire _06695_;
  wire _06696_;
  wire _06697_;
  wire _06698_;
  wire _06699_;
  wire _06700_;
  wire _06701_;
  wire _06702_;
  wire _06703_;
  wire _06704_;
  wire _06705_;
  wire _06706_;
  wire _06707_;
  wire _06708_;
  wire _06709_;
  wire _06710_;
  wire _06711_;
  wire _06712_;
  wire _06713_;
  wire _06714_;
  wire _06715_;
  wire _06716_;
  wire _06717_;
  wire _06718_;
  wire _06719_;
  wire _06720_;
  wire _06721_;
  wire _06722_;
  wire _06723_;
  wire _06724_;
  wire _06725_;
  wire _06726_;
  wire _06727_;
  wire _06728_;
  wire _06729_;
  wire _06730_;
  wire _06731_;
  wire _06732_;
  wire _06733_;
  wire _06734_;
  wire _06735_;
  wire _06736_;
  wire _06737_;
  wire _06738_;
  wire _06739_;
  wire _06740_;
  wire _06741_;
  wire _06742_;
  wire _06743_;
  wire _06744_;
  wire _06745_;
  wire _06746_;
  wire _06747_;
  wire _06748_;
  wire _06749_;
  wire _06750_;
  wire _06751_;
  wire _06752_;
  wire _06753_;
  wire _06754_;
  wire _06755_;
  wire _06756_;
  wire _06757_;
  wire _06758_;
  wire _06759_;
  wire _06760_;
  wire _06761_;
  wire _06762_;
  wire _06763_;
  wire _06764_;
  wire _06765_;
  wire _06766_;
  wire _06767_;
  wire _06768_;
  wire _06769_;
  wire _06770_;
  wire _06771_;
  wire _06772_;
  wire _06773_;
  wire _06774_;
  wire _06775_;
  wire _06776_;
  wire _06777_;
  wire _06778_;
  wire _06779_;
  wire _06780_;
  wire _06781_;
  wire _06782_;
  wire _06783_;
  wire _06784_;
  wire _06785_;
  wire _06786_;
  wire _06787_;
  wire _06788_;
  wire _06789_;
  wire _06790_;
  wire _06791_;
  wire _06792_;
  wire _06793_;
  wire _06794_;
  wire _06795_;
  wire _06796_;
  wire _06797_;
  wire _06798_;
  wire _06799_;
  wire _06800_;
  wire _06801_;
  wire _06802_;
  wire _06803_;
  wire _06804_;
  wire _06805_;
  wire _06806_;
  wire _06807_;
  wire _06808_;
  wire _06809_;
  wire _06810_;
  wire _06811_;
  wire _06812_;
  wire _06813_;
  wire _06814_;
  wire _06815_;
  wire _06816_;
  wire _06817_;
  wire _06818_;
  wire _06819_;
  wire _06820_;
  wire _06821_;
  wire _06822_;
  wire _06823_;
  wire _06824_;
  wire _06825_;
  wire _06826_;
  wire _06827_;
  wire _06828_;
  wire _06829_;
  wire _06830_;
  wire _06831_;
  wire _06832_;
  wire _06833_;
  wire _06834_;
  wire _06835_;
  wire _06836_;
  wire _06837_;
  wire _06838_;
  wire _06839_;
  wire _06840_;
  wire _06841_;
  wire _06842_;
  wire _06843_;
  wire _06844_;
  wire _06845_;
  wire _06846_;
  wire _06847_;
  wire _06848_;
  wire _06849_;
  wire _06850_;
  wire _06851_;
  wire _06852_;
  wire _06853_;
  wire _06854_;
  wire _06855_;
  wire _06856_;
  wire _06857_;
  wire _06858_;
  wire _06859_;
  wire _06860_;
  wire _06861_;
  wire _06862_;
  wire _06863_;
  wire _06864_;
  wire _06865_;
  wire _06866_;
  wire _06867_;
  wire _06868_;
  wire _06869_;
  wire _06870_;
  wire _06871_;
  wire _06872_;
  wire _06873_;
  wire _06874_;
  wire _06875_;
  wire _06876_;
  wire _06877_;
  wire _06878_;
  wire _06879_;
  wire _06880_;
  wire _06881_;
  wire _06882_;
  wire _06883_;
  wire _06884_;
  wire _06885_;
  wire _06886_;
  wire _06887_;
  wire _06888_;
  wire _06889_;
  wire _06890_;
  wire _06891_;
  wire _06892_;
  wire _06893_;
  wire _06894_;
  wire _06895_;
  wire _06896_;
  wire _06897_;
  wire _06898_;
  wire _06899_;
  wire _06900_;
  wire _06901_;
  wire _06902_;
  wire _06903_;
  wire _06904_;
  wire _06905_;
  wire _06906_;
  wire _06907_;
  wire _06908_;
  wire _06909_;
  wire _06910_;
  wire _06911_;
  wire _06912_;
  wire _06913_;
  wire _06914_;
  wire _06915_;
  wire _06916_;
  wire _06917_;
  wire _06918_;
  wire _06919_;
  wire _06920_;
  wire _06921_;
  wire _06922_;
  wire _06923_;
  wire _06924_;
  wire _06925_;
  wire _06926_;
  wire _06927_;
  wire _06928_;
  wire _06929_;
  wire _06930_;
  wire _06931_;
  wire _06932_;
  wire _06933_;
  wire _06934_;
  wire _06935_;
  wire _06936_;
  wire _06937_;
  wire _06938_;
  wire _06939_;
  wire _06940_;
  wire _06941_;
  wire _06942_;
  wire _06943_;
  wire _06944_;
  wire _06945_;
  wire _06946_;
  wire _06947_;
  wire _06948_;
  wire _06949_;
  wire _06950_;
  wire _06951_;
  wire _06952_;
  wire _06953_;
  wire _06954_;
  wire _06955_;
  wire _06956_;
  wire _06957_;
  wire _06958_;
  wire _06959_;
  wire _06960_;
  wire _06961_;
  wire _06962_;
  wire _06963_;
  wire _06964_;
  wire _06965_;
  wire _06966_;
  wire _06967_;
  wire _06968_;
  wire _06969_;
  wire _06970_;
  wire _06971_;
  wire _06972_;
  wire _06973_;
  wire _06974_;
  wire _06975_;
  wire _06976_;
  wire _06977_;
  wire _06978_;
  wire _06979_;
  wire _06980_;
  wire _06981_;
  wire _06982_;
  wire _06983_;
  wire _06984_;
  wire _06985_;
  wire _06986_;
  wire _06987_;
  wire _06988_;
  wire _06989_;
  wire _06990_;
  wire _06991_;
  wire _06992_;
  wire _06993_;
  wire _06994_;
  wire _06995_;
  wire _06996_;
  wire _06997_;
  wire _06998_;
  wire _06999_;
  wire _07000_;
  wire _07001_;
  wire _07002_;
  wire _07003_;
  wire _07004_;
  wire _07005_;
  wire _07006_;
  wire _07007_;
  wire _07008_;
  wire _07009_;
  wire _07010_;
  wire _07011_;
  wire _07012_;
  wire _07013_;
  wire _07014_;
  wire _07015_;
  wire _07016_;
  wire _07017_;
  wire _07018_;
  wire _07019_;
  wire _07020_;
  wire _07021_;
  wire _07022_;
  wire _07023_;
  wire _07024_;
  wire _07025_;
  wire _07026_;
  wire _07027_;
  wire _07028_;
  wire _07029_;
  wire _07030_;
  wire _07031_;
  wire _07032_;
  wire _07033_;
  wire _07034_;
  wire _07035_;
  wire _07036_;
  wire _07037_;
  wire _07038_;
  wire _07039_;
  wire _07040_;
  wire _07041_;
  wire _07042_;
  wire _07043_;
  wire _07044_;
  wire _07045_;
  wire _07046_;
  wire _07047_;
  wire _07048_;
  wire _07049_;
  wire _07050_;
  wire _07051_;
  wire _07052_;
  wire _07053_;
  wire _07054_;
  wire _07055_;
  wire _07056_;
  wire _07057_;
  wire _07058_;
  wire _07059_;
  wire _07060_;
  wire _07061_;
  wire _07062_;
  wire _07063_;
  wire _07064_;
  wire _07065_;
  wire _07066_;
  wire _07067_;
  wire _07068_;
  wire _07069_;
  wire _07070_;
  wire _07071_;
  wire _07072_;
  wire _07073_;
  wire _07074_;
  wire _07075_;
  wire _07076_;
  wire _07077_;
  wire _07078_;
  wire _07079_;
  wire _07080_;
  wire _07081_;
  wire _07082_;
  wire _07083_;
  wire _07084_;
  wire _07085_;
  wire _07086_;
  wire _07087_;
  wire _07088_;
  wire _07089_;
  wire _07090_;
  wire _07091_;
  wire _07092_;
  wire _07093_;
  wire _07094_;
  wire _07095_;
  wire _07096_;
  wire _07097_;
  wire _07098_;
  wire _07099_;
  wire _07100_;
  wire _07101_;
  wire _07102_;
  wire _07103_;
  wire _07104_;
  wire _07105_;
  wire _07106_;
  wire _07107_;
  wire _07108_;
  wire _07109_;
  wire _07110_;
  wire _07111_;
  wire _07112_;
  wire _07113_;
  wire _07114_;
  wire _07115_;
  wire _07116_;
  wire _07117_;
  wire _07118_;
  wire _07119_;
  wire _07120_;
  wire _07121_;
  wire _07122_;
  wire _07123_;
  wire _07124_;
  wire _07125_;
  wire _07126_;
  wire _07127_;
  wire _07128_;
  wire _07129_;
  wire _07130_;
  wire _07131_;
  wire _07132_;
  wire _07133_;
  wire _07134_;
  wire _07135_;
  wire _07136_;
  wire _07137_;
  wire _07138_;
  wire _07139_;
  wire _07140_;
  wire _07141_;
  wire _07142_;
  wire _07143_;
  wire _07144_;
  wire _07145_;
  wire _07146_;
  wire _07147_;
  wire _07148_;
  wire _07149_;
  wire _07150_;
  wire _07151_;
  wire _07152_;
  wire _07153_;
  wire _07154_;
  wire _07155_;
  wire _07156_;
  wire _07157_;
  wire _07158_;
  wire _07159_;
  wire _07160_;
  wire _07161_;
  wire _07162_;
  wire _07163_;
  wire _07164_;
  wire _07165_;
  wire _07166_;
  wire _07167_;
  wire _07168_;
  wire _07169_;
  wire _07170_;
  wire _07171_;
  wire _07172_;
  wire _07173_;
  wire _07174_;
  wire _07175_;
  wire _07176_;
  wire _07177_;
  wire _07178_;
  wire _07179_;
  wire _07180_;
  wire _07181_;
  wire _07182_;
  wire _07183_;
  wire _07184_;
  wire _07185_;
  wire _07186_;
  wire _07187_;
  wire _07188_;
  wire _07189_;
  wire _07190_;
  wire _07191_;
  wire _07192_;
  wire _07193_;
  wire _07194_;
  wire _07195_;
  wire _07196_;
  wire _07197_;
  wire _07198_;
  wire _07199_;
  wire _07200_;
  wire _07201_;
  wire _07202_;
  wire _07203_;
  wire _07204_;
  wire _07205_;
  wire _07206_;
  wire _07207_;
  wire _07208_;
  wire _07209_;
  wire _07210_;
  wire _07211_;
  wire _07212_;
  wire _07213_;
  wire _07214_;
  wire _07215_;
  wire _07216_;
  wire _07217_;
  wire _07218_;
  wire _07219_;
  wire _07220_;
  wire _07221_;
  wire _07222_;
  wire _07223_;
  wire _07224_;
  wire _07225_;
  wire _07226_;
  wire _07227_;
  wire _07228_;
  wire _07229_;
  wire _07230_;
  wire _07231_;
  wire _07232_;
  wire _07233_;
  wire _07234_;
  wire _07235_;
  wire _07236_;
  wire _07237_;
  wire _07238_;
  wire _07239_;
  wire _07240_;
  wire _07241_;
  wire _07242_;
  wire _07243_;
  wire _07244_;
  wire _07245_;
  wire _07246_;
  wire _07247_;
  wire _07248_;
  wire _07249_;
  wire _07250_;
  wire _07251_;
  wire _07252_;
  wire _07253_;
  wire _07254_;
  wire _07255_;
  wire _07256_;
  wire _07257_;
  wire _07258_;
  wire _07259_;
  wire _07260_;
  wire _07261_;
  wire _07262_;
  wire _07263_;
  wire _07264_;
  wire _07265_;
  wire _07266_;
  wire _07267_;
  wire _07268_;
  wire _07269_;
  wire _07270_;
  wire _07271_;
  wire _07272_;
  wire _07273_;
  wire _07274_;
  wire _07275_;
  wire _07276_;
  wire _07277_;
  wire _07278_;
  wire _07279_;
  wire _07280_;
  wire _07281_;
  wire _07282_;
  wire _07283_;
  wire _07284_;
  wire _07285_;
  wire _07286_;
  wire _07287_;
  wire _07288_;
  wire _07289_;
  wire _07290_;
  wire _07291_;
  wire _07292_;
  wire _07293_;
  wire _07294_;
  wire _07295_;
  wire _07296_;
  wire _07297_;
  wire _07298_;
  wire _07299_;
  wire _07300_;
  wire _07301_;
  wire _07302_;
  wire _07303_;
  wire _07304_;
  wire _07305_;
  wire _07306_;
  wire _07307_;
  wire _07308_;
  wire _07309_;
  wire _07310_;
  wire _07311_;
  wire _07312_;
  wire _07313_;
  wire _07314_;
  wire _07315_;
  wire _07316_;
  wire _07317_;
  wire _07318_;
  wire _07319_;
  wire _07320_;
  wire _07321_;
  wire _07322_;
  wire _07323_;
  wire _07324_;
  wire _07325_;
  wire _07326_;
  wire _07327_;
  wire _07328_;
  wire _07329_;
  wire _07330_;
  wire _07331_;
  wire _07332_;
  wire _07333_;
  wire _07334_;
  wire _07335_;
  wire _07336_;
  wire _07337_;
  wire _07338_;
  wire _07339_;
  wire _07340_;
  wire _07341_;
  wire _07342_;
  wire _07343_;
  wire _07344_;
  wire _07345_;
  wire _07346_;
  wire _07347_;
  wire _07348_;
  wire _07349_;
  wire _07350_;
  wire _07351_;
  wire _07352_;
  wire _07353_;
  wire _07354_;
  wire _07355_;
  wire _07356_;
  wire _07357_;
  wire _07358_;
  wire _07359_;
  wire _07360_;
  wire _07361_;
  wire _07362_;
  wire _07363_;
  wire _07364_;
  wire _07365_;
  wire _07366_;
  wire _07367_;
  wire _07368_;
  wire _07369_;
  wire _07370_;
  wire _07371_;
  wire _07372_;
  wire _07373_;
  wire _07374_;
  wire _07375_;
  wire _07376_;
  wire _07377_;
  wire _07378_;
  wire _07379_;
  wire _07380_;
  wire _07381_;
  wire _07382_;
  wire _07383_;
  wire _07384_;
  wire _07385_;
  wire _07386_;
  wire _07387_;
  wire _07388_;
  wire _07389_;
  wire _07390_;
  wire _07391_;
  wire _07392_;
  wire _07393_;
  wire _07394_;
  wire _07395_;
  wire _07396_;
  wire _07397_;
  wire _07398_;
  wire _07399_;
  wire _07400_;
  wire _07401_;
  wire _07402_;
  wire _07403_;
  wire _07404_;
  wire _07405_;
  wire _07406_;
  wire _07407_;
  wire _07408_;
  wire _07409_;
  wire _07410_;
  wire _07411_;
  wire _07412_;
  wire _07413_;
  wire _07414_;
  wire _07415_;
  wire _07416_;
  wire _07417_;
  wire _07418_;
  wire _07419_;
  wire _07420_;
  wire _07421_;
  wire _07422_;
  wire _07423_;
  wire _07424_;
  wire _07425_;
  wire _07426_;
  wire _07427_;
  wire _07428_;
  wire _07429_;
  wire _07430_;
  wire _07431_;
  wire _07432_;
  wire _07433_;
  wire _07434_;
  wire _07435_;
  wire _07436_;
  wire _07437_;
  wire _07438_;
  wire _07439_;
  wire _07440_;
  wire _07441_;
  wire _07442_;
  wire _07443_;
  wire _07444_;
  wire _07445_;
  wire _07446_;
  wire _07447_;
  wire _07448_;
  wire _07449_;
  wire _07450_;
  wire _07451_;
  wire _07452_;
  wire _07453_;
  wire _07454_;
  wire _07455_;
  wire _07456_;
  wire _07457_;
  wire _07458_;
  wire _07459_;
  wire _07460_;
  wire _07461_;
  wire _07462_;
  wire _07463_;
  wire _07464_;
  wire _07465_;
  wire _07466_;
  wire _07467_;
  wire _07468_;
  wire _07469_;
  wire _07470_;
  wire _07471_;
  wire _07472_;
  wire _07473_;
  wire _07474_;
  wire _07475_;
  wire _07476_;
  wire _07477_;
  wire _07478_;
  wire _07479_;
  wire _07480_;
  wire _07481_;
  wire _07482_;
  wire _07483_;
  wire _07484_;
  wire _07485_;
  wire _07486_;
  wire _07487_;
  wire _07488_;
  wire _07489_;
  wire _07490_;
  wire _07491_;
  wire _07492_;
  wire _07493_;
  wire _07494_;
  wire _07495_;
  wire _07496_;
  wire _07497_;
  wire _07498_;
  wire _07499_;
  wire _07500_;
  wire _07501_;
  wire _07502_;
  wire _07503_;
  wire _07504_;
  wire _07505_;
  wire _07506_;
  wire _07507_;
  wire _07508_;
  wire _07509_;
  wire _07510_;
  wire _07511_;
  wire _07512_;
  wire _07513_;
  wire _07514_;
  wire _07515_;
  wire _07516_;
  wire _07517_;
  wire _07518_;
  wire _07519_;
  wire _07520_;
  wire _07521_;
  wire _07522_;
  wire _07523_;
  wire _07524_;
  wire _07525_;
  wire _07526_;
  wire _07527_;
  wire _07528_;
  wire _07529_;
  wire _07530_;
  wire _07531_;
  wire _07532_;
  wire _07533_;
  wire _07534_;
  wire _07535_;
  wire _07536_;
  wire _07537_;
  wire _07538_;
  wire _07539_;
  wire _07540_;
  wire _07541_;
  wire _07542_;
  wire _07543_;
  wire _07544_;
  wire _07545_;
  wire _07546_;
  wire _07547_;
  wire _07548_;
  wire _07549_;
  wire _07550_;
  wire _07551_;
  wire _07552_;
  wire _07553_;
  wire _07554_;
  wire _07555_;
  wire _07556_;
  wire _07557_;
  wire _07558_;
  wire _07559_;
  wire _07560_;
  wire _07561_;
  wire _07562_;
  wire _07563_;
  wire _07564_;
  wire _07565_;
  wire _07566_;
  wire _07567_;
  wire _07568_;
  wire _07569_;
  wire _07570_;
  wire _07571_;
  wire _07572_;
  wire _07573_;
  wire _07574_;
  wire _07575_;
  wire _07576_;
  wire _07577_;
  wire _07578_;
  wire _07579_;
  wire _07580_;
  wire _07581_;
  wire _07582_;
  wire _07583_;
  wire _07584_;
  wire _07585_;
  wire _07586_;
  wire _07587_;
  wire _07588_;
  wire _07589_;
  wire _07590_;
  wire _07591_;
  wire _07592_;
  wire _07593_;
  wire _07594_;
  wire _07595_;
  wire _07596_;
  wire _07597_;
  wire _07598_;
  wire _07599_;
  wire _07600_;
  wire _07601_;
  wire _07602_;
  wire _07603_;
  wire _07604_;
  wire _07605_;
  wire _07606_;
  wire _07607_;
  wire _07608_;
  wire _07609_;
  wire _07610_;
  wire _07611_;
  wire _07612_;
  wire _07613_;
  wire _07614_;
  wire _07615_;
  wire _07616_;
  wire _07617_;
  wire _07618_;
  wire _07619_;
  wire _07620_;
  wire _07621_;
  wire _07622_;
  wire _07623_;
  wire _07624_;
  wire _07625_;
  wire _07626_;
  wire _07627_;
  wire _07628_;
  wire _07629_;
  wire _07630_;
  wire _07631_;
  wire _07632_;
  wire _07633_;
  wire _07634_;
  wire _07635_;
  wire _07636_;
  wire _07637_;
  wire _07638_;
  wire _07639_;
  wire _07640_;
  wire _07641_;
  wire _07642_;
  wire _07643_;
  wire _07644_;
  wire _07645_;
  wire _07646_;
  wire _07647_;
  wire _07648_;
  wire _07649_;
  wire _07650_;
  wire _07651_;
  wire _07652_;
  wire _07653_;
  wire _07654_;
  wire _07655_;
  wire _07656_;
  wire _07657_;
  wire _07658_;
  wire _07659_;
  wire _07660_;
  wire _07661_;
  wire _07662_;
  wire _07663_;
  wire _07664_;
  wire _07665_;
  wire _07666_;
  wire _07667_;
  wire _07668_;
  wire _07669_;
  wire _07670_;
  wire _07671_;
  wire _07672_;
  wire _07673_;
  wire _07674_;
  wire _07675_;
  wire _07676_;
  wire _07677_;
  wire _07678_;
  wire _07679_;
  wire _07680_;
  wire _07681_;
  wire _07682_;
  wire _07683_;
  wire _07684_;
  wire _07685_;
  wire _07686_;
  wire _07687_;
  wire _07688_;
  wire _07689_;
  wire _07690_;
  wire _07691_;
  wire _07692_;
  wire _07693_;
  wire _07694_;
  wire _07695_;
  wire _07696_;
  wire _07697_;
  wire _07698_;
  wire _07699_;
  wire _07700_;
  wire _07701_;
  wire _07702_;
  wire _07703_;
  wire _07704_;
  wire _07705_;
  wire _07706_;
  wire _07707_;
  wire _07708_;
  wire _07709_;
  wire _07710_;
  wire _07711_;
  wire _07712_;
  wire _07713_;
  wire _07714_;
  wire _07715_;
  wire _07716_;
  wire _07717_;
  wire _07718_;
  wire _07719_;
  wire _07720_;
  wire _07721_;
  wire _07722_;
  wire _07723_;
  wire _07724_;
  wire _07725_;
  wire _07726_;
  wire _07727_;
  wire _07728_;
  wire _07729_;
  wire _07730_;
  wire _07731_;
  wire _07732_;
  wire _07733_;
  wire _07734_;
  wire _07735_;
  wire _07736_;
  wire _07737_;
  wire _07738_;
  wire _07739_;
  wire _07740_;
  wire _07741_;
  wire _07742_;
  wire _07743_;
  wire _07744_;
  wire _07745_;
  wire _07746_;
  wire _07747_;
  wire _07748_;
  wire _07749_;
  wire _07750_;
  wire _07751_;
  wire _07752_;
  wire _07753_;
  wire _07754_;
  wire _07755_;
  wire _07756_;
  wire _07757_;
  wire _07758_;
  wire _07759_;
  wire _07760_;
  wire _07761_;
  wire _07762_;
  wire _07763_;
  wire _07764_;
  wire _07765_;
  wire _07766_;
  wire _07767_;
  wire _07768_;
  wire _07769_;
  wire _07770_;
  wire _07771_;
  wire _07772_;
  wire _07773_;
  wire _07774_;
  wire _07775_;
  wire _07776_;
  wire _07777_;
  wire _07778_;
  wire _07779_;
  wire _07780_;
  wire _07781_;
  wire _07782_;
  wire _07783_;
  wire _07784_;
  wire _07785_;
  wire _07786_;
  wire _07787_;
  wire _07788_;
  wire _07789_;
  wire _07790_;
  wire _07791_;
  wire _07792_;
  wire _07793_;
  wire _07794_;
  wire _07795_;
  wire _07796_;
  wire _07797_;
  wire _07798_;
  wire _07799_;
  wire _07800_;
  wire _07801_;
  wire _07802_;
  wire _07803_;
  wire _07804_;
  wire _07805_;
  wire _07806_;
  wire _07807_;
  wire _07808_;
  wire _07809_;
  wire _07810_;
  wire _07811_;
  wire _07812_;
  wire _07813_;
  wire _07814_;
  wire _07815_;
  wire _07816_;
  wire _07817_;
  wire _07818_;
  wire _07819_;
  wire _07820_;
  wire _07821_;
  wire _07822_;
  wire _07823_;
  wire _07824_;
  wire _07825_;
  wire _07826_;
  wire _07827_;
  wire _07828_;
  wire _07829_;
  wire _07830_;
  wire _07831_;
  wire _07832_;
  wire _07833_;
  wire _07834_;
  wire _07835_;
  wire _07836_;
  wire _07837_;
  wire _07838_;
  wire _07839_;
  wire _07840_;
  wire _07841_;
  wire _07842_;
  wire _07843_;
  wire _07844_;
  wire _07845_;
  wire _07846_;
  wire _07847_;
  wire _07848_;
  wire _07849_;
  wire _07850_;
  wire _07851_;
  wire _07852_;
  wire _07853_;
  wire _07854_;
  wire _07855_;
  wire _07856_;
  wire _07857_;
  wire _07858_;
  wire _07859_;
  wire _07860_;
  wire _07861_;
  wire _07862_;
  wire _07863_;
  wire _07864_;
  wire _07865_;
  wire _07866_;
  wire _07867_;
  wire _07868_;
  wire _07869_;
  wire _07870_;
  wire _07871_;
  wire _07872_;
  wire _07873_;
  wire _07874_;
  wire _07875_;
  wire _07876_;
  wire _07877_;
  wire _07878_;
  wire _07879_;
  wire _07880_;
  wire _07881_;
  wire _07882_;
  wire _07883_;
  wire _07884_;
  wire _07885_;
  wire _07886_;
  wire _07887_;
  wire _07888_;
  wire _07889_;
  wire _07890_;
  wire _07891_;
  wire _07892_;
  wire _07893_;
  wire _07894_;
  wire _07895_;
  wire _07896_;
  wire _07897_;
  wire _07898_;
  wire _07899_;
  wire _07900_;
  wire _07901_;
  wire _07902_;
  wire _07903_;
  wire _07904_;
  wire _07905_;
  wire _07906_;
  wire _07907_;
  wire _07908_;
  wire _07909_;
  wire _07910_;
  wire _07911_;
  wire _07912_;
  wire _07913_;
  wire _07914_;
  wire _07915_;
  wire _07916_;
  wire _07917_;
  wire _07918_;
  wire _07919_;
  wire _07920_;
  wire _07921_;
  wire _07922_;
  wire _07923_;
  wire _07924_;
  wire _07925_;
  wire _07926_;
  wire _07927_;
  wire _07928_;
  wire _07929_;
  wire _07930_;
  wire _07931_;
  wire _07932_;
  wire _07933_;
  wire _07934_;
  wire _07935_;
  wire _07936_;
  wire _07937_;
  wire _07938_;
  wire _07939_;
  wire _07940_;
  wire _07941_;
  wire _07942_;
  wire _07943_;
  wire _07944_;
  wire _07945_;
  wire _07946_;
  wire _07947_;
  wire _07948_;
  wire _07949_;
  wire _07950_;
  wire _07951_;
  wire _07952_;
  wire _07953_;
  wire _07954_;
  wire _07955_;
  wire _07956_;
  wire _07957_;
  wire _07958_;
  wire _07959_;
  wire _07960_;
  wire _07961_;
  wire _07962_;
  wire _07963_;
  wire _07964_;
  wire _07965_;
  wire _07966_;
  wire _07967_;
  wire _07968_;
  wire _07969_;
  wire _07970_;
  wire _07971_;
  wire _07972_;
  wire _07973_;
  wire _07974_;
  wire _07975_;
  wire _07976_;
  wire _07977_;
  wire _07978_;
  wire _07979_;
  wire _07980_;
  wire _07981_;
  wire _07982_;
  wire _07983_;
  wire _07984_;
  wire _07985_;
  wire _07986_;
  wire _07987_;
  wire _07988_;
  wire _07989_;
  wire _07990_;
  wire _07991_;
  wire _07992_;
  wire _07993_;
  wire _07994_;
  wire _07995_;
  wire _07996_;
  wire _07997_;
  wire _07998_;
  wire _07999_;
  wire _08000_;
  wire _08001_;
  wire _08002_;
  wire _08003_;
  wire _08004_;
  wire _08005_;
  wire _08006_;
  wire _08007_;
  wire _08008_;
  wire _08009_;
  wire _08010_;
  wire _08011_;
  wire _08012_;
  wire _08013_;
  wire _08014_;
  wire _08015_;
  wire _08016_;
  wire _08017_;
  wire _08018_;
  wire _08019_;
  wire _08020_;
  wire _08021_;
  wire _08022_;
  wire _08023_;
  wire _08024_;
  wire _08025_;
  wire _08026_;
  wire _08027_;
  wire _08028_;
  wire _08029_;
  wire _08030_;
  wire _08031_;
  wire _08032_;
  wire _08033_;
  wire _08034_;
  wire _08035_;
  wire _08036_;
  wire _08037_;
  wire _08038_;
  wire _08039_;
  wire _08040_;
  wire _08041_;
  wire _08042_;
  wire _08043_;
  wire _08044_;
  wire _08045_;
  wire _08046_;
  wire _08047_;
  wire _08048_;
  wire _08049_;
  wire _08050_;
  wire _08051_;
  wire _08052_;
  wire _08053_;
  wire _08054_;
  wire _08055_;
  wire _08056_;
  wire _08057_;
  wire _08058_;
  wire _08059_;
  wire _08060_;
  wire _08061_;
  wire _08062_;
  wire _08063_;
  wire _08064_;
  wire _08065_;
  wire _08066_;
  wire _08067_;
  wire _08068_;
  wire _08069_;
  wire _08070_;
  wire _08071_;
  wire _08072_;
  wire _08073_;
  wire _08074_;
  wire _08075_;
  wire _08076_;
  wire _08077_;
  wire _08078_;
  wire _08079_;
  wire _08080_;
  wire _08081_;
  wire _08082_;
  wire _08083_;
  wire _08084_;
  wire _08085_;
  wire _08086_;
  wire _08087_;
  wire _08088_;
  wire _08089_;
  wire _08090_;
  wire _08091_;
  wire _08092_;
  wire _08093_;
  wire _08094_;
  wire _08095_;
  wire _08096_;
  wire _08097_;
  wire _08098_;
  wire _08099_;
  wire _08100_;
  wire _08101_;
  wire _08102_;
  wire _08103_;
  wire _08104_;
  wire _08105_;
  wire _08106_;
  wire _08107_;
  wire _08108_;
  wire _08109_;
  wire _08110_;
  wire _08111_;
  wire _08112_;
  wire _08113_;
  wire _08114_;
  wire _08115_;
  wire _08116_;
  wire _08117_;
  wire _08118_;
  wire _08119_;
  wire _08120_;
  wire _08121_;
  wire _08122_;
  wire _08123_;
  wire _08124_;
  wire _08125_;
  wire _08126_;
  wire _08127_;
  wire _08128_;
  wire _08129_;
  wire _08130_;
  wire _08131_;
  wire _08132_;
  wire _08133_;
  wire _08134_;
  wire _08135_;
  wire _08136_;
  wire _08137_;
  wire _08138_;
  wire _08139_;
  wire _08140_;
  wire _08141_;
  wire _08142_;
  wire _08143_;
  wire _08144_;
  wire _08145_;
  wire _08146_;
  wire _08147_;
  wire _08148_;
  wire _08149_;
  wire _08150_;
  wire _08151_;
  wire _08152_;
  wire _08153_;
  wire _08154_;
  wire _08155_;
  wire _08156_;
  wire _08157_;
  wire _08158_;
  wire _08159_;
  wire _08160_;
  wire _08161_;
  wire _08162_;
  wire _08163_;
  wire _08164_;
  wire _08165_;
  wire _08166_;
  wire _08167_;
  wire _08168_;
  wire _08169_;
  wire _08170_;
  wire _08171_;
  wire _08172_;
  wire _08173_;
  wire _08174_;
  wire _08175_;
  wire _08176_;
  wire _08177_;
  wire _08178_;
  wire _08179_;
  wire _08180_;
  wire _08181_;
  wire _08182_;
  wire _08183_;
  wire _08184_;
  wire _08185_;
  wire _08186_;
  wire _08187_;
  wire _08188_;
  wire _08189_;
  wire _08190_;
  wire _08191_;
  wire _08192_;
  wire _08193_;
  wire _08194_;
  wire _08195_;
  wire _08196_;
  wire _08197_;
  wire _08198_;
  wire _08199_;
  wire _08200_;
  wire _08201_;
  wire _08202_;
  wire _08203_;
  wire _08204_;
  wire _08205_;
  wire _08206_;
  wire _08207_;
  wire _08208_;
  wire _08209_;
  wire _08210_;
  wire _08211_;
  wire _08212_;
  wire _08213_;
  wire _08214_;
  wire _08215_;
  wire _08216_;
  wire _08217_;
  wire _08218_;
  wire _08219_;
  wire _08220_;
  wire _08221_;
  wire _08222_;
  wire _08223_;
  wire _08224_;
  wire _08225_;
  wire _08226_;
  wire _08227_;
  wire _08228_;
  wire _08229_;
  wire _08230_;
  wire _08231_;
  wire _08232_;
  wire _08233_;
  wire _08234_;
  wire _08235_;
  wire _08236_;
  wire _08237_;
  wire _08238_;
  wire _08239_;
  wire _08240_;
  wire _08241_;
  wire _08242_;
  wire _08243_;
  wire _08244_;
  wire _08245_;
  wire _08246_;
  wire _08247_;
  wire _08248_;
  wire _08249_;
  wire _08250_;
  wire _08251_;
  wire _08252_;
  wire _08253_;
  wire _08254_;
  wire _08255_;
  wire _08256_;
  wire _08257_;
  wire _08258_;
  wire _08259_;
  wire _08260_;
  wire _08261_;
  wire _08262_;
  wire _08263_;
  wire _08264_;
  wire _08265_;
  wire _08266_;
  wire _08267_;
  wire _08268_;
  wire _08269_;
  wire _08270_;
  wire _08271_;
  wire _08272_;
  wire _08273_;
  wire _08274_;
  wire _08275_;
  wire _08276_;
  wire _08277_;
  wire _08278_;
  wire _08279_;
  wire _08280_;
  wire _08281_;
  wire _08282_;
  wire _08283_;
  wire _08284_;
  wire _08285_;
  wire _08286_;
  wire _08287_;
  wire _08288_;
  wire _08289_;
  wire _08290_;
  wire _08291_;
  wire _08292_;
  wire _08293_;
  wire _08294_;
  wire _08295_;
  wire _08296_;
  wire _08297_;
  wire _08298_;
  wire _08299_;
  wire _08300_;
  wire _08301_;
  wire _08302_;
  wire _08303_;
  wire _08304_;
  wire _08305_;
  wire _08306_;
  wire _08307_;
  wire _08308_;
  wire _08309_;
  wire _08310_;
  wire _08311_;
  wire _08312_;
  wire _08313_;
  wire _08314_;
  wire _08315_;
  wire _08316_;
  wire _08317_;
  wire _08318_;
  wire _08319_;
  wire _08320_;
  wire _08321_;
  wire _08322_;
  wire _08323_;
  wire _08324_;
  wire _08325_;
  wire _08326_;
  wire _08327_;
  wire _08328_;
  wire _08329_;
  wire _08330_;
  wire _08331_;
  wire _08332_;
  wire _08333_;
  wire _08334_;
  wire _08335_;
  wire _08336_;
  wire _08337_;
  wire _08338_;
  wire _08339_;
  wire _08340_;
  wire _08341_;
  wire _08342_;
  wire _08343_;
  wire _08344_;
  wire _08345_;
  wire _08346_;
  wire _08347_;
  wire _08348_;
  wire _08349_;
  wire _08350_;
  wire _08351_;
  wire _08352_;
  wire _08353_;
  wire _08354_;
  wire _08355_;
  wire _08356_;
  wire _08357_;
  wire _08358_;
  wire _08359_;
  wire _08360_;
  wire _08361_;
  wire _08362_;
  wire _08363_;
  wire _08364_;
  wire _08365_;
  wire _08366_;
  wire _08367_;
  wire _08368_;
  wire _08369_;
  wire _08370_;
  wire _08371_;
  wire _08372_;
  wire _08373_;
  wire _08374_;
  wire _08375_;
  wire _08376_;
  wire _08377_;
  wire _08378_;
  wire _08379_;
  wire _08380_;
  wire _08381_;
  wire _08382_;
  wire _08383_;
  wire _08384_;
  wire _08385_;
  wire _08386_;
  wire _08387_;
  wire _08388_;
  wire _08389_;
  wire _08390_;
  wire _08391_;
  wire _08392_;
  wire _08393_;
  wire _08394_;
  wire _08395_;
  wire _08396_;
  wire _08397_;
  wire _08398_;
  wire _08399_;
  wire _08400_;
  wire _08401_;
  wire _08402_;
  wire _08403_;
  wire _08404_;
  wire _08405_;
  wire _08406_;
  wire _08407_;
  wire _08408_;
  wire _08409_;
  wire _08410_;
  wire _08411_;
  wire _08412_;
  wire _08413_;
  wire _08414_;
  wire _08415_;
  wire _08416_;
  wire _08417_;
  wire _08418_;
  wire _08419_;
  wire _08420_;
  wire _08421_;
  wire _08422_;
  wire _08423_;
  wire _08424_;
  wire _08425_;
  wire _08426_;
  wire _08427_;
  wire _08428_;
  wire _08429_;
  wire _08430_;
  wire _08431_;
  wire _08432_;
  wire _08433_;
  wire _08434_;
  wire _08435_;
  wire _08436_;
  wire _08437_;
  wire _08438_;
  wire _08439_;
  wire _08440_;
  wire _08441_;
  wire _08442_;
  wire _08443_;
  wire _08444_;
  wire _08445_;
  wire _08446_;
  wire _08447_;
  wire _08448_;
  wire _08449_;
  wire _08450_;
  wire _08451_;
  wire _08452_;
  wire _08453_;
  wire _08454_;
  wire _08455_;
  wire _08456_;
  wire _08457_;
  wire _08458_;
  wire _08459_;
  wire _08460_;
  wire _08461_;
  wire _08462_;
  wire _08463_;
  wire _08464_;
  wire _08465_;
  wire _08466_;
  wire _08467_;
  wire _08468_;
  wire _08469_;
  wire _08470_;
  wire _08471_;
  wire _08472_;
  wire _08473_;
  wire _08474_;
  wire _08475_;
  wire _08476_;
  wire _08477_;
  wire _08478_;
  wire _08479_;
  wire _08480_;
  wire _08481_;
  wire _08482_;
  wire _08483_;
  wire _08484_;
  wire _08485_;
  wire _08486_;
  wire _08487_;
  wire _08488_;
  wire _08489_;
  wire _08490_;
  wire _08491_;
  wire _08492_;
  wire _08493_;
  wire _08494_;
  wire _08495_;
  wire _08496_;
  wire _08497_;
  wire _08498_;
  wire _08499_;
  wire _08500_;
  wire _08501_;
  wire _08502_;
  wire _08503_;
  wire _08504_;
  wire _08505_;
  wire _08506_;
  wire _08507_;
  wire _08508_;
  wire _08509_;
  wire _08510_;
  wire _08511_;
  wire _08512_;
  wire _08513_;
  wire _08514_;
  wire _08515_;
  wire _08516_;
  wire _08517_;
  wire _08518_;
  wire _08519_;
  wire _08520_;
  wire _08521_;
  wire _08522_;
  wire _08523_;
  wire _08524_;
  wire _08525_;
  wire _08526_;
  wire _08527_;
  wire _08528_;
  wire _08529_;
  wire _08530_;
  wire _08531_;
  wire _08532_;
  wire _08533_;
  wire _08534_;
  wire _08535_;
  wire _08536_;
  wire _08537_;
  wire _08538_;
  wire _08539_;
  wire _08540_;
  wire _08541_;
  wire _08542_;
  wire _08543_;
  wire _08544_;
  wire _08545_;
  wire _08546_;
  wire _08547_;
  wire _08548_;
  wire _08549_;
  wire _08550_;
  wire _08551_;
  wire _08552_;
  wire _08553_;
  wire _08554_;
  wire _08555_;
  wire _08556_;
  wire _08557_;
  wire _08558_;
  wire _08559_;
  wire _08560_;
  wire _08561_;
  wire _08562_;
  wire _08563_;
  wire _08564_;
  wire _08565_;
  wire _08566_;
  wire _08567_;
  wire _08568_;
  wire _08569_;
  wire _08570_;
  wire _08571_;
  wire _08572_;
  wire _08573_;
  wire _08574_;
  wire _08575_;
  wire _08576_;
  wire _08577_;
  wire _08578_;
  wire _08579_;
  wire _08580_;
  wire _08581_;
  wire _08582_;
  wire _08583_;
  wire _08584_;
  wire _08585_;
  wire _08586_;
  wire _08587_;
  wire _08588_;
  wire _08589_;
  wire _08590_;
  wire _08591_;
  wire _08592_;
  wire _08593_;
  wire _08594_;
  wire _08595_;
  wire _08596_;
  wire _08597_;
  wire _08598_;
  wire _08599_;
  wire _08600_;
  wire _08601_;
  wire _08602_;
  wire _08603_;
  wire _08604_;
  wire _08605_;
  wire _08606_;
  wire _08607_;
  wire _08608_;
  wire _08609_;
  wire _08610_;
  wire _08611_;
  wire _08612_;
  wire _08613_;
  wire _08614_;
  wire _08615_;
  wire _08616_;
  wire _08617_;
  wire _08618_;
  wire _08619_;
  wire _08620_;
  wire _08621_;
  wire _08622_;
  wire _08623_;
  wire _08624_;
  wire _08625_;
  wire _08626_;
  wire _08627_;
  wire _08628_;
  wire _08629_;
  wire _08630_;
  wire _08631_;
  wire _08632_;
  wire _08633_;
  wire _08634_;
  wire _08635_;
  wire _08636_;
  wire _08637_;
  wire _08638_;
  wire _08639_;
  wire _08640_;
  wire _08641_;
  wire _08642_;
  wire _08643_;
  wire _08644_;
  wire _08645_;
  wire _08646_;
  wire _08647_;
  wire _08648_;
  wire _08649_;
  wire _08650_;
  wire _08651_;
  wire _08652_;
  wire _08653_;
  wire _08654_;
  wire _08655_;
  wire _08656_;
  wire _08657_;
  wire _08658_;
  wire _08659_;
  wire _08660_;
  wire _08661_;
  wire _08662_;
  wire _08663_;
  wire _08664_;
  wire _08665_;
  wire _08666_;
  wire _08667_;
  wire _08668_;
  wire _08669_;
  wire _08670_;
  wire _08671_;
  wire _08672_;
  wire _08673_;
  wire _08674_;
  wire _08675_;
  wire _08676_;
  wire _08677_;
  wire _08678_;
  wire _08679_;
  wire _08680_;
  wire _08681_;
  wire _08682_;
  wire _08683_;
  wire _08684_;
  wire _08685_;
  wire _08686_;
  wire _08687_;
  wire _08688_;
  wire _08689_;
  wire _08690_;
  wire _08691_;
  wire _08692_;
  wire _08693_;
  wire _08694_;
  wire _08695_;
  wire _08696_;
  wire _08697_;
  wire _08698_;
  wire _08699_;
  wire _08700_;
  wire _08701_;
  wire _08702_;
  wire _08703_;
  wire _08704_;
  wire _08705_;
  wire _08706_;
  wire _08707_;
  wire _08708_;
  wire _08709_;
  wire _08710_;
  wire _08711_;
  wire _08712_;
  wire _08713_;
  wire _08714_;
  wire _08715_;
  wire _08716_;
  wire _08717_;
  wire _08718_;
  wire _08719_;
  wire _08720_;
  wire _08721_;
  wire _08722_;
  wire _08723_;
  wire _08724_;
  wire _08725_;
  wire _08726_;
  wire _08727_;
  wire _08728_;
  wire _08729_;
  wire _08730_;
  wire _08731_;
  wire _08732_;
  wire _08733_;
  wire _08734_;
  wire _08735_;
  wire _08736_;
  wire _08737_;
  wire _08738_;
  wire _08739_;
  wire _08740_;
  wire _08741_;
  wire _08742_;
  wire _08743_;
  wire _08744_;
  wire _08745_;
  wire _08746_;
  wire _08747_;
  wire _08748_;
  wire _08749_;
  wire _08750_;
  wire _08751_;
  wire _08752_;
  wire _08753_;
  wire _08754_;
  wire _08755_;
  wire _08756_;
  wire _08757_;
  wire _08758_;
  wire _08759_;
  wire _08760_;
  wire _08761_;
  wire _08762_;
  wire _08763_;
  wire _08764_;
  wire _08765_;
  wire _08766_;
  wire _08767_;
  wire _08768_;
  wire _08769_;
  wire _08770_;
  wire _08771_;
  wire _08772_;
  wire _08773_;
  wire _08774_;
  wire _08775_;
  wire _08776_;
  wire _08777_;
  wire _08778_;
  wire _08779_;
  wire _08780_;
  wire _08781_;
  wire _08782_;
  wire _08783_;
  wire _08784_;
  wire _08785_;
  wire _08786_;
  wire _08787_;
  wire _08788_;
  wire _08789_;
  wire _08790_;
  wire _08791_;
  wire _08792_;
  wire _08793_;
  wire _08794_;
  wire _08795_;
  wire _08796_;
  wire _08797_;
  wire _08798_;
  wire _08799_;
  wire _08800_;
  wire _08801_;
  wire _08802_;
  wire _08803_;
  wire _08804_;
  wire _08805_;
  wire _08806_;
  wire _08807_;
  wire _08808_;
  wire _08809_;
  wire _08810_;
  wire _08811_;
  wire _08812_;
  wire _08813_;
  wire _08814_;
  wire _08815_;
  wire _08816_;
  wire _08817_;
  wire _08818_;
  wire _08819_;
  wire _08820_;
  wire _08821_;
  wire _08822_;
  wire _08823_;
  wire _08824_;
  wire _08825_;
  wire _08826_;
  wire _08827_;
  wire _08828_;
  wire _08829_;
  wire _08830_;
  wire _08831_;
  wire _08832_;
  wire _08833_;
  wire _08834_;
  wire _08835_;
  wire _08836_;
  wire _08837_;
  wire _08838_;
  wire _08839_;
  wire _08840_;
  wire _08841_;
  wire _08842_;
  wire _08843_;
  wire _08844_;
  wire _08845_;
  wire _08846_;
  wire _08847_;
  wire _08848_;
  wire _08849_;
  wire _08850_;
  wire _08851_;
  wire _08852_;
  wire _08853_;
  wire _08854_;
  wire _08855_;
  wire _08856_;
  wire _08857_;
  wire _08858_;
  wire _08859_;
  wire _08860_;
  wire _08861_;
  wire _08862_;
  wire _08863_;
  wire _08864_;
  wire _08865_;
  wire _08866_;
  wire _08867_;
  wire _08868_;
  wire _08869_;
  wire _08870_;
  wire _08871_;
  wire _08872_;
  wire _08873_;
  wire _08874_;
  wire _08875_;
  wire _08876_;
  wire _08877_;
  wire _08878_;
  wire _08879_;
  wire _08880_;
  wire _08881_;
  wire _08882_;
  wire _08883_;
  wire _08884_;
  wire _08885_;
  wire _08886_;
  wire _08887_;
  wire _08888_;
  wire _08889_;
  wire _08890_;
  wire _08891_;
  wire _08892_;
  wire _08893_;
  wire _08894_;
  wire _08895_;
  wire _08896_;
  wire _08897_;
  wire _08898_;
  wire _08899_;
  wire _08900_;
  wire _08901_;
  wire _08902_;
  wire _08903_;
  wire _08904_;
  wire _08905_;
  wire _08906_;
  wire _08907_;
  wire _08908_;
  wire _08909_;
  wire _08910_;
  wire _08911_;
  wire _08912_;
  wire _08913_;
  wire _08914_;
  wire _08915_;
  wire _08916_;
  wire _08917_;
  wire _08918_;
  wire _08919_;
  wire _08920_;
  wire _08921_;
  wire _08922_;
  wire _08923_;
  wire _08924_;
  wire _08925_;
  wire _08926_;
  wire _08927_;
  wire _08928_;
  wire _08929_;
  wire _08930_;
  wire _08931_;
  wire _08932_;
  wire _08933_;
  wire _08934_;
  wire _08935_;
  wire _08936_;
  wire _08937_;
  wire _08938_;
  wire _08939_;
  wire _08940_;
  wire _08941_;
  wire _08942_;
  wire _08943_;
  wire _08944_;
  wire _08945_;
  wire _08946_;
  wire _08947_;
  wire _08948_;
  wire _08949_;
  wire _08950_;
  wire _08951_;
  wire _08952_;
  wire _08953_;
  wire _08954_;
  wire _08955_;
  wire _08956_;
  wire _08957_;
  wire _08958_;
  wire _08959_;
  wire _08960_;
  wire _08961_;
  wire _08962_;
  wire _08963_;
  wire _08964_;
  wire _08965_;
  wire _08966_;
  wire _08967_;
  wire _08968_;
  wire _08969_;
  wire _08970_;
  wire _08971_;
  wire _08972_;
  wire _08973_;
  wire _08974_;
  wire _08975_;
  wire _08976_;
  wire _08977_;
  wire _08978_;
  wire _08979_;
  wire _08980_;
  wire _08981_;
  wire _08982_;
  wire _08983_;
  wire _08984_;
  wire _08985_;
  wire _08986_;
  wire _08987_;
  wire _08988_;
  wire _08989_;
  wire _08990_;
  wire _08991_;
  wire _08992_;
  wire _08993_;
  wire _08994_;
  wire _08995_;
  wire _08996_;
  wire _08997_;
  wire _08998_;
  wire _08999_;
  wire _09000_;
  wire _09001_;
  wire _09002_;
  wire _09003_;
  wire _09004_;
  wire _09005_;
  wire _09006_;
  wire _09007_;
  wire _09008_;
  wire _09009_;
  wire _09010_;
  wire _09011_;
  wire _09012_;
  wire _09013_;
  wire _09014_;
  wire _09015_;
  wire _09016_;
  wire _09017_;
  wire _09018_;
  wire _09019_;
  wire _09020_;
  wire _09021_;
  wire _09022_;
  wire _09023_;
  wire _09024_;
  wire _09025_;
  wire _09026_;
  wire _09027_;
  wire _09028_;
  wire _09029_;
  wire _09030_;
  wire _09031_;
  wire _09032_;
  wire _09033_;
  wire _09034_;
  wire _09035_;
  wire _09036_;
  wire _09037_;
  wire _09038_;
  wire _09039_;
  wire _09040_;
  wire _09041_;
  wire _09042_;
  wire _09043_;
  wire _09044_;
  wire _09045_;
  wire _09046_;
  wire _09047_;
  wire _09048_;
  wire _09049_;
  wire _09050_;
  wire _09051_;
  wire _09052_;
  wire _09053_;
  wire _09054_;
  wire _09055_;
  wire _09056_;
  wire _09057_;
  wire _09058_;
  wire _09059_;
  wire _09060_;
  wire _09061_;
  wire _09062_;
  wire _09063_;
  wire _09064_;
  wire _09065_;
  wire _09066_;
  wire _09067_;
  wire _09068_;
  wire _09069_;
  wire _09070_;
  wire _09071_;
  wire _09072_;
  wire _09073_;
  wire _09074_;
  wire _09075_;
  wire _09076_;
  wire _09077_;
  wire _09078_;
  wire _09079_;
  wire _09080_;
  wire _09081_;
  wire _09082_;
  wire _09083_;
  wire _09084_;
  wire _09085_;
  wire _09086_;
  wire _09087_;
  wire _09088_;
  wire _09089_;
  wire _09090_;
  wire _09091_;
  wire _09092_;
  wire _09093_;
  wire _09094_;
  wire _09095_;
  wire _09096_;
  wire _09097_;
  wire _09098_;
  wire _09099_;
  wire _09100_;
  wire _09101_;
  wire _09102_;
  wire _09103_;
  wire _09104_;
  wire _09105_;
  wire _09106_;
  wire _09107_;
  wire _09108_;
  wire _09109_;
  wire _09110_;
  wire _09111_;
  wire _09112_;
  wire _09113_;
  wire _09114_;
  wire _09115_;
  wire _09116_;
  wire _09117_;
  wire _09118_;
  wire _09119_;
  wire _09120_;
  wire _09121_;
  wire _09122_;
  wire _09123_;
  wire _09124_;
  wire _09125_;
  wire _09126_;
  wire _09127_;
  wire _09128_;
  wire _09129_;
  wire _09130_;
  wire _09131_;
  wire _09132_;
  wire _09133_;
  wire _09134_;
  wire _09135_;
  wire _09136_;
  wire _09137_;
  wire _09138_;
  wire _09139_;
  wire _09140_;
  wire _09141_;
  wire _09142_;
  wire _09143_;
  wire _09144_;
  wire _09145_;
  wire _09146_;
  wire _09147_;
  wire _09148_;
  wire _09149_;
  wire _09150_;
  wire _09151_;
  wire _09152_;
  wire _09153_;
  wire _09154_;
  wire _09155_;
  wire _09156_;
  wire _09157_;
  wire _09158_;
  wire _09159_;
  wire _09160_;
  wire _09161_;
  wire _09162_;
  wire _09163_;
  wire _09164_;
  wire _09165_;
  wire _09166_;
  wire _09167_;
  wire _09168_;
  wire _09169_;
  wire _09170_;
  wire _09171_;
  wire _09172_;
  wire _09173_;
  wire _09174_;
  wire _09175_;
  wire _09176_;
  wire _09177_;
  wire _09178_;
  wire _09179_;
  wire _09180_;
  wire _09181_;
  wire _09182_;
  wire _09183_;
  wire _09184_;
  wire _09185_;
  wire _09186_;
  wire _09187_;
  wire _09188_;
  wire _09189_;
  wire _09190_;
  wire _09191_;
  wire _09192_;
  wire _09193_;
  wire _09194_;
  wire _09195_;
  wire _09196_;
  wire _09197_;
  wire _09198_;
  wire _09199_;
  wire _09200_;
  wire _09201_;
  wire _09202_;
  wire _09203_;
  wire _09204_;
  wire _09205_;
  wire _09206_;
  wire _09207_;
  wire _09208_;
  wire _09209_;
  wire _09210_;
  wire _09211_;
  wire _09212_;
  wire _09213_;
  wire _09214_;
  wire _09215_;
  wire _09216_;
  wire _09217_;
  wire _09218_;
  wire _09219_;
  wire _09220_;
  wire _09221_;
  wire _09222_;
  wire _09223_;
  wire _09224_;
  wire _09225_;
  wire _09226_;
  wire _09227_;
  wire _09228_;
  wire _09229_;
  wire _09230_;
  wire _09231_;
  wire _09232_;
  wire _09233_;
  wire _09234_;
  wire _09235_;
  wire _09236_;
  wire _09237_;
  wire _09238_;
  wire _09239_;
  wire _09240_;
  wire _09241_;
  wire _09242_;
  wire _09243_;
  wire _09244_;
  wire _09245_;
  wire _09246_;
  wire _09247_;
  wire _09248_;
  wire _09249_;
  wire _09250_;
  wire _09251_;
  wire _09252_;
  wire _09253_;
  wire _09254_;
  wire _09255_;
  wire _09256_;
  wire _09257_;
  wire _09258_;
  wire _09259_;
  wire _09260_;
  wire _09261_;
  wire _09262_;
  wire _09263_;
  wire _09264_;
  wire _09265_;
  wire _09266_;
  wire _09267_;
  wire _09268_;
  wire _09269_;
  wire _09270_;
  wire _09271_;
  wire _09272_;
  wire _09273_;
  wire _09274_;
  wire _09275_;
  wire _09276_;
  wire _09277_;
  wire _09278_;
  wire _09279_;
  wire _09280_;
  wire _09281_;
  wire _09282_;
  wire _09283_;
  wire _09284_;
  wire _09285_;
  wire _09286_;
  wire _09287_;
  wire _09288_;
  wire _09289_;
  wire _09290_;
  wire _09291_;
  wire _09292_;
  wire _09293_;
  wire _09294_;
  wire _09295_;
  wire _09296_;
  wire _09297_;
  wire _09298_;
  wire _09299_;
  wire _09300_;
  wire _09301_;
  wire _09302_;
  wire _09303_;
  wire _09304_;
  wire _09305_;
  wire _09306_;
  wire _09307_;
  wire _09308_;
  wire _09309_;
  wire _09310_;
  wire _09311_;
  wire _09312_;
  wire _09313_;
  wire _09314_;
  wire _09315_;
  wire _09316_;
  wire _09317_;
  wire _09318_;
  wire _09319_;
  wire _09320_;
  wire _09321_;
  wire _09322_;
  wire _09323_;
  wire _09324_;
  wire _09325_;
  wire _09326_;
  wire _09327_;
  wire _09328_;
  wire _09329_;
  wire _09330_;
  wire _09331_;
  wire _09332_;
  wire _09333_;
  wire _09334_;
  wire _09335_;
  wire _09336_;
  wire _09337_;
  wire _09338_;
  wire _09339_;
  wire _09340_;
  wire _09341_;
  wire _09342_;
  wire _09343_;
  wire _09344_;
  wire _09345_;
  wire _09346_;
  wire _09347_;
  wire _09348_;
  wire _09349_;
  wire _09350_;
  wire _09351_;
  wire _09352_;
  wire _09353_;
  wire _09354_;
  wire _09355_;
  wire _09356_;
  wire _09357_;
  wire _09358_;
  wire _09359_;
  wire _09360_;
  wire _09361_;
  wire _09362_;
  wire _09363_;
  wire _09364_;
  wire _09365_;
  wire _09366_;
  wire _09367_;
  wire _09368_;
  wire _09369_;
  wire _09370_;
  wire _09371_;
  wire _09372_;
  wire _09373_;
  wire _09374_;
  wire _09375_;
  wire _09376_;
  wire _09377_;
  wire _09378_;
  wire _09379_;
  wire _09380_;
  wire _09381_;
  wire _09382_;
  wire _09383_;
  wire _09384_;
  wire _09385_;
  wire _09386_;
  wire _09387_;
  wire _09388_;
  wire _09389_;
  wire _09390_;
  wire _09391_;
  wire _09392_;
  wire _09393_;
  wire _09394_;
  wire _09395_;
  wire _09396_;
  wire _09397_;
  wire _09398_;
  wire _09399_;
  wire _09400_;
  wire _09401_;
  wire _09402_;
  wire _09403_;
  wire _09404_;
  wire _09405_;
  wire _09406_;
  wire _09407_;
  wire _09408_;
  wire _09409_;
  wire _09410_;
  wire _09411_;
  wire _09412_;
  wire _09413_;
  wire _09414_;
  wire _09415_;
  wire _09416_;
  wire _09417_;
  wire _09418_;
  wire _09419_;
  wire _09420_;
  wire _09421_;
  wire _09422_;
  wire _09423_;
  wire _09424_;
  wire _09425_;
  wire _09426_;
  wire _09427_;
  wire _09428_;
  wire _09429_;
  wire _09430_;
  wire _09431_;
  wire _09432_;
  wire _09433_;
  wire _09434_;
  wire _09435_;
  wire _09436_;
  wire _09437_;
  wire _09438_;
  wire _09439_;
  wire _09440_;
  wire _09441_;
  wire _09442_;
  wire _09443_;
  wire _09444_;
  wire _09445_;
  wire _09446_;
  wire _09447_;
  wire _09448_;
  wire _09449_;
  wire _09450_;
  wire _09451_;
  wire _09452_;
  wire _09453_;
  wire _09454_;
  wire _09455_;
  wire _09456_;
  wire _09457_;
  wire _09458_;
  wire _09459_;
  wire _09460_;
  wire _09461_;
  wire _09462_;
  wire _09463_;
  wire _09464_;
  wire _09465_;
  wire _09466_;
  wire _09467_;
  wire _09468_;
  wire _09469_;
  wire _09470_;
  wire _09471_;
  wire _09472_;
  wire _09473_;
  wire _09474_;
  wire _09475_;
  wire _09476_;
  wire _09477_;
  wire _09478_;
  wire _09479_;
  wire _09480_;
  wire _09481_;
  wire _09482_;
  wire _09483_;
  wire _09484_;
  wire _09485_;
  wire _09486_;
  wire _09487_;
  wire _09488_;
  wire _09489_;
  wire _09490_;
  wire _09491_;
  wire _09492_;
  wire _09493_;
  wire _09494_;
  wire _09495_;
  wire _09496_;
  wire _09497_;
  wire _09498_;
  wire _09499_;
  wire _09500_;
  wire _09501_;
  wire _09502_;
  wire _09503_;
  wire _09504_;
  wire _09505_;
  wire _09506_;
  wire _09507_;
  wire _09508_;
  wire _09509_;
  wire _09510_;
  wire _09511_;
  wire _09512_;
  wire _09513_;
  wire _09514_;
  wire _09515_;
  wire _09516_;
  wire _09517_;
  wire _09518_;
  wire _09519_;
  wire _09520_;
  wire _09521_;
  wire _09522_;
  wire _09523_;
  wire _09524_;
  wire _09525_;
  wire _09526_;
  wire _09527_;
  wire _09528_;
  wire _09529_;
  wire _09530_;
  wire _09531_;
  wire _09532_;
  wire _09533_;
  wire _09534_;
  wire _09535_;
  wire _09536_;
  wire _09537_;
  wire _09538_;
  wire _09539_;
  wire _09540_;
  wire _09541_;
  wire _09542_;
  wire _09543_;
  wire _09544_;
  wire _09545_;
  wire _09546_;
  wire _09547_;
  wire _09548_;
  wire _09549_;
  wire _09550_;
  wire _09551_;
  wire _09552_;
  wire _09553_;
  wire _09554_;
  wire _09555_;
  wire _09556_;
  wire _09557_;
  wire _09558_;
  wire _09559_;
  wire _09560_;
  wire _09561_;
  wire _09562_;
  wire _09563_;
  wire _09564_;
  wire _09565_;
  wire _09566_;
  wire _09567_;
  wire _09568_;
  wire _09569_;
  wire _09570_;
  wire _09571_;
  wire _09572_;
  wire _09573_;
  wire _09574_;
  wire _09575_;
  wire _09576_;
  wire _09577_;
  wire _09578_;
  wire _09579_;
  wire _09580_;
  wire _09581_;
  wire _09582_;
  wire _09583_;
  wire _09584_;
  wire _09585_;
  wire _09586_;
  wire _09587_;
  wire _09588_;
  wire _09589_;
  wire _09590_;
  wire _09591_;
  wire _09592_;
  wire _09593_;
  wire _09594_;
  wire _09595_;
  wire _09596_;
  wire _09597_;
  wire _09598_;
  wire _09599_;
  wire _09600_;
  wire _09601_;
  wire _09602_;
  wire _09603_;
  wire _09604_;
  wire _09605_;
  wire _09606_;
  wire _09607_;
  wire _09608_;
  wire _09609_;
  wire _09610_;
  wire _09611_;
  wire _09612_;
  wire _09613_;
  wire _09614_;
  wire _09615_;
  wire _09616_;
  wire _09617_;
  wire _09618_;
  wire _09619_;
  wire _09620_;
  wire _09621_;
  wire _09622_;
  wire _09623_;
  wire _09624_;
  wire _09625_;
  wire _09626_;
  wire _09627_;
  wire _09628_;
  wire _09629_;
  wire _09630_;
  wire _09631_;
  wire _09632_;
  wire _09633_;
  wire _09634_;
  wire _09635_;
  wire _09636_;
  wire _09637_;
  wire _09638_;
  wire _09639_;
  wire _09640_;
  wire _09641_;
  wire _09642_;
  wire _09643_;
  wire _09644_;
  wire _09645_;
  wire _09646_;
  wire _09647_;
  wire _09648_;
  wire _09649_;
  wire _09650_;
  wire _09651_;
  wire _09652_;
  wire _09653_;
  wire _09654_;
  wire _09655_;
  wire _09656_;
  wire _09657_;
  wire _09658_;
  wire _09659_;
  wire _09660_;
  wire _09661_;
  wire _09662_;
  wire _09663_;
  wire _09664_;
  wire _09665_;
  wire _09666_;
  wire _09667_;
  wire _09668_;
  wire _09669_;
  wire _09670_;
  wire _09671_;
  wire _09672_;
  wire _09673_;
  wire _09674_;
  wire _09675_;
  wire _09676_;
  wire _09677_;
  wire _09678_;
  wire _09679_;
  wire _09680_;
  wire _09681_;
  wire _09682_;
  wire _09683_;
  wire _09684_;
  wire _09685_;
  wire _09686_;
  wire _09687_;
  wire _09688_;
  wire _09689_;
  wire _09690_;
  wire _09691_;
  wire _09692_;
  wire _09693_;
  wire _09694_;
  wire _09695_;
  wire _09696_;
  wire _09697_;
  wire _09698_;
  wire _09699_;
  wire _09700_;
  wire _09701_;
  wire _09702_;
  wire _09703_;
  wire _09704_;
  wire _09705_;
  wire _09706_;
  wire _09707_;
  wire _09708_;
  wire _09709_;
  wire _09710_;
  wire _09711_;
  wire _09712_;
  wire _09713_;
  wire _09714_;
  wire _09715_;
  wire _09716_;
  wire _09717_;
  wire _09718_;
  wire _09719_;
  wire _09720_;
  wire _09721_;
  wire _09722_;
  wire _09723_;
  wire _09724_;
  wire _09725_;
  wire _09726_;
  wire _09727_;
  wire _09728_;
  wire _09729_;
  wire _09730_;
  wire _09731_;
  wire _09732_;
  wire _09733_;
  wire _09734_;
  wire _09735_;
  wire _09736_;
  wire _09737_;
  wire _09738_;
  wire _09739_;
  wire _09740_;
  wire _09741_;
  wire _09742_;
  wire _09743_;
  wire _09744_;
  wire _09745_;
  wire _09746_;
  wire _09747_;
  wire _09748_;
  wire _09749_;
  wire _09750_;
  wire _09751_;
  wire _09752_;
  wire _09753_;
  wire _09754_;
  wire _09755_;
  wire _09756_;
  wire _09757_;
  wire _09758_;
  wire _09759_;
  wire _09760_;
  wire _09761_;
  wire _09762_;
  wire _09763_;
  wire _09764_;
  wire _09765_;
  wire _09766_;
  wire _09767_;
  wire _09768_;
  wire _09769_;
  wire _09770_;
  wire _09771_;
  wire _09772_;
  wire _09773_;
  wire _09774_;
  wire _09775_;
  wire _09776_;
  wire _09777_;
  wire _09778_;
  wire _09779_;
  wire _09780_;
  wire _09781_;
  wire _09782_;
  wire _09783_;
  wire _09784_;
  wire _09785_;
  wire _09786_;
  wire _09787_;
  wire _09788_;
  wire _09789_;
  wire _09790_;
  wire _09791_;
  wire _09792_;
  wire _09793_;
  wire _09794_;
  wire _09795_;
  wire _09796_;
  wire _09797_;
  wire _09798_;
  wire _09799_;
  wire _09800_;
  wire _09801_;
  wire _09802_;
  wire _09803_;
  wire _09804_;
  wire _09805_;
  wire _09806_;
  wire _09807_;
  wire _09808_;
  wire _09809_;
  wire _09810_;
  wire _09811_;
  wire _09812_;
  wire _09813_;
  wire _09814_;
  wire _09815_;
  wire _09816_;
  wire _09817_;
  wire _09818_;
  wire _09819_;
  wire _09820_;
  wire _09821_;
  wire _09822_;
  wire _09823_;
  wire _09824_;
  wire _09825_;
  wire _09826_;
  wire _09827_;
  wire _09828_;
  wire _09829_;
  wire _09830_;
  wire _09831_;
  wire _09832_;
  wire _09833_;
  wire _09834_;
  wire _09835_;
  wire _09836_;
  wire _09837_;
  wire _09838_;
  wire _09839_;
  wire _09840_;
  wire _09841_;
  wire _09842_;
  wire _09843_;
  wire _09844_;
  wire _09845_;
  wire _09846_;
  wire _09847_;
  wire _09848_;
  wire _09849_;
  wire _09850_;
  wire _09851_;
  wire _09852_;
  wire _09853_;
  wire _09854_;
  wire _09855_;
  wire _09856_;
  wire _09857_;
  wire _09858_;
  wire _09859_;
  wire _09860_;
  wire _09861_;
  wire _09862_;
  wire _09863_;
  wire _09864_;
  wire _09865_;
  wire _09866_;
  wire _09867_;
  wire _09868_;
  wire _09869_;
  wire _09870_;
  wire _09871_;
  wire _09872_;
  wire _09873_;
  wire _09874_;
  wire _09875_;
  wire _09876_;
  wire _09877_;
  wire _09878_;
  wire _09879_;
  wire _09880_;
  wire _09881_;
  wire _09882_;
  wire _09883_;
  wire _09884_;
  wire _09885_;
  wire _09886_;
  wire _09887_;
  wire _09888_;
  wire _09889_;
  wire _09890_;
  wire _09891_;
  wire _09892_;
  wire _09893_;
  wire _09894_;
  wire _09895_;
  wire _09896_;
  wire _09897_;
  wire _09898_;
  wire _09899_;
  wire _09900_;
  wire _09901_;
  wire _09902_;
  wire _09903_;
  wire _09904_;
  wire _09905_;
  wire _09906_;
  wire _09907_;
  wire _09908_;
  wire _09909_;
  wire _09910_;
  wire _09911_;
  wire _09912_;
  wire _09913_;
  wire _09914_;
  wire _09915_;
  wire _09916_;
  wire _09917_;
  wire _09918_;
  wire _09919_;
  wire _09920_;
  wire _09921_;
  wire _09922_;
  wire _09923_;
  wire _09924_;
  wire _09925_;
  wire _09926_;
  wire _09927_;
  wire _09928_;
  wire _09929_;
  wire _09930_;
  wire _09931_;
  wire _09932_;
  wire _09933_;
  wire _09934_;
  wire _09935_;
  wire _09936_;
  wire _09937_;
  wire _09938_;
  wire _09939_;
  wire _09940_;
  wire _09941_;
  wire _09942_;
  wire _09943_;
  wire _09944_;
  wire _09945_;
  wire _09946_;
  wire _09947_;
  wire _09948_;
  wire _09949_;
  wire _09950_;
  wire _09951_;
  wire _09952_;
  wire _09953_;
  wire _09954_;
  wire _09955_;
  wire _09956_;
  wire _09957_;
  wire _09958_;
  wire _09959_;
  wire _09960_;
  wire _09961_;
  wire _09962_;
  wire _09963_;
  wire _09964_;
  wire _09965_;
  wire _09966_;
  wire _09967_;
  wire _09968_;
  wire _09969_;
  wire _09970_;
  wire _09971_;
  wire _09972_;
  wire _09973_;
  wire _09974_;
  wire _09975_;
  wire _09976_;
  wire _09977_;
  wire _09978_;
  wire _09979_;
  wire _09980_;
  wire _09981_;
  wire _09982_;
  wire _09983_;
  wire _09984_;
  wire _09985_;
  wire _09986_;
  wire _09987_;
  wire _09988_;
  wire _09989_;
  wire _09990_;
  wire _09991_;
  wire _09992_;
  wire _09993_;
  wire _09994_;
  wire _09995_;
  wire _09996_;
  wire _09997_;
  wire _09998_;
  wire _09999_;
  wire _10000_;
  wire _10001_;
  wire _10002_;
  wire _10003_;
  wire _10004_;
  wire _10005_;
  wire _10006_;
  wire _10007_;
  wire _10008_;
  wire _10009_;
  wire _10010_;
  wire _10011_;
  wire _10012_;
  wire _10013_;
  wire _10014_;
  wire _10015_;
  wire _10016_;
  wire _10017_;
  wire _10018_;
  wire _10019_;
  wire _10020_;
  wire _10021_;
  wire _10022_;
  wire _10023_;
  wire _10024_;
  wire _10025_;
  wire _10026_;
  wire _10027_;
  wire _10028_;
  wire _10029_;
  wire _10030_;
  wire _10031_;
  wire _10032_;
  wire _10033_;
  wire _10034_;
  wire _10035_;
  wire _10036_;
  wire _10037_;
  wire _10038_;
  wire _10039_;
  wire _10040_;
  wire _10041_;
  wire _10042_;
  wire _10043_;
  wire _10044_;
  wire _10045_;
  wire _10046_;
  wire _10047_;
  wire _10048_;
  wire _10049_;
  wire _10050_;
  wire _10051_;
  wire _10052_;
  wire _10053_;
  wire _10054_;
  wire _10055_;
  wire _10056_;
  wire _10057_;
  wire _10058_;
  wire _10059_;
  wire _10060_;
  wire _10061_;
  wire _10062_;
  wire _10063_;
  wire _10064_;
  wire _10065_;
  wire _10066_;
  wire _10067_;
  wire _10068_;
  wire _10069_;
  wire _10070_;
  wire _10071_;
  wire _10072_;
  wire _10073_;
  wire _10074_;
  wire _10075_;
  wire _10076_;
  wire _10077_;
  wire _10078_;
  wire _10079_;
  wire _10080_;
  wire _10081_;
  wire _10082_;
  wire _10083_;
  wire _10084_;
  wire _10085_;
  wire _10086_;
  wire _10087_;
  wire _10088_;
  wire _10089_;
  wire _10090_;
  wire _10091_;
  wire _10092_;
  wire _10093_;
  wire _10094_;
  wire _10095_;
  wire _10096_;
  wire _10097_;
  wire _10098_;
  wire _10099_;
  wire _10100_;
  wire _10101_;
  wire _10102_;
  wire _10103_;
  wire _10104_;
  wire _10105_;
  wire _10106_;
  wire _10107_;
  wire _10108_;
  wire _10109_;
  wire _10110_;
  wire _10111_;
  wire _10112_;
  wire _10113_;
  wire _10114_;
  wire _10115_;
  wire _10116_;
  wire _10117_;
  wire _10118_;
  wire _10119_;
  wire _10120_;
  wire _10121_;
  wire _10122_;
  wire _10123_;
  wire _10124_;
  wire _10125_;
  wire _10126_;
  wire _10127_;
  wire _10128_;
  wire _10129_;
  wire _10130_;
  wire _10131_;
  wire _10132_;
  wire _10133_;
  wire _10134_;
  wire _10135_;
  wire _10136_;
  wire _10137_;
  wire _10138_;
  wire _10139_;
  wire _10140_;
  wire _10141_;
  wire _10142_;
  wire _10143_;
  wire _10144_;
  wire _10145_;
  wire _10146_;
  wire _10147_;
  wire _10148_;
  wire _10149_;
  wire _10150_;
  wire _10151_;
  wire _10152_;
  wire _10153_;
  wire _10154_;
  wire _10155_;
  wire _10156_;
  wire _10157_;
  wire _10158_;
  wire _10159_;
  wire _10160_;
  wire _10161_;
  wire _10162_;
  wire _10163_;
  wire _10164_;
  wire _10165_;
  wire _10166_;
  wire _10167_;
  wire _10168_;
  wire _10169_;
  wire _10170_;
  wire _10171_;
  wire _10172_;
  wire _10173_;
  wire _10174_;
  wire _10175_;
  wire _10176_;
  wire _10177_;
  wire _10178_;
  wire _10179_;
  wire _10180_;
  wire _10181_;
  wire _10182_;
  wire _10183_;
  wire _10184_;
  wire _10185_;
  wire _10186_;
  wire _10187_;
  wire _10188_;
  wire _10189_;
  wire _10190_;
  wire _10191_;
  wire _10192_;
  wire _10193_;
  wire _10194_;
  wire _10195_;
  wire _10196_;
  wire _10197_;
  wire _10198_;
  wire _10199_;
  wire _10200_;
  wire _10201_;
  wire _10202_;
  wire _10203_;
  wire _10204_;
  wire _10205_;
  wire _10206_;
  wire _10207_;
  wire _10208_;
  wire _10209_;
  wire _10210_;
  wire _10211_;
  wire _10212_;
  wire _10213_;
  wire _10214_;
  wire _10215_;
  wire _10216_;
  wire _10217_;
  wire _10218_;
  wire _10219_;
  wire _10220_;
  wire _10221_;
  wire _10222_;
  wire _10223_;
  wire _10224_;
  wire _10225_;
  wire _10226_;
  wire _10227_;
  wire _10228_;
  wire _10229_;
  wire _10230_;
  wire _10231_;
  wire _10232_;
  wire _10233_;
  wire _10234_;
  wire _10235_;
  wire _10236_;
  wire _10237_;
  wire _10238_;
  wire _10239_;
  wire _10240_;
  wire _10241_;
  wire _10242_;
  wire _10243_;
  wire _10244_;
  wire _10245_;
  wire _10246_;
  wire _10247_;
  wire _10248_;
  wire _10249_;
  wire _10250_;
  wire _10251_;
  wire _10252_;
  wire _10253_;
  wire _10254_;
  wire _10255_;
  wire _10256_;
  wire _10257_;
  wire _10258_;
  wire _10259_;
  wire _10260_;
  wire _10261_;
  wire _10262_;
  wire _10263_;
  wire _10264_;
  wire _10265_;
  wire _10266_;
  wire _10267_;
  wire _10268_;
  wire _10269_;
  wire _10270_;
  wire _10271_;
  wire _10272_;
  wire _10273_;
  wire _10274_;
  wire _10275_;
  wire _10276_;
  wire _10277_;
  wire _10278_;
  wire _10279_;
  wire _10280_;
  wire _10281_;
  wire _10282_;
  wire _10283_;
  wire _10284_;
  wire _10285_;
  wire _10286_;
  wire _10287_;
  wire _10288_;
  wire _10289_;
  wire _10290_;
  wire _10291_;
  wire _10292_;
  wire _10293_;
  wire _10294_;
  wire _10295_;
  wire _10296_;
  wire _10297_;
  wire _10298_;
  wire _10299_;
  wire _10300_;
  wire _10301_;
  wire _10302_;
  wire _10303_;
  wire _10304_;
  wire _10305_;
  wire _10306_;
  wire _10307_;
  wire _10308_;
  wire _10309_;
  wire _10310_;
  wire _10311_;
  wire _10312_;
  wire _10313_;
  wire _10314_;
  wire _10315_;
  wire _10316_;
  wire _10317_;
  wire _10318_;
  wire _10319_;
  wire _10320_;
  wire _10321_;
  wire _10322_;
  wire _10323_;
  wire _10324_;
  wire _10325_;
  wire _10326_;
  wire _10327_;
  wire _10328_;
  wire _10329_;
  wire _10330_;
  wire _10331_;
  wire _10332_;
  wire _10333_;
  wire _10334_;
  wire _10335_;
  wire _10336_;
  wire _10337_;
  wire _10338_;
  wire _10339_;
  wire _10340_;
  wire _10341_;
  wire _10342_;
  wire _10343_;
  wire _10344_;
  wire _10345_;
  wire _10346_;
  wire _10347_;
  wire _10348_;
  wire _10349_;
  wire _10350_;
  wire _10351_;
  wire _10352_;
  wire _10353_;
  wire _10354_;
  wire _10355_;
  wire _10356_;
  wire _10357_;
  wire _10358_;
  wire _10359_;
  wire _10360_;
  wire _10361_;
  wire _10362_;
  wire _10363_;
  wire _10364_;
  wire _10365_;
  wire _10366_;
  wire _10367_;
  wire _10368_;
  wire _10369_;
  wire _10370_;
  wire _10371_;
  wire _10372_;
  wire _10373_;
  wire _10374_;
  wire _10375_;
  wire _10376_;
  wire _10377_;
  wire _10378_;
  wire _10379_;
  wire _10380_;
  wire _10381_;
  wire _10382_;
  wire _10383_;
  wire _10384_;
  wire _10385_;
  wire _10386_;
  wire _10387_;
  wire _10388_;
  wire _10389_;
  wire _10390_;
  wire _10391_;
  wire _10392_;
  wire _10393_;
  wire _10394_;
  wire _10395_;
  wire _10396_;
  wire _10397_;
  wire _10398_;
  wire _10399_;
  wire _10400_;
  wire _10401_;
  wire _10402_;
  wire _10403_;
  wire _10404_;
  wire _10405_;
  wire _10406_;
  wire _10407_;
  wire _10408_;
  wire _10409_;
  wire _10410_;
  wire _10411_;
  wire _10412_;
  wire _10413_;
  wire _10414_;
  wire _10415_;
  wire _10416_;
  wire _10417_;
  wire _10418_;
  wire _10419_;
  wire _10420_;
  wire _10421_;
  wire _10422_;
  wire _10423_;
  wire _10424_;
  wire _10425_;
  wire _10426_;
  wire _10427_;
  wire _10428_;
  wire _10429_;
  wire _10430_;
  wire _10431_;
  wire _10432_;
  wire _10433_;
  wire _10434_;
  wire _10435_;
  wire _10436_;
  wire _10437_;
  wire _10438_;
  wire _10439_;
  wire _10440_;
  wire _10441_;
  wire _10442_;
  wire _10443_;
  wire _10444_;
  wire _10445_;
  wire _10446_;
  wire _10447_;
  wire _10448_;
  wire _10449_;
  wire _10450_;
  wire _10451_;
  wire _10452_;
  wire _10453_;
  wire _10454_;
  wire _10455_;
  wire _10456_;
  wire _10457_;
  wire _10458_;
  wire _10459_;
  wire _10460_;
  wire _10461_;
  wire _10462_;
  wire _10463_;
  wire _10464_;
  wire _10465_;
  wire _10466_;
  wire _10467_;
  wire _10468_;
  wire _10469_;
  wire _10470_;
  wire _10471_;
  wire _10472_;
  wire _10473_;
  wire _10474_;
  wire _10475_;
  wire _10476_;
  wire _10477_;
  wire _10478_;
  wire _10479_;
  wire _10480_;
  wire _10481_;
  wire _10482_;
  wire _10483_;
  wire _10484_;
  wire _10485_;
  wire _10486_;
  wire _10487_;
  wire _10488_;
  wire _10489_;
  wire _10490_;
  wire _10491_;
  wire _10492_;
  wire _10493_;
  wire _10494_;
  wire _10495_;
  wire _10496_;
  wire _10497_;
  wire _10498_;
  wire _10499_;
  wire _10500_;
  wire _10501_;
  wire _10502_;
  wire _10503_;
  wire _10504_;
  wire _10505_;
  wire _10506_;
  wire _10507_;
  wire _10508_;
  wire _10509_;
  wire _10510_;
  wire _10511_;
  wire _10512_;
  wire _10513_;
  wire _10514_;
  wire _10515_;
  wire _10516_;
  wire _10517_;
  wire _10518_;
  wire _10519_;
  wire _10520_;
  wire _10521_;
  wire _10522_;
  wire _10523_;
  wire _10524_;
  wire _10525_;
  wire _10526_;
  wire _10527_;
  wire _10528_;
  wire _10529_;
  wire _10530_;
  wire _10531_;
  wire _10532_;
  wire _10533_;
  wire _10534_;
  wire _10535_;
  wire _10536_;
  wire _10537_;
  wire _10538_;
  wire _10539_;
  wire _10540_;
  wire _10541_;
  wire _10542_;
  wire _10543_;
  wire _10544_;
  wire _10545_;
  wire _10546_;
  wire _10547_;
  wire _10548_;
  wire _10549_;
  wire _10550_;
  wire _10551_;
  wire _10552_;
  wire _10553_;
  wire _10554_;
  wire _10555_;
  wire _10556_;
  wire _10557_;
  wire _10558_;
  wire _10559_;
  wire _10560_;
  wire _10561_;
  wire _10562_;
  wire _10563_;
  wire _10564_;
  wire _10565_;
  wire _10566_;
  wire _10567_;
  wire _10568_;
  wire _10569_;
  wire _10570_;
  wire _10571_;
  wire _10572_;
  wire _10573_;
  wire _10574_;
  wire _10575_;
  wire _10576_;
  wire _10577_;
  wire _10578_;
  wire _10579_;
  wire _10580_;
  wire _10581_;
  wire _10582_;
  wire _10583_;
  wire _10584_;
  wire _10585_;
  wire _10586_;
  wire _10587_;
  wire _10588_;
  wire _10589_;
  wire _10590_;
  wire _10591_;
  wire _10592_;
  wire _10593_;
  wire _10594_;
  wire _10595_;
  wire _10596_;
  wire _10597_;
  wire _10598_;
  wire _10599_;
  wire _10600_;
  wire _10601_;
  wire _10602_;
  wire _10603_;
  wire _10604_;
  wire _10605_;
  wire _10606_;
  wire _10607_;
  wire _10608_;
  wire _10609_;
  wire _10610_;
  wire _10611_;
  wire _10612_;
  wire _10613_;
  wire _10614_;
  wire _10615_;
  wire _10616_;
  wire _10617_;
  wire _10618_;
  wire _10619_;
  wire _10620_;
  wire _10621_;
  wire _10622_;
  wire _10623_;
  wire _10624_;
  wire _10625_;
  wire _10626_;
  wire _10627_;
  wire _10628_;
  wire _10629_;
  wire _10630_;
  wire _10631_;
  wire _10632_;
  wire _10633_;
  wire _10634_;
  wire _10635_;
  wire _10636_;
  wire _10637_;
  wire _10638_;
  wire _10639_;
  wire _10640_;
  wire _10641_;
  wire _10642_;
  wire _10643_;
  wire _10644_;
  wire _10645_;
  wire _10646_;
  wire _10647_;
  wire _10648_;
  wire _10649_;
  wire _10650_;
  wire _10651_;
  wire _10652_;
  wire _10653_;
  wire _10654_;
  wire _10655_;
  wire _10656_;
  wire _10657_;
  wire _10658_;
  wire _10659_;
  wire _10660_;
  wire _10661_;
  wire _10662_;
  wire _10663_;
  wire _10664_;
  wire _10665_;
  wire _10666_;
  wire _10667_;
  wire _10668_;
  wire _10669_;
  wire _10670_;
  wire _10671_;
  wire _10672_;
  wire _10673_;
  wire _10674_;
  wire _10675_;
  wire _10676_;
  wire _10677_;
  wire _10678_;
  wire _10679_;
  wire _10680_;
  wire _10681_;
  wire _10682_;
  wire _10683_;
  wire _10684_;
  wire _10685_;
  wire _10686_;
  wire _10687_;
  wire _10688_;
  wire _10689_;
  wire _10690_;
  wire _10691_;
  wire _10692_;
  wire _10693_;
  wire _10694_;
  wire _10695_;
  wire _10696_;
  wire _10697_;
  wire _10698_;
  wire _10699_;
  wire _10700_;
  wire _10701_;
  wire _10702_;
  wire _10703_;
  wire _10704_;
  wire _10705_;
  wire _10706_;
  wire _10707_;
  wire _10708_;
  wire _10709_;
  wire _10710_;
  wire _10711_;
  wire _10712_;
  wire _10713_;
  wire _10714_;
  wire _10715_;
  wire _10716_;
  wire _10717_;
  wire _10718_;
  wire _10719_;
  wire _10720_;
  wire _10721_;
  wire _10722_;
  wire _10723_;
  wire _10724_;
  wire _10725_;
  wire _10726_;
  wire _10727_;
  wire _10728_;
  wire _10729_;
  wire _10730_;
  wire _10731_;
  wire _10732_;
  wire _10733_;
  wire _10734_;
  wire _10735_;
  wire _10736_;
  wire _10737_;
  wire _10738_;
  wire _10739_;
  wire _10740_;
  wire _10741_;
  wire _10742_;
  wire _10743_;
  wire _10744_;
  wire _10745_;
  wire _10746_;
  wire _10747_;
  wire _10748_;
  wire _10749_;
  wire _10750_;
  wire _10751_;
  wire _10752_;
  wire _10753_;
  wire _10754_;
  wire _10755_;
  wire _10756_;
  wire _10757_;
  wire _10758_;
  wire _10759_;
  wire _10760_;
  wire _10761_;
  wire _10762_;
  wire _10763_;
  wire _10764_;
  wire _10765_;
  wire _10766_;
  wire _10767_;
  wire _10768_;
  wire _10769_;
  wire _10770_;
  wire _10771_;
  wire _10772_;
  wire _10773_;
  wire _10774_;
  wire _10775_;
  wire _10776_;
  wire _10777_;
  wire _10778_;
  wire _10779_;
  wire _10780_;
  wire _10781_;
  wire _10782_;
  wire _10783_;
  wire _10784_;
  wire _10785_;
  wire _10786_;
  wire _10787_;
  wire _10788_;
  wire _10789_;
  wire _10790_;
  wire _10791_;
  wire _10792_;
  wire _10793_;
  wire _10794_;
  wire _10795_;
  wire _10796_;
  wire _10797_;
  wire _10798_;
  wire _10799_;
  wire _10800_;
  wire _10801_;
  wire _10802_;
  wire _10803_;
  wire _10804_;
  wire _10805_;
  wire _10806_;
  wire _10807_;
  wire _10808_;
  wire _10809_;
  wire _10810_;
  wire _10811_;
  wire _10812_;
  wire _10813_;
  wire _10814_;
  wire _10815_;
  wire _10816_;
  wire _10817_;
  wire _10818_;
  wire _10819_;
  wire _10820_;
  wire _10821_;
  wire _10822_;
  wire _10823_;
  wire _10824_;
  wire _10825_;
  wire _10826_;
  wire _10827_;
  wire _10828_;
  wire _10829_;
  wire _10830_;
  wire _10831_;
  wire _10832_;
  wire _10833_;
  wire _10834_;
  wire _10835_;
  wire _10836_;
  wire _10837_;
  wire _10838_;
  wire _10839_;
  wire _10840_;
  wire _10841_;
  wire _10842_;
  wire _10843_;
  wire _10844_;
  wire _10845_;
  wire _10846_;
  wire _10847_;
  wire _10848_;
  wire _10849_;
  wire _10850_;
  wire _10851_;
  wire _10852_;
  wire _10853_;
  wire _10854_;
  wire _10855_;
  wire _10856_;
  wire _10857_;
  wire _10858_;
  wire _10859_;
  wire _10860_;
  wire _10861_;
  wire _10862_;
  wire _10863_;
  wire _10864_;
  wire _10865_;
  wire _10866_;
  wire _10867_;
  wire _10868_;
  wire _10869_;
  wire _10870_;
  wire _10871_;
  wire _10872_;
  wire _10873_;
  wire _10874_;
  wire _10875_;
  wire _10876_;
  wire _10877_;
  wire _10878_;
  wire _10879_;
  wire _10880_;
  wire _10881_;
  wire _10882_;
  wire _10883_;
  wire _10884_;
  wire _10885_;
  wire _10886_;
  wire _10887_;
  wire _10888_;
  wire _10889_;
  wire _10890_;
  wire _10891_;
  wire _10892_;
  wire _10893_;
  wire _10894_;
  wire _10895_;
  wire _10896_;
  wire _10897_;
  wire _10898_;
  wire _10899_;
  wire _10900_;
  wire _10901_;
  wire _10902_;
  wire _10903_;
  wire _10904_;
  wire _10905_;
  wire _10906_;
  wire _10907_;
  wire _10908_;
  wire _10909_;
  wire _10910_;
  wire _10911_;
  wire _10912_;
  wire _10913_;
  wire _10914_;
  wire _10915_;
  wire _10916_;
  wire _10917_;
  wire _10918_;
  wire _10919_;
  wire _10920_;
  wire _10921_;
  wire _10922_;
  wire _10923_;
  wire _10924_;
  wire _10925_;
  wire _10926_;
  wire _10927_;
  wire _10928_;
  wire _10929_;
  wire _10930_;
  wire _10931_;
  wire _10932_;
  wire _10933_;
  wire _10934_;
  wire _10935_;
  wire _10936_;
  wire _10937_;
  wire _10938_;
  wire _10939_;
  wire _10940_;
  wire _10941_;
  wire _10942_;
  wire _10943_;
  wire _10944_;
  wire _10945_;
  wire _10946_;
  wire _10947_;
  wire _10948_;
  wire _10949_;
  wire _10950_;
  wire _10951_;
  wire _10952_;
  wire _10953_;
  wire _10954_;
  wire _10955_;
  wire _10956_;
  wire _10957_;
  wire _10958_;
  wire _10959_;
  wire _10960_;
  wire _10961_;
  wire _10962_;
  wire _10963_;
  wire _10964_;
  wire _10965_;
  wire _10966_;
  wire _10967_;
  wire _10968_;
  wire _10969_;
  wire _10970_;
  wire _10971_;
  wire _10972_;
  wire _10973_;
  wire _10974_;
  wire _10975_;
  wire _10976_;
  wire _10977_;
  wire _10978_;
  wire _10979_;
  wire _10980_;
  wire _10981_;
  wire _10982_;
  wire _10983_;
  wire _10984_;
  wire _10985_;
  wire _10986_;
  wire _10987_;
  wire _10988_;
  wire _10989_;
  wire _10990_;
  wire _10991_;
  wire _10992_;
  wire _10993_;
  wire _10994_;
  wire _10995_;
  wire _10996_;
  wire _10997_;
  wire _10998_;
  wire _10999_;
  wire _11000_;
  wire _11001_;
  wire _11002_;
  wire _11003_;
  wire _11004_;
  wire _11005_;
  wire _11006_;
  wire _11007_;
  wire _11008_;
  wire _11009_;
  wire _11010_;
  wire _11011_;
  wire _11012_;
  wire _11013_;
  wire _11014_;
  wire _11015_;
  wire _11016_;
  wire _11017_;
  wire _11018_;
  wire _11019_;
  wire _11020_;
  wire _11021_;
  wire _11022_;
  wire _11023_;
  wire _11024_;
  wire _11025_;
  wire _11026_;
  wire _11027_;
  wire _11028_;
  wire _11029_;
  wire _11030_;
  wire _11031_;
  wire _11032_;
  wire _11033_;
  wire _11034_;
  wire _11035_;
  wire _11036_;
  wire _11037_;
  wire _11038_;
  wire _11039_;
  wire _11040_;
  wire _11041_;
  wire _11042_;
  wire _11043_;
  wire _11044_;
  wire _11045_;
  wire _11046_;
  wire _11047_;
  wire _11048_;
  wire _11049_;
  wire _11050_;
  wire _11051_;
  wire _11052_;
  wire _11053_;
  wire _11054_;
  wire _11055_;
  wire _11056_;
  wire _11057_;
  wire _11058_;
  wire _11059_;
  wire _11060_;
  wire _11061_;
  wire _11062_;
  wire _11063_;
  wire _11064_;
  wire _11065_;
  wire _11066_;
  wire _11067_;
  wire _11068_;
  wire _11069_;
  wire _11070_;
  wire _11071_;
  wire _11072_;
  wire _11073_;
  wire _11074_;
  wire _11075_;
  wire _11076_;
  wire _11077_;
  wire _11078_;
  wire _11079_;
  wire _11080_;
  wire _11081_;
  wire _11082_;
  wire _11083_;
  wire _11084_;
  wire _11085_;
  wire _11086_;
  wire _11087_;
  wire _11088_;
  wire _11089_;
  wire _11090_;
  wire _11091_;
  wire _11092_;
  wire _11093_;
  wire _11094_;
  wire _11095_;
  wire _11096_;
  wire _11097_;
  wire _11098_;
  wire _11099_;
  wire _11100_;
  wire _11101_;
  wire _11102_;
  wire _11103_;
  wire _11104_;
  wire _11105_;
  wire _11106_;
  wire _11107_;
  wire _11108_;
  wire _11109_;
  wire _11110_;
  wire _11111_;
  wire _11112_;
  wire _11113_;
  wire _11114_;
  wire _11115_;
  wire _11116_;
  wire _11117_;
  wire _11118_;
  wire _11119_;
  wire _11120_;
  wire _11121_;
  wire _11122_;
  wire _11123_;
  wire _11124_;
  wire _11125_;
  wire _11126_;
  wire _11127_;
  wire _11128_;
  wire _11129_;
  wire _11130_;
  wire _11131_;
  wire _11132_;
  wire _11133_;
  wire _11134_;
  wire _11135_;
  wire _11136_;
  wire _11137_;
  wire _11138_;
  wire _11139_;
  wire _11140_;
  wire _11141_;
  wire _11142_;
  wire _11143_;
  wire _11144_;
  wire _11145_;
  wire _11146_;
  wire _11147_;
  wire _11148_;
  wire _11149_;
  wire _11150_;
  wire _11151_;
  wire _11152_;
  wire _11153_;
  wire _11154_;
  wire _11155_;
  wire _11156_;
  wire _11157_;
  wire _11158_;
  wire _11159_;
  wire _11160_;
  wire _11161_;
  wire _11162_;
  wire _11163_;
  wire _11164_;
  wire _11165_;
  wire _11166_;
  wire _11167_;
  wire _11168_;
  wire _11169_;
  wire _11170_;
  wire _11171_;
  wire _11172_;
  wire _11173_;
  wire _11174_;
  wire _11175_;
  wire _11176_;
  wire _11177_;
  wire _11178_;
  wire _11179_;
  wire _11180_;
  wire _11181_;
  wire _11182_;
  wire _11183_;
  wire _11184_;
  wire _11185_;
  wire _11186_;
  wire _11187_;
  wire _11188_;
  wire _11189_;
  wire _11190_;
  wire _11191_;
  wire _11192_;
  wire _11193_;
  wire _11194_;
  wire _11195_;
  wire _11196_;
  wire _11197_;
  wire _11198_;
  wire _11199_;
  wire _11200_;
  wire _11201_;
  wire _11202_;
  wire _11203_;
  wire _11204_;
  wire _11205_;
  wire _11206_;
  wire _11207_;
  wire _11208_;
  wire _11209_;
  wire _11210_;
  wire _11211_;
  wire _11212_;
  wire _11213_;
  wire _11214_;
  wire _11215_;
  wire _11216_;
  wire _11217_;
  wire _11218_;
  wire _11219_;
  wire _11220_;
  wire _11221_;
  wire _11222_;
  wire _11223_;
  wire _11224_;
  wire _11225_;
  wire _11226_;
  wire _11227_;
  wire _11228_;
  wire _11229_;
  wire _11230_;
  wire _11231_;
  wire _11232_;
  wire _11233_;
  wire _11234_;
  wire _11235_;
  wire _11236_;
  wire _11237_;
  wire _11238_;
  wire _11239_;
  wire _11240_;
  wire _11241_;
  wire _11242_;
  wire _11243_;
  wire _11244_;
  wire _11245_;
  wire _11246_;
  wire _11247_;
  wire _11248_;
  wire _11249_;
  wire _11250_;
  wire _11251_;
  wire _11252_;
  wire _11253_;
  wire _11254_;
  wire _11255_;
  wire _11256_;
  wire _11257_;
  wire _11258_;
  wire _11259_;
  wire _11260_;
  wire _11261_;
  wire _11262_;
  wire _11263_;
  wire _11264_;
  wire _11265_;
  wire _11266_;
  wire _11267_;
  wire _11268_;
  wire _11269_;
  wire _11270_;
  wire _11271_;
  wire _11272_;
  wire _11273_;
  wire _11274_;
  wire _11275_;
  wire _11276_;
  wire _11277_;
  wire _11278_;
  wire _11279_;
  wire _11280_;
  wire _11281_;
  wire _11282_;
  wire _11283_;
  wire _11284_;
  wire _11285_;
  wire _11286_;
  wire _11287_;
  wire _11288_;
  wire _11289_;
  wire _11290_;
  wire _11291_;
  wire _11292_;
  wire _11293_;
  wire _11294_;
  wire _11295_;
  wire _11296_;
  wire _11297_;
  wire _11298_;
  wire _11299_;
  wire _11300_;
  wire _11301_;
  wire _11302_;
  wire _11303_;
  wire _11304_;
  wire _11305_;
  wire _11306_;
  wire _11307_;
  wire _11308_;
  wire _11309_;
  wire _11310_;
  wire _11311_;
  wire _11312_;
  wire _11313_;
  wire _11314_;
  wire _11315_;
  wire _11316_;
  wire _11317_;
  wire _11318_;
  wire _11319_;
  wire _11320_;
  wire _11321_;
  wire _11322_;
  wire _11323_;
  wire _11324_;
  wire _11325_;
  wire _11326_;
  wire _11327_;
  wire _11328_;
  wire _11329_;
  wire _11330_;
  wire _11331_;
  wire _11332_;
  wire _11333_;
  wire _11334_;
  wire _11335_;
  wire _11336_;
  wire _11337_;
  wire _11338_;
  wire _11339_;
  wire _11340_;
  wire _11341_;
  wire _11342_;
  wire _11343_;
  wire _11344_;
  wire _11345_;
  wire _11346_;
  wire _11347_;
  wire _11348_;
  wire _11349_;
  wire _11350_;
  wire _11351_;
  wire _11352_;
  wire _11353_;
  wire _11354_;
  wire _11355_;
  wire _11356_;
  wire _11357_;
  wire _11358_;
  wire _11359_;
  wire _11360_;
  wire _11361_;
  wire _11362_;
  wire _11363_;
  wire _11364_;
  wire _11365_;
  wire _11366_;
  wire _11367_;
  wire _11368_;
  wire _11369_;
  wire _11370_;
  wire _11371_;
  wire _11372_;
  wire _11373_;
  wire _11374_;
  wire _11375_;
  wire _11376_;
  wire _11377_;
  wire _11378_;
  wire _11379_;
  wire _11380_;
  wire _11381_;
  wire _11382_;
  wire _11383_;
  wire _11384_;
  wire _11385_;
  wire _11386_;
  wire _11387_;
  wire _11388_;
  wire _11389_;
  wire _11390_;
  wire _11391_;
  wire _11392_;
  wire _11393_;
  wire _11394_;
  wire _11395_;
  wire _11396_;
  wire _11397_;
  wire _11398_;
  wire _11399_;
  wire _11400_;
  wire _11401_;
  wire _11402_;
  wire _11403_;
  wire _11404_;
  wire _11405_;
  wire _11406_;
  wire _11407_;
  wire _11408_;
  wire _11409_;
  wire _11410_;
  wire _11411_;
  wire _11412_;
  wire _11413_;
  wire _11414_;
  wire _11415_;
  wire _11416_;
  wire _11417_;
  wire _11418_;
  wire _11419_;
  wire _11420_;
  wire _11421_;
  wire _11422_;
  wire _11423_;
  wire _11424_;
  wire _11425_;
  wire _11426_;
  wire _11427_;
  wire _11428_;
  wire _11429_;
  wire _11430_;
  wire _11431_;
  wire _11432_;
  wire _11433_;
  wire _11434_;
  wire _11435_;
  wire _11436_;
  wire _11437_;
  wire _11438_;
  wire _11439_;
  wire _11440_;
  wire _11441_;
  wire _11442_;
  wire _11443_;
  wire _11444_;
  wire _11445_;
  wire _11446_;
  wire _11447_;
  wire _11448_;
  wire _11449_;
  wire _11450_;
  wire _11451_;
  wire _11452_;
  wire _11453_;
  wire _11454_;
  wire _11455_;
  wire _11456_;
  wire _11457_;
  wire _11458_;
  wire _11459_;
  wire _11460_;
  wire _11461_;
  wire _11462_;
  wire _11463_;
  wire _11464_;
  wire _11465_;
  wire _11466_;
  wire _11467_;
  wire _11468_;
  wire _11469_;
  wire _11470_;
  wire _11471_;
  wire _11472_;
  wire _11473_;
  wire _11474_;
  wire _11475_;
  wire _11476_;
  wire _11477_;
  wire _11478_;
  wire _11479_;
  wire _11480_;
  wire _11481_;
  wire _11482_;
  wire _11483_;
  wire _11484_;
  wire _11485_;
  wire _11486_;
  wire _11487_;
  wire _11488_;
  wire _11489_;
  wire _11490_;
  wire _11491_;
  wire _11492_;
  wire _11493_;
  wire _11494_;
  wire _11495_;
  wire _11496_;
  wire _11497_;
  wire _11498_;
  wire _11499_;
  wire _11500_;
  wire _11501_;
  wire _11502_;
  wire _11503_;
  wire _11504_;
  wire _11505_;
  wire _11506_;
  wire _11507_;
  wire _11508_;
  wire _11509_;
  wire _11510_;
  wire _11511_;
  wire _11512_;
  wire _11513_;
  wire _11514_;
  wire _11515_;
  wire _11516_;
  wire _11517_;
  wire _11518_;
  wire _11519_;
  wire _11520_;
  wire _11521_;
  wire _11522_;
  wire _11523_;
  wire _11524_;
  wire _11525_;
  wire _11526_;
  wire _11527_;
  wire _11528_;
  wire _11529_;
  wire _11530_;
  wire _11531_;
  wire _11532_;
  wire _11533_;
  wire _11534_;
  wire _11535_;
  wire _11536_;
  wire _11537_;
  wire _11538_;
  wire _11539_;
  wire _11540_;
  wire _11541_;
  wire _11542_;
  wire _11543_;
  wire _11544_;
  wire _11545_;
  wire _11546_;
  wire _11547_;
  wire _11548_;
  wire _11549_;
  wire _11550_;
  wire _11551_;
  wire _11552_;
  wire _11553_;
  wire _11554_;
  wire _11555_;
  wire _11556_;
  wire _11557_;
  wire _11558_;
  wire _11559_;
  wire _11560_;
  wire _11561_;
  wire _11562_;
  wire _11563_;
  wire _11564_;
  wire _11565_;
  wire _11566_;
  wire _11567_;
  wire _11568_;
  wire _11569_;
  wire _11570_;
  wire _11571_;
  wire _11572_;
  wire _11573_;
  wire _11574_;
  wire _11575_;
  wire _11576_;
  wire _11577_;
  wire _11578_;
  wire _11579_;
  wire _11580_;
  wire _11581_;
  wire _11582_;
  wire _11583_;
  wire _11584_;
  wire _11585_;
  wire _11586_;
  wire _11587_;
  wire _11588_;
  wire _11589_;
  wire _11590_;
  wire _11591_;
  wire _11592_;
  wire _11593_;
  wire _11594_;
  wire _11595_;
  wire _11596_;
  wire _11597_;
  wire _11598_;
  wire _11599_;
  wire _11600_;
  wire _11601_;
  wire _11602_;
  wire _11603_;
  wire _11604_;
  wire _11605_;
  wire _11606_;
  wire _11607_;
  wire _11608_;
  wire _11609_;
  wire _11610_;
  wire _11611_;
  wire _11612_;
  wire _11613_;
  wire _11614_;
  wire _11615_;
  wire _11616_;
  wire _11617_;
  wire _11618_;
  wire _11619_;
  wire _11620_;
  wire _11621_;
  wire _11622_;
  wire _11623_;
  wire _11624_;
  wire _11625_;
  wire _11626_;
  wire _11627_;
  wire _11628_;
  wire _11629_;
  wire _11630_;
  wire _11631_;
  wire _11632_;
  wire _11633_;
  wire _11634_;
  wire _11635_;
  wire _11636_;
  wire _11637_;
  wire _11638_;
  wire _11639_;
  wire _11640_;
  wire _11641_;
  wire _11642_;
  wire _11643_;
  wire _11644_;
  wire _11645_;
  wire _11646_;
  wire _11647_;
  wire _11648_;
  wire _11649_;
  wire _11650_;
  wire _11651_;
  wire _11652_;
  wire _11653_;
  wire _11654_;
  wire _11655_;
  wire _11656_;
  wire _11657_;
  wire _11658_;
  wire _11659_;
  wire _11660_;
  wire _11661_;
  wire _11662_;
  wire _11663_;
  wire _11664_;
  wire _11665_;
  wire _11666_;
  wire _11667_;
  wire _11668_;
  wire _11669_;
  wire _11670_;
  wire _11671_;
  wire _11672_;
  wire _11673_;
  wire _11674_;
  wire _11675_;
  wire _11676_;
  wire _11677_;
  wire _11678_;
  wire _11679_;
  wire _11680_;
  wire _11681_;
  wire _11682_;
  wire _11683_;
  wire _11684_;
  wire _11685_;
  wire _11686_;
  wire _11687_;
  wire _11688_;
  wire _11689_;
  wire _11690_;
  wire _11691_;
  wire _11692_;
  wire _11693_;
  wire _11694_;
  wire _11695_;
  wire _11696_;
  wire _11697_;
  wire _11698_;
  wire _11699_;
  wire _11700_;
  wire _11701_;
  wire _11702_;
  wire _11703_;
  wire _11704_;
  wire _11705_;
  wire _11706_;
  wire _11707_;
  wire _11708_;
  wire _11709_;
  wire _11710_;
  wire _11711_;
  wire _11712_;
  wire _11713_;
  wire _11714_;
  wire _11715_;
  wire _11716_;
  wire _11717_;
  wire _11718_;
  wire _11719_;
  wire _11720_;
  wire _11721_;
  wire _11722_;
  wire _11723_;
  wire _11724_;
  wire _11725_;
  wire _11726_;
  wire _11727_;
  wire _11728_;
  wire _11729_;
  wire _11730_;
  wire _11731_;
  wire _11732_;
  wire _11733_;
  wire _11734_;
  wire _11735_;
  wire _11736_;
  wire _11737_;
  wire _11738_;
  wire _11739_;
  wire _11740_;
  wire _11741_;
  wire _11742_;
  wire _11743_;
  wire _11744_;
  wire _11745_;
  wire _11746_;
  wire _11747_;
  wire _11748_;
  wire _11749_;
  wire _11750_;
  wire _11751_;
  wire _11752_;
  wire _11753_;
  wire _11754_;
  wire _11755_;
  wire _11756_;
  wire _11757_;
  wire _11758_;
  wire _11759_;
  wire _11760_;
  wire _11761_;
  wire _11762_;
  wire _11763_;
  wire _11764_;
  wire _11765_;
  wire _11766_;
  wire _11767_;
  wire _11768_;
  wire _11769_;
  wire _11770_;
  wire _11771_;
  wire _11772_;
  wire _11773_;
  wire _11774_;
  wire _11775_;
  wire _11776_;
  wire _11777_;
  wire _11778_;
  wire _11779_;
  wire _11780_;
  wire _11781_;
  wire _11782_;
  wire _11783_;
  wire _11784_;
  wire _11785_;
  wire _11786_;
  wire _11787_;
  wire _11788_;
  wire _11789_;
  wire _11790_;
  wire _11791_;
  wire _11792_;
  wire _11793_;
  wire _11794_;
  wire _11795_;
  wire _11796_;
  wire _11797_;
  wire _11798_;
  wire _11799_;
  wire _11800_;
  wire _11801_;
  wire _11802_;
  wire _11803_;
  wire _11804_;
  wire _11805_;
  wire _11806_;
  wire _11807_;
  wire _11808_;
  wire _11809_;
  wire _11810_;
  wire _11811_;
  wire _11812_;
  wire _11813_;
  wire _11814_;
  wire _11815_;
  wire _11816_;
  wire _11817_;
  wire _11818_;
  wire _11819_;
  wire _11820_;
  wire _11821_;
  wire _11822_;
  wire _11823_;
  wire _11824_;
  wire _11825_;
  wire _11826_;
  wire _11827_;
  wire _11828_;
  wire _11829_;
  wire _11830_;
  wire _11831_;
  wire _11832_;
  wire _11833_;
  wire _11834_;
  wire _11835_;
  wire _11836_;
  wire _11837_;
  wire _11838_;
  wire _11839_;
  wire _11840_;
  wire _11841_;
  wire _11842_;
  wire _11843_;
  wire _11844_;
  wire _11845_;
  wire _11846_;
  wire _11847_;
  wire _11848_;
  wire _11849_;
  wire _11850_;
  wire _11851_;
  wire _11852_;
  wire _11853_;
  wire _11854_;
  wire _11855_;
  wire _11856_;
  wire _11857_;
  wire _11858_;
  wire _11859_;
  wire _11860_;
  wire _11861_;
  wire _11862_;
  wire _11863_;
  wire _11864_;
  wire _11865_;
  wire _11866_;
  wire _11867_;
  wire _11868_;
  wire _11869_;
  wire _11870_;
  wire _11871_;
  wire _11872_;
  wire _11873_;
  wire _11874_;
  wire _11875_;
  wire _11876_;
  wire _11877_;
  wire _11878_;
  wire _11879_;
  wire _11880_;
  wire _11881_;
  wire _11882_;
  wire _11883_;
  wire _11884_;
  wire _11885_;
  wire _11886_;
  wire _11887_;
  wire _11888_;
  wire _11889_;
  wire _11890_;
  wire _11891_;
  wire _11892_;
  wire _11893_;
  wire _11894_;
  wire _11895_;
  wire _11896_;
  wire _11897_;
  wire _11898_;
  wire _11899_;
  wire _11900_;
  wire _11901_;
  wire _11902_;
  wire _11903_;
  wire _11904_;
  wire _11905_;
  wire _11906_;
  wire _11907_;
  wire _11908_;
  wire _11909_;
  wire _11910_;
  wire _11911_;
  wire _11912_;
  wire _11913_;
  wire _11914_;
  wire _11915_;
  wire _11916_;
  wire _11917_;
  wire _11918_;
  wire _11919_;
  wire _11920_;
  wire _11921_;
  wire _11922_;
  wire _11923_;
  wire _11924_;
  wire _11925_;
  wire _11926_;
  wire _11927_;
  wire _11928_;
  wire _11929_;
  wire _11930_;
  wire _11931_;
  wire _11932_;
  wire _11933_;
  wire _11934_;
  wire _11935_;
  wire _11936_;
  wire _11937_;
  wire _11938_;
  wire _11939_;
  wire _11940_;
  wire _11941_;
  wire _11942_;
  wire _11943_;
  wire _11944_;
  wire _11945_;
  wire _11946_;
  wire _11947_;
  wire _11948_;
  wire _11949_;
  wire _11950_;
  wire _11951_;
  wire _11952_;
  wire _11953_;
  wire _11954_;
  wire _11955_;
  wire _11956_;
  wire _11957_;
  wire _11958_;
  wire _11959_;
  wire _11960_;
  wire _11961_;
  wire _11962_;
  wire _11963_;
  wire _11964_;
  wire _11965_;
  wire _11966_;
  wire _11967_;
  wire _11968_;
  wire _11969_;
  wire _11970_;
  wire _11971_;
  wire _11972_;
  wire _11973_;
  wire _11974_;
  wire _11975_;
  wire _11976_;
  wire _11977_;
  wire _11978_;
  wire _11979_;
  wire _11980_;
  wire _11981_;
  wire _11982_;
  wire _11983_;
  wire _11984_;
  wire _11985_;
  wire _11986_;
  wire _11987_;
  wire _11988_;
  wire _11989_;
  wire _11990_;
  wire _11991_;
  wire _11992_;
  wire _11993_;
  wire _11994_;
  wire _11995_;
  wire _11996_;
  wire _11997_;
  wire _11998_;
  wire _11999_;
  wire _12000_;
  wire _12001_;
  wire _12002_;
  wire _12003_;
  wire _12004_;
  wire _12005_;
  wire _12006_;
  wire _12007_;
  wire _12008_;
  wire _12009_;
  wire _12010_;
  wire _12011_;
  wire _12012_;
  wire _12013_;
  wire _12014_;
  wire _12015_;
  wire _12016_;
  wire _12017_;
  wire _12018_;
  wire _12019_;
  wire _12020_;
  wire _12021_;
  wire _12022_;
  wire _12023_;
  wire _12024_;
  wire _12025_;
  wire _12026_;
  wire _12027_;
  wire _12028_;
  wire _12029_;
  wire _12030_;
  wire _12031_;
  wire _12032_;
  wire _12033_;
  wire _12034_;
  wire _12035_;
  wire _12036_;
  wire _12037_;
  wire _12038_;
  wire _12039_;
  wire _12040_;
  wire _12041_;
  wire _12042_;
  wire _12043_;
  wire _12044_;
  wire _12045_;
  wire _12046_;
  wire _12047_;
  wire _12048_;
  wire _12049_;
  wire _12050_;
  wire _12051_;
  wire _12052_;
  wire _12053_;
  wire _12054_;
  wire _12055_;
  wire _12056_;
  wire _12057_;
  wire _12058_;
  wire _12059_;
  wire _12060_;
  wire _12061_;
  wire _12062_;
  wire _12063_;
  wire _12064_;
  wire _12065_;
  wire _12066_;
  wire _12067_;
  wire _12068_;
  wire _12069_;
  wire _12070_;
  wire _12071_;
  wire _12072_;
  wire _12073_;
  wire _12074_;
  wire _12075_;
  wire _12076_;
  wire _12077_;
  wire _12078_;
  wire _12079_;
  wire _12080_;
  wire _12081_;
  wire _12082_;
  wire _12083_;
  wire _12084_;
  wire _12085_;
  wire _12086_;
  wire _12087_;
  wire _12088_;
  wire _12089_;
  wire _12090_;
  wire _12091_;
  wire _12092_;
  wire _12093_;
  wire _12094_;
  wire _12095_;
  wire _12096_;
  wire _12097_;
  wire _12098_;
  wire _12099_;
  wire _12100_;
  wire _12101_;
  wire _12102_;
  wire _12103_;
  wire _12104_;
  wire _12105_;
  wire _12106_;
  wire _12107_;
  wire _12108_;
  wire _12109_;
  wire _12110_;
  wire _12111_;
  wire _12112_;
  wire _12113_;
  wire _12114_;
  wire _12115_;
  wire _12116_;
  wire _12117_;
  wire _12118_;
  wire _12119_;
  wire _12120_;
  wire _12121_;
  wire _12122_;
  wire _12123_;
  wire _12124_;
  wire _12125_;
  wire _12126_;
  wire _12127_;
  wire _12128_;
  wire _12129_;
  wire _12130_;
  wire _12131_;
  wire _12132_;
  wire _12133_;
  wire _12134_;
  wire _12135_;
  wire _12136_;
  wire _12137_;
  wire _12138_;
  wire _12139_;
  wire _12140_;
  wire _12141_;
  wire _12142_;
  wire _12143_;
  wire _12144_;
  wire _12145_;
  wire _12146_;
  wire _12147_;
  wire _12148_;
  wire _12149_;
  wire _12150_;
  wire _12151_;
  wire _12152_;
  wire _12153_;
  wire _12154_;
  wire _12155_;
  wire _12156_;
  wire _12157_;
  wire _12158_;
  wire _12159_;
  wire _12160_;
  wire _12161_;
  wire _12162_;
  wire _12163_;
  wire _12164_;
  wire _12165_;
  wire _12166_;
  wire _12167_;
  wire _12168_;
  wire _12169_;
  wire _12170_;
  wire _12171_;
  wire _12172_;
  wire _12173_;
  wire _12174_;
  wire _12175_;
  wire _12176_;
  wire _12177_;
  wire _12178_;
  wire _12179_;
  wire _12180_;
  wire _12181_;
  wire _12182_;
  wire _12183_;
  wire _12184_;
  wire _12185_;
  wire _12186_;
  wire _12187_;
  wire _12188_;
  wire _12189_;
  wire _12190_;
  wire _12191_;
  wire _12192_;
  wire _12193_;
  wire _12194_;
  wire _12195_;
  wire _12196_;
  wire _12197_;
  wire _12198_;
  wire _12199_;
  wire _12200_;
  wire _12201_;
  wire _12202_;
  wire _12203_;
  wire _12204_;
  wire _12205_;
  wire _12206_;
  wire _12207_;
  wire _12208_;
  wire _12209_;
  wire _12210_;
  wire _12211_;
  wire _12212_;
  wire _12213_;
  wire _12214_;
  wire _12215_;
  wire _12216_;
  wire _12217_;
  wire _12218_;
  wire _12219_;
  wire _12220_;
  wire _12221_;
  wire _12222_;
  wire _12223_;
  wire _12224_;
  wire _12225_;
  wire _12226_;
  wire _12227_;
  wire _12228_;
  wire _12229_;
  wire _12230_;
  wire _12231_;
  wire _12232_;
  wire _12233_;
  wire _12234_;
  wire _12235_;
  wire _12236_;
  wire _12237_;
  wire _12238_;
  wire _12239_;
  wire _12240_;
  wire _12241_;
  wire _12242_;
  wire _12243_;
  wire _12244_;
  wire _12245_;
  wire _12246_;
  wire _12247_;
  wire _12248_;
  wire _12249_;
  wire _12250_;
  wire _12251_;
  wire _12252_;
  wire _12253_;
  wire _12254_;
  wire _12255_;
  wire _12256_;
  wire _12257_;
  wire _12258_;
  wire _12259_;
  wire _12260_;
  wire _12261_;
  wire _12262_;
  wire _12263_;
  wire _12264_;
  wire _12265_;
  wire _12266_;
  wire _12267_;
  wire _12268_;
  wire _12269_;
  wire _12270_;
  wire _12271_;
  wire _12272_;
  wire _12273_;
  wire _12274_;
  wire _12275_;
  wire _12276_;
  wire _12277_;
  wire _12278_;
  wire _12279_;
  wire _12280_;
  wire _12281_;
  wire _12282_;
  wire _12283_;
  wire _12284_;
  wire _12285_;
  wire _12286_;
  wire _12287_;
  wire _12288_;
  wire _12289_;
  wire _12290_;
  wire _12291_;
  wire _12292_;
  wire _12293_;
  wire _12294_;
  wire _12295_;
  wire _12296_;
  wire _12297_;
  wire _12298_;
  wire _12299_;
  wire _12300_;
  wire _12301_;
  wire _12302_;
  wire _12303_;
  wire _12304_;
  wire _12305_;
  wire _12306_;
  wire _12307_;
  wire _12308_;
  wire _12309_;
  wire _12310_;
  wire _12311_;
  wire _12312_;
  wire _12313_;
  wire _12314_;
  wire _12315_;
  wire _12316_;
  wire _12317_;
  wire _12318_;
  wire _12319_;
  wire _12320_;
  wire _12321_;
  wire _12322_;
  wire _12323_;
  wire _12324_;
  wire _12325_;
  wire _12326_;
  wire _12327_;
  wire _12328_;
  wire _12329_;
  wire _12330_;
  wire _12331_;
  wire _12332_;
  wire _12333_;
  wire _12334_;
  wire _12335_;
  wire _12336_;
  wire _12337_;
  wire _12338_;
  wire _12339_;
  wire _12340_;
  wire _12341_;
  wire _12342_;
  wire _12343_;
  wire _12344_;
  wire _12345_;
  wire _12346_;
  wire _12347_;
  wire _12348_;
  wire _12349_;
  wire _12350_;
  wire _12351_;
  wire _12352_;
  wire _12353_;
  wire _12354_;
  wire _12355_;
  wire _12356_;
  wire _12357_;
  wire _12358_;
  wire _12359_;
  wire _12360_;
  wire _12361_;
  wire _12362_;
  wire _12363_;
  wire _12364_;
  wire _12365_;
  wire _12366_;
  wire _12367_;
  wire _12368_;
  wire _12369_;
  wire _12370_;
  wire _12371_;
  wire _12372_;
  wire _12373_;
  wire _12374_;
  wire _12375_;
  wire _12376_;
  wire _12377_;
  wire _12378_;
  wire _12379_;
  wire _12380_;
  wire _12381_;
  wire _12382_;
  wire _12383_;
  wire _12384_;
  wire _12385_;
  wire _12386_;
  wire _12387_;
  wire _12388_;
  wire _12389_;
  wire _12390_;
  wire _12391_;
  wire _12392_;
  wire _12393_;
  wire _12394_;
  wire _12395_;
  wire _12396_;
  wire _12397_;
  wire _12398_;
  wire _12399_;
  wire _12400_;
  wire _12401_;
  wire _12402_;
  wire _12403_;
  wire _12404_;
  wire _12405_;
  wire _12406_;
  wire _12407_;
  wire _12408_;
  wire _12409_;
  wire _12410_;
  wire _12411_;
  wire _12412_;
  wire _12413_;
  wire _12414_;
  wire _12415_;
  wire _12416_;
  wire _12417_;
  wire _12418_;
  wire _12419_;
  wire _12420_;
  wire _12421_;
  wire _12422_;
  wire _12423_;
  wire _12424_;
  wire _12425_;
  wire _12426_;
  wire _12427_;
  wire _12428_;
  wire _12429_;
  wire _12430_;
  wire _12431_;
  wire _12432_;
  wire _12433_;
  wire _12434_;
  wire _12435_;
  wire _12436_;
  wire _12437_;
  wire _12438_;
  wire _12439_;
  wire _12440_;
  wire _12441_;
  wire _12442_;
  wire _12443_;
  wire _12444_;
  wire _12445_;
  wire _12446_;
  wire _12447_;
  wire _12448_;
  wire _12449_;
  wire _12450_;
  wire _12451_;
  wire _12452_;
  wire _12453_;
  wire _12454_;
  wire _12455_;
  wire _12456_;
  wire _12457_;
  wire _12458_;
  wire _12459_;
  wire _12460_;
  wire _12461_;
  wire _12462_;
  wire _12463_;
  wire _12464_;
  wire _12465_;
  wire _12466_;
  wire _12467_;
  wire _12468_;
  wire _12469_;
  wire _12470_;
  wire _12471_;
  wire _12472_;
  wire _12473_;
  wire _12474_;
  wire _12475_;
  wire _12476_;
  wire _12477_;
  wire _12478_;
  wire _12479_;
  wire _12480_;
  wire _12481_;
  wire _12482_;
  wire _12483_;
  wire _12484_;
  wire _12485_;
  wire _12486_;
  wire _12487_;
  wire _12488_;
  wire _12489_;
  wire _12490_;
  wire _12491_;
  wire _12492_;
  wire _12493_;
  wire _12494_;
  wire _12495_;
  wire _12496_;
  wire _12497_;
  wire _12498_;
  wire _12499_;
  wire _12500_;
  wire _12501_;
  wire _12502_;
  wire _12503_;
  wire _12504_;
  wire _12505_;
  wire _12506_;
  wire _12507_;
  wire _12508_;
  wire _12509_;
  wire _12510_;
  wire _12511_;
  wire _12512_;
  wire _12513_;
  wire _12514_;
  wire _12515_;
  wire _12516_;
  wire _12517_;
  wire _12518_;
  wire _12519_;
  wire _12520_;
  wire _12521_;
  wire _12522_;
  wire _12523_;
  wire _12524_;
  wire _12525_;
  wire _12526_;
  wire _12527_;
  wire _12528_;
  wire _12529_;
  wire _12530_;
  wire _12531_;
  wire _12532_;
  wire _12533_;
  wire _12534_;
  wire _12535_;
  wire _12536_;
  wire _12537_;
  wire _12538_;
  wire _12539_;
  wire _12540_;
  wire _12541_;
  wire _12542_;
  wire _12543_;
  wire _12544_;
  wire _12545_;
  wire _12546_;
  wire _12547_;
  wire _12548_;
  wire _12549_;
  wire _12550_;
  wire _12551_;
  wire _12552_;
  wire _12553_;
  wire _12554_;
  wire _12555_;
  wire _12556_;
  wire _12557_;
  wire _12558_;
  wire _12559_;
  wire _12560_;
  wire _12561_;
  wire _12562_;
  wire _12563_;
  wire _12564_;
  wire _12565_;
  wire _12566_;
  wire _12567_;
  wire _12568_;
  wire _12569_;
  wire _12570_;
  wire _12571_;
  wire _12572_;
  wire _12573_;
  wire _12574_;
  wire _12575_;
  wire _12576_;
  wire _12577_;
  wire _12578_;
  wire _12579_;
  wire _12580_;
  wire _12581_;
  wire _12582_;
  wire _12583_;
  wire _12584_;
  wire _12585_;
  wire _12586_;
  wire _12587_;
  wire _12588_;
  wire _12589_;
  wire _12590_;
  wire _12591_;
  wire _12592_;
  wire _12593_;
  wire _12594_;
  wire _12595_;
  wire _12596_;
  wire _12597_;
  wire _12598_;
  wire _12599_;
  wire _12600_;
  wire _12601_;
  wire _12602_;
  wire _12603_;
  wire _12604_;
  wire _12605_;
  wire _12606_;
  wire _12607_;
  wire _12608_;
  wire _12609_;
  wire _12610_;
  wire _12611_;
  wire _12612_;
  wire _12613_;
  wire _12614_;
  wire _12615_;
  wire _12616_;
  wire _12617_;
  wire _12618_;
  wire _12619_;
  wire _12620_;
  wire _12621_;
  wire _12622_;
  wire _12623_;
  wire _12624_;
  wire _12625_;
  wire _12626_;
  wire _12627_;
  wire _12628_;
  wire _12629_;
  wire _12630_;
  wire _12631_;
  wire _12632_;
  wire _12633_;
  wire _12634_;
  wire _12635_;
  wire _12636_;
  wire _12637_;
  wire _12638_;
  wire _12639_;
  wire _12640_;
  wire _12641_;
  wire _12642_;
  wire _12643_;
  wire _12644_;
  wire _12645_;
  wire _12646_;
  wire _12647_;
  wire _12648_;
  wire _12649_;
  wire _12650_;
  wire _12651_;
  wire _12652_;
  wire _12653_;
  wire _12654_;
  wire _12655_;
  wire _12656_;
  wire _12657_;
  wire _12658_;
  wire _12659_;
  wire _12660_;
  wire _12661_;
  wire _12662_;
  wire _12663_;
  wire _12664_;
  wire _12665_;
  wire _12666_;
  wire _12667_;
  wire _12668_;
  wire _12669_;
  wire _12670_;
  wire _12671_;
  wire _12672_;
  wire _12673_;
  wire _12674_;
  wire _12675_;
  wire _12676_;
  wire _12677_;
  wire _12678_;
  wire _12679_;
  wire _12680_;
  wire _12681_;
  wire _12682_;
  wire _12683_;
  wire _12684_;
  wire _12685_;
  wire _12686_;
  wire _12687_;
  wire _12688_;
  wire _12689_;
  wire _12690_;
  wire _12691_;
  wire _12692_;
  wire _12693_;
  wire _12694_;
  wire _12695_;
  wire _12696_;
  wire _12697_;
  wire _12698_;
  wire _12699_;
  wire _12700_;
  wire _12701_;
  wire _12702_;
  wire _12703_;
  wire _12704_;
  wire _12705_;
  wire _12706_;
  wire _12707_;
  wire _12708_;
  wire _12709_;
  wire _12710_;
  wire _12711_;
  wire _12712_;
  wire _12713_;
  wire _12714_;
  wire _12715_;
  wire _12716_;
  wire _12717_;
  wire _12718_;
  wire _12719_;
  wire _12720_;
  wire _12721_;
  wire _12722_;
  wire _12723_;
  wire _12724_;
  wire _12725_;
  wire _12726_;
  wire _12727_;
  wire _12728_;
  wire _12729_;
  wire _12730_;
  wire _12731_;
  wire _12732_;
  wire _12733_;
  wire _12734_;
  wire _12735_;
  wire _12736_;
  wire _12737_;
  wire _12738_;
  wire _12739_;
  wire _12740_;
  wire _12741_;
  wire _12742_;
  wire _12743_;
  wire _12744_;
  wire _12745_;
  wire _12746_;
  wire _12747_;
  wire _12748_;
  wire _12749_;
  wire _12750_;
  wire _12751_;
  wire _12752_;
  wire _12753_;
  wire _12754_;
  wire _12755_;
  wire _12756_;
  wire _12757_;
  wire _12758_;
  wire _12759_;
  wire _12760_;
  wire _12761_;
  wire _12762_;
  wire _12763_;
  wire _12764_;
  wire _12765_;
  wire _12766_;
  wire _12767_;
  wire _12768_;
  wire _12769_;
  wire _12770_;
  wire _12771_;
  wire _12772_;
  wire _12773_;
  wire _12774_;
  wire _12775_;
  wire _12776_;
  wire _12777_;
  wire _12778_;
  wire _12779_;
  wire _12780_;
  wire _12781_;
  wire _12782_;
  wire _12783_;
  wire _12784_;
  wire _12785_;
  wire _12786_;
  wire _12787_;
  wire _12788_;
  wire _12789_;
  wire _12790_;
  wire _12791_;
  wire _12792_;
  wire _12793_;
  wire _12794_;
  wire _12795_;
  wire _12796_;
  wire _12797_;
  wire _12798_;
  wire _12799_;
  wire _12800_;
  wire _12801_;
  wire _12802_;
  wire _12803_;
  wire _12804_;
  wire _12805_;
  wire _12806_;
  wire _12807_;
  wire _12808_;
  wire _12809_;
  wire _12810_;
  wire _12811_;
  wire _12812_;
  wire _12813_;
  wire _12814_;
  wire _12815_;
  wire _12816_;
  wire _12817_;
  wire _12818_;
  wire _12819_;
  wire _12820_;
  wire _12821_;
  wire _12822_;
  wire _12823_;
  wire _12824_;
  wire _12825_;
  wire _12826_;
  wire _12827_;
  wire _12828_;
  wire _12829_;
  wire _12830_;
  wire _12831_;
  wire _12832_;
  wire _12833_;
  wire _12834_;
  wire _12835_;
  wire _12836_;
  wire _12837_;
  wire _12838_;
  wire _12839_;
  wire _12840_;
  wire _12841_;
  wire _12842_;
  wire _12843_;
  wire _12844_;
  wire _12845_;
  wire _12846_;
  wire _12847_;
  wire _12848_;
  wire _12849_;
  wire _12850_;
  wire _12851_;
  wire _12852_;
  wire _12853_;
  wire _12854_;
  wire _12855_;
  wire _12856_;
  wire _12857_;
  wire _12858_;
  wire _12859_;
  wire _12860_;
  wire _12861_;
  wire _12862_;
  wire _12863_;
  wire _12864_;
  wire _12865_;
  wire _12866_;
  wire _12867_;
  wire _12868_;
  wire _12869_;
  wire _12870_;
  wire _12871_;
  wire _12872_;
  wire _12873_;
  wire _12874_;
  wire _12875_;
  wire _12876_;
  wire _12877_;
  wire _12878_;
  wire _12879_;
  wire _12880_;
  wire _12881_;
  wire _12882_;
  wire _12883_;
  wire _12884_;
  wire _12885_;
  wire _12886_;
  wire _12887_;
  wire _12888_;
  wire _12889_;
  wire _12890_;
  wire _12891_;
  wire _12892_;
  wire _12893_;
  wire _12894_;
  wire _12895_;
  wire _12896_;
  wire _12897_;
  wire _12898_;
  wire _12899_;
  wire _12900_;
  wire _12901_;
  wire _12902_;
  wire _12903_;
  wire _12904_;
  wire _12905_;
  wire _12906_;
  wire _12907_;
  wire _12908_;
  wire _12909_;
  wire _12910_;
  wire _12911_;
  wire _12912_;
  wire _12913_;
  wire _12914_;
  wire _12915_;
  wire _12916_;
  wire _12917_;
  wire _12918_;
  wire _12919_;
  wire _12920_;
  wire _12921_;
  wire _12922_;
  wire _12923_;
  wire _12924_;
  wire _12925_;
  wire _12926_;
  wire _12927_;
  wire _12928_;
  wire _12929_;
  wire _12930_;
  wire _12931_;
  wire _12932_;
  wire _12933_;
  wire _12934_;
  wire _12935_;
  wire _12936_;
  wire _12937_;
  wire _12938_;
  wire _12939_;
  wire _12940_;
  wire _12941_;
  wire _12942_;
  wire _12943_;
  wire _12944_;
  wire _12945_;
  wire _12946_;
  wire _12947_;
  wire _12948_;
  wire _12949_;
  wire _12950_;
  wire _12951_;
  wire _12952_;
  wire _12953_;
  wire _12954_;
  wire _12955_;
  wire _12956_;
  wire _12957_;
  wire _12958_;
  wire _12959_;
  wire _12960_;
  wire _12961_;
  wire _12962_;
  wire _12963_;
  wire _12964_;
  wire _12965_;
  wire _12966_;
  wire _12967_;
  wire _12968_;
  wire _12969_;
  wire _12970_;
  wire _12971_;
  wire _12972_;
  wire _12973_;
  wire _12974_;
  wire _12975_;
  wire _12976_;
  wire _12977_;
  wire _12978_;
  wire _12979_;
  wire _12980_;
  wire _12981_;
  wire _12982_;
  wire _12983_;
  wire _12984_;
  wire _12985_;
  wire _12986_;
  wire _12987_;
  wire _12988_;
  wire _12989_;
  wire _12990_;
  wire _12991_;
  wire _12992_;
  wire _12993_;
  wire _12994_;
  wire _12995_;
  wire _12996_;
  wire _12997_;
  wire _12998_;
  wire _12999_;
  wire _13000_;
  wire _13001_;
  wire _13002_;
  wire _13003_;
  wire _13004_;
  wire _13005_;
  wire _13006_;
  wire _13007_;
  wire _13008_;
  wire _13009_;
  wire _13010_;
  wire _13011_;
  wire _13012_;
  wire _13013_;
  wire _13014_;
  wire _13015_;
  wire _13016_;
  wire _13017_;
  wire _13018_;
  wire _13019_;
  wire _13020_;
  wire _13021_;
  wire _13022_;
  wire _13023_;
  wire _13024_;
  wire _13025_;
  wire _13026_;
  wire _13027_;
  wire _13028_;
  wire _13029_;
  wire _13030_;
  wire _13031_;
  wire _13032_;
  wire _13033_;
  wire _13034_;
  wire _13035_;
  wire _13036_;
  wire _13037_;
  wire _13038_;
  wire _13039_;
  wire _13040_;
  wire _13041_;
  wire _13042_;
  wire _13043_;
  wire _13044_;
  wire _13045_;
  wire _13046_;
  wire _13047_;
  wire _13048_;
  wire _13049_;
  wire _13050_;
  wire _13051_;
  wire _13052_;
  wire _13053_;
  wire _13054_;
  wire _13055_;
  wire _13056_;
  wire _13057_;
  wire _13058_;
  wire _13059_;
  wire _13060_;
  wire _13061_;
  wire _13062_;
  wire _13063_;
  wire _13064_;
  wire _13065_;
  wire _13066_;
  wire _13067_;
  wire _13068_;
  wire _13069_;
  wire _13070_;
  wire _13071_;
  wire _13072_;
  wire _13073_;
  wire _13074_;
  wire _13075_;
  wire _13076_;
  wire _13077_;
  wire _13078_;
  wire _13079_;
  wire _13080_;
  wire _13081_;
  wire _13082_;
  wire _13083_;
  wire _13084_;
  wire _13085_;
  wire _13086_;
  wire _13087_;
  wire _13088_;
  wire _13089_;
  wire _13090_;
  wire _13091_;
  wire _13092_;
  wire _13093_;
  wire _13094_;
  wire _13095_;
  wire _13096_;
  wire _13097_;
  wire _13098_;
  wire _13099_;
  wire _13100_;
  wire _13101_;
  wire _13102_;
  wire _13103_;
  wire _13104_;
  wire _13105_;
  wire _13106_;
  wire _13107_;
  wire _13108_;
  wire _13109_;
  wire _13110_;
  wire _13111_;
  wire _13112_;
  wire _13113_;
  wire _13114_;
  wire _13115_;
  wire _13116_;
  wire _13117_;
  wire _13118_;
  wire _13119_;
  wire _13120_;
  wire _13121_;
  wire _13122_;
  wire _13123_;
  wire _13124_;
  wire _13125_;
  wire _13126_;
  wire _13127_;
  wire _13128_;
  wire _13129_;
  wire _13130_;
  wire _13131_;
  wire _13132_;
  wire _13133_;
  wire _13134_;
  wire _13135_;
  wire _13136_;
  wire _13137_;
  wire _13138_;
  wire _13139_;
  wire _13140_;
  wire _13141_;
  wire _13142_;
  wire _13143_;
  wire _13144_;
  wire _13145_;
  wire _13146_;
  wire _13147_;
  wire _13148_;
  wire _13149_;
  wire _13150_;
  wire _13151_;
  wire _13152_;
  wire _13153_;
  wire _13154_;
  wire _13155_;
  wire _13156_;
  wire _13157_;
  wire _13158_;
  wire _13159_;
  wire _13160_;
  wire _13161_;
  wire _13162_;
  wire _13163_;
  wire _13164_;
  wire _13165_;
  wire _13166_;
  wire _13167_;
  wire _13168_;
  wire _13169_;
  wire _13170_;
  wire _13171_;
  wire _13172_;
  wire _13173_;
  wire _13174_;
  wire _13175_;
  wire _13176_;
  wire _13177_;
  wire _13178_;
  wire _13179_;
  wire _13180_;
  wire _13181_;
  wire _13182_;
  wire _13183_;
  wire _13184_;
  wire _13185_;
  wire _13186_;
  wire _13187_;
  wire _13188_;
  wire _13189_;
  wire _13190_;
  wire _13191_;
  wire _13192_;
  wire _13193_;
  wire _13194_;
  wire _13195_;
  wire _13196_;
  wire _13197_;
  wire _13198_;
  wire _13199_;
  wire _13200_;
  wire _13201_;
  wire _13202_;
  wire _13203_;
  wire _13204_;
  wire _13205_;
  wire _13206_;
  wire _13207_;
  wire _13208_;
  wire _13209_;
  wire _13210_;
  wire _13211_;
  wire _13212_;
  wire _13213_;
  wire _13214_;
  wire _13215_;
  wire _13216_;
  wire _13217_;
  wire _13218_;
  wire _13219_;
  wire _13220_;
  wire _13221_;
  wire _13222_;
  wire _13223_;
  wire _13224_;
  wire _13225_;
  wire _13226_;
  wire _13227_;
  wire _13228_;
  wire _13229_;
  wire _13230_;
  wire _13231_;
  wire _13232_;
  wire _13233_;
  wire _13234_;
  wire _13235_;
  wire _13236_;
  wire _13237_;
  wire _13238_;
  wire _13239_;
  wire _13240_;
  wire _13241_;
  wire _13242_;
  wire _13243_;
  wire _13244_;
  wire _13245_;
  wire _13246_;
  wire _13247_;
  wire _13248_;
  wire _13249_;
  wire _13250_;
  wire _13251_;
  wire _13252_;
  wire _13253_;
  wire _13254_;
  wire _13255_;
  wire _13256_;
  wire _13257_;
  wire _13258_;
  wire _13259_;
  wire _13260_;
  wire _13261_;
  wire _13262_;
  wire _13263_;
  wire _13264_;
  wire _13265_;
  wire _13266_;
  wire _13267_;
  wire _13268_;
  wire _13269_;
  wire _13270_;
  wire _13271_;
  wire _13272_;
  wire _13273_;
  wire _13274_;
  wire _13275_;
  wire _13276_;
  wire _13277_;
  wire _13278_;
  wire _13279_;
  wire _13280_;
  wire _13281_;
  wire _13282_;
  wire _13283_;
  wire _13284_;
  wire _13285_;
  wire _13286_;
  wire _13287_;
  wire _13288_;
  wire _13289_;
  wire _13290_;
  wire _13291_;
  wire _13292_;
  wire _13293_;
  wire _13294_;
  wire _13295_;
  wire _13296_;
  wire _13297_;
  wire _13298_;
  wire _13299_;
  wire _13300_;
  wire _13301_;
  wire _13302_;
  wire _13303_;
  wire _13304_;
  wire _13305_;
  wire _13306_;
  wire _13307_;
  wire _13308_;
  wire _13309_;
  wire _13310_;
  wire _13311_;
  wire _13312_;
  wire _13313_;
  wire _13314_;
  wire _13315_;
  wire _13316_;
  wire _13317_;
  wire _13318_;
  wire _13319_;
  wire _13320_;
  wire _13321_;
  wire _13322_;
  wire _13323_;
  wire _13324_;
  wire _13325_;
  wire _13326_;
  wire _13327_;
  wire _13328_;
  wire _13329_;
  wire _13330_;
  wire _13331_;
  wire _13332_;
  wire _13333_;
  wire _13334_;
  wire _13335_;
  wire _13336_;
  wire _13337_;
  wire _13338_;
  wire _13339_;
  wire _13340_;
  wire _13341_;
  wire _13342_;
  wire _13343_;
  wire _13344_;
  wire _13345_;
  wire _13346_;
  wire _13347_;
  wire _13348_;
  wire _13349_;
  wire _13350_;
  wire _13351_;
  wire _13352_;
  wire _13353_;
  wire _13354_;
  wire _13355_;
  wire _13356_;
  wire _13357_;
  wire _13358_;
  wire _13359_;
  wire _13360_;
  wire _13361_;
  wire _13362_;
  wire _13363_;
  wire _13364_;
  wire _13365_;
  wire _13366_;
  wire _13367_;
  wire _13368_;
  wire _13369_;
  wire _13370_;
  wire _13371_;
  wire _13372_;
  wire _13373_;
  wire _13374_;
  wire _13375_;
  wire _13376_;
  wire _13377_;
  wire _13378_;
  wire _13379_;
  wire _13380_;
  wire _13381_;
  wire _13382_;
  wire _13383_;
  wire _13384_;
  wire _13385_;
  wire _13386_;
  wire _13387_;
  wire _13388_;
  wire _13389_;
  wire _13390_;
  wire _13391_;
  wire _13392_;
  wire _13393_;
  wire _13394_;
  wire _13395_;
  wire _13396_;
  wire _13397_;
  wire _13398_;
  wire _13399_;
  wire _13400_;
  wire _13401_;
  wire _13402_;
  wire _13403_;
  wire _13404_;
  wire _13405_;
  wire _13406_;
  wire _13407_;
  wire _13408_;
  wire _13409_;
  wire _13410_;
  wire _13411_;
  wire _13412_;
  wire _13413_;
  wire _13414_;
  wire _13415_;
  wire _13416_;
  wire _13417_;
  wire _13418_;
  wire _13419_;
  wire _13420_;
  wire _13421_;
  wire _13422_;
  wire _13423_;
  wire _13424_;
  wire _13425_;
  wire _13426_;
  wire _13427_;
  wire _13428_;
  wire _13429_;
  wire _13430_;
  wire _13431_;
  wire _13432_;
  wire _13433_;
  wire _13434_;
  wire _13435_;
  wire _13436_;
  wire _13437_;
  wire _13438_;
  wire _13439_;
  wire _13440_;
  wire _13441_;
  wire _13442_;
  wire _13443_;
  wire _13444_;
  wire _13445_;
  wire _13446_;
  wire _13447_;
  wire _13448_;
  wire _13449_;
  wire _13450_;
  wire _13451_;
  wire _13452_;
  wire _13453_;
  wire _13454_;
  wire _13455_;
  wire _13456_;
  wire _13457_;
  wire _13458_;
  wire _13459_;
  wire _13460_;
  wire _13461_;
  wire _13462_;
  wire _13463_;
  wire _13464_;
  wire _13465_;
  wire _13466_;
  wire _13467_;
  wire _13468_;
  wire _13469_;
  wire _13470_;
  wire _13471_;
  wire _13472_;
  wire _13473_;
  wire _13474_;
  wire _13475_;
  wire _13476_;
  wire _13477_;
  wire _13478_;
  wire _13479_;
  wire _13480_;
  wire _13481_;
  wire _13482_;
  wire _13483_;
  wire _13484_;
  wire _13485_;
  wire _13486_;
  wire _13487_;
  wire _13488_;
  wire _13489_;
  wire _13490_;
  wire _13491_;
  wire _13492_;
  wire _13493_;
  wire _13494_;
  wire _13495_;
  wire _13496_;
  wire _13497_;
  wire _13498_;
  wire _13499_;
  wire _13500_;
  wire _13501_;
  wire _13502_;
  wire _13503_;
  wire _13504_;
  wire _13505_;
  wire _13506_;
  wire _13507_;
  wire _13508_;
  wire _13509_;
  wire _13510_;
  wire _13511_;
  wire _13512_;
  wire _13513_;
  wire _13514_;
  wire _13515_;
  wire _13516_;
  wire _13517_;
  wire _13518_;
  wire _13519_;
  wire _13520_;
  wire _13521_;
  wire _13522_;
  wire _13523_;
  wire _13524_;
  wire _13525_;
  wire _13526_;
  wire _13527_;
  wire _13528_;
  wire _13529_;
  wire _13530_;
  wire _13531_;
  wire _13532_;
  wire _13533_;
  wire _13534_;
  wire _13535_;
  wire _13536_;
  wire _13537_;
  wire _13538_;
  wire _13539_;
  wire _13540_;
  wire _13541_;
  wire _13542_;
  wire _13543_;
  wire _13544_;
  wire _13545_;
  wire _13546_;
  wire _13547_;
  wire _13548_;
  wire _13549_;
  wire _13550_;
  wire _13551_;
  wire _13552_;
  wire _13553_;
  wire _13554_;
  wire _13555_;
  wire _13556_;
  wire _13557_;
  wire _13558_;
  wire _13559_;
  wire _13560_;
  wire _13561_;
  wire _13562_;
  wire _13563_;
  wire _13564_;
  wire _13565_;
  wire _13566_;
  wire _13567_;
  wire _13568_;
  wire _13569_;
  wire _13570_;
  wire _13571_;
  wire _13572_;
  wire _13573_;
  wire _13574_;
  wire _13575_;
  wire _13576_;
  wire _13577_;
  wire _13578_;
  wire _13579_;
  wire _13580_;
  wire _13581_;
  wire _13582_;
  wire _13583_;
  wire _13584_;
  wire _13585_;
  wire _13586_;
  wire _13587_;
  wire _13588_;
  wire _13589_;
  wire _13590_;
  wire _13591_;
  wire _13592_;
  wire _13593_;
  wire _13594_;
  wire _13595_;
  wire _13596_;
  wire _13597_;
  wire _13598_;
  wire _13599_;
  wire _13600_;
  wire _13601_;
  wire _13602_;
  wire _13603_;
  wire _13604_;
  wire _13605_;
  wire _13606_;
  wire _13607_;
  wire _13608_;
  wire _13609_;
  wire _13610_;
  wire _13611_;
  wire _13612_;
  wire _13613_;
  wire _13614_;
  wire _13615_;
  wire _13616_;
  wire _13617_;
  wire _13618_;
  wire _13619_;
  wire _13620_;
  wire _13621_;
  wire _13622_;
  wire _13623_;
  wire _13624_;
  wire _13625_;
  wire _13626_;
  wire _13627_;
  wire _13628_;
  wire _13629_;
  wire _13630_;
  wire _13631_;
  wire _13632_;
  wire _13633_;
  wire _13634_;
  wire _13635_;
  wire _13636_;
  wire _13637_;
  wire _13638_;
  wire _13639_;
  wire _13640_;
  wire _13641_;
  wire _13642_;
  wire _13643_;
  wire _13644_;
  wire _13645_;
  wire _13646_;
  wire _13647_;
  wire _13648_;
  wire _13649_;
  wire _13650_;
  wire _13651_;
  wire _13652_;
  wire _13653_;
  wire _13654_;
  wire _13655_;
  wire _13656_;
  wire _13657_;
  wire _13658_;
  wire _13659_;
  wire _13660_;
  wire _13661_;
  wire _13662_;
  wire _13663_;
  wire _13664_;
  wire _13665_;
  wire _13666_;
  wire _13667_;
  wire _13668_;
  wire _13669_;
  wire _13670_;
  wire _13671_;
  wire _13672_;
  wire _13673_;
  wire _13674_;
  wire _13675_;
  wire _13676_;
  wire _13677_;
  wire _13678_;
  wire _13679_;
  wire _13680_;
  wire _13681_;
  wire _13682_;
  wire _13683_;
  wire _13684_;
  wire _13685_;
  wire _13686_;
  wire _13687_;
  wire _13688_;
  wire _13689_;
  wire _13690_;
  wire _13691_;
  wire _13692_;
  wire _13693_;
  wire _13694_;
  wire _13695_;
  wire _13696_;
  wire _13697_;
  wire _13698_;
  wire _13699_;
  wire _13700_;
  wire _13701_;
  wire _13702_;
  wire _13703_;
  wire _13704_;
  wire _13705_;
  wire _13706_;
  wire _13707_;
  wire _13708_;
  wire _13709_;
  wire _13710_;
  wire _13711_;
  wire _13712_;
  wire _13713_;
  wire _13714_;
  wire _13715_;
  wire _13716_;
  wire _13717_;
  wire _13718_;
  wire _13719_;
  wire _13720_;
  wire _13721_;
  wire _13722_;
  wire _13723_;
  wire _13724_;
  wire _13725_;
  wire _13726_;
  wire _13727_;
  wire _13728_;
  wire _13729_;
  wire _13730_;
  wire _13731_;
  wire _13732_;
  wire _13733_;
  wire _13734_;
  wire _13735_;
  wire _13736_;
  wire _13737_;
  wire _13738_;
  wire _13739_;
  wire _13740_;
  wire _13741_;
  wire _13742_;
  wire _13743_;
  wire _13744_;
  wire _13745_;
  wire _13746_;
  wire _13747_;
  wire _13748_;
  wire _13749_;
  wire _13750_;
  wire _13751_;
  wire _13752_;
  wire _13753_;
  wire _13754_;
  wire _13755_;
  wire _13756_;
  wire _13757_;
  wire _13758_;
  wire _13759_;
  wire _13760_;
  wire _13761_;
  wire _13762_;
  wire _13763_;
  wire _13764_;
  wire _13765_;
  wire _13766_;
  wire _13767_;
  wire _13768_;
  wire _13769_;
  wire _13770_;
  wire _13771_;
  wire _13772_;
  wire _13773_;
  wire _13774_;
  wire _13775_;
  wire _13776_;
  wire _13777_;
  wire _13778_;
  wire _13779_;
  wire _13780_;
  wire _13781_;
  wire _13782_;
  wire _13783_;
  wire _13784_;
  wire _13785_;
  wire _13786_;
  wire _13787_;
  wire _13788_;
  wire _13789_;
  wire _13790_;
  wire _13791_;
  wire _13792_;
  wire _13793_;
  wire _13794_;
  wire _13795_;
  wire _13796_;
  wire _13797_;
  wire _13798_;
  wire _13799_;
  wire _13800_;
  wire _13801_;
  wire _13802_;
  wire _13803_;
  wire _13804_;
  wire _13805_;
  wire _13806_;
  wire _13807_;
  wire _13808_;
  wire _13809_;
  wire _13810_;
  wire _13811_;
  wire _13812_;
  wire _13813_;
  wire _13814_;
  wire _13815_;
  wire _13816_;
  wire _13817_;
  wire _13818_;
  wire _13819_;
  wire _13820_;
  wire _13821_;
  wire _13822_;
  wire _13823_;
  wire _13824_;
  wire _13825_;
  wire _13826_;
  wire _13827_;
  wire _13828_;
  wire _13829_;
  wire _13830_;
  wire _13831_;
  wire _13832_;
  wire _13833_;
  wire _13834_;
  wire _13835_;
  wire _13836_;
  wire _13837_;
  wire _13838_;
  wire _13839_;
  wire _13840_;
  wire _13841_;
  wire _13842_;
  wire _13843_;
  wire _13844_;
  wire _13845_;
  wire _13846_;
  wire _13847_;
  wire _13848_;
  wire _13849_;
  wire _13850_;
  wire _13851_;
  wire _13852_;
  wire _13853_;
  wire _13854_;
  wire _13855_;
  wire _13856_;
  wire _13857_;
  wire _13858_;
  wire _13859_;
  wire _13860_;
  wire _13861_;
  wire _13862_;
  wire _13863_;
  wire _13864_;
  wire _13865_;
  wire _13866_;
  wire _13867_;
  wire _13868_;
  wire _13869_;
  wire _13870_;
  wire _13871_;
  wire _13872_;
  wire _13873_;
  wire _13874_;
  wire _13875_;
  wire _13876_;
  wire _13877_;
  wire _13878_;
  wire _13879_;
  wire _13880_;
  wire _13881_;
  wire _13882_;
  wire _13883_;
  wire _13884_;
  wire _13885_;
  wire _13886_;
  wire _13887_;
  wire _13888_;
  wire _13889_;
  wire _13890_;
  wire _13891_;
  wire _13892_;
  wire _13893_;
  wire _13894_;
  wire _13895_;
  wire _13896_;
  wire _13897_;
  wire _13898_;
  wire _13899_;
  wire _13900_;
  wire _13901_;
  wire _13902_;
  wire _13903_;
  wire _13904_;
  wire _13905_;
  wire _13906_;
  wire _13907_;
  wire _13908_;
  wire _13909_;
  wire _13910_;
  wire _13911_;
  wire _13912_;
  wire _13913_;
  wire _13914_;
  wire _13915_;
  wire _13916_;
  wire _13917_;
  wire _13918_;
  wire _13919_;
  wire _13920_;
  wire _13921_;
  wire _13922_;
  wire _13923_;
  wire _13924_;
  wire _13925_;
  wire _13926_;
  wire _13927_;
  wire _13928_;
  wire _13929_;
  wire _13930_;
  wire _13931_;
  wire _13932_;
  wire _13933_;
  wire _13934_;
  wire _13935_;
  wire _13936_;
  wire _13937_;
  wire _13938_;
  wire _13939_;
  wire _13940_;
  wire _13941_;
  wire _13942_;
  wire _13943_;
  wire _13944_;
  wire _13945_;
  wire _13946_;
  wire _13947_;
  wire _13948_;
  wire _13949_;
  wire _13950_;
  wire _13951_;
  wire _13952_;
  wire _13953_;
  wire _13954_;
  wire _13955_;
  wire _13956_;
  wire _13957_;
  wire _13958_;
  wire _13959_;
  wire _13960_;
  wire _13961_;
  wire _13962_;
  wire _13963_;
  wire _13964_;
  wire _13965_;
  wire _13966_;
  wire _13967_;
  wire _13968_;
  wire _13969_;
  wire _13970_;
  wire _13971_;
  wire _13972_;
  wire _13973_;
  wire _13974_;
  wire _13975_;
  wire _13976_;
  wire _13977_;
  wire _13978_;
  wire _13979_;
  wire _13980_;
  wire _13981_;
  wire _13982_;
  wire _13983_;
  wire _13984_;
  wire _13985_;
  wire _13986_;
  wire _13987_;
  wire _13988_;
  wire _13989_;
  wire _13990_;
  wire _13991_;
  wire _13992_;
  wire _13993_;
  wire _13994_;
  wire _13995_;
  wire _13996_;
  wire _13997_;
  wire _13998_;
  wire _13999_;
  wire _14000_;
  wire _14001_;
  wire _14002_;
  wire _14003_;
  wire _14004_;
  wire _14005_;
  wire _14006_;
  wire _14007_;
  wire _14008_;
  wire _14009_;
  wire _14010_;
  wire _14011_;
  wire _14012_;
  wire _14013_;
  wire _14014_;
  wire _14015_;
  wire _14016_;
  wire _14017_;
  wire _14018_;
  wire _14019_;
  wire _14020_;
  wire _14021_;
  wire _14022_;
  wire _14023_;
  wire _14024_;
  wire _14025_;
  wire _14026_;
  wire _14027_;
  wire _14028_;
  wire _14029_;
  wire _14030_;
  wire _14031_;
  wire _14032_;
  wire _14033_;
  wire _14034_;
  wire _14035_;
  wire _14036_;
  wire _14037_;
  wire _14038_;
  wire _14039_;
  wire _14040_;
  wire _14041_;
  wire _14042_;
  wire _14043_;
  wire _14044_;
  wire _14045_;
  wire _14046_;
  wire _14047_;
  wire _14048_;
  wire _14049_;
  wire _14050_;
  wire _14051_;
  wire _14052_;
  wire _14053_;
  wire _14054_;
  wire _14055_;
  wire _14056_;
  wire _14057_;
  wire _14058_;
  wire _14059_;
  wire _14060_;
  wire _14061_;
  wire _14062_;
  wire _14063_;
  wire _14064_;
  wire _14065_;
  wire _14066_;
  wire _14067_;
  wire _14068_;
  wire _14069_;
  wire _14070_;
  wire _14071_;
  wire _14072_;
  wire _14073_;
  wire _14074_;
  wire _14075_;
  wire _14076_;
  wire _14077_;
  wire _14078_;
  wire _14079_;
  wire _14080_;
  wire _14081_;
  wire _14082_;
  wire _14083_;
  wire _14084_;
  wire _14085_;
  wire _14086_;
  wire _14087_;
  wire _14088_;
  wire _14089_;
  wire _14090_;
  wire _14091_;
  wire _14092_;
  wire _14093_;
  wire _14094_;
  wire _14095_;
  wire _14096_;
  wire _14097_;
  wire _14098_;
  wire _14099_;
  wire _14100_;
  wire _14101_;
  wire _14102_;
  wire _14103_;
  wire _14104_;
  wire _14105_;
  wire _14106_;
  wire _14107_;
  wire _14108_;
  wire _14109_;
  wire _14110_;
  wire _14111_;
  wire _14112_;
  wire _14113_;
  wire _14114_;
  wire _14115_;
  wire _14116_;
  wire _14117_;
  wire _14118_;
  wire _14119_;
  wire _14120_;
  wire _14121_;
  wire _14122_;
  wire _14123_;
  wire _14124_;
  wire _14125_;
  wire _14126_;
  wire _14127_;
  wire _14128_;
  wire _14129_;
  wire _14130_;
  wire _14131_;
  wire _14132_;
  wire _14133_;
  wire _14134_;
  wire _14135_;
  wire _14136_;
  wire _14137_;
  wire _14138_;
  wire _14139_;
  wire _14140_;
  wire _14141_;
  wire _14142_;
  wire _14143_;
  wire _14144_;
  wire _14145_;
  wire _14146_;
  wire _14147_;
  wire _14148_;
  wire _14149_;
  wire _14150_;
  wire _14151_;
  wire _14152_;
  wire _14153_;
  wire _14154_;
  wire _14155_;
  wire _14156_;
  wire _14157_;
  wire _14158_;
  wire _14159_;
  wire _14160_;
  wire _14161_;
  wire _14162_;
  wire _14163_;
  wire _14164_;
  wire _14165_;
  wire _14166_;
  wire _14167_;
  wire _14168_;
  wire _14169_;
  wire _14170_;
  wire _14171_;
  wire _14172_;
  wire _14173_;
  wire _14174_;
  wire _14175_;
  wire _14176_;
  wire _14177_;
  wire _14178_;
  wire _14179_;
  wire _14180_;
  wire _14181_;
  wire _14182_;
  wire _14183_;
  wire _14184_;
  wire _14185_;
  wire _14186_;
  wire _14187_;
  wire _14188_;
  wire _14189_;
  wire _14190_;
  wire _14191_;
  wire _14192_;
  wire _14193_;
  wire _14194_;
  wire _14195_;
  wire _14196_;
  wire _14197_;
  wire _14198_;
  wire _14199_;
  wire _14200_;
  wire _14201_;
  wire _14202_;
  wire _14203_;
  wire _14204_;
  wire _14205_;
  wire _14206_;
  wire _14207_;
  wire _14208_;
  wire _14209_;
  wire _14210_;
  wire _14211_;
  wire _14212_;
  wire _14213_;
  wire _14214_;
  wire _14215_;
  wire _14216_;
  wire _14217_;
  wire _14218_;
  wire _14219_;
  wire _14220_;
  wire _14221_;
  wire _14222_;
  wire _14223_;
  wire _14224_;
  wire _14225_;
  wire _14226_;
  wire _14227_;
  wire _14228_;
  wire _14229_;
  wire _14230_;
  wire _14231_;
  wire _14232_;
  wire _14233_;
  wire _14234_;
  wire _14235_;
  wire _14236_;
  wire _14237_;
  wire _14238_;
  wire _14239_;
  wire _14240_;
  wire _14241_;
  wire _14242_;
  wire _14243_;
  wire _14244_;
  wire _14245_;
  wire _14246_;
  wire _14247_;
  wire _14248_;
  wire _14249_;
  wire _14250_;
  wire _14251_;
  wire _14252_;
  wire _14253_;
  wire _14254_;
  wire _14255_;
  wire _14256_;
  wire _14257_;
  wire _14258_;
  wire _14259_;
  wire _14260_;
  wire _14261_;
  wire _14262_;
  wire _14263_;
  wire _14264_;
  wire _14265_;
  wire _14266_;
  wire _14267_;
  wire _14268_;
  wire _14269_;
  wire _14270_;
  wire _14271_;
  wire _14272_;
  wire _14273_;
  wire _14274_;
  wire _14275_;
  wire _14276_;
  wire _14277_;
  wire _14278_;
  wire _14279_;
  wire _14280_;
  wire _14281_;
  wire _14282_;
  wire _14283_;
  wire _14284_;
  wire _14285_;
  wire _14286_;
  wire _14287_;
  wire _14288_;
  wire _14289_;
  wire _14290_;
  wire _14291_;
  wire _14292_;
  wire _14293_;
  wire _14294_;
  wire _14295_;
  wire _14296_;
  wire _14297_;
  wire _14298_;
  wire _14299_;
  wire _14300_;
  wire _14301_;
  wire _14302_;
  wire _14303_;
  wire _14304_;
  wire _14305_;
  wire _14306_;
  wire _14307_;
  wire _14308_;
  wire _14309_;
  wire _14310_;
  wire _14311_;
  wire _14312_;
  wire _14313_;
  wire _14314_;
  wire _14315_;
  wire _14316_;
  wire _14317_;
  wire _14318_;
  wire _14319_;
  wire _14320_;
  wire _14321_;
  wire _14322_;
  wire _14323_;
  wire _14324_;
  wire _14325_;
  wire _14326_;
  wire _14327_;
  wire _14328_;
  wire _14329_;
  wire _14330_;
  wire _14331_;
  wire _14332_;
  wire _14333_;
  wire _14334_;
  wire _14335_;
  wire _14336_;
  wire _14337_;
  wire _14338_;
  wire _14339_;
  wire _14340_;
  wire _14341_;
  wire _14342_;
  wire _14343_;
  wire _14344_;
  wire _14345_;
  wire _14346_;
  wire _14347_;
  wire _14348_;
  wire _14349_;
  wire _14350_;
  wire _14351_;
  wire _14352_;
  wire _14353_;
  wire _14354_;
  wire _14355_;
  wire _14356_;
  wire _14357_;
  wire _14358_;
  wire _14359_;
  wire _14360_;
  wire _14361_;
  wire _14362_;
  wire _14363_;
  wire _14364_;
  wire _14365_;
  wire _14366_;
  wire _14367_;
  wire _14368_;
  wire _14369_;
  wire _14370_;
  wire _14371_;
  wire _14372_;
  wire _14373_;
  wire _14374_;
  wire _14375_;
  wire _14376_;
  wire _14377_;
  wire _14378_;
  wire _14379_;
  wire _14380_;
  wire _14381_;
  wire _14382_;
  wire _14383_;
  wire _14384_;
  wire _14385_;
  wire _14386_;
  wire _14387_;
  wire _14388_;
  wire _14389_;
  wire _14390_;
  wire _14391_;
  wire _14392_;
  wire _14393_;
  wire _14394_;
  wire _14395_;
  wire _14396_;
  wire _14397_;
  wire _14398_;
  wire _14399_;
  wire _14400_;
  wire _14401_;
  wire _14402_;
  wire _14403_;
  wire _14404_;
  wire _14405_;
  wire _14406_;
  wire _14407_;
  wire _14408_;
  wire _14409_;
  wire _14410_;
  wire _14411_;
  wire _14412_;
  wire _14413_;
  wire _14414_;
  wire _14415_;
  wire _14416_;
  wire _14417_;
  wire _14418_;
  wire _14419_;
  wire _14420_;
  wire _14421_;
  wire _14422_;
  wire _14423_;
  wire _14424_;
  wire _14425_;
  wire _14426_;
  wire _14427_;
  wire _14428_;
  wire _14429_;
  wire _14430_;
  wire _14431_;
  wire _14432_;
  wire _14433_;
  wire _14434_;
  wire _14435_;
  wire _14436_;
  wire _14437_;
  wire _14438_;
  wire _14439_;
  wire _14440_;
  wire _14441_;
  wire _14442_;
  wire _14443_;
  wire _14444_;
  wire _14445_;
  wire _14446_;
  wire _14447_;
  wire _14448_;
  wire _14449_;
  wire _14450_;
  wire _14451_;
  wire _14452_;
  wire _14453_;
  wire _14454_;
  wire _14455_;
  wire _14456_;
  wire _14457_;
  wire _14458_;
  wire _14459_;
  wire _14460_;
  wire _14461_;
  wire _14462_;
  wire _14463_;
  wire _14464_;
  wire _14465_;
  wire _14466_;
  wire _14467_;
  wire _14468_;
  wire _14469_;
  wire _14470_;
  wire _14471_;
  wire _14472_;
  wire _14473_;
  wire _14474_;
  wire _14475_;
  wire _14476_;
  wire _14477_;
  wire _14478_;
  wire _14479_;
  wire _14480_;
  wire _14481_;
  wire _14482_;
  wire _14483_;
  wire _14484_;
  wire _14485_;
  wire _14486_;
  wire _14487_;
  wire _14488_;
  wire _14489_;
  wire _14490_;
  wire _14491_;
  wire _14492_;
  wire _14493_;
  wire _14494_;
  wire _14495_;
  wire _14496_;
  wire _14497_;
  wire _14498_;
  wire _14499_;
  wire _14500_;
  wire _14501_;
  wire _14502_;
  wire _14503_;
  wire _14504_;
  wire _14505_;
  wire _14506_;
  wire _14507_;
  wire _14508_;
  wire _14509_;
  wire _14510_;
  wire _14511_;
  wire _14512_;
  wire _14513_;
  wire _14514_;
  wire _14515_;
  wire _14516_;
  wire _14517_;
  wire _14518_;
  wire _14519_;
  wire _14520_;
  wire _14521_;
  wire _14522_;
  wire _14523_;
  wire _14524_;
  wire _14525_;
  wire _14526_;
  wire _14527_;
  wire _14528_;
  wire _14529_;
  wire _14530_;
  wire _14531_;
  wire _14532_;
  wire _14533_;
  wire _14534_;
  wire _14535_;
  wire _14536_;
  wire _14537_;
  wire _14538_;
  wire _14539_;
  wire _14540_;
  wire _14541_;
  wire _14542_;
  wire _14543_;
  wire _14544_;
  wire _14545_;
  wire _14546_;
  wire _14547_;
  wire _14548_;
  wire _14549_;
  wire _14550_;
  wire _14551_;
  wire _14552_;
  wire _14553_;
  wire _14554_;
  wire _14555_;
  wire _14556_;
  wire _14557_;
  wire _14558_;
  wire _14559_;
  wire _14560_;
  wire _14561_;
  wire _14562_;
  wire _14563_;
  wire _14564_;
  wire _14565_;
  wire _14566_;
  wire _14567_;
  wire _14568_;
  wire _14569_;
  wire _14570_;
  wire _14571_;
  wire _14572_;
  wire _14573_;
  wire _14574_;
  wire _14575_;
  wire _14576_;
  wire _14577_;
  wire _14578_;
  wire _14579_;
  wire _14580_;
  wire _14581_;
  wire _14582_;
  wire _14583_;
  wire _14584_;
  wire _14585_;
  wire _14586_;
  wire _14587_;
  wire _14588_;
  wire _14589_;
  wire _14590_;
  wire _14591_;
  wire _14592_;
  wire _14593_;
  wire _14594_;
  wire _14595_;
  wire _14596_;
  wire _14597_;
  wire _14598_;
  wire _14599_;
  wire _14600_;
  wire _14601_;
  wire _14602_;
  wire _14603_;
  wire _14604_;
  wire _14605_;
  wire _14606_;
  wire _14607_;
  input [8:0] ABINPUT;
  input clk;
  wire [31:0] cxrom_data_out;
  wire first_instr;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.bytein3 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout0 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout1 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout2 ;
  wire [7:0] \oc8051_symbolic_cxrom1.byteout3 ;
  wire \oc8051_symbolic_cxrom1.clk ;
  wire [31:0] \oc8051_symbolic_cxrom1.cxrom_data_out ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc1 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc10 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc12 ;
  wire [15:0] \oc8051_symbolic_cxrom1.pc2 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc20 ;
  wire [3:0] \oc8051_symbolic_cxrom1.pc22 ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[0] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[10] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[11] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[12] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[13] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[14] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[15] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[1] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[2] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[3] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[4] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[5] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[6] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[7] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[8] ;
  wire [7:0] \oc8051_symbolic_cxrom1.regarray[9] ;
  wire [15:0] \oc8051_symbolic_cxrom1.regvalid ;
  wire \oc8051_symbolic_cxrom1.rst ;
  wire [31:0] \oc8051_symbolic_cxrom1.word_in ;
  wire [8:0] \oc8051_top_1.ABINPUT ;
  wire [7:0] \oc8051_top_1.acc ;
  wire \oc8051_top_1.bit_data ;
  wire [31:0] \oc8051_top_1.cxrom_data_out ;
  wire \oc8051_top_1.cy ;
  wire [1:0] \oc8051_top_1.cy_sel ;
  wire [7:0] \oc8051_top_1.dptr_hi ;
  wire [7:0] \oc8051_top_1.dptr_lo ;
  wire [31:0] \oc8051_top_1.idat_onchip ;
  wire \oc8051_top_1.int_ack ;
  wire [7:0] \oc8051_top_1.int_src ;
  wire \oc8051_top_1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.mem_act ;
  wire \oc8051_top_1.oc8051_alu1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.divsrc2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.des2 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div0 ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.div1 ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.div_out ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_div1.rst ;
  wire [5:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div ;
  wire [7:0] \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle ;
  wire \oc8051_top_1.oc8051_alu1.oc8051_mul1.rst ;
  wire [15:0] \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul ;
  wire \oc8051_top_1.oc8051_alu1.rst ;
  wire \oc8051_top_1.oc8051_alu1.srcAc ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.acc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.clk ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.dptr ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op1_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op2_r ;
  wire [7:0] \oc8051_top_1.oc8051_alu_src_sel1.op3_r ;
  wire [15:0] \oc8051_top_1.oc8051_alu_src_sel1.pc ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_alu_src_sel1.sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_alu_src_sel1.sel2 ;
  wire \oc8051_top_1.oc8051_alu_src_sel1.sel3 ;
  wire [7:0] \oc8051_top_1.oc8051_comp1.acc ;
  wire \oc8051_top_1.oc8051_comp1.cy ;
  wire \oc8051_top_1.oc8051_cy_select1.cy_in ;
  wire [1:0] \oc8051_top_1.oc8051_cy_select1.cy_sel ;
  wire [3:0] \oc8051_top_1.oc8051_decoder1.alu_op ;
  wire \oc8051_top_1.oc8051_decoder1.clk ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.cy_sel ;
  wire \oc8051_top_1.oc8051_decoder1.irom_out_of_rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_decoder1.op ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.psw_set ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.ram_wr_sel ;
  wire \oc8051_top_1.oc8051_decoder1.rst ;
  wire [2:0] \oc8051_top_1.oc8051_decoder1.src_sel1 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.src_sel2 ;
  wire \oc8051_top_1.oc8051_decoder1.src_sel3 ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.state ;
  wire \oc8051_top_1.oc8051_decoder1.wait_data ;
  wire \oc8051_top_1.oc8051_decoder1.wr ;
  wire [1:0] \oc8051_top_1.oc8051_decoder1.wr_sfr ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[0] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[1] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[2] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[3] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[4] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[5] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[6] ;
  wire [7:0] \oc8051_top_1.oc8051_indi_addr1.buff[7] ;
  wire \oc8051_top_1.oc8051_indi_addr1.clk ;
  wire \oc8051_top_1.oc8051_indi_addr1.rst ;
  wire \oc8051_top_1.oc8051_indi_addr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.acc ;
  wire \oc8051_top_1.oc8051_memory_interface1.bit_in ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.cdata ;
  wire \oc8051_top_1.oc8051_memory_interface1.cdone ;
  wire \oc8051_top_1.oc8051_memory_interface1.clk ;
  wire \oc8051_top_1.oc8051_memory_interface1.dmem_wait ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.dptr ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.iadr_t ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_cur ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_old ;
  wire [31:0] \oc8051_top_1.oc8051_memory_interface1.idat_onchip ;
  wire \oc8051_top_1.oc8051_memory_interface1.imem_wait ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm2_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.imm_r ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.in_ram ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.int_ack_t ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_v ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.int_vec_buff ;
  wire \oc8051_top_1.oc8051_memory_interface1.istb_t ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.mem_act ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op2_buff ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.op3_buff ;
  wire [2:0] \oc8051_top_1.oc8051_memory_interface1.op_pos ;
  wire \oc8051_top_1.oc8051_memory_interface1.out_of_rst ;
  wire [3:0] \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_buf ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_log_prev ;
  wire [15:0] \oc8051_top_1.oc8051_memory_interface1.pc_out ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_addr_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rd_ind ;
  wire \oc8051_top_1.oc8051_memory_interface1.reti ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.ri_r ;
  wire [4:0] \oc8051_top_1.oc8051_memory_interface1.rn_r ;
  wire \oc8051_top_1.oc8051_memory_interface1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_memory_interface1.sfr ;
  wire \oc8051_top_1.oc8051_memory_interface1.sfr_bit ;
  wire \oc8051_top_1.oc8051_rom1.clk ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.cxrom_data_out ;
  wire [31:0] \oc8051_top_1.oc8051_rom1.data_o ;
  wire \oc8051_top_1.oc8051_rom1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.acc ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.b_reg ;
  wire \oc8051_top_1.oc8051_sfr1.bit_out ;
  wire \oc8051_top_1.oc8051_sfr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.cy ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dat0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.dptr_lo ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ie ;
  wire \oc8051_top_1.oc8051_sfr1.int_ack ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.ip ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.ack ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip ;
  wire [5:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] ;
  wire [2:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk ;
  wire [7:1] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.p ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_psw1.set ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd ;
  wire [11:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp ;
  wire [10:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done ;
  wire \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p0_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p1_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p2_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_in ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.p3_out ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.pcon ;
  wire \oc8051_top_1.oc8051_sfr1.pres_ow ;
  wire [3:0] \oc8051_top_1.oc8051_sfr1.prescaler ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.psw ;
  wire [1:0] \oc8051_top_1.oc8051_sfr1.psw_set ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2h ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.rcap2l ;
  wire \oc8051_top_1.oc8051_sfr1.rclk ;
  wire \oc8051_top_1.oc8051_sfr1.reti ;
  wire \oc8051_top_1.oc8051_sfr1.rst ;
  wire \oc8051_top_1.oc8051_sfr1.rxd ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.sbuf ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.scon ;
  wire \oc8051_top_1.oc8051_sfr1.srcAc ;
  wire \oc8051_top_1.oc8051_sfr1.t0 ;
  wire \oc8051_top_1.oc8051_sfr1.t1 ;
  wire \oc8051_top_1.oc8051_sfr1.t2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.t2con ;
  wire \oc8051_top_1.oc8051_sfr1.t2ex ;
  wire \oc8051_top_1.oc8051_sfr1.tc2_int ;
  wire \oc8051_top_1.oc8051_sfr1.tclk ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tcon ;
  wire \oc8051_top_1.oc8051_sfr1.tf0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.th2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl0 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl1 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tl2 ;
  wire [7:0] \oc8051_top_1.oc8051_sfr1.tmod ;
  wire \oc8051_top_1.oc8051_sfr1.tr0 ;
  wire \oc8051_top_1.oc8051_sfr1.tr1 ;
  wire \oc8051_top_1.oc8051_sfr1.uart_int ;
  wire \oc8051_top_1.oc8051_sfr1.wait_data ;
  wire \oc8051_top_1.oc8051_sfr1.wr_bit_r ;
  wire [7:0] \oc8051_top_1.p0_i ;
  wire [7:0] \oc8051_top_1.p0_o ;
  wire [7:0] \oc8051_top_1.p1_i ;
  wire [7:0] \oc8051_top_1.p1_o ;
  wire [7:0] \oc8051_top_1.p2_i ;
  wire [7:0] \oc8051_top_1.p2_o ;
  wire [7:0] \oc8051_top_1.p3_i ;
  wire [7:0] \oc8051_top_1.p3_o ;
  wire [15:0] \oc8051_top_1.pc ;
  wire [15:0] \oc8051_top_1.pc_log ;
  wire [15:0] \oc8051_top_1.pc_log_prev ;
  wire [1:0] \oc8051_top_1.psw_set ;
  wire [7:0] \oc8051_top_1.ram_data ;
  wire \oc8051_top_1.rd_ind ;
  wire \oc8051_top_1.reti ;
  wire \oc8051_top_1.rxd_i ;
  wire \oc8051_top_1.sfr_bit ;
  wire [7:0] \oc8051_top_1.sfr_out ;
  wire \oc8051_top_1.srcAc ;
  wire [2:0] \oc8051_top_1.src_sel1 ;
  wire [1:0] \oc8051_top_1.src_sel2 ;
  wire \oc8051_top_1.src_sel3 ;
  wire \oc8051_top_1.t0_i ;
  wire \oc8051_top_1.t1_i ;
  wire \oc8051_top_1.t2_i ;
  wire \oc8051_top_1.t2ex_i ;
  wire \oc8051_top_1.wait_data ;
  wire \oc8051_top_1.wb_clk_i ;
  wire \oc8051_top_1.wb_rst_i ;
  input [7:0] p0_in;
  wire [7:0] p0_out;
  input [7:0] p1_in;
  wire [7:0] p1_out;
  input [7:0] p2_in;
  wire [7:0] p2_out;
  input [7:0] p3_in;
  wire [7:0] p3_out;
  wire [15:0] pc1;
  wire [15:0] pc1_plus_2;
  wire [15:0] pc2;
  output property_invalid;
  input rst;
  input rxd_i;
  input t0_i;
  input t1_i;
  input t2_i;
  input t2ex_i;
  input [31:0] word_in;
  nor (_06295_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  not (_06296_, _06295_);
  and (_06297_, _06296_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr );
  and (_06298_, _06297_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  and (_06299_, _06298_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_06300_, _06298_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  nor (_06301_, _06300_, _06299_);
  and (_06302_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_06303_, _06302_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  and (_06304_, _06303_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  and (_06305_, _06304_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  not (_06306_, _06305_);
  not (_06307_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  not (_06308_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06309_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _06308_);
  and (_06310_, _06309_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0]);
  and (_06311_, _06310_, _06307_);
  not (_06312_, _06311_);
  nor (_06313_, _06304_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_06314_, _06313_, _06312_);
  and (_06315_, _06314_, _06306_);
  not (_06316_, _06315_);
  not (_06317_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1]);
  and (_06318_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _06308_);
  and (_06319_, _06318_, _06317_);
  and (_06320_, _06319_, _06307_);
  and (_06321_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  nor (_06322_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_06323_, _06322_, _06317_);
  or (_06324_, _06323_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_06325_, _06324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [4]);
  nor (_06326_, _06325_, _06321_);
  and (_06327_, _06319_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_06328_, _06327_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  not (_06329_, _06328_);
  and (_06330_, _06310_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2]);
  and (_06331_, _06322_, _06309_);
  and (_06332_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [4]);
  nor (_06333_, _06332_, _06330_);
  and (_06334_, _06333_, _06329_);
  and (_06335_, _06334_, _06326_);
  and (_06336_, _06335_, _06316_);
  not (_06337_, _06336_);
  and (_06338_, _06305_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  not (_06339_, _06338_);
  nor (_06340_, _06305_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_06341_, _06340_, _06312_);
  and (_06342_, _06341_, _06339_);
  not (_06343_, _06342_);
  and (_06344_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [5]);
  and (_06345_, _06327_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  and (_06346_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  or (_06347_, _06346_, _06345_);
  or (_06348_, _06347_, _06330_);
  nor (_06349_, _06348_, _06344_);
  and (_06350_, _06349_, _06343_);
  and (_06351_, _06350_, _06337_);
  and (_06352_, _06338_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  not (_06353_, _06352_);
  nor (_06354_, _06338_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_06355_, _06354_, _06312_);
  and (_06356_, _06355_, _06353_);
  not (_06357_, _06356_);
  and (_06358_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [6]);
  and (_06359_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  and (_06360_, _06327_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or (_06361_, _06360_, _06359_);
  or (_06362_, _06361_, _06330_);
  nor (_06363_, _06362_, _06358_);
  and (_06364_, _06363_, _06357_);
  not (_06365_, _06364_);
  not (_06366_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7]);
  nor (_06367_, _06352_, _06366_);
  and (_06368_, _06352_, _06366_);
  nor (_06369_, _06368_, _06367_);
  nor (_06370_, _06369_, _06312_);
  not (_06371_, _06370_);
  and (_06372_, _06320_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  not (_06373_, _06372_);
  and (_06374_, _06327_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  not (_06375_, _06374_);
  and (_06376_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [7]);
  nor (_06377_, _06376_, _06330_);
  and (_06378_, _06377_, _06375_);
  and (_06379_, _06378_, _06373_);
  and (_06380_, _06379_, _06371_);
  nor (_06381_, _06380_, _06365_);
  and (_06382_, _06381_, _06351_);
  and (_06383_, _06327_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_06384_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  nor (_06385_, _06384_, _06383_);
  nor (_06386_, _06303_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_06387_, _06386_, _06304_);
  and (_06388_, _06387_, _06311_);
  not (_06389_, _06388_);
  and (_06390_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [3]);
  and (_06391_, _06324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [3]);
  nor (_06392_, _06391_, _06390_);
  and (_06393_, _06392_, _06389_);
  and (_06394_, _06393_, _06385_);
  not (_06395_, _06394_);
  and (_06396_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  and (_06397_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [0]);
  nor (_06398_, _06397_, _06396_);
  and (_06399_, _06327_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  not (_06400_, _06399_);
  not (_06401_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  and (_06402_, _06311_, _06401_);
  and (_06403_, _06324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [0]);
  nor (_06404_, _06403_, _06402_);
  and (_06405_, _06404_, _06400_);
  and (_06406_, _06405_, _06398_);
  not (_06407_, _06406_);
  nor (_06408_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0]);
  nor (_06409_, _06408_, _06302_);
  and (_06410_, _06409_, _06311_);
  and (_06411_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [1]);
  nor (_06412_, _06411_, _06410_);
  and (_06413_, _06327_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_06414_, _06320_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_06415_, _06324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [1]);
  or (_06416_, _06415_, _06414_);
  nor (_06417_, _06416_, _06413_);
  and (_06418_, _06417_, _06412_);
  nor (_06419_, _06302_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_06420_, _06419_, _06303_);
  and (_06421_, _06420_, _06311_);
  and (_06422_, _06331_, \oc8051_top_1.oc8051_memory_interface1.ri_r [2]);
  nor (_06423_, _06422_, _06421_);
  and (_06424_, _06327_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_06425_, _06320_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and (_06426_, _06324_, \oc8051_top_1.oc8051_memory_interface1.rn_r [2]);
  or (_06427_, _06426_, _06425_);
  nor (_06428_, _06427_, _06424_);
  and (_06430_, _06428_, _06423_);
  and (_06431_, _06430_, _06418_);
  and (_06432_, _06431_, _06407_);
  and (_06434_, _06432_, _06395_);
  and (_06435_, _06309_, _06307_);
  not (_06436_, _06435_);
  not (_06437_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_06438_, \oc8051_top_1.oc8051_decoder1.wr , _06308_);
  and (_06439_, _06438_, _06437_);
  and (_06440_, _06439_, _06436_);
  and (_06441_, _06440_, _06434_);
  and (_06442_, _06441_, _06382_);
  nor (_06443_, _06442_, rst);
  and (_14257_, _06443_, _06301_);
  not (_06444_, rst);
  and (_06445_, _06380_, _06364_);
  and (_06446_, _06445_, _06351_);
  and (_06447_, _06446_, _06434_);
  and (_06448_, _06447_, _06439_);
  not (_06449_, _06448_);
  and (_06450_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_06451_, \oc8051_top_1.oc8051_decoder1.alu_op [1], _06308_);
  and (_06452_, _06451_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_06453_, \oc8051_top_1.oc8051_decoder1.alu_op [3], _06308_);
  and (_06454_, _06453_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_06455_, _06454_, _06452_);
  and (_06456_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_06457_, _06456_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  not (_06458_, \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  and (_06459_, _06458_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  nor (_06460_, _06459_, ABINPUT[0]);
  nand (_06461_, _06458_, \oc8051_top_1.oc8051_memory_interface1.rd_addr_r );
  nor (_06462_, _06461_, \oc8051_top_1.oc8051_sfr1.bit_out );
  nor (_06463_, _06462_, _06460_);
  nor (_06464_, _06463_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  nor (_06465_, _06464_, _06457_);
  or (_06466_, _06459_, ABINPUT[6]);
  or (_06467_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  nand (_06468_, _06467_, _06466_);
  nor (_06469_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  not (_06470_, _06469_);
  or (_06472_, _06470_, _06468_);
  not (_06474_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  nand (_06475_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_06476_, _06475_, _06474_);
  not (_06477_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  not (_06478_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  nand (_06479_, _06478_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_06480_, _06479_, _06477_);
  and (_06481_, _06480_, _06476_);
  and (_06482_, _06481_, _06472_);
  not (_06483_, _06482_);
  and (_06484_, _06483_, _06465_);
  not (_06485_, \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  not (_06486_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  and (_06487_, _06486_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  and (_06488_, _06487_, _06485_);
  nand (_06489_, _06488_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  nor (_06490_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], _06485_);
  and (_06491_, _06490_, _06486_);
  nand (_06492_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  and (_06493_, _06492_, _06489_);
  nor (_06494_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_06495_, _06494_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_06496_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_06497_, _06490_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_06498_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_06499_, _06498_, _06496_);
  and (_06500_, _06499_, _06493_);
  and (_06501_, _06494_, _06486_);
  not (_06502_, _06501_);
  or (_06503_, _06502_, _06468_);
  and (_06504_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  and (_06505_, _06504_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  nand (_06506_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [5]);
  and (_06507_, _06504_, _06486_);
  nand (_06508_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_06509_, _06508_, _06506_);
  and (_06510_, _06509_, _06503_);
  and (_06511_, _06510_, _06500_);
  nor (_06512_, _06511_, _06465_);
  or (_06513_, _06512_, _06484_);
  and (_06514_, _06513_, _06455_);
  not (_06515_, _06465_);
  nand (_06516_, _06488_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  nand (_06518_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  and (_06519_, _06518_, _06516_);
  nand (_06520_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nand (_06521_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_06522_, _06521_, _06520_);
  and (_06523_, _06522_, _06519_);
  or (_06524_, _06459_, ABINPUT[5]);
  or (_06525_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  nand (_06526_, _06525_, _06524_);
  or (_06527_, _06526_, _06502_);
  nand (_06528_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [4]);
  nand (_06529_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  and (_06530_, _06529_, _06528_);
  and (_06531_, _06530_, _06527_);
  and (_06532_, _06531_, _06523_);
  not (_06534_, _06532_);
  nand (_06535_, _06488_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  nand (_06537_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  and (_06538_, _06537_, _06535_);
  and (_06539_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_06540_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_06541_, _06540_, _06539_);
  and (_06542_, _06541_, _06538_);
  or (_06543_, _06459_, ABINPUT[4]);
  or (_06544_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  nand (_06545_, _06544_, _06543_);
  or (_06546_, _06545_, _06502_);
  and (_06547_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [3]);
  and (_06548_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  nor (_06549_, _06548_, _06547_);
  and (_06550_, _06549_, _06546_);
  and (_06551_, _06550_, _06542_);
  not (_06552_, _06551_);
  nand (_06553_, _06488_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  nand (_06554_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  and (_06555_, _06554_, _06553_);
  nand (_06556_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nand (_06557_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_06558_, _06557_, _06556_);
  and (_06559_, _06558_, _06555_);
  or (_06560_, _06459_, ABINPUT[2]);
  or (_06561_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  nand (_06562_, _06561_, _06560_);
  or (_06563_, _06562_, _06502_);
  nand (_06564_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [1]);
  nand (_06565_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_06567_, _06565_, _06564_);
  and (_06568_, _06567_, _06563_);
  and (_06570_, _06568_, _06559_);
  and (_06571_, _06488_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_06572_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  nor (_06573_, _06572_, _06571_);
  and (_06574_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_06575_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_06576_, _06575_, _06574_);
  and (_06577_, _06576_, _06573_);
  or (_06578_, _06459_, ABINPUT[1]);
  or (_06579_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  and (_06580_, _06579_, _06578_);
  and (_06581_, _06580_, _06501_);
  and (_06582_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [0]);
  and (_06583_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  nor (_06584_, _06583_, _06582_);
  not (_06585_, _06584_);
  nor (_06586_, _06585_, _06581_);
  and (_06587_, _06586_, _06577_);
  nor (_06588_, _06587_, _06570_);
  nand (_06589_, _06488_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  nand (_06590_, _06491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  and (_06591_, _06590_, _06589_);
  or (_06592_, _06459_, ABINPUT[3]);
  or (_06593_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  nand (_06594_, _06593_, _06592_);
  or (_06595_, _06594_, _06502_);
  and (_06596_, _06595_, _06591_);
  nand (_06597_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nand (_06598_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_06599_, _06598_, _06597_);
  nand (_06600_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nand (_06601_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [2]);
  and (_06602_, _06601_, _06600_);
  and (_06603_, _06602_, _06599_);
  and (_06604_, _06603_, _06596_);
  not (_06605_, _06604_);
  and (_06606_, _06605_, _06588_);
  and (_06607_, _06606_, _06552_);
  and (_06608_, _06607_, _06534_);
  and (_06609_, _06608_, _06515_);
  and (_06610_, _06604_, _06570_);
  and (_06611_, _06610_, _06587_);
  and (_06612_, _06611_, _06551_);
  and (_06613_, _06612_, _06532_);
  and (_06614_, _06613_, _06465_);
  nor (_06615_, _06614_, _06609_);
  nor (_06616_, _06615_, _06511_);
  not (_06617_, _06616_);
  not (_06618_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  and (_06619_, _06451_, _06618_);
  and (_06620_, _06619_, _06454_);
  not (_06621_, _06620_);
  and (_06622_, _06615_, _06511_);
  nor (_06623_, _06622_, _06621_);
  and (_06624_, _06623_, _06617_);
  nor (_06625_, _06624_, _06514_);
  and (_06626_, \oc8051_top_1.oc8051_decoder1.alu_op [0], _06308_);
  and (_06627_, \oc8051_top_1.oc8051_decoder1.alu_op [2], _06308_);
  nor (_06628_, _06627_, _06453_);
  and (_06629_, _06628_, _06626_);
  not (_06630_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  not (_06631_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  and (_06632_, _06627_, _06631_);
  and (_06633_, _06632_, _06630_);
  nor (_06634_, _06633_, _06629_);
  not (_06635_, \oc8051_top_1.oc8051_decoder1.alu_op [2]);
  and (_06636_, _06453_, _06635_);
  and (_06637_, _06636_, _06451_);
  not (_06638_, _06637_);
  nor (_06639_, _06626_, _06451_);
  and (_06640_, _06639_, _06628_);
  and (_06641_, _06454_, _06630_);
  nor (_06642_, _06641_, _06640_);
  and (_06643_, _06642_, _06638_);
  and (_06644_, _06643_, _06634_);
  nor (_06645_, _06644_, _06511_);
  not (_06646_, _06645_);
  and (_06647_, _06639_, _06636_);
  nor (_06648_, _06511_, _06482_);
  and (_06649_, _06511_, _06482_);
  nor (_06650_, _06649_, _06648_);
  and (_06651_, _06650_, _06647_);
  not (_06652_, _06651_);
  and (_06653_, _06626_, _06630_);
  and (_06654_, _06653_, _06636_);
  not (_06655_, _06654_);
  nor (_06656_, _06655_, _06649_);
  not (_06657_, _06656_);
  and (_06658_, _06632_, _06452_);
  and (_06659_, _06658_, _06648_);
  and (_06660_, _06632_, _06619_);
  and (_06661_, _06660_, _06511_);
  nor (_06662_, _06661_, _06659_);
  and (_06663_, _06662_, _06657_);
  and (_06664_, _06663_, _06652_);
  and (_06665_, _06664_, _06646_);
  and (_06666_, _06665_, _06625_);
  nor (_06667_, _06666_, _06449_);
  or (_06668_, _06667_, _06450_);
  and (_06471_, _06668_, _06444_);
  or (_06669_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_06670_, _06395_, _06336_);
  not (_06671_, _06350_);
  nor (_06672_, _06364_, _06671_);
  and (_06673_, _06438_, _06436_);
  and (_06674_, _06673_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  not (_06675_, _06674_);
  nor (_06676_, _06675_, _06380_);
  and (_06677_, _06676_, _06672_);
  and (_06678_, _06677_, _06670_);
  or (_06679_, _06678_, _06669_);
  and (_06680_, _06628_, _06619_);
  not (_06681_, _06680_);
  nand (_06682_, _06491_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  nand (_06683_, _06488_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_06684_, _06683_, _06682_);
  and (_06685_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_06686_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  nor (_06687_, _06686_, _06685_);
  and (_06688_, _06687_, _06684_);
  or (_06689_, _06459_, ABINPUT[8]);
  or (_06690_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  nand (_06691_, _06690_, _06689_);
  or (_06692_, _06691_, _06502_);
  and (_06693_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [7]);
  and (_06694_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  nor (_06695_, _06694_, _06693_);
  and (_06696_, _06695_, _06692_);
  and (_06697_, _06696_, _06688_);
  or (_06698_, _06691_, _06470_);
  not (_06699_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  or (_06700_, _06475_, _06699_);
  not (_06701_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_06702_, _06479_, _06701_);
  and (_06703_, _06702_, _06700_);
  and (_06704_, _06703_, _06698_);
  not (_06705_, _06704_);
  and (_06706_, _06705_, _06697_);
  nor (_06707_, _06704_, _06697_);
  and (_06708_, _06704_, _06697_);
  nor (_06709_, _06708_, _06707_);
  nand (_06710_, _06488_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  nand (_06711_, _06491_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  and (_06712_, _06711_, _06710_);
  and (_06714_, _06497_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_06716_, _06495_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_06718_, _06716_, _06714_);
  and (_06720_, _06718_, _06712_);
  or (_06722_, _06459_, ABINPUT[7]);
  or (_06723_, _06461_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  nand (_06725_, _06723_, _06722_);
  or (_06727_, _06725_, _06502_);
  and (_06728_, _06505_, \oc8051_top_1.oc8051_alu_src_sel1.op1_r [6]);
  and (_06729_, _06507_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  nor (_06730_, _06729_, _06728_);
  and (_06731_, _06730_, _06727_);
  and (_06732_, _06731_, _06720_);
  or (_06733_, _06725_, _06470_);
  not (_06734_, \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  or (_06735_, _06475_, _06734_);
  not (_06736_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_06737_, _06479_, _06736_);
  and (_06738_, _06737_, _06735_);
  and (_06739_, _06738_, _06733_);
  not (_06740_, _06739_);
  nor (_06741_, _06740_, _06732_);
  nor (_06742_, _06739_, _06732_);
  and (_06743_, _06739_, _06732_);
  nor (_06744_, _06743_, _06742_);
  nor (_06745_, _06511_, _06483_);
  or (_06746_, _06526_, _06470_);
  not (_06747_, \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  or (_06748_, _06475_, _06747_);
  not (_06749_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_06750_, _06479_, _06749_);
  and (_06751_, _06750_, _06748_);
  and (_06752_, _06751_, _06746_);
  not (_06753_, _06752_);
  and (_06754_, _06753_, _06532_);
  nor (_06755_, _06754_, _06650_);
  nor (_06756_, _06755_, _06745_);
  nor (_06757_, _06756_, _06744_);
  nor (_06758_, _06757_, _06741_);
  and (_06759_, _06756_, _06744_);
  nor (_06760_, _06759_, _06757_);
  not (_06761_, _06760_);
  and (_06762_, _06754_, _06650_);
  nor (_06763_, _06762_, _06755_);
  not (_06764_, _06763_);
  nor (_06765_, _06752_, _06532_);
  and (_06766_, _06752_, _06532_);
  nor (_06767_, _06766_, _06765_);
  not (_06768_, _06767_);
  or (_06769_, _06545_, _06470_);
  not (_06770_, \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  or (_06771_, _06475_, _06770_);
  not (_06772_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_06773_, _06479_, _06772_);
  and (_06774_, _06773_, _06771_);
  and (_06775_, _06774_, _06769_);
  and (_06776_, _06775_, _06551_);
  nor (_06777_, _06775_, _06551_);
  nor (_06778_, _06777_, _06776_);
  or (_06779_, _06594_, _06470_);
  not (_06780_, \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  or (_06781_, _06475_, _06780_);
  not (_06782_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_06783_, _06479_, _06782_);
  and (_06784_, _06783_, _06781_);
  and (_06785_, _06784_, _06779_);
  nor (_06786_, _06785_, _06604_);
  and (_06787_, _06785_, _06604_);
  nor (_06788_, _06787_, _06786_);
  or (_06789_, _06562_, _06470_);
  not (_06790_, \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  or (_06791_, _06475_, _06790_);
  not (_06792_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_06793_, _06479_, _06792_);
  and (_06794_, _06793_, _06791_);
  nand (_06795_, _06794_, _06789_);
  not (_06796_, _06795_);
  nor (_06797_, _06796_, _06570_);
  and (_06798_, _06796_, _06570_);
  nor (_06799_, _06798_, _06797_);
  nand (_06800_, _06580_, _06469_);
  not (_06801_, \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  or (_06802_, _06475_, _06801_);
  not (_06803_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_06804_, _06479_, _06803_);
  and (_06805_, _06804_, _06802_);
  nand (_06806_, _06805_, _06800_);
  and (_06807_, _06806_, _06587_);
  nor (_06808_, _06807_, _06799_);
  nor (_06809_, _06795_, _06570_);
  nor (_06810_, _06809_, _06808_);
  nor (_06811_, _06810_, _06788_);
  not (_06812_, _06785_);
  nor (_06813_, _06812_, _06604_);
  nor (_06814_, _06813_, _06811_);
  nor (_06815_, _06814_, _06778_);
  and (_06816_, _06814_, _06778_);
  nor (_06817_, _06816_, _06815_);
  and (_06818_, _06810_, _06788_);
  nor (_06819_, _06818_, _06811_);
  not (_06820_, _06819_);
  and (_06821_, _06807_, _06799_);
  nor (_06822_, _06821_, _06808_);
  not (_06823_, _06822_);
  not (_06824_, _06806_);
  nor (_06825_, _06824_, _06587_);
  and (_06826_, _06824_, _06587_);
  nor (_06827_, _06826_, _06825_);
  nor (_06828_, _06827_, _06515_);
  and (_06829_, _06828_, _06823_);
  and (_06830_, _06829_, _06820_);
  not (_06831_, _06830_);
  nor (_06832_, _06831_, _06817_);
  not (_06833_, _06775_);
  or (_06834_, _06833_, _06551_);
  and (_06835_, _06833_, _06551_);
  or (_06836_, _06814_, _06835_);
  and (_06837_, _06836_, _06834_);
  or (_06838_, _06837_, _06832_);
  and (_06839_, _06838_, _06768_);
  and (_06840_, _06839_, _06764_);
  and (_06841_, _06840_, _06761_);
  nor (_06842_, _06841_, _06758_);
  nor (_06843_, _06842_, _06709_);
  nor (_06844_, _06843_, _06706_);
  nor (_06845_, _06844_, _06681_);
  not (_06846_, _06845_);
  and (_06847_, _06653_, _06628_);
  not (_06848_, _06847_);
  not (_06849_, _06744_);
  and (_06850_, _06765_, _06650_);
  nor (_06851_, _06850_, _06648_);
  nor (_06852_, _06851_, _06849_);
  not (_06853_, _06788_);
  and (_06854_, _06825_, _06799_);
  nor (_06855_, _06854_, _06797_);
  nor (_06856_, _06855_, _06853_);
  nor (_06857_, _06856_, _06786_);
  nor (_06858_, _06857_, _06778_);
  and (_06859_, _06857_, _06778_);
  nor (_06860_, _06859_, _06858_);
  and (_06861_, _06827_, _06465_);
  and (_06862_, _06861_, _06799_);
  and (_06863_, _06855_, _06853_);
  nor (_06864_, _06863_, _06856_);
  and (_06865_, _06864_, _06862_);
  not (_06866_, _06865_);
  nor (_06867_, _06866_, _06860_);
  nor (_06868_, _06857_, _06776_);
  or (_06869_, _06868_, _06777_);
  or (_06870_, _06869_, _06867_);
  and (_06871_, _06870_, _06767_);
  and (_06872_, _06871_, _06650_);
  and (_06873_, _06851_, _06849_);
  nor (_06874_, _06873_, _06852_);
  and (_06875_, _06874_, _06872_);
  or (_06876_, _06875_, _06742_);
  nor (_06877_, _06876_, _06852_);
  nor (_06878_, _06877_, _06708_);
  nor (_06879_, _06878_, _06707_);
  nor (_06880_, _06879_, _06848_);
  and (_06881_, _06732_, _06511_);
  not (_06882_, _06881_);
  and (_06883_, _06653_, _06632_);
  nor (_06884_, _06610_, _06551_);
  and (_06885_, _06884_, _06883_);
  and (_06886_, _06885_, _06534_);
  nor (_06887_, _06886_, _06882_);
  nor (_06888_, _06887_, _06697_);
  nor (_06889_, _06888_, _06465_);
  not (_06890_, _06889_);
  not (_06891_, _06883_);
  nor (_06892_, _06697_, _06515_);
  not (_06893_, _06892_);
  nor (_06894_, _06893_, _06887_);
  nor (_06895_, _06894_, _06891_);
  and (_06896_, _06895_, _06890_);
  nor (_06897_, _06465_, _06463_);
  not (_06898_, _06647_);
  and (_06899_, _06465_, _06463_);
  or (_06900_, _06899_, _06898_);
  and (_06901_, _06900_, _06655_);
  or (_06902_, _06901_, _06897_);
  not (_06903_, _06587_);
  and (_06904_, _06653_, _06454_);
  and (_06905_, _06904_, _06903_);
  and (_06906_, _06463_, _06457_);
  and (_06907_, _06636_, _06619_);
  and (_06908_, _06658_, _06463_);
  nor (_06909_, _06908_, _06907_);
  nor (_06910_, _06909_, _06906_);
  nor (_06911_, _06910_, _06905_);
  and (_06912_, _06911_, _06902_);
  and (_06913_, _06636_, _06452_);
  not (_06914_, _06697_);
  and (_06915_, _06914_, _06913_);
  nor (_06916_, _06660_, _06465_);
  not (_06917_, _06463_);
  and (_06918_, _06639_, _06454_);
  and (_06919_, _06918_, _06917_);
  nor (_06920_, _06919_, _06640_);
  and (_06921_, _06920_, _06465_);
  nor (_06922_, _06921_, _06916_);
  or (_06923_, _06922_, _06885_);
  nor (_06924_, _06923_, _06915_);
  and (_06925_, _06924_, _06912_);
  not (_06926_, _06925_);
  nor (_06927_, _06926_, _06896_);
  not (_06928_, _06927_);
  nor (_06929_, _06928_, _06880_);
  and (_06930_, _06929_, _06846_);
  not (_06931_, _06430_);
  nor (_06932_, _06418_, _06406_);
  and (_06933_, _06932_, _06931_);
  not (_06934_, _06933_);
  nor (_06935_, _06934_, _06930_);
  nand (_06936_, _06934_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  nand (_06937_, _06936_, _06678_);
  or (_06938_, _06937_, _06935_);
  and (_06939_, _06938_, _06679_);
  nor (_06940_, _06380_, _06337_);
  and (_06941_, _06940_, _06672_);
  and (_06942_, _06431_, _06406_);
  not (_06943_, _06440_);
  nor (_06944_, _06943_, _06394_);
  and (_06945_, _06944_, _06942_);
  and (_06946_, _06945_, _06941_);
  or (_06947_, _06946_, _06939_);
  and (_06948_, _06697_, _06515_);
  not (_06949_, _06948_);
  not (_06951_, _06455_);
  and (_06952_, _06704_, _06465_);
  nor (_06953_, _06952_, _06951_);
  and (_06954_, _06953_, _06949_);
  and (_06955_, _06881_, _06613_);
  nor (_06956_, _06955_, _06515_);
  not (_06957_, _06732_);
  not (_06958_, _06511_);
  and (_06959_, _06608_, _06958_);
  and (_06960_, _06959_, _06957_);
  nor (_06961_, _06960_, _06465_);
  nor (_06962_, _06961_, _06956_);
  and (_06963_, _06962_, _06914_);
  nor (_06964_, _06962_, _06914_);
  nor (_06965_, _06964_, _06963_);
  and (_06966_, _06965_, _06620_);
  nor (_06967_, _06966_, _06954_);
  and (_06968_, _06709_, _06647_);
  and (_06969_, _06707_, _06658_);
  nor (_06970_, _06708_, _06655_);
  and (_06971_, _06697_, _06660_);
  or (_06972_, _06971_, _06970_);
  or (_06973_, _06972_, _06969_);
  nor (_06974_, _06973_, _06968_);
  nor (_06975_, _06697_, _06644_);
  not (_06976_, _06975_);
  and (_06977_, _06976_, _06974_);
  and (_06978_, _06977_, _06967_);
  nand (_06979_, _06978_, _06946_);
  and (_06980_, _06979_, _06444_);
  and (_09333_, _06980_, _06947_);
  not (_06981_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set );
  and (_06982_, _06418_, _06406_);
  and (_06983_, _06982_, _06931_);
  and (_06984_, _06944_, _06983_);
  and (_06985_, _06984_, _06941_);
  and (_06986_, _06418_, _06407_);
  and (_06987_, _06986_, _06931_);
  and (_06988_, _06944_, _06987_);
  and (_06989_, _06988_, _06941_);
  nor (_06990_, _06989_, _06985_);
  nor (_06991_, _06990_, _06981_);
  and (_06992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_06993_, _06992_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_06994_, _06993_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_06995_, _06994_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_06996_, _06995_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  and (_06997_, _06996_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_06998_, _06997_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_06999_, _06998_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_07000_, _06999_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_07001_, _07000_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_07002_, _07001_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_07003_, _07002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_07004_, _07003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  and (_07005_, _07004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_07006_, _07005_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_07007_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  not (_07008_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_07009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _07008_);
  and (_07010_, _07009_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  and (_07011_, _07010_, _07007_);
  nor (_07012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not (_07013_, _07012_);
  not (_07014_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_07015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_07016_, _07015_, _07012_);
  and (_07017_, _07016_, _07014_);
  nor (_07018_, _07017_, _07013_);
  and (_07019_, _07018_, _07011_);
  and (_07020_, _07019_, _06990_);
  and (_07021_, _07020_, _07006_);
  or (_07022_, _07021_, _06991_);
  and (_09435_, _07022_, _06444_);
  nand (_07023_, _06989_, _06978_);
  and (_07024_, _07011_, _07005_);
  nor (_07025_, _07024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_07026_, _07011_, _07006_);
  nor (_07027_, _07026_, _07025_);
  and (_07028_, _07012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  not (_07029_, _07028_);
  and (_07030_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_07031_, _07030_, _07011_);
  and (_07032_, _07031_, _07006_);
  or (_07033_, _07032_, _07017_);
  or (_07034_, _07033_, _07027_);
  not (_07035_, _07017_);
  nor (_07036_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  nor (_07037_, _07036_, _06985_);
  and (_07038_, _07037_, _07034_);
  and (_07039_, _06985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_07040_, _07039_, _06989_);
  or (_07041_, _07040_, _07038_);
  and (_07042_, _07041_, _06444_);
  and (_11388_, _07042_, _07023_);
  and (_07043_, _06432_, _06394_);
  and (_07044_, _07043_, _06446_);
  and (_07045_, _07044_, _06439_);
  not (_07046_, _07045_);
  and (_07047_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  and (_07048_, _06795_, _06455_);
  and (_07049_, _06587_, _06570_);
  nor (_07050_, _07049_, _06588_);
  and (_07052_, _07050_, _06465_);
  nor (_07053_, _07050_, _06465_);
  or (_07054_, _07053_, _06621_);
  nor (_07055_, _07054_, _07052_);
  nor (_07056_, _07055_, _07048_);
  nor (_07057_, _06644_, _06570_);
  not (_07058_, _07057_);
  and (_07059_, _06799_, _06647_);
  not (_07060_, _07059_);
  nor (_07061_, _06798_, _06655_);
  not (_07062_, _07061_);
  and (_07063_, _06797_, _06658_);
  and (_07064_, _06660_, _06570_);
  nor (_07065_, _07064_, _07063_);
  and (_07066_, _07065_, _07062_);
  and (_07067_, _07066_, _07060_);
  and (_07068_, _07067_, _07058_);
  and (_07069_, _07068_, _07056_);
  not (_07070_, _07069_);
  and (_07071_, _07070_, _07045_);
  or (_07072_, _07071_, _07047_);
  and (_11722_, _07072_, _06444_);
  and (_07073_, \oc8051_top_1.oc8051_memory_interface1.reti , \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  and (_07074_, _06444_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_12487_, _07074_, _07073_);
  not (_07075_, _07073_);
  not (_07076_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc );
  not (_07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  and (_07078_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _07077_);
  and (_07079_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_07080_, _07079_, _07078_);
  and (_07081_, _07080_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  nor (_07082_, _07081_, _07076_);
  and (_07083_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_07084_, _07083_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  not (_07085_, _07084_);
  and (_07086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_07087_, _07086_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_07088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_07089_, _07088_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  nor (_07090_, _07089_, _07087_);
  and (_07091_, _07090_, _07085_);
  not (_07092_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  nor (_07093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nor (_07094_, _07093_, _07092_);
  and (_07095_, _07094_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  not (_07096_, _07095_);
  not (_07098_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  nor (_07099_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nor (_07100_, _07099_, _07098_);
  nand (_07101_, _07100_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_07102_, _07101_, _07096_);
  and (_07103_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_07104_, _07103_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  not (_07105_, _07104_);
  and (_07106_, _07105_, _07102_);
  and (_07107_, _07106_, _07091_);
  nor (_07108_, _07107_, _07082_);
  and (_07109_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _07076_);
  not (_07110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_07111_, _07094_, _07110_);
  not (_07112_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_07113_, _07100_, _07112_);
  nor (_07114_, _07113_, _07111_);
  not (_07115_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_07116_, _07103_, _07115_);
  not (_07117_, _07116_);
  not (_07118_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_07119_, _07083_, _07118_);
  not (_07120_, _07119_);
  not (_07121_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_07122_, _07086_, _07121_);
  not (_07123_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  and (_07124_, _07088_, _07123_);
  nor (_07125_, _07124_, _07122_);
  and (_07126_, _07125_, _07120_);
  and (_07127_, _07126_, _07117_);
  nand (_07128_, _07127_, _07114_);
  nand (_07130_, _07128_, _07109_);
  not (_07131_, _07130_);
  nor (_07132_, _07131_, _07108_);
  and (_07133_, _07132_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  not (_07134_, _07108_);
  nor (_07135_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  and (_07136_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1]);
  nor (_07137_, _07136_, _07135_);
  nor (_07138_, _07137_, _07134_);
  or (_07139_, _07138_, _07133_);
  and (_07140_, _07139_, _07075_);
  and (_07141_, _07137_, _07073_);
  or (_07142_, _07141_, _07140_);
  and (_12749_, _07142_, _06444_);
  nand (_07143_, _07130_, _07076_);
  or (_07144_, _07143_, _07108_);
  nand (_07145_, _07135_, _07073_);
  and (_07146_, _07145_, _06444_);
  and (_12769_, _07146_, _07144_);
  and (_07147_, _06942_, _06395_);
  and (_07148_, _07147_, _06446_);
  not (_07149_, _07044_);
  and (_07150_, _06942_, _06394_);
  and (_07151_, _07150_, _06446_);
  and (_07152_, _06350_, _06336_);
  and (_07153_, _07152_, _06445_);
  and (_07154_, _07153_, _06434_);
  nor (_07155_, _07154_, _07151_);
  nand (_07156_, _07155_, _07149_);
  nor (_07157_, _07156_, _07148_);
  not (_07158_, _06439_);
  and (_07159_, _07153_, _07150_);
  or (_07160_, _07159_, _07158_);
  or (_07161_, _07160_, _07157_);
  and (_07162_, _07161_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_07163_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_07164_, _07163_, _07156_);
  nor (_07166_, _06532_, _06465_);
  and (_07167_, _06753_, _06465_);
  or (_07168_, _07167_, _07166_);
  and (_07169_, _07168_, _06455_);
  nor (_07170_, _06607_, _06465_);
  nor (_07171_, _06612_, _06515_);
  nor (_07172_, _07171_, _07170_);
  nor (_07173_, _07172_, _06534_);
  and (_07174_, _07172_, _06534_);
  nor (_07175_, _07174_, _07173_);
  and (_07176_, _07175_, _06620_);
  nor (_07177_, _07176_, _07169_);
  nor (_07178_, _06644_, _06532_);
  not (_07179_, _07178_);
  and (_07180_, _06767_, _06647_);
  and (_07181_, _06765_, _06658_);
  nor (_07182_, _06766_, _06655_);
  and (_07183_, _06660_, _06532_);
  or (_07184_, _07183_, _07182_);
  or (_07185_, _07184_, _07181_);
  nor (_07186_, _07185_, _07180_);
  and (_07187_, _07186_, _07179_);
  and (_07188_, _07187_, _07177_);
  and (_07189_, _07148_, _06439_);
  not (_07190_, _07189_);
  nor (_07191_, _07190_, _07188_);
  or (_07192_, _07191_, _07164_);
  or (_07193_, _07192_, _07162_);
  and (_13150_, _07193_, _06444_);
  or (_07194_, _07091_, _07082_);
  nor (_07195_, _07130_, _07108_);
  not (_07196_, _07195_);
  or (_07197_, _07196_, _07126_);
  and (_07198_, _07197_, _07194_);
  nor (_07199_, _07073_, _07077_);
  not (_07200_, _07199_);
  or (_07201_, _07200_, _07198_);
  not (_07202_, _07114_);
  and (_07203_, _07202_, _07109_);
  and (_07204_, _07116_, _07109_);
  or (_07205_, _07204_, _07203_);
  or (_07206_, _07205_, _07108_);
  not (_07207_, _07106_);
  or (_07208_, _07194_, _07207_);
  and (_07209_, _07208_, _07199_);
  and (_07210_, _07209_, _07206_);
  or (_07211_, _07210_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2]);
  and (_07213_, _07211_, _06444_);
  and (_13339_, _07213_, _07201_);
  and (_07214_, _06440_, _06394_);
  and (_07215_, _07214_, _06942_);
  nor (_07216_, _06380_, _06364_);
  and (_07217_, _07216_, _06351_);
  and (_07218_, _07217_, _07215_);
  not (_07219_, _07218_);
  and (_07220_, _07219_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  nor (_07221_, _07219_, _07188_);
  nor (_07222_, _07221_, _07220_);
  nor (_07223_, _07222_, _06337_);
  and (_07224_, _07222_, _06337_);
  nor (_07225_, _07224_, _07223_);
  not (_07226_, \oc8051_top_1.oc8051_memory_interface1.dmem_wait );
  nor (_07227_, \oc8051_top_1.oc8051_memory_interface1.imem_wait , \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_07228_, _07227_, _07226_);
  nor (_07229_, \oc8051_top_1.oc8051_decoder1.state [1], \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_07230_, _07229_, _06308_);
  and (_07231_, _07230_, _07228_);
  not (_07232_, _07231_);
  not (_07233_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_07234_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  not (_07235_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  not (_07236_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  nor (_07237_, _07236_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_07238_, _07237_, _07235_);
  nand (_07239_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  and (_07240_, _07236_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nand (_07241_, _07240_, _07235_);
  not (_07242_, _07241_);
  nand (_07243_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_07244_, _07243_, _07239_);
  nor (_07245_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_07246_, _07245_, _07235_);
  nand (_07247_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  and (_07248_, _07245_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nand (_07249_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_07250_, _07249_, _07247_);
  and (_07251_, _07245_, _07235_);
  nand (_07252_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  and (_07253_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_07254_, _07253_, _07235_);
  nand (_07255_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  and (_07256_, _07255_, _07252_);
  and (_07257_, _07256_, _07250_);
  nand (_07258_, _07257_, _07244_);
  nand (_07259_, _07258_, _07234_);
  nand (_07260_, _07259_, _07233_);
  nor (_07261_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _07233_);
  not (_07262_, _07261_);
  and (_07263_, _07262_, _07260_);
  or (_07264_, _07263_, _07232_);
  not (_07265_, _07228_);
  nor (_07266_, _07230_, \oc8051_top_1.oc8051_decoder1.op [0]);
  nor (_07267_, _07266_, _07265_);
  and (_07268_, _07267_, _07264_);
  and (_07269_, _07268_, _06406_);
  not (_07270_, _07269_);
  and (_07271_, _06439_, _06431_);
  and (_07272_, _07271_, _06350_);
  and (_07273_, _07272_, _06445_);
  nor (_07274_, _07268_, _06406_);
  not (_07275_, _07274_);
  and (_07276_, _07275_, _07273_);
  and (_07277_, _07276_, _07270_);
  and (_07278_, _07219_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  nor (_07280_, _06775_, _06951_);
  nor (_07281_, _06611_, _06515_);
  nor (_07282_, _06606_, _06465_);
  nor (_07283_, _07282_, _07281_);
  and (_07284_, _07283_, _06552_);
  not (_07285_, _07284_);
  nor (_07286_, _07283_, _06552_);
  nor (_07287_, _07286_, _06621_);
  and (_07288_, _07287_, _07285_);
  nor (_07289_, _07288_, _07280_);
  nor (_07290_, _06776_, _06655_);
  and (_07291_, _06778_, _06647_);
  nor (_07292_, _07291_, _07290_);
  and (_07293_, _06777_, _06658_);
  and (_07294_, _06660_, _06551_);
  nor (_07295_, _07294_, _07293_);
  nor (_07296_, _06644_, _06551_);
  not (_07297_, _07296_);
  and (_07298_, _07297_, _07295_);
  and (_07299_, _07298_, _07292_);
  and (_07300_, _07299_, _07289_);
  nor (_07301_, _07300_, _07219_);
  nor (_07302_, _07301_, _07278_);
  and (_07303_, _07302_, _06395_);
  nor (_07304_, _07302_, _06395_);
  nor (_07305_, _07304_, _07303_);
  and (_07306_, _07305_, _07277_);
  and (_07307_, _07306_, _07225_);
  nor (_07308_, _07268_, _07302_);
  and (_07309_, _07308_, _07222_);
  and (_07310_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  not (_07311_, _07268_);
  and (_07312_, _07311_, _07302_);
  and (_07313_, _07312_, _07222_);
  and (_07314_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  nor (_07315_, _07314_, _07310_);
  not (_07316_, _07222_);
  and (_07317_, _07268_, _07302_);
  and (_07318_, _07317_, _07316_);
  and (_07319_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor (_07320_, _07311_, _07302_);
  and (_07321_, _07320_, _07316_);
  and (_07322_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  nor (_07323_, _07322_, _07319_);
  and (_07324_, _07323_, _07315_);
  and (_07325_, _07308_, _07316_);
  and (_07326_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  and (_07327_, _07312_, _07316_);
  and (_07329_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  nor (_07330_, _07329_, _07326_);
  and (_07331_, _07320_, _07222_);
  and (_07332_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  and (_07333_, _07317_, _07222_);
  and (_07334_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  nor (_07335_, _07334_, _07332_);
  and (_07336_, _07335_, _07330_);
  and (_07338_, _07336_, _07324_);
  nor (_07339_, _07338_, _07307_);
  not (_07340_, _07300_);
  and (_07341_, _07307_, _07340_);
  nor (_07342_, _07341_, _07339_);
  nor (_14055_, _07342_, rst);
  and (_07343_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  and (_07344_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  nor (_07345_, _07344_, _07343_);
  and (_07346_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_07347_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  nor (_07348_, _07347_, _07346_);
  and (_07349_, _07348_, _07345_);
  and (_07350_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [4]);
  and (_07351_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_07352_, _07351_, _07350_);
  and (_07353_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  and (_07354_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  nor (_07355_, _07354_, _07353_);
  and (_07356_, _07355_, _07352_);
  and (_07357_, _07356_, _07349_);
  nor (_07358_, _07357_, _07307_);
  not (_07359_, _07188_);
  and (_07360_, _07307_, _07359_);
  nor (_07361_, _07360_, _07358_);
  nor (_14295_, _07361_, rst);
  and (_07362_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [5]);
  and (_07363_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  nor (_07364_, _07363_, _07362_);
  and (_07365_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  and (_07366_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  nor (_07367_, _07366_, _07365_);
  and (_07368_, _07367_, _07364_);
  and (_07369_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_07370_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  nor (_07371_, _07370_, _07369_);
  and (_07372_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  and (_07373_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_07374_, _07373_, _07372_);
  and (_07375_, _07374_, _07371_);
  and (_07376_, _07375_, _07368_);
  nor (_07377_, _07376_, _07307_);
  not (_07378_, _06666_);
  and (_07379_, _07307_, _07378_);
  nor (_07380_, _07379_, _07377_);
  nor (_01145_, _07380_, rst);
  nor (_07381_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_07382_, _07381_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  not (_07383_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  and (_07384_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_07385_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  nor (_07386_, _07385_, _07384_);
  nor (_07387_, _07386_, _07076_);
  or (_07388_, _07387_, _07383_);
  and (_07389_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _07077_);
  and (_07390_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  nor (_07391_, _07390_, _07389_);
  nor (_07392_, _07391_, _07076_);
  and (_07393_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_07394_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor (_07396_, _07394_, _07393_);
  nand (_07397_, _07396_, _07392_);
  or (_07398_, _07397_, _07388_);
  and (_07399_, _07398_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_07400_, _07399_, _07382_);
  and (_07401_, _06364_, _06350_);
  and (_07402_, _07401_, _06940_);
  nor (_07403_, _06675_, _06394_);
  and (_07404_, _07403_, _06933_);
  and (_07405_, _07404_, _07402_);
  or (_07406_, _07405_, _07400_);
  and (_07407_, _07402_, _06945_);
  not (_07408_, _07407_);
  and (_07409_, _07408_, _07406_);
  nand (_07410_, _07405_, _06930_);
  and (_07411_, _07410_, _07409_);
  nor (_07412_, _07408_, _06978_);
  or (_07413_, _07412_, _07411_);
  and (_01342_, _07413_, _06444_);
  and (_07414_, _07153_, _07043_);
  nor (_07415_, _07159_, _07414_);
  and (_07416_, _07153_, _07147_);
  not (_07417_, _07416_);
  and (_07418_, _07155_, _07417_);
  and (_07419_, _07418_, _07415_);
  or (_07420_, _07419_, _07158_);
  and (_07421_, _07420_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_07422_, _07153_, _06431_);
  and (_07423_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [3]);
  and (_07424_, _07423_, _07422_);
  and (_07425_, _07151_, _06439_);
  and (_07426_, _07425_, _07340_);
  or (_07427_, _07426_, _07424_);
  or (_07428_, _07427_, _07421_);
  and (_01560_, _07428_, _06444_);
  not (_07429_, _07230_);
  nor (_07430_, _07253_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  nor (_07431_, _07430_, _07429_);
  nor (_07432_, _07431_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  and (_07433_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  not (_07434_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  nor (_07435_, _07432_, _07434_);
  or (_07436_, _07435_, _07433_);
  and (_01936_, _07436_, _06444_);
  not (_07437_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0]);
  and (_07438_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], _06308_);
  and (_07439_, _07438_, _07437_);
  and (_07440_, _06795_, _06640_);
  and (_07441_, _06913_, _06958_);
  and (_07442_, _06955_, _06697_);
  and (_07443_, _07442_, _06824_);
  and (_07444_, _07443_, _06465_);
  nor (_07445_, _06824_, _06697_);
  and (_07446_, _07445_, _06960_);
  and (_07447_, _07446_, _06515_);
  nor (_07448_, _07447_, _07444_);
  nor (_07450_, _07448_, _06795_);
  and (_07451_, _07448_, _06795_);
  nor (_07453_, _07451_, _07450_);
  nor (_07454_, _07453_, _06621_);
  nor (_07456_, _06570_, _06951_);
  or (_07457_, _07456_, _07454_);
  or (_07458_, _07457_, _07441_);
  and (_07459_, _06639_, _06632_);
  nor (_07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07461_, _07460_, _06697_);
  nor (_07462_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7]);
  not (_07463_, _07462_);
  and (_07464_, _07463_, _07461_);
  not (_07465_, _07464_);
  or (_07466_, _06806_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07467_, _06785_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_07468_, _07467_, _07466_);
  or (_07470_, _07468_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07471_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07472_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07473_, _06752_, _07472_);
  nand (_07474_, _06739_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_07475_, _07474_, _07473_);
  or (_07476_, _07475_, _07471_);
  and (_07477_, _07476_, _07470_);
  nor (_07478_, _07477_, _07465_);
  and (_07479_, _07477_, _07465_);
  nand (_07480_, _07460_, _06732_);
  nor (_07481_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6]);
  not (_07482_, _07481_);
  and (_07483_, _07482_, _07480_);
  not (_07484_, _07483_);
  and (_07486_, _06795_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07487_, _07486_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07488_, _06775_, _07472_);
  nand (_07489_, _06482_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_07490_, _07489_, _07488_);
  or (_07491_, _07490_, _07471_);
  and (_07492_, _07491_, _07487_);
  or (_07493_, _07492_, _07484_);
  nor (_07495_, _07493_, _07479_);
  nor (_07496_, _07495_, _07478_);
  nor (_07497_, _07479_, _07478_);
  nand (_07499_, _07492_, _07484_);
  and (_07500_, _07499_, _07493_);
  and (_07501_, _07500_, _07497_);
  nand (_07502_, _07460_, _06511_);
  nor (_07503_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5]);
  not (_07504_, _07503_);
  and (_07505_, _07504_, _07502_);
  not (_07506_, _07505_);
  and (_07507_, _06806_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_07508_, _07507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nand (_07509_, _06785_, _07472_);
  nand (_07510_, _06752_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_07511_, _07510_, _07509_);
  or (_07512_, _07511_, _07471_);
  and (_07513_, _07512_, _07508_);
  nor (_07515_, _07513_, _07506_);
  not (_07516_, _07515_);
  or (_07517_, _06795_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_07518_, _06775_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  and (_07519_, _07518_, _07517_);
  and (_07520_, _07519_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07521_, _07520_);
  nor (_07522_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4]);
  not (_07523_, _07522_);
  nand (_07524_, _07460_, _06532_);
  and (_07525_, _07524_, _07523_);
  and (_07526_, _07525_, _07521_);
  and (_07527_, _07513_, _07506_);
  nor (_07528_, _07527_, _07515_);
  nand (_07529_, _07528_, _07526_);
  nand (_07530_, _07529_, _07516_);
  nand (_07531_, _07530_, _07501_);
  and (_07532_, _07531_, _07496_);
  and (_07533_, _07468_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_07534_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3]);
  not (_07535_, _07534_);
  nand (_07536_, _07460_, _06551_);
  and (_07537_, _07536_, _07535_);
  not (_07538_, _07537_);
  or (_07539_, _07538_, _07533_);
  not (_07540_, _07533_);
  or (_07541_, _07537_, _07540_);
  nand (_07542_, _07541_, _07539_);
  and (_07543_, _07486_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07544_, _07543_);
  nand (_07545_, _07460_, _06604_);
  nor (_07546_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2]);
  not (_07547_, _07546_);
  and (_07548_, _07547_, _07545_);
  nand (_07549_, _07548_, _07544_);
  and (_07550_, _07507_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  not (_07551_, _07550_);
  nand (_07552_, _07460_, _06570_);
  nor (_07553_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1]);
  not (_07554_, _07553_);
  and (_07555_, _07554_, _07552_);
  nor (_07556_, _07555_, _07551_);
  or (_07557_, _07548_, _07544_);
  nand (_07558_, _07557_, _07549_);
  or (_07559_, _07558_, _07556_);
  and (_07560_, _07559_, _07549_);
  or (_07561_, _07560_, _07542_);
  nand (_07562_, _07561_, _07539_);
  not (_07564_, _07525_);
  and (_07565_, _07564_, _07520_);
  nor (_07566_, _07565_, _07526_);
  and (_07567_, _07528_, _07566_);
  and (_07568_, _07567_, _07501_);
  nand (_07569_, _07568_, _07562_);
  nand (_07570_, _07569_, _07532_);
  nor (_07571_, _07519_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  and (_07572_, _06482_, _07472_);
  and (_07573_, _06704_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_07574_, _07573_, _07572_);
  nor (_07575_, _07574_, _07471_);
  nor (_07576_, _07575_, _07571_);
  not (_07577_, _07576_);
  and (_07578_, _06739_, _06704_);
  nor (_07579_, _07578_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nor (_07580_, _07490_, _07475_);
  nor (_07581_, _07574_, _07511_);
  and (_07582_, _07581_, _07580_);
  nor (_07583_, _07582_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1]);
  nor (_07584_, _07583_, _07579_);
  and (_07585_, _07584_, _07577_);
  and (_07586_, _07585_, _07570_);
  and (_07587_, _07586_, _07459_);
  nor (_07588_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  not (_07589_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_07590_, _07589_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07591_, _07590_, _07588_);
  not (_07592_, _07591_);
  nor (_07593_, _07592_, _06879_);
  nor (_07594_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_07595_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_07596_, _07595_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_07597_, _07596_, _07594_);
  nor (_07598_, _07597_, _07593_);
  and (_07599_, _07597_, _07593_);
  nor (_07600_, _07599_, _07598_);
  and (_07601_, _07600_, _06847_);
  and (_07602_, _06628_, _06452_);
  not (_07603_, _06570_);
  nor (_07604_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  nand (_07605_, _07604_, _06704_);
  not (_07606_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0]);
  or (_07607_, _07606_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  or (_07608_, _07607_, _06482_);
  not (_07609_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  or (_07610_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _07609_);
  or (_07611_, _07610_, _06775_);
  and (_07612_, _07611_, _07608_);
  and (_07613_, _07610_, _07607_);
  or (_07614_, _06795_, _07609_);
  nand (_07615_, _07614_, _07613_);
  nand (_07616_, _07615_, _07612_);
  and (_07617_, _07616_, _07605_);
  and (_07618_, _07617_, _07603_);
  nand (_07619_, _07604_, _06739_);
  or (_07620_, _07607_, _06752_);
  or (_07621_, _07610_, _06785_);
  and (_07622_, _07621_, _07620_);
  or (_07624_, _06806_, _07609_);
  nand (_07625_, _07624_, _07613_);
  nand (_07626_, _07625_, _07622_);
  and (_07627_, _07626_, _07619_);
  and (_07628_, _07627_, _06903_);
  and (_07629_, _07628_, _07618_);
  nand (_07630_, _07626_, _07619_);
  or (_07631_, _07630_, _06570_);
  and (_07632_, _07617_, _06903_);
  not (_07633_, _07632_);
  and (_07634_, _07633_, _07631_);
  nor (_07635_, _07634_, _07629_);
  and (_07636_, _07635_, _07602_);
  or (_07637_, _07636_, _07601_);
  or (_07638_, _07637_, _07587_);
  or (_07639_, _07638_, _07458_);
  nor (_07640_, _07639_, _07440_);
  and (_07641_, _07640_, _07439_);
  not (_07642_, _07641_);
  not (_07643_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  and (_07644_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], _06308_);
  and (_07646_, _07644_, _07643_);
  and (_07647_, _06671_, _06336_);
  and (_07649_, _07647_, _07216_);
  and (_07650_, _07649_, _07150_);
  and (_07651_, _07650_, _06440_);
  nor (_07652_, _07651_, _07646_);
  not (_07653_, _07652_);
  nor (_07654_, _07586_, _07465_);
  not (_07655_, _07654_);
  not (_07656_, _07500_);
  and (_07657_, _07566_, _07562_);
  nor (_07659_, _07657_, _07526_);
  or (_07660_, _07659_, _07527_);
  and (_07661_, _07660_, _07516_);
  or (_07662_, _07661_, _07656_);
  and (_07664_, _07662_, _07493_);
  nand (_07665_, _07664_, _07497_);
  or (_07666_, _07664_, _07497_);
  nand (_07667_, _07666_, _07665_);
  nand (_07668_, _07667_, _07586_);
  and (_07669_, _07668_, _07655_);
  or (_07670_, _07669_, _07576_);
  nand (_07671_, _07669_, _07576_);
  not (_07672_, _07477_);
  not (_07673_, _07586_);
  and (_07674_, _07661_, _07656_);
  not (_07675_, _07674_);
  and (_07676_, _07675_, _07662_);
  nor (_07677_, _07676_, _07673_);
  nor (_07679_, _07586_, _07483_);
  nor (_07680_, _07679_, _07677_);
  and (_07681_, _07680_, _07672_);
  nand (_07682_, _07681_, _07671_);
  and (_07683_, _07682_, _07670_);
  and (_07684_, _07671_, _07670_);
  nor (_07685_, _07680_, _07672_);
  nor (_07686_, _07685_, _07681_);
  and (_07687_, _07686_, _07684_);
  not (_07688_, _07492_);
  nor (_07689_, _07528_, _07659_);
  and (_07690_, _07528_, _07659_);
  or (_07691_, _07690_, _07689_);
  nor (_07692_, _07691_, _07673_);
  nor (_07693_, _07586_, _07505_);
  nor (_07694_, _07693_, _07692_);
  and (_07695_, _07694_, _07688_);
  not (_07696_, _07513_);
  nor (_07697_, _07566_, _07562_);
  or (_07698_, _07697_, _07657_);
  and (_07699_, _07698_, _07586_);
  nor (_07700_, _07586_, _07525_);
  nor (_07701_, _07700_, _07699_);
  and (_07703_, _07701_, _07696_);
  not (_07704_, _07703_);
  nor (_07706_, _07694_, _07688_);
  or (_07707_, _07695_, _07706_);
  nor (_07708_, _07707_, _07704_);
  nor (_07709_, _07708_, _07695_);
  not (_07711_, _07709_);
  nor (_07712_, _07586_, _07538_);
  and (_07713_, _07560_, _07542_);
  not (_07714_, _07713_);
  and (_07715_, _07714_, _07561_);
  and (_07716_, _07715_, _07586_);
  or (_07717_, _07716_, _07712_);
  nor (_07718_, _07717_, _07521_);
  not (_07719_, _07718_);
  nand (_07720_, _07673_, _07555_);
  nor (_07721_, _07555_, _07550_);
  and (_07722_, _07555_, _07550_);
  nor (_07723_, _07722_, _07721_);
  nand (_07724_, _07586_, _07723_);
  nand (_07725_, _07724_, _07720_);
  nand (_07726_, _07725_, _07544_);
  or (_07727_, _07725_, _07544_);
  nand (_07728_, _07727_, _07726_);
  nor (_07729_, _07460_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0]);
  and (_07730_, _07460_, _06587_);
  nor (_07731_, _07730_, _07729_);
  nor (_07732_, _07731_, _07551_);
  or (_07733_, _07732_, _07728_);
  and (_07734_, _07733_, _07726_);
  or (_07735_, _07586_, _07548_);
  and (_07736_, _07558_, _07556_);
  not (_07737_, _07736_);
  and (_07738_, _07737_, _07559_);
  or (_07739_, _07738_, _07673_);
  and (_07740_, _07739_, _07735_);
  and (_07741_, _07740_, _07540_);
  nor (_07742_, _07740_, _07540_);
  or (_07743_, _07742_, _07741_);
  or (_07744_, _07743_, _07734_);
  and (_07745_, _07717_, _07521_);
  nor (_07746_, _07745_, _07741_);
  nand (_07747_, _07746_, _07744_);
  and (_07748_, _07747_, _07719_);
  nor (_07749_, _07701_, _07696_);
  nor (_07750_, _07749_, _07703_);
  not (_07751_, _07750_);
  nor (_07752_, _07707_, _07751_);
  and (_07753_, _07752_, _07748_);
  or (_07754_, _07753_, _07711_);
  nand (_07755_, _07754_, _07687_);
  nand (_07756_, _07755_, _07683_);
  and (_07757_, _07756_, _07584_);
  not (_07758_, _07757_);
  and (_07760_, _07732_, _07728_);
  not (_07761_, _07760_);
  and (_07762_, _07761_, _07733_);
  or (_07763_, _07762_, _07758_);
  or (_07764_, _07757_, _07725_);
  and (_07765_, _07764_, _07763_);
  nand (_07766_, _07765_, _07459_);
  not (_07767_, _07604_);
  and (_07768_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6]);
  and (_07769_, _07617_, _06534_);
  and (_07770_, _07627_, _06552_);
  and (_07771_, _07770_, _07769_);
  and (_07772_, _07627_, _06534_);
  and (_07773_, _07617_, _06958_);
  nand (_07774_, _07773_, _07772_);
  and (_07775_, _07627_, _06958_);
  or (_07776_, _07775_, _07769_);
  and (_07777_, _07776_, _07774_);
  and (_07778_, _07777_, _07771_);
  or (_07779_, _07774_, _06732_);
  and (_07780_, _07627_, _06957_);
  not (_07781_, _07780_);
  nand (_07782_, _07781_, _07774_);
  and (_07783_, _07782_, _07779_);
  nand (_07784_, _07783_, _07773_);
  or (_07785_, _07780_, _07773_);
  and (_07786_, _07785_, _07784_);
  nand (_07787_, _07786_, _07778_);
  not (_07788_, _07787_);
  not (_07789_, _07779_);
  and (_07790_, _07783_, _07773_);
  or (_07791_, _07630_, _06697_);
  nand (_07792_, _07616_, _07605_);
  or (_07793_, _07792_, _06732_);
  or (_07794_, _07793_, _07791_);
  nand (_07795_, _07793_, _07791_);
  and (_07796_, _07795_, _07794_);
  nand (_07797_, _07796_, _07790_);
  or (_07798_, _07796_, _07790_);
  and (_07799_, _07798_, _07797_);
  nand (_07800_, _07799_, _07789_);
  or (_07801_, _07799_, _07789_);
  and (_07802_, _07801_, _07800_);
  nand (_07803_, _07802_, _07788_);
  or (_07804_, _07802_, _07788_);
  nand (_07805_, _07804_, _07803_);
  not (_07806_, _07805_);
  and (_07807_, _07627_, _06605_);
  nand (_07808_, _07807_, _07618_);
  and (_07810_, _07617_, _06605_);
  and (_07811_, _07810_, _07631_);
  nand (_07812_, _07811_, _07770_);
  nand (_07813_, _07812_, _07808_);
  not (_07814_, _07771_);
  and (_07815_, _07617_, _06552_);
  or (_07816_, _07815_, _07772_);
  and (_07817_, _07816_, _07814_);
  nand (_07818_, _07817_, _07813_);
  not (_07819_, _07818_);
  not (_07820_, _07778_);
  or (_07821_, _07777_, _07771_);
  and (_07822_, _07821_, _07820_);
  and (_07823_, _07822_, _07819_);
  or (_07825_, _07786_, _07778_);
  and (_07826_, _07825_, _07787_);
  nand (_07827_, _07826_, _07823_);
  or (_07828_, _07807_, _07618_);
  and (_07829_, _07828_, _07808_);
  and (_07830_, _07829_, _07629_);
  or (_07831_, _07811_, _07770_);
  and (_07832_, _07831_, _07812_);
  nand (_07833_, _07832_, _07830_);
  not (_07834_, _07833_);
  or (_07835_, _07817_, _07813_);
  and (_07836_, _07835_, _07818_);
  nand (_07837_, _07836_, _07834_);
  not (_07838_, _07837_);
  nand (_07839_, _07822_, _07819_);
  or (_07840_, _07822_, _07819_);
  and (_07841_, _07840_, _07839_);
  nand (_07842_, _07841_, _07838_);
  not (_07843_, _07842_);
  or (_07844_, _07826_, _07823_);
  and (_07845_, _07844_, _07827_);
  nand (_07846_, _07845_, _07843_);
  nand (_07847_, _07846_, _07827_);
  nand (_07848_, _07847_, _07806_);
  nand (_07850_, _07848_, _07803_);
  and (_07851_, _07617_, _06914_);
  and (_07853_, _07851_, _07781_);
  and (_07854_, _07800_, _07797_);
  not (_07856_, _07854_);
  nand (_07857_, _07856_, _07853_);
  or (_07858_, _07856_, _07853_);
  and (_07859_, _07858_, _07857_);
  nand (_07861_, _07859_, _07850_);
  or (_07862_, _07859_, _07850_);
  and (_07864_, _07862_, _07861_);
  nand (_07865_, _07864_, _07768_);
  and (_07866_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5]);
  or (_07868_, _07847_, _07806_);
  and (_07869_, _07868_, _07848_);
  nand (_07870_, _07869_, _07866_);
  or (_07871_, _07869_, _07866_);
  nand (_07872_, _07871_, _07870_);
  and (_07873_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4]);
  or (_07874_, _07845_, _07843_);
  and (_07875_, _07874_, _07846_);
  nand (_07877_, _07875_, _07873_);
  or (_07879_, _07875_, _07873_);
  nand (_07880_, _07879_, _07877_);
  and (_07881_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3]);
  or (_07882_, _07841_, _07838_);
  and (_07883_, _07882_, _07842_);
  nand (_07884_, _07883_, _07881_);
  or (_07885_, _07883_, _07881_);
  and (_07886_, _07885_, _07884_);
  and (_07887_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2]);
  or (_07888_, _07836_, _07834_);
  and (_07889_, _07888_, _07837_);
  nand (_07890_, _07889_, _07887_);
  and (_07891_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1]);
  or (_07892_, _07832_, _07830_);
  and (_07893_, _07892_, _07833_);
  nand (_07894_, _07893_, _07891_);
  and (_07895_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0]);
  nand (_07896_, _07829_, _07629_);
  or (_07897_, _07829_, _07629_);
  and (_07898_, _07897_, _07896_);
  and (_07899_, _07898_, _07895_);
  or (_07900_, _07893_, _07891_);
  and (_07901_, _07900_, _07894_);
  nand (_07902_, _07901_, _07899_);
  nand (_07903_, _07902_, _07894_);
  or (_07904_, _07889_, _07887_);
  and (_07905_, _07904_, _07890_);
  nand (_07906_, _07905_, _07903_);
  nand (_07907_, _07906_, _07890_);
  nand (_07908_, _07907_, _07886_);
  and (_07910_, _07908_, _07884_);
  or (_07911_, _07910_, _07880_);
  and (_07912_, _07911_, _07877_);
  or (_07913_, _07912_, _07872_);
  and (_07914_, _07913_, _07870_);
  or (_07915_, _07864_, _07768_);
  nand (_07916_, _07915_, _07865_);
  or (_07917_, _07916_, _07914_);
  and (_07918_, _07917_, _07865_);
  and (_07919_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7]);
  and (_07920_, _07857_, _07794_);
  nand (_07921_, _07920_, _07861_);
  nand (_07922_, _07921_, _07919_);
  or (_07923_, _07921_, _07919_);
  nand (_07924_, _07923_, _07922_);
  or (_07925_, _07924_, _07918_);
  nand (_07926_, _07924_, _07918_);
  and (_07927_, _07926_, _07925_);
  nand (_07928_, _07927_, _07602_);
  nor (_07929_, _06828_, _06823_);
  nor (_07930_, _07929_, _06829_);
  nor (_07931_, _07930_, _06681_);
  not (_07932_, _07931_);
  not (_07933_, _06641_);
  nor (_07935_, _07933_, _06604_);
  not (_07936_, _07935_);
  and (_07937_, _06640_, _07603_);
  nor (_07938_, _06638_, _06587_);
  nor (_07939_, _07938_, _07937_);
  and (_07940_, _07939_, _07936_);
  and (_07941_, _07940_, _07067_);
  and (_07942_, _07941_, _07056_);
  nor (_07943_, _06884_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_07944_, _07943_, _07603_);
  nor (_07945_, _07943_, _07603_);
  nor (_07946_, _07945_, _07944_);
  nor (_07947_, _07946_, _06891_);
  nor (_07948_, _06825_, _06799_);
  or (_07949_, _07948_, _06854_);
  and (_07950_, _07949_, _06861_);
  nor (_07951_, _07949_, _06861_);
  or (_07952_, _07951_, _07950_);
  and (_07953_, _07952_, _06847_);
  nor (_07955_, _07953_, _07947_);
  and (_07956_, _07955_, _07942_);
  and (_07957_, _07956_, _07932_);
  and (_07958_, _07957_, _07928_);
  nand (_07959_, _07958_, _07766_);
  nand (_07960_, _07959_, _07653_);
  not (_07961_, _07439_);
  and (_07962_, _06940_, _06394_);
  nor (_07963_, _06364_, _06350_);
  and (_07965_, _07963_, _06674_);
  and (_07966_, _07965_, _07962_);
  and (_07967_, _07966_, _06432_);
  and (_07968_, _07967_, _06930_);
  nor (_07969_, _07967_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  or (_07971_, _07969_, _07653_);
  or (_07972_, _07971_, _07968_);
  and (_07974_, _07972_, _07961_);
  nand (_07975_, _07974_, _07960_);
  and (_07976_, _07975_, _07642_);
  and (_06429_, _07976_, _06444_);
  not (_07978_, _07731_);
  and (_07979_, _07757_, _07550_);
  nor (_07980_, _07979_, _07978_);
  and (_07981_, _07979_, _07978_);
  or (_07982_, _07981_, _07980_);
  nand (_07984_, _07982_, _07459_);
  not (_07985_, _07917_);
  and (_07986_, _07916_, _07914_);
  nor (_07987_, _07986_, _07985_);
  and (_07988_, _07987_, _07602_);
  nor (_07989_, _06827_, _06465_);
  nor (_07990_, _07989_, _06861_);
  not (_07991_, _07990_);
  nor (_07993_, _06847_, _06680_);
  nor (_07994_, _07993_, _07991_);
  not (_07995_, _07994_);
  nor (_07996_, _06825_, _06898_);
  nor (_07997_, _07996_, _06654_);
  or (_07998_, _07997_, _06826_);
  and (_07999_, _06825_, _06658_);
  and (_08000_, _06806_, _06455_);
  or (_08001_, _06660_, _06620_);
  and (_08002_, _08001_, _06587_);
  or (_08003_, _08002_, _08000_);
  nor (_08004_, _08003_, _07999_);
  and (_08005_, _06914_, _06907_);
  and (_08006_, _06913_, _06465_);
  nor (_08007_, _08006_, _08005_);
  or (_08008_, _07933_, _06570_);
  nor (_08009_, _06883_, _06640_);
  nor (_08010_, _08009_, _06587_);
  not (_08011_, _08010_);
  and (_08012_, _08011_, _08008_);
  and (_08013_, _08012_, _08007_);
  and (_08014_, _08013_, _08004_);
  and (_08015_, _08014_, _07998_);
  and (_08016_, _08015_, _07995_);
  not (_08017_, _08016_);
  nor (_08018_, _08017_, _07988_);
  nand (_08019_, _08018_, _07984_);
  nand (_08020_, _08019_, _07653_);
  not (_08021_, _06942_);
  nor (_08022_, _06930_, _08021_);
  nor (_08023_, _06942_, _06803_);
  nor (_08024_, _08023_, _08022_);
  or (_08025_, _07646_, _07439_);
  nor (_08026_, _08025_, _07651_);
  and (_08027_, _08026_, _07966_);
  not (_08028_, _08027_);
  nor (_08029_, _08028_, _08024_);
  not (_08030_, _06380_);
  and (_08031_, _06394_, _06336_);
  and (_08032_, _08031_, _07963_);
  and (_08033_, _08032_, _08030_);
  and (_08034_, _08033_, _06674_);
  not (_08035_, _08034_);
  and (_08036_, _08035_, _08026_);
  and (_08037_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_08038_, _08037_, _07439_);
  nor (_08039_, _08038_, _08029_);
  nand (_08040_, _08039_, _08020_);
  and (_08041_, _06806_, _06640_);
  and (_08042_, _06913_, _06534_);
  nor (_08043_, _06948_, _06892_);
  and (_08044_, _08043_, _06962_);
  nor (_08045_, _08044_, _06806_);
  and (_08046_, _08044_, _06806_);
  nor (_08047_, _08046_, _08045_);
  and (_08048_, _08047_, _06620_);
  nor (_08049_, _06587_, _06951_);
  or (_08050_, _08049_, _08048_);
  or (_08051_, _08050_, _08042_);
  and (_08052_, _07757_, _07459_);
  and (_08053_, _07592_, _06879_);
  nor (_08054_, _08053_, _07593_);
  and (_08055_, _08054_, _06847_);
  and (_08056_, _07628_, _07602_);
  or (_08057_, _08056_, _08055_);
  or (_08058_, _08057_, _08052_);
  or (_08059_, _08058_, _08051_);
  nor (_08060_, _08059_, _08041_);
  and (_08061_, _08060_, _07439_);
  not (_08062_, _08061_);
  and (_08063_, _08062_, _08040_);
  and (_06433_, _08063_, _06444_);
  and (_08064_, _07231_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  and (_08065_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  not (_08066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_08067_, _08064_, _08066_);
  or (_08069_, _08067_, _08065_);
  and (_06473_, _08069_, _06444_);
  and (_08070_, _07758_, _07694_);
  nand (_08071_, _07750_, _07748_);
  nand (_08072_, _08071_, _07704_);
  nor (_08073_, _08072_, _07707_);
  and (_08074_, _08072_, _07707_);
  or (_08076_, _08074_, _08073_);
  and (_08077_, _08076_, _07757_);
  or (_08078_, _08077_, _08070_);
  and (_08079_, _08078_, _07459_);
  or (_08080_, _07924_, _07865_);
  nand (_08081_, _08080_, _07922_);
  and (_08082_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8]);
  and (_08083_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9]);
  and (_08084_, _08083_, _08082_);
  and (_08085_, _08084_, _08081_);
  nor (_08086_, _07924_, _07916_);
  nand (_08087_, _08084_, _08086_);
  nor (_08088_, _08087_, _07914_);
  or (_08089_, _08088_, _08085_);
  and (_08090_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10]);
  and (_08091_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11]);
  and (_08092_, _08091_, _08090_);
  nand (_08093_, _08092_, _08089_);
  nand (_08094_, _08089_, _08090_);
  not (_08095_, _08091_);
  nand (_08096_, _08095_, _08094_);
  and (_08097_, _08096_, _08093_);
  and (_08098_, _08097_, _07602_);
  nor (_08099_, _06765_, _06650_);
  nor (_08100_, _08099_, _06850_);
  or (_08101_, _08100_, _06871_);
  nor (_08102_, _06872_, _06848_);
  and (_08103_, _08102_, _08101_);
  nor (_08104_, _06839_, _06764_);
  or (_08105_, _08104_, _06840_);
  and (_08106_, _08105_, _06680_);
  nor (_08107_, _06881_, _06697_);
  or (_08108_, _06885_, _06465_);
  nor (_08109_, _08108_, _08107_);
  nor (_08110_, _08109_, _06886_);
  and (_08111_, _08110_, _06511_);
  nor (_08112_, _08110_, _06511_);
  or (_08113_, _08112_, _08111_);
  and (_08114_, _08113_, _06883_);
  and (_08115_, _06640_, _06958_);
  nor (_08116_, _06638_, _06532_);
  nor (_08117_, _06732_, _07933_);
  or (_08119_, _08117_, _08116_);
  nor (_08120_, _08119_, _08115_);
  nand (_08121_, _08120_, _06664_);
  nor (_08122_, _08121_, _08114_);
  nand (_08123_, _08122_, _06625_);
  or (_08124_, _08123_, _08106_);
  or (_08125_, _08124_, _08103_);
  or (_08126_, _08125_, _08098_);
  or (_08127_, _08126_, _08079_);
  and (_08128_, _08127_, _07653_);
  nand (_08129_, _06987_, _06930_);
  or (_08130_, _06987_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_08131_, _08130_, _08027_);
  and (_08132_, _08131_, _08129_);
  and (_08133_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  or (_08134_, _08133_, _07439_);
  or (_08135_, _08134_, _08132_);
  or (_08136_, _08135_, _08128_);
  nor (_08137_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_08138_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_08139_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08138_);
  nor (_08141_, _08139_, _08137_);
  nor (_08142_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_08143_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_08144_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08143_);
  nor (_08145_, _08144_, _08142_);
  and (_08146_, _08145_, _07599_);
  and (_08147_, _08146_, _08141_);
  nor (_08148_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], \oc8051_top_1.oc8051_decoder1.src_sel3 );
  not (_08150_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_08151_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _08150_);
  nor (_08152_, _08151_, _08148_);
  and (_08153_, _08152_, _08147_);
  nor (_08154_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  not (_08155_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_08156_, _08155_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_08157_, _08156_, _08154_);
  or (_08158_, _08157_, _08153_);
  and (_08159_, _08157_, _08153_);
  nor (_08160_, _08159_, _06848_);
  and (_08161_, _08160_, _08158_);
  or (_08162_, _07907_, _07886_);
  and (_08163_, _08162_, _07908_);
  and (_08164_, _08163_, _07602_);
  nor (_08165_, _06806_, _06795_);
  and (_08166_, _06785_, _06775_);
  and (_08167_, _08166_, _08165_);
  and (_08168_, _08167_, _07442_);
  and (_08169_, _08168_, _06752_);
  nor (_08170_, _08169_, _06515_);
  and (_08171_, _07446_, _06795_);
  and (_08172_, _08171_, _06812_);
  nand (_08173_, _08172_, _06833_);
  nor (_08174_, _08173_, _06752_);
  nor (_08175_, _08174_, _06465_);
  nor (_08176_, _08175_, _08170_);
  or (_08177_, _08176_, _06483_);
  nand (_08178_, _08176_, _06483_);
  and (_08179_, _08178_, _06620_);
  and (_08180_, _08179_, _08177_);
  and (_08181_, _06913_, _07603_);
  nor (_08182_, _06465_, _06951_);
  nor (_08183_, _08182_, _06640_);
  nor (_08184_, _08183_, _06482_);
  and (_08185_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  nand (_08186_, _06465_, _06455_);
  nor (_08187_, _08186_, _06511_);
  or (_08188_, _08187_, _08185_);
  or (_08190_, _08188_, _08184_);
  or (_08191_, _08190_, _08181_);
  or (_08192_, _08191_, _08180_);
  or (_08193_, _08192_, _08164_);
  or (_08194_, _08193_, _08161_);
  or (_08195_, _08194_, _07961_);
  and (_08196_, _08195_, _08136_);
  and (_06517_, _08196_, _06444_);
  or (_08197_, _07750_, _07748_);
  nand (_08198_, _08197_, _08071_);
  nand (_08199_, _08198_, _07757_);
  or (_08200_, _07757_, _07701_);
  and (_08201_, _08200_, _08199_);
  and (_08202_, _08201_, _07459_);
  or (_08203_, _08089_, _08090_);
  and (_08205_, _08203_, _08094_);
  and (_08206_, _08205_, _07602_);
  nor (_08207_, _06838_, _06767_);
  and (_08208_, _06838_, _06767_);
  nor (_08209_, _08208_, _08207_);
  and (_08210_, _08209_, _06680_);
  or (_08211_, _06870_, _06767_);
  nor (_08212_, _06871_, _06848_);
  and (_08213_, _08212_, _08211_);
  nor (_08214_, _06884_, _06891_);
  and (_08215_, _08214_, _06534_);
  and (_08216_, _06885_, _06532_);
  and (_08217_, _06640_, _06534_);
  nor (_08218_, _07933_, _06511_);
  nor (_08220_, _06638_, _06551_);
  or (_08221_, _08220_, _08218_);
  or (_08222_, _08221_, _08217_);
  or (_08223_, _08222_, _08216_);
  nor (_08224_, _08223_, _08215_);
  and (_08225_, _08224_, _07186_);
  nand (_08226_, _08225_, _07177_);
  or (_08227_, _08226_, _08213_);
  or (_08228_, _08227_, _08210_);
  or (_08229_, _08228_, _08206_);
  or (_08230_, _08229_, _08202_);
  and (_08231_, _08230_, _07653_);
  not (_08232_, _06930_);
  and (_08233_, _06983_, _08232_);
  nor (_08234_, _06983_, _06749_);
  or (_08235_, _08234_, _08233_);
  and (_08236_, _08235_, _08027_);
  and (_08237_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_08238_, _08237_, _07439_);
  or (_08239_, _08238_, _08236_);
  or (_08241_, _08239_, _08231_);
  or (_08242_, _08152_, _08147_);
  nor (_08243_, _08153_, _06848_);
  and (_08244_, _08243_, _08242_);
  or (_08245_, _07905_, _07903_);
  and (_08246_, _08245_, _07906_);
  and (_08247_, _08246_, _07602_);
  and (_08248_, _08173_, _06515_);
  nor (_08249_, _08168_, _06515_);
  or (_08250_, _08249_, _08248_);
  nand (_08251_, _08250_, _06752_);
  or (_08252_, _08250_, _06752_);
  and (_08253_, _08252_, _06620_);
  and (_08254_, _08253_, _08251_);
  and (_08255_, _06913_, _06903_);
  nand (_08256_, _06532_, _06465_);
  or (_08257_, _06753_, _06465_);
  and (_08258_, _08257_, _06455_);
  and (_08259_, _08258_, _08256_);
  and (_08260_, _06753_, _06640_);
  and (_08261_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  or (_08262_, _08261_, _08260_);
  or (_08263_, _08262_, _08259_);
  or (_08264_, _08263_, _08255_);
  or (_08265_, _08264_, _08254_);
  or (_08266_, _08265_, _08247_);
  or (_08267_, _08266_, _08244_);
  or (_08268_, _08267_, _07961_);
  and (_08269_, _08268_, _08241_);
  and (_06533_, _08269_, _06444_);
  and (_08270_, _07758_, _07717_);
  or (_08271_, _07745_, _07718_);
  not (_08272_, _07741_);
  and (_08273_, _07744_, _08272_);
  nand (_08274_, _08273_, _08271_);
  or (_08275_, _08273_, _08271_);
  and (_08276_, _08275_, _08274_);
  and (_08277_, _08276_, _07757_);
  or (_08278_, _08277_, _08270_);
  and (_08279_, _08278_, _07459_);
  nand (_08280_, _07925_, _07922_);
  nand (_08281_, _08280_, _08082_);
  not (_08282_, _08083_);
  and (_08283_, _08282_, _08281_);
  nor (_08284_, _08283_, _08089_);
  and (_08285_, _08284_, _07602_);
  and (_08286_, _06831_, _06817_);
  nor (_08287_, _08286_, _06832_);
  nor (_08288_, _08287_, _06681_);
  nand (_08289_, _06866_, _06860_);
  nor (_08290_, _06867_, _06848_);
  and (_08291_, _08290_, _08289_);
  or (_08292_, _08214_, _06640_);
  and (_08293_, _08292_, _06552_);
  not (_08294_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_08295_, _06610_, _08294_);
  and (_08296_, _08295_, _08214_);
  nor (_08297_, _07933_, _06532_);
  nor (_08298_, _06638_, _06604_);
  nor (_08299_, _08298_, _08297_);
  and (_08300_, _08299_, _07295_);
  nand (_08301_, _08300_, _07292_);
  or (_08302_, _08301_, _08296_);
  nor (_08303_, _08302_, _08293_);
  nand (_08304_, _08303_, _07289_);
  or (_08305_, _08304_, _08291_);
  or (_08306_, _08305_, _08288_);
  or (_08307_, _08306_, _08285_);
  or (_08308_, _08307_, _08279_);
  and (_08309_, _08308_, _07653_);
  and (_08310_, _06932_, _06430_);
  nand (_08311_, _08310_, _06930_);
  or (_08312_, _08310_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_08313_, _08312_, _08027_);
  and (_08314_, _08313_, _08311_);
  and (_08315_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_08316_, _08315_, _07439_);
  or (_08317_, _08316_, _08314_);
  or (_08318_, _08317_, _08309_);
  or (_08319_, _08146_, _08141_);
  nor (_08320_, _08147_, _06848_);
  and (_08321_, _08320_, _08319_);
  and (_08322_, _08165_, _07442_);
  and (_08323_, _08322_, _06785_);
  nor (_08324_, _08323_, _06515_);
  nor (_08325_, _08172_, _06465_);
  nor (_08326_, _08325_, _08324_);
  nand (_08327_, _08326_, _06833_);
  or (_08328_, _08326_, _06833_);
  and (_08329_, _08328_, _06620_);
  and (_08330_, _08329_, _08327_);
  or (_08331_, _07901_, _07899_);
  and (_08332_, _08331_, _07902_);
  and (_08333_, _08332_, _07602_);
  nor (_08334_, _06551_, _06951_);
  and (_08335_, _06833_, _06640_);
  and (_08336_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  or (_08337_, _08336_, _08335_);
  or (_08338_, _08337_, _06915_);
  or (_08339_, _08338_, _08334_);
  or (_08340_, _08339_, _08333_);
  or (_08341_, _08340_, _08330_);
  or (_08342_, _08341_, _08321_);
  or (_08343_, _08342_, _07961_);
  and (_08344_, _08343_, _08318_);
  and (_06536_, _08344_, _06444_);
  nand (_08345_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  nand (_08346_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  and (_08347_, _08346_, _08345_);
  nand (_08348_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nand (_08349_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_08350_, _08349_, _08348_);
  nand (_08351_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nand (_08352_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_08353_, _08352_, _08351_);
  and (_08354_, _08353_, _08350_);
  nand (_08355_, _08354_, _08347_);
  nand (_08356_, _08355_, _07234_);
  nand (_08357_, _08356_, _07233_);
  nor (_08358_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _07233_);
  not (_08359_, _08358_);
  and (_08360_, _08359_, _08357_);
  and (_06566_, _08360_, _06444_);
  nor (_08361_, _07230_, _06699_);
  and (_08362_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  and (_08363_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_08364_, _08363_, _08362_);
  and (_08365_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_08366_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_08367_, _08366_, _08365_);
  and (_08368_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  and (_08369_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_08370_, _08369_, _08368_);
  and (_08371_, _08370_, _08367_);
  and (_08372_, _08371_, _08364_);
  and (_08373_, _07230_, _07234_);
  not (_08374_, _08373_);
  nor (_08375_, _08374_, _08372_);
  nor (_08376_, _08375_, _08361_);
  nor (_06569_, _08376_, rst);
  and (_06713_, _07263_, _06444_);
  nand (_08377_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nand (_08378_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  and (_08379_, _08378_, _08377_);
  nand (_08380_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_08381_, _08380_, _08379_);
  nand (_08382_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  and (_08383_, _08382_, _07234_);
  nand (_08384_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nand (_08385_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  and (_08386_, _08385_, _08384_);
  and (_08387_, _08386_, _08383_);
  nand (_08388_, _08387_, _08381_);
  or (_08389_, _08388_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_08390_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _07233_);
  not (_08391_, _08390_);
  and (_08392_, _08391_, _08389_);
  and (_06715_, _08392_, _06444_);
  and (_08393_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_08394_, _08393_);
  nand (_08395_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nand (_08396_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  and (_08397_, _08396_, _08395_);
  nand (_08398_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nand (_08399_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and (_08400_, _08399_, _08398_);
  and (_08401_, _08400_, _08397_);
  nand (_08402_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nand (_08403_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  and (_08404_, _08403_, _08402_);
  and (_08405_, _08404_, _08401_);
  or (_08406_, \oc8051_top_1.oc8051_memory_interface1.cdone , \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_08407_, _08406_, _08405_);
  and (_08408_, _08407_, _08394_);
  nor (_06717_, _08408_, rst);
  nand (_08410_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nand (_08411_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  and (_08412_, _08411_, _08410_);
  nand (_08413_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nand (_08414_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_08415_, _08414_, _08413_);
  nand (_08416_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nand (_08417_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_08418_, _08417_, _08416_);
  and (_08419_, _08418_, _08415_);
  nand (_08420_, _08419_, _08412_);
  nand (_08421_, _08420_, _07234_);
  nand (_08422_, _08421_, _07233_);
  nor (_08423_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _07233_);
  not (_08424_, _08423_);
  and (_08425_, _08424_, _08422_);
  and (_06719_, _08425_, _06444_);
  and (_08426_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_08427_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  and (_08428_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_08429_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_08430_, _08429_, _08428_);
  and (_08431_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_08432_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_08433_, _08432_, _08431_);
  nand (_08434_, _08433_, _08430_);
  or (_08435_, _08434_, _08427_);
  or (_08436_, _08435_, _08426_);
  or (_08437_, _08436_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_08438_, _08437_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_08439_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _07233_);
  not (_08440_, _08439_);
  and (_08441_, _08440_, _08438_);
  and (_06721_, _08441_, _06444_);
  nand (_08442_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  nand (_08443_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  and (_08444_, _08443_, _08442_);
  nand (_08445_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nand (_08446_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_08447_, _08446_, _08445_);
  nand (_08448_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nand (_08449_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  and (_08450_, _08449_, _08448_);
  and (_08451_, _08450_, _08447_);
  nand (_08452_, _08451_, _08444_);
  and (_08453_, _08452_, _07234_);
  or (_08454_, _08453_, \oc8051_top_1.oc8051_memory_interface1.cdone );
  nor (_08455_, _07233_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  not (_08456_, _08455_);
  and (_08457_, _08456_, _08454_);
  and (_06724_, _08457_, _06444_);
  nand (_08458_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nand (_08459_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_08460_, _08459_, _08458_);
  nand (_08461_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nand (_08462_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_08463_, _08462_, _08461_);
  nand (_08464_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  nand (_08465_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  and (_08466_, _08465_, _08464_);
  and (_08467_, _08466_, _08463_);
  and (_08468_, _08467_, _08460_);
  or (_08469_, _08468_, _08406_);
  and (_08470_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], \oc8051_top_1.oc8051_memory_interface1.cdone );
  not (_08471_, _08470_);
  and (_08472_, _08471_, _08469_);
  nor (_06726_, _08472_, rst);
  and (_08473_, _06299_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  and (_08474_, _08473_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_08475_, _08473_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_08476_, _08475_, _08474_);
  and (_06950_, _08476_, _06443_);
  nor (_08477_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  not (_08478_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08479_, _08478_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  nor (_08480_, _08479_, _08477_);
  not (_08481_, \oc8051_symbolic_cxrom1.regvalid [13]);
  not (_08482_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_08483_, _07432_, _08482_);
  and (_08484_, _08483_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_08485_, _08483_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_08486_, _08485_, _08484_);
  nor (_08487_, _08486_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08488_, _08478_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  nor (_08489_, _08488_, _08487_);
  and (_08490_, _08489_, _08481_);
  nor (_08491_, _08489_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08492_, _08491_, _08490_);
  not (_08493_, _08492_);
  nor (_08494_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_08495_, _08478_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  nor (_08496_, _08495_, _08494_);
  not (_08497_, _08496_);
  and (_08498_, _07432_, _08482_);
  nor (_08499_, _08498_, _08483_);
  nor (_08500_, _08499_, \oc8051_top_1.oc8051_memory_interface1.istb_t );
  nor (_08501_, _08478_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  nor (_08502_, _08501_, _08500_);
  and (_08503_, _08502_, _08497_);
  nand (_08504_, _08503_, _08493_);
  and (_08505_, _08504_, _08480_);
  nor (_08506_, _08502_, _08497_);
  not (_08507_, _08506_);
  not (_08508_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_08509_, _08489_, _08508_);
  and (_08510_, _08489_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08511_, _08510_, _08509_);
  nor (_08512_, _08511_, _08507_);
  and (_08513_, _08502_, _08496_);
  not (_08514_, _08513_);
  not (_08515_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_08516_, _08489_, _08515_);
  nor (_08517_, _08489_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_08518_, _08517_, _08516_);
  nor (_08519_, _08518_, _08514_);
  nor (_08520_, _08519_, _08512_);
  not (_08521_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08522_, _08489_, _08521_);
  nor (_08523_, _08502_, _08496_);
  not (_08524_, _08523_);
  nor (_08525_, _08489_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08526_, _08525_, _08524_);
  or (_08527_, _08526_, _08522_);
  and (_08528_, _08527_, _08520_);
  and (_08529_, _08528_, _08505_);
  not (_08530_, _08502_);
  and (_08531_, _08489_, \oc8051_symbolic_cxrom1.regvalid [12]);
  not (_08532_, _08489_);
  and (_08533_, _08532_, \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_08534_, _08533_, _08531_);
  nor (_08535_, _08534_, _08530_);
  nor (_08536_, _08502_, _08489_);
  and (_08537_, _08536_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_08538_, _08530_, _08489_);
  and (_08539_, _08538_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_08540_, _08539_, _08537_);
  not (_08541_, _08540_);
  nor (_08542_, _08541_, _08535_);
  nor (_08543_, _08542_, _08496_);
  and (_08544_, _08536_, _08496_);
  and (_08545_, _08544_, \oc8051_symbolic_cxrom1.regvalid [2]);
  not (_08546_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_08547_, _08489_, _08546_);
  nor (_08548_, _08489_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08549_, _08548_, _08547_);
  nor (_08550_, _08549_, _08514_);
  and (_08551_, _08489_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08552_, _08551_, _08506_);
  or (_08553_, _08552_, _08480_);
  or (_08554_, _08553_, _08550_);
  or (_08555_, _08554_, _08545_);
  nor (_08556_, _08555_, _08543_);
  nor (_08557_, _08556_, _08529_);
  not (_08558_, _08557_);
  and (_08559_, _08558_, word_in[7]);
  not (_08560_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  nand (_08561_, _08480_, _08560_);
  or (_08562_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_08563_, _08562_, _08561_);
  and (_08564_, _08563_, _08513_);
  not (_08565_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nand (_08566_, _08480_, _08565_);
  or (_08567_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_08568_, _08567_, _08566_);
  and (_08569_, _08568_, _08506_);
  or (_08570_, _08569_, _08564_);
  not (_08571_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nand (_08572_, _08480_, _08571_);
  or (_08573_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_08574_, _08573_, _08572_);
  and (_08575_, _08574_, _08503_);
  not (_08576_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  nand (_08577_, _08480_, _08576_);
  or (_08578_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_08579_, _08578_, _08577_);
  and (_08580_, _08579_, _08523_);
  or (_08581_, _08580_, _08575_);
  or (_08582_, _08581_, _08570_);
  and (_08583_, _08582_, _08489_);
  not (_08584_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  nand (_08585_, _08480_, _08584_);
  or (_08586_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_08587_, _08586_, _08585_);
  and (_08588_, _08587_, _08544_);
  and (_08589_, _08513_, _08532_);
  not (_08590_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  nand (_08591_, _08480_, _08590_);
  or (_08592_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_08593_, _08592_, _08591_);
  and (_08594_, _08593_, _08589_);
  not (_08595_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nand (_08596_, _08480_, _08595_);
  or (_08597_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_08598_, _08597_, _08596_);
  and (_08599_, _08598_, _08503_);
  not (_08600_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nand (_08601_, _08480_, _08600_);
  or (_08602_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_08603_, _08602_, _08601_);
  and (_08604_, _08603_, _08523_);
  or (_08605_, _08604_, _08599_);
  and (_08606_, _08605_, _08532_);
  or (_08607_, _08606_, _08594_);
  or (_08608_, _08607_, _08588_);
  or (_08609_, _08608_, _08583_);
  and (_08610_, _08609_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [7], _08610_, _08559_);
  nor (_08611_, _08496_, _08480_);
  not (_08612_, _08611_);
  and (_08613_, _08496_, _08480_);
  nor (_08614_, _08613_, _08502_);
  and (_08615_, _08613_, _08502_);
  nor (_08616_, _08615_, _08614_);
  not (_08617_, _08616_);
  nor (_08618_, _08617_, _08492_);
  nor (_08619_, _08615_, _08532_);
  and (_08620_, _08615_, _08532_);
  nor (_08622_, _08620_, _08619_);
  nor (_08623_, _08622_, _08616_);
  and (_08624_, _08623_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_08626_, _08622_, _08617_);
  and (_08627_, _08626_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08628_, _08627_, _08624_);
  nor (_08630_, _08628_, _08618_);
  nor (_08631_, _08630_, _08612_);
  not (_08632_, _08631_);
  not (_08634_, _08613_);
  nor (_08635_, _08617_, _08534_);
  and (_08636_, _08626_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_08638_, _08636_, _08635_);
  or (_08639_, _08638_, _08634_);
  nand (_08640_, _08620_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_08642_, _08640_, _08639_);
  and (_08643_, _08642_, _08632_);
  and (_08644_, _08497_, _08480_);
  not (_08645_, _08644_);
  nor (_08646_, _08617_, _08549_);
  and (_08648_, _08623_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08649_, _08626_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08651_, _08649_, _08648_);
  nor (_08652_, _08651_, _08646_);
  nor (_08653_, _08652_, _08645_);
  not (_08654_, _08480_);
  and (_08655_, _08496_, _08654_);
  not (_08656_, _08655_);
  nor (_08657_, _08617_, _08518_);
  and (_08658_, _08623_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_08659_, _08626_, \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_08660_, _08659_, _08658_);
  nor (_08661_, _08660_, _08657_);
  nor (_08662_, _08661_, _08656_);
  nor (_08663_, _08662_, _08653_);
  and (_08664_, _08663_, _08643_);
  or (_08665_, _08613_, _08611_);
  not (_08666_, _08665_);
  not (_08667_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  nand (_08668_, _08480_, _08667_);
  or (_08669_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  and (_08670_, _08669_, _08668_);
  and (_08671_, _08670_, _08666_);
  not (_08672_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nand (_08673_, _08480_, _08672_);
  or (_08674_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_08675_, _08674_, _08673_);
  and (_08676_, _08675_, _08665_);
  or (_08677_, _08676_, _08671_);
  and (_08678_, _08677_, _08623_);
  and (_08679_, _08616_, _08489_);
  not (_08680_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  nand (_08681_, _08480_, _08680_);
  or (_08682_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_08683_, _08682_, _08681_);
  and (_08684_, _08683_, _08666_);
  not (_08685_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nand (_08686_, _08480_, _08685_);
  or (_08687_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  and (_08688_, _08687_, _08686_);
  and (_08689_, _08688_, _08665_);
  or (_08691_, _08689_, _08684_);
  and (_08692_, _08691_, _08679_);
  or (_08693_, _08692_, _08678_);
  not (_08695_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nand (_08696_, _08480_, _08695_);
  or (_08697_, _08480_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  and (_08698_, _08697_, _08696_);
  and (_08699_, _08698_, _08665_);
  not (_08700_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  nand (_08702_, _08480_, _08700_);
  or (_08703_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_08704_, _08703_, _08702_);
  and (_08705_, _08704_, _08666_);
  or (_08706_, _08705_, _08699_);
  and (_08707_, _08706_, _08626_);
  and (_08708_, _08616_, _08532_);
  not (_08709_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nand (_08710_, _08480_, _08709_);
  or (_08711_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  and (_08712_, _08711_, _08710_);
  and (_08713_, _08712_, _08665_);
  not (_08714_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  nand (_08715_, _08480_, _08714_);
  or (_08716_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_08717_, _08716_, _08715_);
  and (_08718_, _08717_, _08666_);
  or (_08720_, _08718_, _08713_);
  and (_08721_, _08720_, _08708_);
  or (_08722_, _08721_, _08707_);
  nor (_08723_, _08722_, _08693_);
  nor (_08724_, _08723_, _08664_);
  and (_08725_, _08664_, word_in[15]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [15], _08725_, _08724_);
  nor (_08726_, _08513_, _08523_);
  not (_08727_, _08726_);
  nor (_08728_, _08727_, _08492_);
  and (_08729_, _08513_, _08489_);
  nor (_08730_, _08513_, _08489_);
  nor (_08731_, _08730_, _08729_);
  nor (_08732_, _08726_, _08731_);
  and (_08733_, _08732_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_08734_, _08727_, _08731_);
  and (_08735_, _08734_, \oc8051_symbolic_cxrom1.regvalid [9]);
  or (_08736_, _08735_, _08733_);
  nor (_08737_, _08736_, _08728_);
  nor (_08738_, _08737_, _08634_);
  and (_08739_, _08732_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_08740_, _08739_);
  nor (_08742_, _08727_, _08518_);
  and (_08744_, _08734_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08746_, _08744_, _08742_);
  and (_08747_, _08746_, _08740_);
  nor (_08748_, _08747_, _08645_);
  nor (_08749_, _08748_, _08738_);
  nor (_08751_, _08727_, _08549_);
  and (_08752_, _08734_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_08753_, _08732_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08754_, _08753_, _08752_);
  nor (_08756_, _08754_, _08751_);
  nor (_08758_, _08756_, _08612_);
  and (_08759_, _08732_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not (_08760_, _08759_);
  nor (_08761_, _08727_, _08534_);
  and (_08763_, _08734_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_08764_, _08763_, _08761_);
  and (_08765_, _08764_, _08760_);
  nor (_08766_, _08765_, _08656_);
  nor (_08768_, _08766_, _08758_);
  and (_08769_, _08768_, _08749_);
  not (_08770_, _08731_);
  and (_08771_, _08593_, _08503_);
  and (_08772_, _08603_, _08489_);
  or (_08773_, _08772_, _08771_);
  and (_08774_, _08598_, _08506_);
  and (_08775_, _08587_, _08523_);
  or (_08776_, _08775_, _08774_);
  or (_08777_, _08776_, _08773_);
  and (_08778_, _08777_, _08770_);
  and (_08779_, _08574_, _08506_);
  and (_08780_, _08568_, _08523_);
  or (_08781_, _08780_, _08779_);
  and (_08782_, _08563_, _08503_);
  and (_08783_, _08579_, _08513_);
  or (_08784_, _08783_, _08782_);
  or (_08785_, _08784_, _08781_);
  and (_08786_, _08785_, _08731_);
  nor (_08787_, _08786_, _08778_);
  nor (_08788_, _08787_, _08769_);
  and (_08789_, _08769_, word_in[23]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [23], _08789_, _08788_);
  and (_08790_, _08729_, _08654_);
  and (_08791_, _08790_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_08792_, _08612_, _08502_);
  nor (_08793_, _08612_, _08502_);
  nor (_08794_, _08793_, _08792_);
  not (_08795_, _08794_);
  nor (_08796_, _08795_, _08518_);
  and (_08797_, _08792_, _08489_);
  nor (_08798_, _08792_, _08489_);
  nor (_08799_, _08798_, _08797_);
  and (_08800_, _08799_, _08795_);
  and (_08801_, _08800_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_08802_, _08801_, _08796_);
  nor (_08803_, _08802_, _08612_);
  nor (_08804_, _08803_, _08791_);
  nor (_08805_, _08795_, _08492_);
  and (_08806_, _08800_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_08807_, _08806_, _08805_);
  nor (_08808_, _08807_, _08656_);
  and (_08809_, _08793_, _08509_);
  nor (_08810_, _08809_, _08808_);
  and (_08811_, _08810_, _08804_);
  nor (_08812_, _08549_, _08795_);
  and (_08813_, _08800_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_08814_, _08799_, _08794_);
  and (_08815_, _08814_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_08816_, _08815_, _08813_);
  nor (_08817_, _08816_, _08812_);
  nor (_08818_, _08817_, _08634_);
  and (_08819_, _08502_, _08489_);
  and (_08820_, _08644_, _08819_);
  and (_08821_, _08820_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_08822_, _08795_, _08534_);
  and (_08823_, _08800_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_08824_, _08823_, _08822_);
  nor (_08825_, _08824_, _08645_);
  or (_08826_, _08825_, _08821_);
  nor (_08827_, _08826_, _08818_);
  and (_08828_, _08827_, _08811_);
  and (_08829_, _08675_, _08666_);
  and (_08830_, _08670_, _08665_);
  or (_08831_, _08830_, _08829_);
  and (_08832_, _08831_, _08800_);
  and (_08833_, _08698_, _08666_);
  and (_08834_, _08704_, _08665_);
  or (_08835_, _08834_, _08833_);
  and (_08836_, _08835_, _08814_);
  and (_08837_, _08794_, _08532_);
  and (_08838_, _08712_, _08666_);
  and (_08839_, _08717_, _08665_);
  or (_08840_, _08839_, _08838_);
  and (_08841_, _08840_, _08837_);
  and (_08842_, _08794_, _08489_);
  and (_08843_, _08688_, _08666_);
  and (_08844_, _08683_, _08665_);
  or (_08845_, _08844_, _08843_);
  and (_08846_, _08845_, _08842_);
  or (_08847_, _08846_, _08841_);
  or (_08848_, _08847_, _08836_);
  nor (_08849_, _08848_, _08832_);
  nor (_08850_, _08849_, _08828_);
  and (_08852_, _08828_, word_in[31]);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [31], _08852_, _08850_);
  or (_08853_, _08819_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_07051_, _08853_, _06444_);
  and (_08855_, _08828_, _06444_);
  and (_08856_, _08855_, word_in[31]);
  and (_08857_, _08819_, _08611_);
  and (_08859_, _08855_, _08857_);
  and (_08860_, _08859_, _08856_);
  not (_08862_, _08859_);
  and (_08863_, _08769_, _06444_);
  and (_08865_, _08863_, _08726_);
  and (_08866_, _08865_, _08731_);
  and (_08867_, _08866_, _08644_);
  not (_08868_, _08867_);
  and (_08869_, _08664_, _06444_);
  and (_08870_, _08869_, _08655_);
  and (_08871_, _08870_, _08679_);
  and (_08872_, _08529_, _06444_);
  and (_08874_, _08872_, _08496_);
  nor (_08875_, _08557_, rst);
  and (_08877_, _08875_, _08819_);
  and (_08878_, _08877_, _08874_);
  and (_08879_, _08878_, word_in[7]);
  nor (_08880_, _08878_, _08560_);
  nor (_08881_, _08880_, _08879_);
  nor (_08882_, _08881_, _08871_);
  and (_08883_, _08871_, word_in[15]);
  or (_08884_, _08883_, _08882_);
  and (_08885_, _08884_, _08868_);
  and (_08886_, _08863_, word_in[23]);
  and (_08887_, _08886_, _08867_);
  or (_08888_, _08887_, _08885_);
  and (_08889_, _08888_, _08862_);
  or (_14579_, _08889_, _08860_);
  or (_08890_, _08814_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_07097_, _08890_, _06444_);
  and (_08891_, _08523_, _08532_);
  or (_08892_, _08891_, \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_08893_, _08892_, _08729_);
  and (_07129_, _08893_, _06444_);
  and (_08894_, _08615_, _08489_);
  or (_08895_, _08894_, _08891_);
  or (_08896_, _08645_, _08502_);
  nor (_08897_, _08896_, _08489_);
  and (_08898_, _08837_, _08655_);
  nor (_08899_, _08898_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_08900_, _08899_, _08897_);
  or (_08901_, _08900_, _08895_);
  and (_07165_, _08901_, _06444_);
  or (_08902_, _08536_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_07212_, _08902_, _06444_);
  not (_08903_, _08536_);
  nor (_08904_, _08530_, _08489_);
  and (_08905_, _08904_, _08611_);
  or (_08906_, _08905_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_08907_, _08906_, _08903_);
  and (_08908_, _08793_, _08533_);
  or (_08909_, _08897_, _08544_);
  or (_08910_, _08909_, _08908_);
  or (_08911_, _08910_, _08907_);
  and (_07279_, _08911_, _06444_);
  and (_08912_, _06364_, _06671_);
  and (_08913_, _08912_, _07962_);
  and (_08914_, _08913_, _06933_);
  nand (_08915_, _08914_, _06930_);
  or (_08916_, _08914_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_08917_, _08916_, _06674_);
  and (_08918_, _08917_, _08915_);
  and (_08919_, _08913_, _06942_);
  not (_08920_, _08919_);
  nor (_08921_, _08920_, _06978_);
  and (_08922_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_08923_, _08922_, _08921_);
  and (_08924_, _08923_, _06440_);
  not (_08925_, _06673_);
  and (_08926_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  or (_08927_, _08926_, rst);
  or (_08928_, _08927_, _08924_);
  or (_07328_, _08928_, _08918_);
  not (_08929_, _08730_);
  and (_08930_, _08613_, _08536_);
  or (_08931_, _08905_, _08930_);
  or (_08932_, _08931_, _08929_);
  and (_08933_, _08932_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_08934_, _08904_, _08644_);
  and (_08935_, _08898_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08936_, _08935_, _08934_);
  nor (_08937_, _08936_, _08933_);
  nor (_08938_, _08937_, _08798_);
  and (_08939_, _08891_, \oc8051_symbolic_cxrom1.regvalid [5]);
  or (_08940_, _08939_, _08898_);
  or (_08941_, _08940_, _08905_);
  or (_08942_, _08941_, _08930_);
  or (_08944_, _08942_, _08938_);
  and (_07337_, _08944_, _06444_);
  and (_08946_, _08792_, _08532_);
  or (_08947_, _08619_, _08946_);
  or (_08949_, _08790_, _08731_);
  or (_08950_, _08489_, _08480_);
  nor (_08952_, _08950_, _08514_);
  and (_08953_, _08931_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08955_, _08953_, _08952_);
  and (_08956_, _08903_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08958_, _08956_, _08950_);
  and (_08959_, _08898_, \oc8051_symbolic_cxrom1.regvalid [6]);
  and (_08961_, _08891_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_08962_, _08961_, _08959_);
  or (_08963_, _08962_, _08958_);
  or (_08964_, _08963_, _08955_);
  and (_08965_, _08964_, _08949_);
  or (_08966_, _08953_, _08934_);
  or (_08967_, _08966_, _08965_);
  and (_08968_, _08967_, _08947_);
  and (_08969_, _08964_, _08894_);
  or (_08970_, _08961_, _08930_);
  or (_08971_, _08970_, _08959_);
  or (_08972_, _08971_, _08905_);
  or (_08973_, _08972_, _08969_);
  or (_08974_, _08973_, _08968_);
  and (_07395_, _08974_, _06444_);
  and (_08975_, _07644_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1]);
  nor (_08976_, _06418_, _06407_);
  and (_08977_, _08976_, _06430_);
  and (_08978_, _07402_, _07214_);
  and (_08979_, _08978_, _08977_);
  nor (_08980_, _08979_, _08975_);
  or (_08981_, _08980_, _08019_);
  not (_08982_, _08980_);
  or (_08983_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_08984_, _08983_, _06444_);
  and (_07449_, _08984_, _08981_);
  nand (_08985_, _07754_, _07686_);
  or (_08986_, _07754_, _07686_);
  nand (_08987_, _08986_, _08985_);
  nand (_08988_, _08987_, _07757_);
  or (_08989_, _07757_, _07680_);
  and (_08990_, _08989_, _08988_);
  nand (_08991_, _08990_, _07459_);
  and (_08992_, _08092_, _08089_);
  and (_08993_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12]);
  nand (_08994_, _08993_, _08992_);
  or (_08995_, _08993_, _08992_);
  and (_08996_, _08995_, _08994_);
  nand (_08997_, _08996_, _07602_);
  nor (_08998_, _06840_, _06761_);
  nor (_08999_, _08998_, _06841_);
  nor (_09000_, _08999_, _06681_);
  not (_09001_, _09000_);
  nor (_09002_, _06874_, _06872_);
  not (_09003_, _09002_);
  nor (_09004_, _06875_, _06848_);
  and (_09005_, _09004_, _09003_);
  and (_09006_, _06740_, _06465_);
  nor (_09007_, _06732_, _06465_);
  or (_09008_, _09007_, _09006_);
  and (_09009_, _09008_, _06455_);
  nor (_09010_, _06959_, _06957_);
  not (_09011_, _09010_);
  and (_09012_, _09011_, _06961_);
  and (_09013_, _06613_, _06511_);
  nor (_09014_, _06732_, _09013_);
  nor (_09015_, _09014_, _06955_);
  nor (_09016_, _09015_, _06515_);
  nor (_09017_, _09016_, _09012_);
  nor (_09018_, _09017_, _06621_);
  nor (_09019_, _09018_, _09009_);
  nor (_09020_, _08111_, _06732_);
  and (_09021_, _08111_, _06732_);
  nor (_09022_, _09021_, _09020_);
  nor (_09023_, _09022_, _06891_);
  and (_09024_, _06744_, _06647_);
  and (_09025_, _06742_, _06658_);
  nor (_09026_, _06743_, _06655_);
  and (_09027_, _06732_, _06660_);
  or (_09028_, _09027_, _09026_);
  or (_09029_, _09028_, _09025_);
  nor (_09030_, _09029_, _09024_);
  or (_09031_, _06697_, _07933_);
  nor (_09032_, _06638_, _06511_);
  and (_09033_, _06957_, _06640_);
  nor (_09034_, _09033_, _09032_);
  and (_09035_, _09034_, _09031_);
  and (_09036_, _09035_, _09030_);
  not (_09037_, _09036_);
  nor (_09038_, _09037_, _09023_);
  and (_09039_, _09038_, _09019_);
  not (_09040_, _09039_);
  nor (_09041_, _09040_, _09005_);
  and (_09042_, _09041_, _09001_);
  and (_09043_, _09042_, _08997_);
  and (_09045_, _09043_, _08991_);
  nand (_09046_, _09045_, _08982_);
  or (_09048_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_09049_, _09048_, _06444_);
  and (_07452_, _09049_, _09046_);
  or (_09051_, _08980_, _08127_);
  or (_09052_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_09053_, _09052_, _06444_);
  and (_07455_, _09053_, _09051_);
  or (_09054_, _08980_, _08230_);
  or (_09055_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_09056_, _09055_, _06444_);
  and (_07469_, _09056_, _09054_);
  not (_09057_, _08622_);
  and (_09059_, _08536_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_09060_, _08952_, _08489_);
  and (_09062_, _09060_, \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_09063_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_09064_, _08496_, _09063_);
  and (_09065_, _09064_, _08904_);
  or (_09066_, _09065_, _08620_);
  or (_09067_, _09066_, _09062_);
  or (_09068_, _09067_, _09059_);
  and (_09069_, _09068_, _09057_);
  and (_09070_, _08837_, \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_09071_, _09070_, _08480_);
  and (_09072_, _08898_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_09073_, _09065_, _08952_);
  or (_09074_, _09073_, _09072_);
  or (_09075_, _09074_, _09071_);
  or (_09076_, _09075_, _09069_);
  and (_09077_, _09076_, _08949_);
  and (_09078_, _09068_, _08894_);
  or (_09079_, _09059_, _08905_);
  or (_09080_, _09079_, _08934_);
  or (_09081_, _09080_, _09078_);
  or (_09082_, _09081_, _09077_);
  and (_07485_, _09082_, _06444_);
  or (_09083_, _08980_, _08308_);
  or (_09084_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_09085_, _09084_, _06444_);
  and (_07494_, _09085_, _09083_);
  not (_09086_, _07459_);
  and (_09087_, _07743_, _07734_);
  not (_09088_, _09087_);
  and (_09089_, _09088_, _07744_);
  nor (_09090_, _09089_, _07758_);
  nor (_09091_, _07757_, _07740_);
  or (_09092_, _09091_, _09090_);
  or (_09093_, _09092_, _09086_);
  or (_09094_, _08280_, _08082_);
  and (_09095_, _09094_, _08281_);
  nand (_09096_, _09095_, _07602_);
  nor (_09097_, _06829_, _06820_);
  nor (_09098_, _09097_, _06830_);
  nor (_09099_, _09098_, _06681_);
  not (_09100_, _09099_);
  nor (_09101_, _06864_, _06862_);
  not (_09102_, _09101_);
  nor (_09103_, _06865_, _06848_);
  and (_09104_, _09103_, _09102_);
  not (_09105_, _09104_);
  nor (_09106_, _06785_, _06951_);
  and (_09107_, _07049_, _06465_);
  and (_09108_, _06588_, _06515_);
  nor (_09109_, _09108_, _09107_);
  nor (_09110_, _09109_, _06605_);
  and (_09111_, _09109_, _06605_);
  or (_09112_, _09111_, _09110_);
  and (_09113_, _09112_, _06620_);
  nor (_09114_, _09113_, _09106_);
  and (_09115_, _06610_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nor (_09116_, _07945_, _06604_);
  nor (_09117_, _09116_, _09115_);
  nor (_09118_, _09117_, _06891_);
  nor (_09119_, _06787_, _06655_);
  and (_09120_, _06788_, _06647_);
  nor (_09121_, _09120_, _09119_);
  and (_09122_, _06786_, _06658_);
  and (_09123_, _06660_, _06604_);
  nor (_09124_, _09123_, _09122_);
  or (_09125_, _07933_, _06551_);
  nor (_09126_, _06638_, _06570_);
  and (_09127_, _06640_, _06605_);
  nor (_09128_, _09127_, _09126_);
  and (_09129_, _09128_, _09125_);
  and (_09130_, _09129_, _09124_);
  and (_09131_, _09130_, _09121_);
  not (_09132_, _09131_);
  nor (_09133_, _09132_, _09118_);
  and (_09134_, _09133_, _09114_);
  and (_09135_, _09134_, _09105_);
  and (_09136_, _09135_, _09100_);
  and (_09137_, _09136_, _09096_);
  and (_09138_, _09137_, _09093_);
  nand (_09139_, _09138_, _08982_);
  or (_09140_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_09141_, _09140_, _06444_);
  and (_07498_, _09141_, _09139_);
  or (_09142_, _08980_, _07959_);
  or (_09143_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_09144_, _09143_, _06444_);
  and (_07514_, _09144_, _09142_);
  or (_09145_, _08800_, \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_07563_, _09145_, _06444_);
  not (_09146_, _07414_);
  nor (_09147_, _09146_, _06666_);
  and (_09149_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  or (_09151_, _09149_, _07158_);
  or (_09152_, _09151_, _09147_);
  or (_09154_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [5]);
  and (_09155_, _09154_, _06444_);
  and (_07623_, _09155_, _09152_);
  and (_09157_, _08978_, _08310_);
  not (_09158_, _09157_);
  nor (_09160_, _09158_, _09045_);
  and (_09161_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_09163_, _09161_, _08975_);
  or (_09164_, _09163_, _09160_);
  and (_09165_, _06740_, _06640_);
  and (_09167_, _06913_, _06605_);
  or (_09168_, _06752_, _06482_);
  and (_09169_, _09168_, _06515_);
  or (_09171_, _09169_, _06484_);
  or (_09172_, _09171_, _08170_);
  nor (_09173_, _09172_, _08248_);
  and (_09174_, _09173_, _06739_);
  nor (_09175_, _09173_, _06739_);
  or (_09176_, _09175_, _09174_);
  and (_09177_, _09176_, _06620_);
  nor (_09178_, _06739_, _06465_);
  nor (_09179_, _06732_, _06515_);
  or (_09180_, _09179_, _09178_);
  and (_09181_, _09180_, _06455_);
  or (_09182_, _09181_, _09177_);
  or (_09183_, _09182_, _09167_);
  and (_09184_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  nor (_09185_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  not (_09186_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_09187_, _09186_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  nor (_09188_, _09187_, _09185_);
  nor (_09189_, _09188_, _08159_);
  not (_09190_, _09189_);
  and (_09191_, _09188_, _08159_);
  nor (_09192_, _09191_, _06848_);
  and (_09193_, _09192_, _09190_);
  and (_09194_, _07910_, _07880_);
  not (_09195_, _09194_);
  and (_09196_, _09195_, _07911_);
  and (_09197_, _09196_, _07602_);
  or (_09198_, _09197_, _09193_);
  or (_09199_, _09198_, _09184_);
  or (_09200_, _09199_, _09183_);
  nor (_09201_, _09200_, _09165_);
  nand (_09202_, _09201_, _08975_);
  and (_09203_, _09202_, _06444_);
  and (_07645_, _09203_, _09164_);
  and (_09204_, _09157_, _08127_);
  and (_09205_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_09206_, _09205_, _08975_);
  or (_09207_, _09206_, _09204_);
  not (_09208_, _08975_);
  or (_09209_, _09208_, _08194_);
  and (_09210_, _09209_, _06444_);
  and (_07648_, _09210_, _09207_);
  and (_09211_, _09157_, _08230_);
  and (_09212_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_09213_, _09212_, _08975_);
  or (_09214_, _09213_, _09211_);
  or (_09215_, _09208_, _08267_);
  and (_09216_, _09215_, _06444_);
  and (_07658_, _09216_, _09214_);
  not (_09217_, _08793_);
  and (_09218_, _08619_, _09217_);
  nor (_09219_, _08896_, _08532_);
  nor (_09220_, _08730_, _08521_);
  or (_09221_, _09220_, _09219_);
  and (_09222_, _09221_, _09218_);
  and (_09223_, _08793_, _08489_);
  nor (_09224_, _08489_, _08521_);
  and (_09225_, _09224_, _08513_);
  or (_09226_, _09225_, _09223_);
  or (_09227_, _09226_, _09222_);
  and (_09228_, _09227_, _08619_);
  or (_09229_, _08934_, _08837_);
  and (_09230_, _09229_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_09231_, _09221_, _08894_);
  and (_09232_, _09224_, _08793_);
  or (_09233_, _09232_, _08952_);
  or (_09235_, _09233_, _09231_);
  or (_09236_, _09235_, _09230_);
  or (_09237_, _09236_, _08620_);
  or (_09238_, _09237_, _09228_);
  and (_07663_, _09238_, _06444_);
  and (_09239_, _09157_, _08308_);
  and (_09241_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_09242_, _09241_, _08975_);
  or (_09243_, _09242_, _09239_);
  or (_09244_, _09208_, _08342_);
  and (_09246_, _09244_, _06444_);
  and (_07678_, _09246_, _09243_);
  nor (_09247_, _09158_, _09138_);
  and (_09249_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_09250_, _09249_, _08975_);
  or (_09251_, _09250_, _09247_);
  and (_09252_, _06812_, _06640_);
  and (_09254_, _06957_, _06913_);
  nor (_09255_, _06604_, _06951_);
  nor (_09256_, _08171_, _06465_);
  nor (_09257_, _08322_, _06515_);
  or (_09259_, _09257_, _09256_);
  and (_09260_, _09259_, _06785_);
  nor (_09262_, _09259_, _06785_);
  nor (_09263_, _09262_, _09260_);
  and (_09264_, _09263_, _06620_);
  or (_09266_, _09264_, _09255_);
  or (_09267_, _09266_, _09254_);
  and (_09268_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  nor (_09269_, _08145_, _07599_);
  not (_09271_, _09269_);
  nor (_09272_, _08146_, _06848_);
  and (_09273_, _09272_, _09271_);
  nor (_09274_, _07898_, _07895_);
  nor (_09275_, _09274_, _07899_);
  and (_09276_, _09275_, _07602_);
  or (_09277_, _09276_, _09273_);
  or (_09278_, _09277_, _09268_);
  or (_09279_, _09278_, _09267_);
  nor (_09280_, _09279_, _09252_);
  nand (_09281_, _09280_, _08975_);
  and (_09282_, _09281_, _06444_);
  and (_07702_, _09282_, _09251_);
  and (_09283_, _09157_, _07959_);
  and (_09284_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_09285_, _09284_, _08975_);
  or (_09286_, _09285_, _09283_);
  nand (_09287_, _08975_, _07640_);
  and (_09288_, _09287_, _06444_);
  and (_07705_, _09288_, _09286_);
  and (_09289_, _09157_, _08019_);
  and (_09290_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_09291_, _09290_, _08975_);
  or (_09292_, _09291_, _09289_);
  nand (_09293_, _08975_, _08060_);
  and (_09294_, _09293_, _06444_);
  and (_07710_, _09294_, _09292_);
  and (_09295_, _08619_, _08524_);
  or (_09296_, _09295_, _08894_);
  and (_09297_, _08655_, _08842_);
  nand (_09298_, _08614_, _08896_);
  and (_09299_, _09298_, _08551_);
  or (_09300_, _09299_, _09297_);
  and (_09301_, _08708_, \oc8051_symbolic_cxrom1.regvalid [10]);
  not (_09302_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_09303_, _08665_, _09302_);
  and (_09304_, _09303_, _08837_);
  or (_09305_, _09304_, _09301_);
  or (_09306_, _09305_, _09300_);
  or (_09307_, _08620_, _09223_);
  and (_09308_, _09307_, \oc8051_symbolic_cxrom1.regvalid [10]);
  nor (_09309_, _08950_, _08524_);
  and (_09310_, _09309_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_09311_, _09310_, _09308_);
  or (_09312_, _09311_, _09306_);
  and (_09313_, _09312_, _09296_);
  and (_09314_, _08523_, _08489_);
  and (_09315_, _08730_, _08524_);
  and (_09316_, _09315_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_09317_, _08952_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_09318_, _08891_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_09319_, _09318_, _08620_);
  or (_09320_, _09319_, _09317_);
  or (_09321_, _09320_, _09316_);
  or (_09322_, _09321_, _09314_);
  or (_09323_, _09322_, _09313_);
  and (_07759_, _09323_, _06444_);
  nand (_09324_, _08408_, _07231_);
  nor (_09325_, _07230_, \oc8051_top_1.oc8051_decoder1.op [2]);
  nor (_09326_, _09325_, _07265_);
  and (_09327_, _09326_, _09324_);
  and (_07809_, _09327_, _06444_);
  or (_09328_, _07420_, _07159_);
  and (_09329_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  not (_09330_, _07154_);
  nor (_09331_, _07414_, _07416_);
  nand (_09332_, _09331_, _09330_);
  and (_09334_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  and (_09335_, _09334_, _09332_);
  and (_09336_, _07425_, _07070_);
  or (_09337_, _09336_, _09335_);
  or (_09338_, _09337_, _09329_);
  and (_07824_, _09338_, _06444_);
  not (_09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_09340_, _06295_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  and (_09341_, _09340_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_09342_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive );
  nor (_09343_, _06295_, _09342_);
  and (_09344_, _09343_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re );
  not (_09345_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  nor (_09346_, _09345_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  not (_09347_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  nor (_09348_, _09347_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_09349_, _09348_, _09346_);
  and (_09350_, _09349_, _09344_);
  nor (_09351_, _09350_, _09341_);
  not (_09352_, _09351_);
  and (_09353_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_09354_, _09353_, _06296_);
  not (_09355_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  nor (_09356_, _09355_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_09357_, _09356_, _09342_);
  and (_09358_, _09357_, _06295_);
  nor (_09359_, _09358_, _09354_);
  nor (_09360_, _09359_, _09344_);
  nor (_09361_, _09360_, _09352_);
  nor (_09362_, _09361_, _09339_);
  or (_09363_, _09362_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_09364_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  or (_09365_, _09364_, _09351_);
  and (_09366_, _09365_, _06444_);
  and (_07849_, _09366_, _09363_);
  and (_09367_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_09368_, _09367_, _06444_);
  or (_09369_, _09360_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  and (_09370_, _09369_, _09351_);
  and (_09371_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  or (_09372_, _09371_, _09370_);
  and (_09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _06444_);
  and (_09374_, _09373_, _09372_);
  or (_07852_, _09374_, _09368_);
  and (_09375_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_09376_, _09375_, _06444_);
  or (_09377_, _09360_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_09378_, _09377_, _09351_);
  and (_09379_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6]);
  or (_09380_, _09379_, _09378_);
  and (_09381_, _09380_, _09373_);
  or (_07855_, _09381_, _09376_);
  and (_09382_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  and (_09383_, _09382_, _06444_);
  or (_09384_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_09385_, _09384_, _09360_);
  or (_09386_, _09351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5]);
  and (_09387_, _09386_, _09373_);
  and (_09388_, _09387_, _09385_);
  or (_07860_, _09388_, _09383_);
  and (_09389_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_09390_, _09389_, _06444_);
  or (_09391_, _09360_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3]);
  and (_09392_, _09391_, _09351_);
  and (_09393_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4]);
  or (_09394_, _09393_, _09392_);
  and (_09395_, _09394_, _09373_);
  or (_07863_, _09395_, _09390_);
  or (_09396_, _08620_, _09309_);
  and (_09397_, _08666_, _08536_);
  or (_09398_, _09397_, _09396_);
  and (_09399_, _09398_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_09400_, _08613_, _08842_);
  and (_09401_, _08819_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_09402_, _09401_, _09400_);
  and (_09403_, _08708_, \oc8051_symbolic_cxrom1.regvalid [11]);
  or (_09404_, _09403_, _09223_);
  or (_09405_, _09404_, _09297_);
  or (_09406_, _09405_, _09402_);
  or (_09407_, _09406_, _09219_);
  or (_09408_, _09407_, _09399_);
  and (_07867_, _09408_, _06444_);
  or (_09409_, _09362_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_09411_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2]);
  or (_09412_, _09411_, _09351_);
  and (_09413_, _09412_, _06444_);
  and (_07876_, _09413_, _09409_);
  and (_09414_, _07912_, _07872_);
  not (_09415_, _09414_);
  and (_09416_, _09415_, _07913_);
  and (_07878_, _09416_, _06444_);
  and (_09417_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_09418_, _09417_, _06444_);
  or (_09419_, _09360_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7]);
  and (_09420_, _09419_, _09351_);
  and (_09421_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  or (_09422_, _09421_, _09420_);
  and (_09423_, _09422_, _09373_);
  or (_07909_, _09423_, _09418_);
  and (_09424_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  and (_09425_, _09424_, _06444_);
  and (_09426_, _09352_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  nor (_09427_, _09358_, _09344_);
  and (_09428_, _09427_, _09354_);
  or (_09429_, _09428_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8]);
  not (_09430_, _09341_);
  not (_09431_, _09349_);
  and (_09432_, _09431_, _09344_);
  or (_09433_, _09427_, _09432_);
  and (_09434_, _09433_, _09430_);
  and (_09436_, _09434_, _09429_);
  or (_09437_, _09436_, _09426_);
  and (_09438_, _09437_, _09373_);
  or (_07934_, _09438_, _09425_);
  nor (_09439_, _07188_, _06449_);
  and (_09440_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [4]);
  or (_09441_, _09440_, _09439_);
  and (_07954_, _09441_, _06444_);
  nor (_07964_, _07302_, rst);
  or (_09442_, _09362_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_09443_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1]);
  or (_09444_, _09443_, _09351_);
  and (_09445_, _09444_, _06444_);
  and (_07970_, _09445_, _09442_);
  and (_09447_, _09349_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_09448_, _09447_, _09359_);
  or (_09450_, _09448_, _09361_);
  and (_09451_, _09450_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_09452_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  nand (_09453_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  nor (_09454_, _09453_, _09351_);
  or (_09455_, _09454_, _09452_);
  or (_09456_, _09455_, _09451_);
  and (_07973_, _09456_, _06444_);
  and (_09457_, _08797_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_09458_, _08544_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_09459_, _08897_, _08793_);
  and (_09460_, _09459_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_09461_, _08904_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_09462_, _09461_, _08842_);
  or (_09463_, _09462_, _09460_);
  or (_09464_, _09463_, _09458_);
  or (_09465_, _09464_, _09457_);
  and (_07977_, _09465_, _06444_);
  not (_09466_, _09362_);
  and (_09467_, _06444_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_09468_, _09467_, _09466_);
  and (_09469_, _09349_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9]);
  and (_09470_, _09469_, _09359_);
  or (_09471_, _09470_, _09352_);
  and (_09472_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10]);
  and (_09473_, _09472_, _09471_);
  or (_07983_, _09473_, _09468_);
  or (_09474_, _08392_, _07232_);
  nor (_09475_, _07230_, \oc8051_top_1.oc8051_decoder1.op [1]);
  nor (_09476_, _09475_, _07265_);
  and (_09477_, _09476_, _09474_);
  and (_07992_, _09477_, _06444_);
  and (_09478_, _06944_, _08310_);
  and (_09479_, _09478_, _06941_);
  nand (_09480_, _09479_, _06978_);
  and (_09481_, _07028_, _07015_);
  not (_09482_, _09481_);
  and (_09483_, _06944_, _08977_);
  and (_09484_, _09483_, _06941_);
  nor (_09485_, _09484_, _09482_);
  not (_09486_, _09485_);
  and (_09487_, _09486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  and (_09488_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  or (_09489_, _09488_, _09487_);
  or (_09490_, _09489_, _09479_);
  and (_09491_, _09490_, _06444_);
  and (_08068_, _09491_, _09480_);
  and (_08075_, _07268_, _06444_);
  and (_09492_, _08726_, _08731_);
  or (_09493_, _09492_, \oc8051_symbolic_cxrom1.regvalid [13]);
  and (_08118_, _09493_, _06444_);
  nor (_09494_, t2_i, rst);
  and (_08140_, _09494_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r );
  not (_09495_, _07006_);
  and (_09496_, _07013_, _07011_);
  and (_09497_, _09496_, _06990_);
  nand (_09498_, _09497_, _09495_);
  or (_09499_, _09497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  and (_09500_, _09499_, _06444_);
  and (_08149_, _09500_, _09498_);
  nand (_09501_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _06444_);
  nor (_08189_, _09501_, t2ex_i);
  and (_08204_, t2ex_i, _06444_);
  nand (_09502_, _06985_, _06978_);
  not (_09503_, _06989_);
  and (_09504_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_09505_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_09506_, _09505_, _07026_);
  and (_09507_, _07011_, _06997_);
  or (_09508_, _09507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  nand (_09509_, _09507_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  and (_09510_, _09509_, _09508_);
  or (_09511_, _09510_, _09506_);
  and (_09512_, _09511_, _07035_);
  or (_09513_, _09512_, _09504_);
  or (_09514_, _09513_, _06985_);
  and (_09515_, _09514_, _09503_);
  and (_09516_, _09515_, _09502_);
  and (_09517_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_09518_, _09517_, _09516_);
  and (_08219_, _09518_, _06444_);
  or (_09519_, _08679_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_08240_, _09519_, _06444_);
  and (_09520_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_09521_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  and (_09522_, _09521_, _09332_);
  nor (_09523_, _06644_, _06587_);
  not (_09524_, _09523_);
  and (_09525_, _09524_, _08004_);
  and (_09526_, _09525_, _07998_);
  not (_09527_, _09526_);
  and (_09528_, _09527_, _07425_);
  or (_09529_, _09528_, _09522_);
  or (_09530_, _09529_, _09520_);
  and (_08409_, _09530_, _06444_);
  and (_09531_, _08875_, _08496_);
  not (_09532_, _09531_);
  not (_09533_, _08872_);
  and (_09534_, _08875_, _09533_);
  and (_09535_, _09534_, _09532_);
  and (_09536_, _09535_, _08536_);
  not (_09537_, _09536_);
  or (_09538_, _09537_, word_in[0]);
  and (_09539_, _08869_, _08894_);
  not (_09540_, _09539_);
  or (_09541_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_09542_, _09541_, _09540_);
  and (_09543_, _09542_, _09538_);
  and (_09544_, _08863_, _08790_);
  and (_09545_, _09539_, word_in[8]);
  or (_09546_, _09545_, _09544_);
  or (_09547_, _09546_, _09543_);
  and (_09548_, _08855_, _08820_);
  not (_09549_, _09548_);
  not (_09550_, _09544_);
  or (_09551_, _09550_, word_in[16]);
  and (_09552_, _09551_, _09549_);
  and (_09553_, _09552_, _09547_);
  and (_09554_, _08855_, word_in[24]);
  and (_09555_, _09554_, _09548_);
  or (_08621_, _09555_, _09553_);
  not (_09556_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_09557_, _09536_, _09556_);
  and (_09558_, _09536_, word_in[1]);
  or (_09559_, _09558_, _09557_);
  and (_09560_, _09559_, _09540_);
  and (_09562_, _09539_, word_in[9]);
  or (_09563_, _09562_, _09560_);
  and (_09564_, _09563_, _09550_);
  and (_09565_, _08863_, word_in[17]);
  and (_09567_, _09565_, _09544_);
  or (_09568_, _09567_, _09564_);
  and (_09569_, _09568_, _09549_);
  and (_09570_, _09548_, word_in[25]);
  or (_08625_, _09570_, _09569_);
  or (_09572_, _09537_, word_in[2]);
  or (_09573_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_09574_, _09573_, _09540_);
  and (_09575_, _09574_, _09572_);
  and (_09576_, _09539_, word_in[10]);
  or (_09577_, _09576_, _09544_);
  or (_09578_, _09577_, _09575_);
  or (_09579_, _09550_, word_in[18]);
  and (_09580_, _09579_, _09549_);
  and (_09581_, _09580_, _09578_);
  and (_09582_, _08855_, word_in[26]);
  and (_09583_, _09582_, _09548_);
  or (_08629_, _09583_, _09581_);
  or (_09584_, _09537_, word_in[3]);
  or (_09585_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_09586_, _09585_, _09540_);
  and (_09587_, _09586_, _09584_);
  and (_09588_, _09539_, word_in[11]);
  or (_09589_, _09588_, _09544_);
  or (_09591_, _09589_, _09587_);
  or (_09592_, _09550_, word_in[19]);
  and (_09593_, _09592_, _09549_);
  and (_09595_, _09593_, _09591_);
  and (_09596_, _08855_, word_in[27]);
  and (_09597_, _09596_, _09548_);
  or (_08633_, _09597_, _09595_);
  or (_09599_, _09537_, word_in[4]);
  or (_09600_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_09601_, _09600_, _09540_);
  and (_09602_, _09601_, _09599_);
  and (_09603_, _09539_, word_in[12]);
  or (_09604_, _09603_, _09544_);
  or (_09605_, _09604_, _09602_);
  or (_09606_, _09550_, word_in[20]);
  and (_09607_, _09606_, _09549_);
  and (_09608_, _09607_, _09605_);
  and (_09609_, _08855_, word_in[28]);
  and (_09611_, _09609_, _09548_);
  or (_08637_, _09611_, _09608_);
  or (_09612_, _09537_, word_in[5]);
  or (_09613_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_09614_, _09613_, _09540_);
  and (_09615_, _09614_, _09612_);
  and (_09616_, _09539_, word_in[13]);
  or (_09617_, _09616_, _09544_);
  or (_09618_, _09617_, _09615_);
  or (_09620_, _09550_, word_in[21]);
  and (_09621_, _09620_, _09549_);
  and (_09622_, _09621_, _09618_);
  and (_09623_, _08855_, word_in[29]);
  and (_09625_, _09623_, _09548_);
  or (_08641_, _09625_, _09622_);
  and (_09626_, _08855_, word_in[30]);
  and (_09627_, _09626_, _09548_);
  or (_09628_, _09537_, word_in[6]);
  or (_09629_, _09536_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_09631_, _09629_, _09540_);
  and (_09632_, _09631_, _09628_);
  and (_09633_, _09539_, word_in[14]);
  or (_09634_, _09633_, _09544_);
  or (_09635_, _09634_, _09632_);
  or (_09636_, _09550_, word_in[22]);
  and (_09637_, _09636_, _09549_);
  and (_09638_, _09637_, _09635_);
  or (_08647_, _09638_, _09627_);
  nor (_09639_, _09536_, _08695_);
  and (_09640_, _08875_, word_in[7]);
  and (_09641_, _09536_, _09640_);
  or (_09642_, _09641_, _09639_);
  and (_09643_, _09642_, _09540_);
  and (_09644_, _09539_, word_in[15]);
  or (_09645_, _09644_, _09544_);
  or (_09646_, _09645_, _09643_);
  or (_09647_, _09550_, word_in[23]);
  and (_09648_, _09647_, _09549_);
  and (_09649_, _09648_, _09646_);
  and (_09650_, _09548_, word_in[31]);
  or (_08650_, _09650_, _09649_);
  nor (_09651_, _07300_, _07190_);
  and (_09652_, _07190_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [3]);
  or (_09653_, _09652_, _09651_);
  and (_08690_, _09653_, _06444_);
  and (_09654_, _07429_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  and (_09655_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_09656_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_09657_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_09658_, _09657_, _09656_);
  and (_09659_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_09660_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_09661_, _09660_, _09659_);
  not (_09662_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_09663_, _07241_, _09662_);
  and (_09664_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_09665_, _09664_, _09663_);
  and (_09666_, _09665_, _09661_);
  and (_09667_, _09666_, _09658_);
  nor (_09669_, _09667_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_09670_, _09669_, _09655_);
  nor (_09671_, _09670_, _07429_);
  nor (_09672_, _09671_, _09654_);
  nor (_08694_, _09672_, rst);
  nor (_09674_, _09354_, _09344_);
  or (_09675_, _09674_, _09339_);
  and (_09676_, _09675_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  and (_09677_, _09344_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_09678_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_09679_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1]);
  nor (_09680_, _09679_, _09678_);
  and (_09681_, _09680_, _09677_);
  or (_09682_, _09681_, _09676_);
  and (_08701_, _09682_, _06444_);
  nand (_09683_, _09484_, _06978_);
  not (_09684_, _09479_);
  and (_09685_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  and (_09686_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_09687_, _09686_, _09685_);
  or (_09688_, _09687_, _09484_);
  and (_09689_, _09688_, _09684_);
  and (_09690_, _09689_, _09683_);
  and (_09691_, _09479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_09692_, _09691_, _09690_);
  and (_08719_, _09692_, _06444_);
  and (_09693_, _08863_, _08613_);
  and (_09694_, _09693_, _08732_);
  and (_09695_, _08869_, _08611_);
  and (_09696_, _09695_, _08626_);
  not (_09697_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  and (_09698_, _08875_, _08903_);
  and (_09699_, _08872_, _08497_);
  not (_09700_, _09699_);
  nor (_09701_, _09700_, _09698_);
  nor (_09702_, _09701_, _09697_);
  and (_09703_, _08875_, word_in[0]);
  and (_09704_, _09701_, _09703_);
  or (_09705_, _09704_, _09702_);
  or (_09706_, _09705_, _09696_);
  not (_09707_, _09696_);
  or (_09709_, _09707_, word_in[8]);
  and (_09710_, _09709_, _09706_);
  or (_09711_, _09710_, _09694_);
  and (_09712_, _08855_, _08790_);
  not (_09713_, _09712_);
  not (_09714_, _09694_);
  or (_09715_, _09714_, word_in[16]);
  and (_09716_, _09715_, _09713_);
  and (_09717_, _09716_, _09711_);
  and (_09718_, _09712_, word_in[24]);
  or (_08741_, _09718_, _09717_);
  and (_09719_, _09712_, word_in[25]);
  not (_09720_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  nor (_09721_, _09701_, _09720_);
  and (_09722_, _08875_, word_in[1]);
  and (_09723_, _09701_, _09722_);
  or (_09724_, _09723_, _09721_);
  or (_09726_, _09724_, _09696_);
  or (_09727_, _09707_, word_in[9]);
  and (_09728_, _09727_, _09726_);
  or (_09729_, _09728_, _09694_);
  or (_09731_, _09714_, word_in[17]);
  and (_09732_, _09731_, _09713_);
  and (_09733_, _09732_, _09729_);
  or (_08743_, _09733_, _09719_);
  not (_09734_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_09735_, _09701_, _09734_);
  and (_09736_, _08875_, word_in[2]);
  and (_09737_, _09701_, _09736_);
  or (_09738_, _09737_, _09735_);
  or (_09739_, _09738_, _09696_);
  or (_09740_, _09707_, word_in[10]);
  and (_09741_, _09740_, _09739_);
  or (_09743_, _09741_, _09694_);
  or (_09744_, _09714_, word_in[18]);
  and (_09745_, _09744_, _09713_);
  and (_09746_, _09745_, _09743_);
  and (_09747_, _09712_, word_in[26]);
  or (_08745_, _09747_, _09746_);
  and (_09748_, _09712_, word_in[27]);
  not (_09749_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_09750_, _09701_, _09749_);
  and (_09751_, _08875_, word_in[3]);
  and (_09752_, _09701_, _09751_);
  or (_09753_, _09752_, _09750_);
  or (_09754_, _09753_, _09696_);
  or (_09755_, _09707_, word_in[11]);
  and (_09756_, _09755_, _09754_);
  or (_09757_, _09756_, _09694_);
  or (_09758_, _09714_, word_in[19]);
  and (_09759_, _09758_, _09713_);
  and (_09760_, _09759_, _09757_);
  or (_08750_, _09760_, _09748_);
  not (_09761_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_09762_, _09701_, _09761_);
  and (_09763_, _08875_, word_in[4]);
  and (_09764_, _09701_, _09763_);
  or (_09765_, _09764_, _09762_);
  or (_09766_, _09765_, _09696_);
  or (_09767_, _09707_, word_in[12]);
  and (_09768_, _09767_, _09766_);
  or (_09769_, _09768_, _09694_);
  or (_09770_, _09714_, word_in[20]);
  and (_09771_, _09770_, _09713_);
  and (_09772_, _09771_, _09769_);
  and (_09773_, _09712_, word_in[28]);
  or (_08755_, _09773_, _09772_);
  and (_09774_, _09712_, word_in[29]);
  not (_09775_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  nor (_09776_, _09701_, _09775_);
  and (_09777_, _08875_, word_in[5]);
  and (_09778_, _09701_, _09777_);
  or (_09779_, _09778_, _09776_);
  or (_09780_, _09779_, _09696_);
  or (_09781_, _09707_, word_in[13]);
  and (_09782_, _09781_, _09780_);
  or (_09783_, _09782_, _09694_);
  or (_09785_, _09714_, word_in[21]);
  and (_09787_, _09785_, _09713_);
  and (_09788_, _09787_, _09783_);
  or (_08757_, _09788_, _09774_);
  and (_09790_, _09712_, word_in[30]);
  not (_09792_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  nor (_09794_, _09701_, _09792_);
  and (_09795_, _08875_, word_in[6]);
  and (_09797_, _09701_, _09795_);
  or (_09798_, _09797_, _09794_);
  or (_09800_, _09798_, _09696_);
  or (_09802_, _09707_, word_in[14]);
  and (_09803_, _09802_, _09800_);
  or (_09804_, _09803_, _09694_);
  or (_09805_, _09714_, word_in[22]);
  and (_09806_, _09805_, _09713_);
  and (_09807_, _09806_, _09804_);
  or (_08762_, _09807_, _09790_);
  nor (_09808_, _09701_, _08600_);
  and (_09809_, _09701_, _09640_);
  or (_09810_, _09809_, _09808_);
  or (_09811_, _09810_, _09696_);
  or (_09812_, _09707_, word_in[15]);
  and (_09813_, _09812_, _09811_);
  or (_09814_, _09813_, _09694_);
  or (_09815_, _09714_, word_in[23]);
  and (_09816_, _09815_, _09713_);
  and (_09817_, _09816_, _09814_);
  and (_09818_, _09712_, word_in[31]);
  or (_08767_, _09818_, _09817_);
  and (_09819_, _08869_, _08644_);
  and (_09820_, _09819_, _08626_);
  not (_09821_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_09822_, _09531_, _09533_);
  and (_09823_, _09822_, _08536_);
  nor (_09824_, _09823_, _09821_);
  and (_09825_, _09823_, _09703_);
  or (_09826_, _09825_, _09824_);
  or (_09827_, _09826_, _09820_);
  and (_09828_, _08863_, _08611_);
  and (_09829_, _09828_, _08732_);
  not (_09830_, _09829_);
  not (_09831_, _09820_);
  or (_09832_, _09831_, word_in[8]);
  and (_09833_, _09832_, _09830_);
  and (_09834_, _09833_, _09827_);
  and (_09835_, _08855_, _08613_);
  and (_09836_, _09835_, _08814_);
  and (_09837_, _08863_, word_in[16]);
  and (_09838_, _09829_, _09837_);
  or (_09839_, _09838_, _09836_);
  or (_09840_, _09839_, _09834_);
  not (_09841_, _09836_);
  or (_09842_, _09841_, word_in[24]);
  and (_08851_, _09842_, _09840_);
  not (_09843_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  nor (_09844_, _09823_, _09843_);
  and (_09845_, _09823_, _09722_);
  or (_09846_, _09845_, _09844_);
  or (_09847_, _09846_, _09820_);
  or (_09848_, _09831_, word_in[9]);
  and (_09850_, _09848_, _09830_);
  and (_09851_, _09850_, _09847_);
  and (_09853_, _09829_, word_in[17]);
  or (_09854_, _09853_, _09836_);
  or (_09855_, _09854_, _09851_);
  or (_09856_, _09841_, word_in[25]);
  and (_08854_, _09856_, _09855_);
  not (_09857_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  nor (_09858_, _09823_, _09857_);
  and (_09860_, _09823_, _09736_);
  or (_09861_, _09860_, _09858_);
  or (_09862_, _09861_, _09820_);
  or (_09864_, _09831_, word_in[10]);
  and (_09865_, _09864_, _09830_);
  and (_09866_, _09865_, _09862_);
  and (_09867_, _09829_, word_in[18]);
  or (_09868_, _09867_, _09866_);
  and (_09869_, _09868_, _09841_);
  and (_09870_, _09836_, word_in[26]);
  or (_08858_, _09870_, _09869_);
  not (_09871_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  nor (_09873_, _09823_, _09871_);
  and (_09874_, _09823_, _09751_);
  or (_09875_, _09874_, _09873_);
  or (_09876_, _09875_, _09820_);
  or (_09878_, _09831_, word_in[11]);
  and (_09879_, _09878_, _09830_);
  and (_09881_, _09879_, _09876_);
  and (_09882_, _09829_, word_in[19]);
  or (_09883_, _09882_, _09836_);
  or (_09885_, _09883_, _09881_);
  or (_09886_, _09841_, word_in[27]);
  and (_08861_, _09886_, _09885_);
  and (_09888_, _09829_, word_in[20]);
  not (_09889_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  nor (_09891_, _09823_, _09889_);
  and (_09892_, _09823_, _09763_);
  or (_09893_, _09892_, _09891_);
  or (_09895_, _09893_, _09820_);
  or (_09896_, _09831_, word_in[12]);
  and (_09897_, _09896_, _09830_);
  and (_09898_, _09897_, _09895_);
  or (_09899_, _09898_, _09888_);
  and (_09900_, _09899_, _09841_);
  and (_09901_, _09836_, word_in[28]);
  or (_08864_, _09901_, _09900_);
  or (_09902_, _09823_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  not (_09903_, _09823_);
  or (_09904_, _09903_, _09777_);
  and (_09905_, _09904_, _09902_);
  or (_09906_, _09905_, _09820_);
  or (_09907_, _09831_, word_in[13]);
  and (_09908_, _09907_, _09906_);
  or (_09909_, _09908_, _09829_);
  or (_09910_, _09830_, word_in[21]);
  and (_09911_, _09910_, _09841_);
  and (_09912_, _09911_, _09909_);
  and (_09913_, _09836_, word_in[29]);
  or (_14580_, _09913_, _09912_);
  and (_09914_, _09829_, word_in[22]);
  not (_09915_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_09916_, _09823_, _09915_);
  and (_09917_, _09823_, _09795_);
  or (_09918_, _09917_, _09916_);
  or (_09919_, _09918_, _09820_);
  or (_09920_, _09831_, word_in[14]);
  and (_09921_, _09920_, _09830_);
  and (_09922_, _09921_, _09919_);
  or (_09923_, _09922_, _09914_);
  and (_09924_, _09923_, _09841_);
  and (_09925_, _09836_, word_in[30]);
  or (_08873_, _09925_, _09924_);
  nor (_09926_, _09823_, _08700_);
  and (_09927_, _09823_, _09640_);
  or (_09928_, _09927_, _09926_);
  or (_09929_, _09928_, _09820_);
  or (_09930_, _09831_, word_in[15]);
  and (_09931_, _09930_, _09830_);
  and (_09932_, _09931_, _09929_);
  and (_09933_, _09829_, word_in[23]);
  or (_09934_, _09933_, _09836_);
  or (_09935_, _09934_, _09932_);
  or (_09936_, _09841_, word_in[31]);
  and (_08876_, _09936_, _09935_);
  and (_09937_, _08855_, _09309_);
  and (_09938_, _09937_, word_in[24]);
  and (_09939_, _08863_, _08644_);
  and (_09940_, _09939_, _08732_);
  not (_09941_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  not (_09942_, _08874_);
  nor (_09943_, _09698_, _09942_);
  nor (_09944_, _09943_, _09941_);
  and (_09945_, _09943_, _09703_);
  or (_09946_, _09945_, _09944_);
  and (_09947_, _08870_, _08626_);
  or (_09948_, _09947_, _09946_);
  not (_09950_, _09947_);
  or (_09951_, _09950_, word_in[8]);
  and (_09952_, _09951_, _09948_);
  or (_09953_, _09952_, _09940_);
  not (_09954_, _09937_);
  not (_09956_, _09940_);
  or (_09957_, _09956_, word_in[16]);
  and (_09959_, _09957_, _09954_);
  and (_09961_, _09959_, _09953_);
  or (_14581_, _09961_, _09938_);
  not (_09963_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_09965_, _09943_, _09963_);
  and (_09966_, _09943_, _09722_);
  or (_09968_, _09966_, _09965_);
  or (_09970_, _09968_, _09947_);
  or (_09971_, _09950_, word_in[9]);
  and (_09973_, _09971_, _09970_);
  or (_09975_, _09973_, _09940_);
  or (_09977_, _09956_, word_in[17]);
  and (_09978_, _09977_, _09954_);
  and (_09980_, _09978_, _09975_);
  and (_09982_, _09937_, word_in[25]);
  or (_08943_, _09982_, _09980_);
  and (_09984_, _09937_, word_in[26]);
  not (_09985_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  nor (_09986_, _09943_, _09985_);
  and (_09987_, _09943_, _09736_);
  or (_09988_, _09987_, _09986_);
  or (_09989_, _09988_, _09947_);
  or (_09990_, _09950_, word_in[10]);
  and (_09991_, _09990_, _09989_);
  or (_09992_, _09991_, _09940_);
  or (_09993_, _09956_, word_in[18]);
  and (_09994_, _09993_, _09954_);
  and (_09995_, _09994_, _09992_);
  or (_08945_, _09995_, _09984_);
  and (_09997_, _09937_, word_in[27]);
  not (_09998_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  nor (_09999_, _09943_, _09998_);
  and (_10000_, _09943_, _09751_);
  or (_10001_, _10000_, _09999_);
  or (_10002_, _10001_, _09947_);
  or (_10003_, _09950_, word_in[11]);
  and (_10004_, _10003_, _10002_);
  or (_10005_, _10004_, _09940_);
  or (_10006_, _09956_, word_in[19]);
  and (_10007_, _10006_, _09954_);
  and (_10008_, _10007_, _10005_);
  or (_08948_, _10008_, _09997_);
  and (_10010_, _09943_, _09763_);
  not (_10011_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  nor (_10013_, _09943_, _10011_);
  nor (_10014_, _10013_, _10010_);
  nor (_10015_, _10014_, _09947_);
  and (_10016_, _09947_, word_in[12]);
  or (_10018_, _10016_, _10015_);
  and (_10019_, _10018_, _09956_);
  and (_10020_, _08863_, word_in[20]);
  and (_10021_, _09940_, _10020_);
  or (_10022_, _10021_, _09937_);
  or (_10023_, _10022_, _10019_);
  or (_10024_, _09954_, word_in[28]);
  and (_08951_, _10024_, _10023_);
  and (_10026_, _09937_, word_in[29]);
  not (_10027_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  nor (_10028_, _09943_, _10027_);
  and (_10030_, _09943_, _09777_);
  or (_10031_, _10030_, _10028_);
  or (_10032_, _10031_, _09947_);
  or (_10033_, _09950_, word_in[13]);
  and (_10034_, _10033_, _10032_);
  or (_10035_, _10034_, _09940_);
  or (_10036_, _09956_, word_in[21]);
  and (_10038_, _10036_, _09954_);
  and (_10039_, _10038_, _10035_);
  or (_08954_, _10039_, _10026_);
  and (_10041_, _09937_, word_in[30]);
  not (_10042_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  nor (_10043_, _09943_, _10042_);
  and (_10044_, _09943_, _09795_);
  or (_10045_, _10044_, _10043_);
  or (_10046_, _10045_, _09947_);
  or (_10047_, _09950_, word_in[14]);
  and (_10048_, _10047_, _10046_);
  or (_10049_, _10048_, _09940_);
  or (_10050_, _09956_, word_in[22]);
  and (_10051_, _10050_, _09954_);
  and (_10052_, _10051_, _10049_);
  or (_08957_, _10052_, _10041_);
  nor (_10054_, _09943_, _08584_);
  and (_10055_, _09943_, _09640_);
  or (_10056_, _10055_, _10054_);
  or (_10057_, _10056_, _09947_);
  or (_10058_, _09950_, word_in[15]);
  and (_10059_, _10058_, _10057_);
  or (_10060_, _10059_, _09940_);
  or (_10061_, _09956_, word_in[23]);
  and (_10062_, _10061_, _09954_);
  and (_10063_, _10062_, _10060_);
  and (_10064_, _09937_, word_in[31]);
  or (_08960_, _10064_, _10063_);
  and (_10065_, _08865_, _08770_);
  and (_10066_, _10065_, _08655_);
  and (_10067_, _08869_, _08930_);
  not (_10068_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_10069_, _09531_, _08872_);
  and (_10070_, _08875_, _08904_);
  and (_10071_, _10070_, _10069_);
  nor (_10072_, _10071_, _10068_);
  and (_10073_, _10071_, word_in[0]);
  or (_10074_, _10073_, _10072_);
  or (_10075_, _10074_, _10067_);
  not (_10076_, _10067_);
  or (_10077_, _10076_, word_in[8]);
  and (_10078_, _10077_, _10075_);
  or (_10079_, _10078_, _10066_);
  and (_10080_, _08855_, _08897_);
  not (_10081_, _10080_);
  not (_10082_, _10066_);
  or (_10083_, _10082_, _09837_);
  and (_10084_, _10083_, _10081_);
  and (_10085_, _10084_, _10079_);
  and (_10086_, _10080_, word_in[24]);
  or (_09044_, _10086_, _10085_);
  not (_10087_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_10088_, _10071_, _10087_);
  and (_10089_, _10071_, word_in[1]);
  or (_10090_, _10089_, _10088_);
  or (_10091_, _10090_, _10067_);
  or (_10092_, _10076_, word_in[9]);
  and (_10093_, _10092_, _10091_);
  or (_10094_, _10093_, _10066_);
  or (_10095_, _10082_, _09565_);
  and (_10096_, _10095_, _10081_);
  and (_10097_, _10096_, _10094_);
  and (_10098_, _10080_, word_in[25]);
  or (_09047_, _10098_, _10097_);
  and (_10099_, _08863_, word_in[18]);
  and (_10100_, _10066_, _10099_);
  not (_10101_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_10102_, _10071_, _10101_);
  and (_10103_, _10071_, word_in[2]);
  or (_10104_, _10103_, _10102_);
  and (_10105_, _10104_, _10076_);
  and (_10106_, _10067_, word_in[10]);
  or (_10107_, _10106_, _10105_);
  and (_10108_, _10107_, _10082_);
  or (_10109_, _10108_, _10100_);
  and (_10110_, _10109_, _10081_);
  and (_10111_, _10080_, word_in[26]);
  or (_14582_, _10111_, _10110_);
  and (_10112_, _07159_, _06439_);
  nand (_10113_, _10112_, _06666_);
  or (_10114_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [5]);
  and (_10115_, _10114_, _06444_);
  and (_09050_, _10115_, _10113_);
  and (_10116_, _08863_, word_in[19]);
  and (_10117_, _10066_, _10116_);
  not (_10118_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_10119_, _10071_, _10118_);
  and (_10120_, _10071_, word_in[3]);
  or (_10121_, _10120_, _10119_);
  and (_10122_, _10121_, _10076_);
  and (_10123_, _10067_, word_in[11]);
  or (_10124_, _10123_, _10122_);
  and (_10125_, _10124_, _10082_);
  or (_10126_, _10125_, _10117_);
  and (_10127_, _10126_, _10081_);
  and (_10128_, _10080_, word_in[27]);
  or (_14583_, _10128_, _10127_);
  not (_10129_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_10130_, _10071_, _10129_);
  and (_10131_, _10071_, word_in[4]);
  or (_10132_, _10131_, _10130_);
  or (_10133_, _10132_, _10067_);
  or (_10134_, _10076_, word_in[12]);
  and (_10135_, _10134_, _10133_);
  or (_10136_, _10135_, _10066_);
  or (_10137_, _10082_, _10020_);
  and (_10138_, _10137_, _10081_);
  and (_10139_, _10138_, _10136_);
  and (_10140_, _10080_, word_in[28]);
  or (_14584_, _10140_, _10139_);
  not (_10141_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_10142_, _10071_, _10141_);
  and (_10143_, _10071_, word_in[5]);
  or (_10144_, _10143_, _10142_);
  or (_10145_, _10144_, _10067_);
  or (_10146_, _10076_, word_in[13]);
  and (_10147_, _10146_, _10145_);
  or (_10148_, _10147_, _10066_);
  and (_10149_, _08863_, word_in[21]);
  or (_10150_, _10082_, _10149_);
  and (_10151_, _10150_, _10081_);
  and (_10152_, _10151_, _10148_);
  and (_10153_, _10080_, word_in[29]);
  or (_14585_, _10153_, _10152_);
  and (_10154_, _08863_, word_in[22]);
  and (_10155_, _10066_, _10154_);
  not (_10156_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_10157_, _10071_, _10156_);
  and (_10158_, _10071_, word_in[6]);
  or (_10159_, _10158_, _10157_);
  and (_10160_, _10159_, _10076_);
  and (_10161_, _10067_, word_in[14]);
  or (_10162_, _10161_, _10160_);
  and (_10163_, _10162_, _10082_);
  or (_10164_, _10163_, _10155_);
  and (_10165_, _10164_, _10081_);
  and (_10166_, _10080_, word_in[30]);
  or (_09058_, _10166_, _10165_);
  nor (_10167_, _10071_, _08709_);
  and (_10168_, _10071_, word_in[7]);
  or (_10169_, _10168_, _10167_);
  or (_10170_, _10169_, _10067_);
  or (_10171_, _10076_, word_in[15]);
  and (_10172_, _10171_, _10170_);
  or (_10173_, _10172_, _10066_);
  or (_10174_, _10082_, _08886_);
  and (_10175_, _10174_, _10081_);
  and (_10176_, _10175_, _10173_);
  and (_10177_, _10080_, word_in[31]);
  or (_09061_, _10177_, _10176_);
  and (_10178_, _10065_, _08613_);
  not (_10179_, _10178_);
  and (_10180_, _09695_, _08708_);
  and (_10181_, _10070_, _09699_);
  and (_10182_, _10181_, word_in[0]);
  not (_10183_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_10184_, _10181_, _10183_);
  nor (_10185_, _10184_, _10182_);
  nor (_10186_, _10185_, _10180_);
  and (_10187_, _10180_, word_in[8]);
  or (_10188_, _10187_, _10186_);
  and (_10189_, _10188_, _10179_);
  and (_10190_, _10178_, _09837_);
  or (_10191_, _10190_, _10189_);
  and (_10192_, _08855_, _08898_);
  not (_10193_, _10192_);
  and (_10194_, _10193_, _10191_);
  and (_10195_, _10192_, word_in[24]);
  or (_09148_, _10195_, _10194_);
  and (_10196_, _10181_, word_in[1]);
  not (_10197_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_10198_, _10181_, _10197_);
  nor (_10199_, _10198_, _10196_);
  nor (_10200_, _10199_, _10180_);
  and (_10201_, _10180_, word_in[9]);
  or (_10202_, _10201_, _10200_);
  and (_10203_, _10202_, _10179_);
  and (_10204_, _10178_, _09565_);
  or (_10205_, _10204_, _10203_);
  and (_10206_, _10205_, _10193_);
  and (_10207_, _10192_, word_in[25]);
  or (_09150_, _10207_, _10206_);
  and (_10208_, _10181_, word_in[2]);
  not (_10209_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_10210_, _10181_, _10209_);
  nor (_10211_, _10210_, _10208_);
  nor (_10212_, _10211_, _10180_);
  and (_10213_, _10180_, word_in[10]);
  or (_10214_, _10213_, _10212_);
  and (_10215_, _10214_, _10179_);
  and (_10216_, _10178_, _10099_);
  or (_10217_, _10216_, _10215_);
  and (_10218_, _10217_, _10193_);
  and (_10219_, _10192_, word_in[26]);
  or (_09153_, _10219_, _10218_);
  and (_10220_, _10181_, word_in[3]);
  not (_10221_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_10222_, _10181_, _10221_);
  nor (_10223_, _10222_, _10220_);
  nor (_10224_, _10223_, _10180_);
  and (_10225_, _10180_, word_in[11]);
  or (_10226_, _10225_, _10224_);
  and (_10227_, _10226_, _10179_);
  and (_10228_, _10178_, _10116_);
  or (_10229_, _10228_, _10227_);
  and (_10230_, _10229_, _10193_);
  and (_10231_, _10192_, word_in[27]);
  or (_09156_, _10231_, _10230_);
  and (_10232_, _10181_, word_in[4]);
  not (_10233_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_10234_, _10181_, _10233_);
  nor (_10235_, _10234_, _10232_);
  nor (_10236_, _10235_, _10180_);
  and (_10237_, _10180_, word_in[12]);
  or (_10238_, _10237_, _10236_);
  and (_10239_, _10238_, _10179_);
  and (_10240_, _10178_, _10020_);
  or (_10241_, _10240_, _10239_);
  and (_10242_, _10241_, _10193_);
  and (_10243_, _10192_, word_in[28]);
  or (_09159_, _10243_, _10242_);
  and (_10244_, _10181_, word_in[5]);
  not (_10245_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_10246_, _10181_, _10245_);
  nor (_10247_, _10246_, _10244_);
  nor (_10248_, _10247_, _10180_);
  and (_10249_, _10180_, word_in[13]);
  or (_10250_, _10249_, _10248_);
  and (_10251_, _10250_, _10179_);
  and (_10252_, _10178_, _10149_);
  or (_10253_, _10252_, _10251_);
  and (_10254_, _10253_, _10193_);
  and (_10255_, _10192_, word_in[29]);
  or (_09162_, _10255_, _10254_);
  and (_10256_, _10178_, _10154_);
  and (_10257_, _10181_, word_in[6]);
  not (_10258_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_10259_, _10181_, _10258_);
  nor (_10260_, _10259_, _10257_);
  nor (_10261_, _10260_, _10180_);
  and (_10262_, _10180_, word_in[14]);
  or (_10263_, _10262_, _10261_);
  and (_10264_, _10263_, _10179_);
  or (_10265_, _10264_, _10256_);
  and (_10266_, _10265_, _10193_);
  and (_10267_, _10192_, word_in[30]);
  or (_09166_, _10267_, _10266_);
  and (_10268_, _10181_, word_in[7]);
  nor (_10269_, _10181_, _08595_);
  nor (_10270_, _10269_, _10268_);
  nor (_10271_, _10270_, _10180_);
  and (_10272_, _10180_, word_in[15]);
  or (_10273_, _10272_, _10271_);
  and (_10274_, _10273_, _10179_);
  and (_10275_, _10178_, _08886_);
  or (_10276_, _10275_, _10274_);
  and (_10277_, _10276_, _10193_);
  and (_10278_, _10192_, word_in[31]);
  or (_09170_, _10278_, _10277_);
  nand (_10279_, _10112_, _07300_);
  or (_10280_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [3]);
  and (_10281_, _10280_, _06444_);
  and (_09234_, _10281_, _10279_);
  and (_10282_, _08855_, _08930_);
  not (_10283_, _10282_);
  and (_10284_, _10065_, _08611_);
  and (_10285_, _10284_, _09837_);
  not (_10286_, _10284_);
  and (_10287_, _09819_, _08708_);
  and (_10288_, _09822_, _08904_);
  and (_10289_, _10288_, word_in[0]);
  not (_10290_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  nor (_10291_, _10288_, _10290_);
  nor (_10292_, _10291_, _10289_);
  nor (_10293_, _10292_, _10287_);
  and (_10294_, _10287_, word_in[8]);
  or (_10295_, _10294_, _10293_);
  and (_10296_, _10295_, _10286_);
  or (_10297_, _10296_, _10285_);
  and (_10298_, _10297_, _10283_);
  and (_10299_, _10282_, word_in[24]);
  or (_09240_, _10299_, _10298_);
  and (_10300_, _10284_, _09565_);
  not (_10301_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  nor (_10302_, _10288_, _10301_);
  and (_10303_, _10288_, word_in[1]);
  nor (_10304_, _10303_, _10302_);
  nor (_10305_, _10304_, _10287_);
  and (_10306_, _10287_, word_in[9]);
  or (_10307_, _10306_, _10305_);
  and (_10308_, _10307_, _10286_);
  or (_10309_, _10308_, _10300_);
  and (_10310_, _10309_, _10283_);
  and (_10311_, _10282_, word_in[25]);
  or (_09245_, _10311_, _10310_);
  and (_10312_, _10284_, _10099_);
  not (_10313_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  nor (_10314_, _10288_, _10313_);
  and (_10315_, _10288_, word_in[2]);
  nor (_10316_, _10315_, _10314_);
  nor (_10317_, _10316_, _10287_);
  and (_10318_, _10287_, word_in[10]);
  or (_10319_, _10318_, _10317_);
  and (_10320_, _10319_, _10286_);
  or (_10321_, _10320_, _10312_);
  and (_10322_, _10321_, _10283_);
  and (_10323_, _10282_, word_in[26]);
  or (_09248_, _10323_, _10322_);
  and (_10324_, _10284_, _10116_);
  not (_10325_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  nor (_10326_, _10288_, _10325_);
  and (_10327_, _10288_, word_in[3]);
  nor (_10328_, _10327_, _10326_);
  nor (_10329_, _10328_, _10287_);
  and (_10330_, _10287_, word_in[11]);
  or (_10331_, _10330_, _10329_);
  and (_10332_, _10331_, _10286_);
  or (_10333_, _10332_, _10324_);
  and (_10334_, _10333_, _10283_);
  and (_10335_, _10282_, word_in[27]);
  or (_09253_, _10335_, _10334_);
  and (_10336_, _10284_, _10020_);
  not (_10337_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  nor (_10338_, _10288_, _10337_);
  and (_10339_, _10288_, word_in[4]);
  nor (_10340_, _10339_, _10338_);
  nor (_10341_, _10340_, _10287_);
  and (_10342_, _10287_, word_in[12]);
  or (_10343_, _10342_, _10341_);
  and (_10344_, _10343_, _10286_);
  or (_10346_, _10344_, _10336_);
  and (_10347_, _10346_, _10283_);
  and (_10348_, _10282_, word_in[28]);
  or (_09258_, _10348_, _10347_);
  and (_10349_, _10284_, _10149_);
  not (_10350_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  nor (_10351_, _10288_, _10350_);
  and (_10352_, _10288_, word_in[5]);
  nor (_10353_, _10352_, _10351_);
  nor (_10355_, _10353_, _10287_);
  and (_10356_, _10287_, word_in[13]);
  or (_10358_, _10356_, _10355_);
  and (_10359_, _10358_, _10286_);
  or (_10360_, _10359_, _10349_);
  and (_10361_, _10360_, _10283_);
  and (_10363_, _10282_, word_in[29]);
  or (_09261_, _10363_, _10361_);
  and (_10365_, _10284_, _10154_);
  not (_10366_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  nor (_10367_, _10288_, _10366_);
  and (_10368_, _10288_, word_in[6]);
  nor (_10369_, _10368_, _10367_);
  nor (_10370_, _10369_, _10287_);
  and (_10371_, _10287_, word_in[14]);
  or (_10372_, _10371_, _10370_);
  and (_10373_, _10372_, _10286_);
  or (_10374_, _10373_, _10365_);
  and (_10375_, _10374_, _10283_);
  and (_10376_, _10282_, word_in[30]);
  or (_09265_, _10376_, _10375_);
  and (_10377_, _10284_, _08886_);
  nor (_10378_, _10288_, _08714_);
  and (_10379_, _10288_, word_in[7]);
  nor (_10380_, _10379_, _10378_);
  nor (_10381_, _10380_, _10287_);
  and (_10382_, _10287_, word_in[15]);
  or (_10383_, _10382_, _10381_);
  and (_10384_, _10383_, _10286_);
  or (_10385_, _10384_, _10377_);
  and (_10386_, _10385_, _10283_);
  and (_10387_, _10282_, word_in[31]);
  or (_09270_, _10387_, _10386_);
  and (_10388_, _08855_, _08905_);
  not (_10389_, _10388_);
  and (_10390_, _10065_, _08644_);
  and (_10391_, _10390_, _09837_);
  not (_10392_, _10390_);
  and (_10393_, _08870_, _08708_);
  and (_10394_, _10070_, _08874_);
  and (_10395_, _10394_, word_in[0]);
  not (_10396_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  nor (_10397_, _10394_, _10396_);
  nor (_10398_, _10397_, _10395_);
  nor (_10399_, _10398_, _10393_);
  and (_10400_, _10393_, word_in[8]);
  or (_10401_, _10400_, _10399_);
  and (_10402_, _10401_, _10392_);
  or (_10403_, _10402_, _10391_);
  and (_10404_, _10403_, _10389_);
  and (_10405_, _10388_, word_in[24]);
  or (_14586_, _10405_, _10404_);
  not (_10406_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  nor (_10407_, _10394_, _10406_);
  and (_10408_, _10394_, word_in[1]);
  nor (_10409_, _10408_, _10407_);
  nor (_10410_, _10409_, _10393_);
  and (_10411_, _10393_, word_in[9]);
  or (_10412_, _10411_, _10410_);
  and (_10413_, _10412_, _10392_);
  and (_10414_, _10390_, _09565_);
  or (_10415_, _10414_, _10413_);
  and (_10416_, _10415_, _10389_);
  and (_10417_, _10388_, word_in[25]);
  or (_14587_, _10417_, _10416_);
  and (_10418_, _10390_, _10099_);
  and (_10419_, _10394_, word_in[2]);
  not (_10420_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  nor (_10421_, _10394_, _10420_);
  nor (_10422_, _10421_, _10419_);
  nor (_10423_, _10422_, _10393_);
  and (_10424_, _10393_, word_in[10]);
  or (_10425_, _10424_, _10423_);
  and (_10426_, _10425_, _10392_);
  or (_10427_, _10426_, _10418_);
  and (_10428_, _10427_, _10389_);
  and (_10429_, _10388_, word_in[26]);
  or (_14588_, _10429_, _10428_);
  and (_10430_, _10394_, word_in[3]);
  not (_10431_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  nor (_10432_, _10394_, _10431_);
  nor (_10433_, _10432_, _10430_);
  nor (_10434_, _10433_, _10393_);
  and (_10435_, _10393_, word_in[11]);
  or (_10436_, _10435_, _10434_);
  and (_10437_, _10436_, _10392_);
  and (_10438_, _10390_, _10116_);
  or (_10439_, _10438_, _10437_);
  and (_10440_, _10439_, _10389_);
  and (_10441_, _10388_, word_in[27]);
  or (_14589_, _10441_, _10440_);
  and (_10442_, _10394_, word_in[4]);
  not (_10443_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  nor (_10444_, _10394_, _10443_);
  nor (_10445_, _10444_, _10442_);
  nor (_10446_, _10445_, _10393_);
  and (_10447_, _10393_, word_in[12]);
  or (_10448_, _10447_, _10446_);
  and (_10449_, _10448_, _10392_);
  and (_10450_, _10390_, _10020_);
  or (_10451_, _10450_, _10449_);
  and (_10452_, _10451_, _10389_);
  and (_10453_, _10388_, word_in[28]);
  or (_14590_, _10453_, _10452_);
  not (_10454_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  nor (_10455_, _10394_, _10454_);
  and (_10456_, _10394_, word_in[5]);
  or (_10457_, _10456_, _10455_);
  or (_10458_, _10457_, _10393_);
  not (_10459_, _10393_);
  or (_10460_, _10459_, word_in[13]);
  and (_10461_, _10460_, _10458_);
  or (_10462_, _10461_, _10390_);
  or (_10463_, _10392_, _10149_);
  and (_10464_, _10463_, _10462_);
  and (_10465_, _10464_, _10389_);
  and (_10466_, _10388_, word_in[29]);
  or (_14591_, _10466_, _10465_);
  and (_10467_, _10394_, word_in[6]);
  not (_10469_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  nor (_10470_, _10394_, _10469_);
  nor (_10471_, _10470_, _10467_);
  nor (_10472_, _10471_, _10393_);
  and (_10473_, _10393_, word_in[14]);
  or (_10474_, _10473_, _10472_);
  and (_10475_, _10474_, _10392_);
  and (_10476_, _10390_, _10154_);
  or (_10477_, _10476_, _10475_);
  and (_10478_, _10477_, _10389_);
  and (_10479_, _10388_, word_in[30]);
  or (_14592_, _10479_, _10478_);
  or (_10480_, _10392_, _08886_);
  nor (_10481_, _10394_, _08590_);
  and (_10482_, _10394_, word_in[7]);
  or (_10483_, _10482_, _10481_);
  or (_10484_, _10483_, _10393_);
  or (_10485_, _10459_, word_in[15]);
  and (_10486_, _10485_, _10484_);
  or (_10487_, _10486_, _10390_);
  and (_10488_, _10487_, _10480_);
  or (_10489_, _10488_, _10388_);
  or (_10490_, _10389_, word_in[31]);
  and (_14593_, _10490_, _10489_);
  nor (_10491_, _06732_, _06644_);
  not (_10492_, _10491_);
  and (_10493_, _10492_, _09030_);
  and (_10494_, _10493_, _09019_);
  nor (_10495_, _10494_, _07190_);
  and (_10496_, _07156_, _06439_);
  or (_10497_, _10496_, _07161_);
  and (_10498_, _10497_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  or (_10499_, _10498_, _10495_);
  and (_09410_, _10499_, _06444_);
  and (_10500_, _08855_, _08800_);
  and (_10501_, _10500_, _08644_);
  and (_10502_, _08863_, _08952_);
  and (_10503_, _08869_, _08620_);
  not (_10504_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_10505_, _08875_, _08538_);
  and (_10506_, _10505_, _10069_);
  nor (_10507_, _10506_, _10504_);
  and (_10508_, _10506_, word_in[0]);
  or (_10509_, _10508_, _10507_);
  or (_10510_, _10509_, _10503_);
  not (_10511_, _10503_);
  or (_10512_, _10511_, word_in[8]);
  and (_10513_, _10512_, _10510_);
  or (_10514_, _10513_, _10502_);
  not (_10515_, _10502_);
  or (_10516_, _10515_, word_in[16]);
  and (_10517_, _10516_, _10514_);
  or (_10518_, _10517_, _10501_);
  not (_10519_, _10501_);
  or (_10520_, _10519_, word_in[24]);
  and (_09446_, _10520_, _10518_);
  and (_10521_, _10502_, word_in[17]);
  not (_10522_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_10523_, _10506_, _10522_);
  and (_10524_, _10506_, word_in[1]);
  or (_10525_, _10524_, _10523_);
  and (_10526_, _10525_, _10511_);
  and (_10527_, _10503_, word_in[9]);
  or (_10528_, _10527_, _10526_);
  and (_10529_, _10528_, _10515_);
  or (_10530_, _10529_, _10521_);
  and (_10531_, _10530_, _10519_);
  and (_10532_, _10501_, word_in[25]);
  or (_09449_, _10532_, _10531_);
  and (_10533_, _10502_, word_in[18]);
  not (_10534_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_10535_, _10506_, _10534_);
  and (_10536_, _10506_, word_in[2]);
  or (_10537_, _10536_, _10535_);
  and (_10538_, _10537_, _10511_);
  and (_10539_, _10503_, word_in[10]);
  or (_10540_, _10539_, _10538_);
  and (_10541_, _10540_, _10515_);
  or (_10542_, _10541_, _10533_);
  and (_10543_, _10542_, _10519_);
  and (_10544_, _10501_, word_in[26]);
  or (_14594_, _10544_, _10543_);
  and (_10545_, _10502_, word_in[19]);
  not (_10546_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_10547_, _10506_, _10546_);
  and (_10548_, _10506_, word_in[3]);
  or (_10549_, _10548_, _10547_);
  and (_10550_, _10549_, _10511_);
  and (_10551_, _10503_, word_in[11]);
  or (_10552_, _10551_, _10550_);
  and (_10553_, _10552_, _10515_);
  or (_10554_, _10553_, _10545_);
  and (_10555_, _10554_, _10519_);
  and (_10556_, _10501_, word_in[27]);
  or (_14595_, _10556_, _10555_);
  and (_10557_, _10502_, word_in[20]);
  not (_10558_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_10559_, _10506_, _10558_);
  and (_10561_, _10506_, word_in[4]);
  or (_10562_, _10561_, _10559_);
  and (_10563_, _10562_, _10511_);
  and (_10564_, _10503_, word_in[12]);
  or (_10565_, _10564_, _10563_);
  and (_10566_, _10565_, _10515_);
  or (_10567_, _10566_, _10557_);
  and (_10568_, _10567_, _10519_);
  and (_10569_, _10501_, word_in[28]);
  or (_14596_, _10569_, _10568_);
  and (_10570_, _10502_, word_in[21]);
  not (_10571_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_10572_, _10506_, _10571_);
  and (_10573_, _10506_, word_in[5]);
  or (_10574_, _10573_, _10572_);
  and (_10575_, _10574_, _10511_);
  and (_10576_, _10503_, word_in[13]);
  or (_10577_, _10576_, _10575_);
  and (_10578_, _10577_, _10515_);
  or (_10579_, _10578_, _10570_);
  and (_10580_, _10579_, _10519_);
  and (_10581_, _10501_, word_in[29]);
  or (_14597_, _10581_, _10580_);
  and (_10582_, _10502_, word_in[22]);
  not (_10583_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_10584_, _10506_, _10583_);
  and (_10585_, _10506_, word_in[6]);
  or (_10586_, _10585_, _10584_);
  and (_10587_, _10586_, _10511_);
  and (_10588_, _10503_, word_in[14]);
  or (_10589_, _10588_, _10587_);
  and (_10590_, _10589_, _10515_);
  or (_10591_, _10590_, _10582_);
  and (_10592_, _10591_, _10519_);
  and (_10593_, _10501_, word_in[30]);
  or (_14598_, _10593_, _10592_);
  and (_10594_, _10502_, word_in[23]);
  nor (_10595_, _10506_, _08672_);
  and (_10596_, _10506_, word_in[7]);
  or (_10597_, _10596_, _10595_);
  and (_10598_, _10597_, _10511_);
  and (_10599_, _10503_, word_in[15]);
  or (_10600_, _10599_, _10598_);
  and (_10601_, _10600_, _10515_);
  or (_10602_, _10601_, _10594_);
  and (_10603_, _10602_, _10519_);
  and (_10604_, _10501_, word_in[31]);
  or (_14599_, _10604_, _10603_);
  and (_10605_, _10500_, _08655_);
  and (_10606_, _09693_, _08734_);
  and (_10607_, _09695_, _08623_);
  not (_10608_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_10609_, _10505_, _09699_);
  nor (_10610_, _10609_, _10608_);
  and (_10611_, _10609_, word_in[0]);
  or (_10612_, _10611_, _10610_);
  or (_10613_, _10612_, _10607_);
  not (_10614_, _10607_);
  or (_10615_, _10614_, word_in[8]);
  and (_10616_, _10615_, _10613_);
  or (_10617_, _10616_, _10606_);
  not (_10618_, _10606_);
  or (_10619_, _10618_, _09837_);
  and (_10620_, _10619_, _10617_);
  or (_10621_, _10620_, _10605_);
  not (_10622_, _10605_);
  or (_10623_, _10622_, word_in[24]);
  and (_14600_, _10623_, _10621_);
  not (_10624_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  nor (_10625_, _10609_, _10624_);
  and (_10626_, _10609_, _09722_);
  or (_10627_, _10626_, _10625_);
  or (_10628_, _10627_, _10607_);
  or (_10629_, _10614_, word_in[9]);
  and (_10630_, _10629_, _10628_);
  or (_10631_, _10630_, _10606_);
  or (_10632_, _10618_, _09565_);
  and (_10633_, _10632_, _10622_);
  and (_10634_, _10633_, _10631_);
  and (_10635_, _10605_, word_in[25]);
  or (_14601_, _10635_, _10634_);
  not (_10636_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  nor (_10637_, _10609_, _10636_);
  and (_10638_, _10609_, word_in[2]);
  or (_10639_, _10638_, _10637_);
  or (_10640_, _10639_, _10607_);
  or (_10641_, _10614_, word_in[10]);
  and (_10642_, _10641_, _10640_);
  or (_10643_, _10642_, _10606_);
  or (_10644_, _10618_, _10099_);
  and (_10645_, _10644_, _10643_);
  or (_10646_, _10645_, _10605_);
  or (_10647_, _10622_, word_in[26]);
  and (_14602_, _10647_, _10646_);
  or (_10648_, _10618_, _10116_);
  not (_10649_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  nor (_10650_, _10609_, _10649_);
  and (_10651_, _10609_, word_in[3]);
  or (_10652_, _10651_, _10650_);
  or (_10653_, _10652_, _10607_);
  or (_10654_, _10614_, word_in[11]);
  and (_10655_, _10654_, _10653_);
  or (_10656_, _10655_, _10606_);
  and (_10657_, _10656_, _10648_);
  or (_10658_, _10657_, _10605_);
  or (_10659_, _10622_, word_in[27]);
  and (_14603_, _10659_, _10658_);
  not (_10660_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  nor (_10661_, _10609_, _10660_);
  and (_10662_, _10609_, word_in[4]);
  or (_10663_, _10662_, _10661_);
  or (_10664_, _10663_, _10607_);
  or (_10665_, _10614_, word_in[12]);
  and (_10666_, _10665_, _10664_);
  or (_10667_, _10666_, _10606_);
  or (_10668_, _10618_, _10020_);
  and (_10669_, _10668_, _10622_);
  and (_10670_, _10669_, _10667_);
  and (_10671_, _10605_, word_in[28]);
  or (_14604_, _10671_, _10670_);
  not (_10672_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_10673_, _10609_, _10672_);
  and (_10674_, _10609_, _09777_);
  or (_10675_, _10674_, _10673_);
  or (_10676_, _10675_, _10607_);
  or (_10677_, _10614_, word_in[13]);
  and (_10678_, _10677_, _10676_);
  or (_10679_, _10678_, _10606_);
  or (_10680_, _10618_, _10149_);
  and (_10681_, _10680_, _10679_);
  or (_10682_, _10681_, _10605_);
  or (_10683_, _10622_, word_in[29]);
  and (_14605_, _10683_, _10682_);
  or (_10684_, _10618_, _10154_);
  not (_10685_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_10686_, _10609_, _10685_);
  and (_10687_, _10609_, word_in[6]);
  or (_10688_, _10687_, _10686_);
  or (_10689_, _10688_, _10607_);
  or (_10690_, _10614_, word_in[14]);
  and (_10691_, _10690_, _10689_);
  or (_10692_, _10691_, _10606_);
  and (_10693_, _10692_, _10684_);
  or (_10694_, _10693_, _10605_);
  or (_10695_, _10622_, word_in[30]);
  and (_14606_, _10695_, _10694_);
  nor (_10696_, _10609_, _08576_);
  and (_10697_, _10609_, word_in[7]);
  or (_10698_, _10697_, _10696_);
  or (_10699_, _10698_, _10607_);
  or (_10700_, _10614_, word_in[15]);
  and (_10701_, _10700_, _10699_);
  or (_10702_, _10701_, _10606_);
  or (_10703_, _10618_, _08886_);
  and (_10704_, _10703_, _10702_);
  or (_10705_, _10704_, _10605_);
  or (_10706_, _10622_, word_in[31]);
  and (_14607_, _10706_, _10705_);
  and (_10707_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  not (_10708_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  nor (_10709_, _07432_, _10708_);
  or (_10710_, _10709_, _10707_);
  and (_09561_, _10710_, _06444_);
  and (_10711_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  not (_10712_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  nor (_10713_, _07432_, _10712_);
  or (_10714_, _10713_, _10711_);
  and (_09566_, _10714_, _06444_);
  and (_10715_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [5]);
  not (_10716_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_10717_, _07432_, _10716_);
  or (_10718_, _10717_, _10715_);
  and (_09571_, _10718_, _06444_);
  nor (_10719_, _07230_, _06734_);
  and (_10720_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  and (_10721_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  nor (_10722_, _10721_, _10720_);
  and (_10723_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_10724_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  nor (_10725_, _10724_, _10723_);
  and (_10726_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  not (_10728_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  nor (_10729_, _07241_, _10728_);
  nor (_10730_, _10729_, _10726_);
  and (_10731_, _10730_, _10725_);
  and (_10732_, _10731_, _10722_);
  nor (_10733_, _10732_, _08374_);
  nor (_10734_, _10733_, _10719_);
  nor (_09590_, _10734_, rst);
  not (_10735_, _08425_);
  and (_10736_, _08472_, _08360_);
  and (_10737_, _10736_, _08457_);
  not (_10738_, _10737_);
  not (_10739_, _08472_);
  and (_10740_, _10739_, _08360_);
  not (_10741_, _08457_);
  and (_10742_, _10741_, _08441_);
  and (_10743_, _10742_, _10740_);
  nor (_10744_, _08472_, _08360_);
  and (_10745_, _08457_, _08441_);
  and (_10746_, _10745_, _10744_);
  nor (_10747_, _10746_, _10743_);
  and (_10748_, _10747_, _10738_);
  nor (_10749_, _10748_, _10735_);
  not (_10750_, _10749_);
  and (_10751_, _08408_, _08392_);
  nor (_10752_, _08425_, _07263_);
  and (_10753_, _10752_, _10751_);
  not (_10754_, _08392_);
  nor (_10755_, _08425_, _08408_);
  and (_10756_, _10755_, _10754_);
  nor (_10757_, _10756_, _10753_);
  nor (_10758_, _08457_, _08441_);
  and (_10759_, _10758_, _10744_);
  and (_10760_, _10754_, _07263_);
  and (_10761_, _10760_, _10755_);
  and (_10762_, _10745_, _10740_);
  and (_10763_, _10762_, _10761_);
  nor (_10764_, _10763_, _10759_);
  nor (_10765_, _10764_, _10757_);
  not (_10766_, _10765_);
  not (_10767_, _08408_);
  nor (_10768_, _08425_, _10767_);
  nor (_10769_, _08392_, _07263_);
  and (_10770_, _10769_, _10768_);
  nor (_10771_, _10739_, _08360_);
  nor (_10772_, _10758_, _10745_);
  and (_10773_, _10772_, _10771_);
  and (_10774_, _10773_, _10770_);
  and (_10775_, _10761_, _10743_);
  nor (_10776_, _10775_, _10774_);
  not (_10777_, _10761_);
  and (_10778_, _10758_, _10736_);
  nor (_10779_, _10778_, _10746_);
  nor (_10780_, _10779_, _10777_);
  and (_10781_, _10745_, _10736_);
  and (_10782_, _10769_, _10755_);
  and (_10783_, _10782_, _10781_);
  and (_10784_, _10771_, _10741_);
  and (_10785_, _10784_, _10753_);
  nor (_10786_, _10785_, _10783_);
  not (_10787_, _10786_);
  nor (_10788_, _10787_, _10780_);
  and (_10789_, _10788_, _10776_);
  and (_10790_, _10789_, _10766_);
  and (_10791_, _10790_, _10750_);
  and (_10792_, _10782_, _10746_);
  and (_10793_, _10771_, _10761_);
  nor (_10794_, _10793_, _10792_);
  and (_10795_, _10767_, _08392_);
  nor (_10796_, _08441_, _08425_);
  and (_10797_, _10796_, _10795_);
  and (_10798_, _10797_, _10736_);
  and (_10799_, _10771_, _08457_);
  and (_10800_, _10799_, _10782_);
  nor (_10801_, _10800_, _10798_);
  and (_10803_, _10801_, _10794_);
  and (_10804_, _10770_, _10781_);
  not (_10805_, _10778_);
  nor (_10806_, _10753_, _08425_);
  nor (_10807_, _10806_, _10805_);
  nor (_10808_, _10807_, _10804_);
  and (_10810_, _10808_, _10803_);
  not (_10811_, _10756_);
  not (_10812_, _08441_);
  and (_10813_, _10744_, _08457_);
  and (_10814_, _10813_, _10812_);
  and (_10815_, _10742_, _10736_);
  nor (_10816_, _10815_, _10814_);
  nor (_10817_, _10816_, _10811_);
  and (_10818_, _10744_, _10742_);
  and (_10819_, _10818_, _10770_);
  and (_10820_, _10771_, _10745_);
  and (_10821_, _10820_, _10770_);
  nor (_10822_, _10821_, _10819_);
  not (_10823_, _10822_);
  nor (_10824_, _10823_, _10817_);
  and (_10825_, _10824_, _10810_);
  and (_10826_, _10770_, _10759_);
  not (_10827_, _10826_);
  and (_10828_, _10768_, _10754_);
  not (_10829_, _10828_);
  nor (_10830_, _10778_, _07263_);
  nor (_10831_, _10830_, _10829_);
  not (_10832_, _10818_);
  nor (_10833_, _10832_, _10757_);
  nor (_10834_, _10833_, _10831_);
  and (_10835_, _10834_, _10827_);
  and (_10836_, _10740_, _08457_);
  and (_10837_, _10836_, _10812_);
  and (_10838_, _10837_, _10761_);
  and (_10839_, _08441_, _10735_);
  and (_10840_, _10839_, _10795_);
  nor (_10841_, _10813_, _10737_);
  not (_10842_, _10841_);
  and (_10843_, _10842_, _10840_);
  nor (_10844_, _10843_, _10838_);
  and (_10845_, _10758_, _10740_);
  and (_10846_, _10845_, _10761_);
  not (_10847_, _10846_);
  and (_10848_, _10761_, _10781_);
  and (_10849_, _08392_, _07263_);
  and (_10850_, _10849_, _10768_);
  and (_10851_, _10850_, _10818_);
  nor (_10852_, _10851_, _10848_);
  and (_10853_, _10852_, _10847_);
  and (_10854_, _10853_, _10844_);
  and (_10855_, _10854_, _10835_);
  and (_10856_, _10855_, _10825_);
  not (_10857_, _10753_);
  and (_10858_, _10737_, _10812_);
  not (_10859_, _10858_);
  not (_10860_, _10845_);
  nor (_10861_, _10815_, _10781_);
  and (_10862_, _10861_, _10860_);
  and (_10863_, _10862_, _10859_);
  and (_10864_, _10863_, _10747_);
  nor (_10865_, _10864_, _10857_);
  and (_10866_, _10850_, _10759_);
  and (_10867_, _10815_, _10770_);
  nor (_10868_, _10867_, _10866_);
  not (_10869_, _10770_);
  and (_10870_, _10740_, _10741_);
  nor (_10871_, _10858_, _10870_);
  nor (_10872_, _10871_, _10869_);
  not (_10873_, _10813_);
  and (_10874_, _10796_, _10751_);
  nor (_10875_, _10874_, _10770_);
  nor (_10876_, _10875_, _10873_);
  nor (_10877_, _10876_, _10872_);
  and (_10878_, _10877_, _10868_);
  not (_10879_, _10878_);
  nor (_10880_, _10879_, _10865_);
  and (_10881_, _10880_, _10856_);
  and (_10882_, _10881_, _10791_);
  or (_10883_, _10795_, _08425_);
  and (_10884_, _10883_, _10781_);
  or (_10885_, _10884_, _10821_);
  nand (_10886_, _10850_, _10814_);
  nand (_10887_, _10886_, _10852_);
  nor (_10888_, _10887_, _10885_);
  and (_10889_, _10888_, _10868_);
  nand (_10890_, _10889_, _10789_);
  or (_10891_, _10890_, _10882_);
  and (_10892_, _10891_, _07230_);
  nand (_10893_, _10892_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_10894_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , rst);
  or (_10895_, _10892_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  and (_10896_, _10895_, _10894_);
  and (_09594_, _10896_, _10893_);
  not (_10897_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_10898_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_10899_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  and (_10900_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_10901_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_10902_, _10901_, _10899_);
  and (_10903_, _10902_, _10900_);
  nor (_10904_, _10903_, _10899_);
  not (_10906_, _10904_);
  nor (_10907_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2], \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  nor (_10908_, _10907_, _10898_);
  and (_10909_, _10908_, _10906_);
  nor (_10910_, _10909_, _10898_);
  not (_10911_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  not (_10912_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_10913_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  and (_10914_, _10913_, _10912_);
  and (_10915_, _10914_, _10911_);
  and (_10916_, _10915_, _10910_);
  nor (_10917_, _10916_, _10897_);
  and (_10918_, _10916_, _10897_);
  nor (_10919_, _10918_, _10917_);
  not (_10920_, _10919_);
  and (_10921_, _10914_, _10910_);
  nor (_10923_, _10921_, _10911_);
  nor (_10924_, _10923_, _10916_);
  not (_10925_, _10924_);
  and (_10926_, _10913_, _10910_);
  nor (_10927_, _10926_, _10912_);
  nor (_10928_, _10927_, _10921_);
  not (_10929_, _10928_);
  nor (_10930_, _10910_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  and (_10931_, _10910_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_10932_, _10931_, _10930_);
  not (_10933_, _10932_);
  not (_10934_, _10882_);
  nor (_10935_, _10902_, _10900_);
  nor (_10936_, _10935_, _10903_);
  nand (_10937_, _10936_, _10934_);
  nor (_10938_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0], \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  nor (_10939_, _10938_, _10900_);
  and (_10940_, _10939_, _10891_);
  or (_10941_, _10936_, _10934_);
  and (_10942_, _10941_, _10937_);
  nand (_10943_, _10942_, _10940_);
  nand (_10944_, _10943_, _10937_);
  nor (_10945_, _10908_, _10906_);
  nor (_10946_, _10945_, _10909_);
  and (_10947_, _10946_, _10944_);
  and (_10948_, _10947_, _10933_);
  and (_10949_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3], \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_10950_, _10949_, _10913_);
  nand (_10951_, _10950_, _10930_);
  or (_10952_, _10950_, _10930_);
  and (_10953_, _10952_, _10951_);
  and (_10954_, _10953_, _10948_);
  and (_10955_, _10954_, _10929_);
  and (_10956_, _10955_, _10925_);
  and (_10957_, _10956_, _10920_);
  not (_10958_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_10959_, _10918_, _10958_);
  and (_10960_, _10915_, _10897_);
  and (_10961_, _10960_, _10958_);
  and (_10962_, _10961_, _10910_);
  or (_10963_, _10962_, _10959_);
  nand (_10964_, _10963_, _10957_);
  not (_10965_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_10966_, _10962_, _10965_);
  and (_10967_, _10962_, _10965_);
  nor (_10968_, _10967_, _10966_);
  and (_10969_, _10968_, _10964_);
  nor (_10970_, _10968_, _10964_);
  nor (_10971_, _10970_, _10969_);
  or (_10972_, _10971_, _08374_);
  or (_10973_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_10974_, _10973_, _10894_);
  and (_10975_, _10974_, _10972_);
  and (_10976_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _06444_);
  and (_10977_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_09598_, _10977_, _10975_);
  and (_10978_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  and (_10979_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  nor (_10980_, _10979_, _10978_);
  and (_10981_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_10982_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [1]);
  nor (_10983_, _10982_, _10981_);
  and (_10984_, _10983_, _10980_);
  and (_10985_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_10986_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  nor (_10987_, _10986_, _10985_);
  and (_10988_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  and (_10989_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [1]);
  nor (_10990_, _10989_, _10988_);
  and (_10991_, _10990_, _10987_);
  and (_10992_, _10991_, _10984_);
  nor (_10993_, _10992_, _07307_);
  and (_10994_, _07307_, _07070_);
  nor (_10995_, _10994_, _10993_);
  nor (_09610_, _10995_, rst);
  and (_10996_, _09828_, _08734_);
  and (_10997_, _09819_, _08623_);
  not (_10998_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_10999_, _09822_, _08538_);
  nor (_11000_, _10999_, _10998_);
  and (_11001_, _10999_, word_in[0]);
  or (_11002_, _11001_, _11000_);
  or (_11003_, _11002_, _10997_);
  not (_11004_, _10997_);
  or (_11005_, _11004_, word_in[8]);
  and (_11006_, _11005_, _11003_);
  or (_11007_, _11006_, _10996_);
  and (_11008_, _10500_, _08613_);
  not (_11009_, _11008_);
  not (_11010_, _10996_);
  or (_11011_, _11010_, _09837_);
  and (_11012_, _11011_, _11009_);
  and (_11013_, _11012_, _11007_);
  and (_11014_, _11008_, word_in[24]);
  or (_14555_, _11014_, _11013_);
  or (_11015_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [23]);
  not (_11016_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  nand (_11017_, _07432_, _11016_);
  and (_11018_, _11017_, _06444_);
  and (_09619_, _11018_, _11015_);
  not (_11019_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  nor (_11020_, _10999_, _11019_);
  and (_11021_, _10999_, word_in[1]);
  or (_11022_, _11021_, _11020_);
  or (_11023_, _11022_, _10997_);
  or (_11024_, _11004_, word_in[9]);
  and (_11025_, _11024_, _11023_);
  or (_11026_, _11025_, _10996_);
  or (_11027_, _11010_, _09565_);
  and (_11028_, _11027_, _11009_);
  and (_11029_, _11028_, _11026_);
  and (_11030_, _11008_, word_in[25]);
  or (_14556_, _11030_, _11029_);
  or (_11031_, _11010_, _10099_);
  not (_11032_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  nor (_11033_, _10999_, _11032_);
  and (_11034_, _10999_, word_in[2]);
  or (_11035_, _11034_, _11033_);
  or (_11036_, _11035_, _10997_);
  or (_11037_, _11004_, word_in[10]);
  and (_11038_, _11037_, _11036_);
  or (_11039_, _11038_, _10996_);
  and (_11040_, _11039_, _11031_);
  or (_11041_, _11040_, _11008_);
  or (_11042_, _11009_, word_in[26]);
  and (_14557_, _11042_, _11041_);
  or (_11043_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [4]);
  not (_11044_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  nand (_11045_, _07432_, _11044_);
  and (_11046_, _11045_, _06444_);
  and (_09624_, _11046_, _11043_);
  not (_11047_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  nor (_11048_, _10999_, _11047_);
  and (_11049_, _10999_, word_in[3]);
  or (_11050_, _11049_, _11048_);
  or (_11051_, _11050_, _10997_);
  or (_11052_, _11004_, word_in[11]);
  and (_11053_, _11052_, _11051_);
  or (_11054_, _11053_, _10996_);
  or (_11055_, _11010_, _10116_);
  and (_11056_, _11055_, _11009_);
  and (_11057_, _11056_, _11054_);
  and (_11058_, _11008_, word_in[27]);
  or (_14558_, _11058_, _11057_);
  not (_11059_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  nor (_11060_, _10999_, _11059_);
  and (_11061_, _10999_, word_in[4]);
  or (_11062_, _11061_, _11060_);
  or (_11063_, _11062_, _10997_);
  or (_11064_, _11004_, word_in[12]);
  and (_11065_, _11064_, _11063_);
  or (_11066_, _11065_, _10996_);
  or (_11067_, _11010_, _10020_);
  and (_11068_, _11067_, _11066_);
  or (_11069_, _11068_, _11008_);
  or (_11070_, _11009_, word_in[28]);
  and (_14559_, _11070_, _11069_);
  not (_11071_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  nor (_11072_, _10999_, _11071_);
  and (_11073_, _10999_, word_in[5]);
  or (_11074_, _11073_, _11072_);
  or (_11075_, _11074_, _10997_);
  or (_11076_, _11004_, word_in[13]);
  and (_11077_, _11076_, _11075_);
  or (_11078_, _11077_, _10996_);
  or (_11079_, _11010_, _10149_);
  and (_11080_, _11079_, _11078_);
  or (_11081_, _11080_, _11008_);
  or (_11082_, _11009_, word_in[29]);
  and (_14560_, _11082_, _11081_);
  or (_11083_, _11010_, _10154_);
  not (_11084_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  nor (_11085_, _10999_, _11084_);
  and (_11086_, _10999_, word_in[6]);
  or (_11087_, _11086_, _11085_);
  or (_11088_, _11087_, _10997_);
  or (_11089_, _11004_, word_in[14]);
  and (_11090_, _11089_, _11088_);
  or (_11091_, _11090_, _10996_);
  and (_11092_, _11091_, _11083_);
  or (_11093_, _11092_, _11008_);
  or (_11094_, _11009_, word_in[30]);
  and (_14561_, _11094_, _11093_);
  or (_11095_, _07757_, _07669_);
  not (_11096_, _07681_);
  and (_11097_, _08985_, _11096_);
  nand (_11098_, _11097_, _07684_);
  or (_11099_, _11097_, _07684_);
  nand (_11100_, _11099_, _11098_);
  nand (_11101_, _11100_, _07757_);
  nand (_11102_, _11101_, _11095_);
  nand (_11103_, _11102_, _07459_);
  and (_11104_, _07767_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_11105_, _11104_, _08994_);
  or (_11106_, _08994_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13]);
  nand (_11107_, _11106_, _11105_);
  nand (_11108_, _11107_, _07602_);
  nor (_11109_, _08109_, _06887_);
  nor (_11110_, _11109_, _06697_);
  and (_11111_, _11109_, _06697_);
  nor (_11112_, _11111_, _11110_);
  nor (_11113_, _11112_, _06891_);
  nor (_11114_, _06732_, _06638_);
  and (_11115_, _06904_, _06465_);
  nor (_11116_, _11115_, _11114_);
  and (_11117_, _06914_, _06640_);
  and (_11118_, _06918_, _06903_);
  nor (_11119_, _11118_, _11117_);
  and (_11120_, _11119_, _11116_);
  and (_11121_, _11120_, _06974_);
  not (_11122_, _11121_);
  nor (_11123_, _11122_, _11113_);
  and (_11124_, _11123_, _06967_);
  not (_11125_, _06709_);
  and (_11126_, _06842_, _11125_);
  nor (_11127_, _06842_, _11125_);
  nor (_11128_, _11127_, _11126_);
  and (_11129_, _11128_, _06680_);
  nor (_11130_, _06877_, _06709_);
  and (_11131_, _06877_, _06709_);
  or (_11132_, _11131_, _11130_);
  and (_11133_, _11132_, _06847_);
  nor (_11134_, _11133_, _11129_);
  and (_11135_, _11134_, _11124_);
  and (_11136_, _11135_, _11108_);
  nand (_11137_, _11136_, _11103_);
  nand (_11138_, _11137_, _07653_);
  nor (_11139_, _06933_, _06701_);
  nor (_11140_, _11139_, _06935_);
  nor (_11142_, _11140_, _08028_);
  and (_11143_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_11144_, _11143_, _07439_);
  nor (_11145_, _11144_, _11142_);
  nand (_11146_, _11145_, _11138_);
  and (_11147_, _06705_, _06640_);
  and (_11148_, _06913_, _06552_);
  nor (_11149_, _06740_, _06465_);
  nor (_11150_, _11149_, _09006_);
  and (_11151_, _11150_, _09173_);
  and (_11152_, _11151_, _06704_);
  nor (_11153_, _11151_, _06704_);
  nor (_11155_, _11153_, _11152_);
  nor (_11156_, _11155_, _06621_);
  nor (_11157_, _06704_, _06465_);
  or (_11158_, _11157_, _06892_);
  and (_11160_, _11158_, _06455_);
  or (_11161_, _11160_, _11156_);
  or (_11162_, _11161_, _11148_);
  and (_11163_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  nor (_11164_, \oc8051_top_1.oc8051_decoder1.src_sel3 , \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  not (_11165_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_11166_, \oc8051_top_1.oc8051_decoder1.src_sel3 , _11165_);
  nor (_11167_, _11166_, _11164_);
  nand (_11168_, _11167_, _09191_);
  or (_11169_, _11167_, _09191_);
  and (_11170_, _11169_, _06847_);
  and (_11171_, _11170_, _11168_);
  and (_11172_, _09416_, _07602_);
  or (_11173_, _11172_, _11171_);
  or (_11174_, _11173_, _11163_);
  or (_11175_, _11174_, _11162_);
  or (_11177_, _11175_, _11147_);
  or (_11178_, _11177_, _07961_);
  and (_11179_, _11178_, _11146_);
  and (_09630_, _11179_, _06444_);
  nor (_11180_, _10999_, _08667_);
  and (_11181_, _10999_, word_in[7]);
  or (_11182_, _11181_, _11180_);
  or (_11183_, _11182_, _10997_);
  or (_11184_, _11004_, word_in[15]);
  and (_11185_, _11184_, _11183_);
  or (_11186_, _11185_, _10996_);
  or (_11187_, _11010_, _08886_);
  and (_11188_, _11187_, _11009_);
  and (_11189_, _11188_, _11186_);
  and (_11190_, _11008_, word_in[31]);
  or (_14562_, _11190_, _11189_);
  and (_11191_, _07429_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  and (_11192_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_11193_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  not (_11194_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_11195_, _07241_, _11194_);
  nor (_11196_, _11195_, _11193_);
  and (_11197_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_11199_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_11200_, _11199_, _11197_);
  and (_11201_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  and (_11202_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_11203_, _11202_, _11201_);
  and (_11204_, _11203_, _11200_);
  and (_11205_, _11204_, _11196_);
  nor (_11206_, _11205_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_11207_, _11206_, _11192_);
  nor (_11208_, _11207_, _07429_);
  nor (_11209_, _11208_, _11191_);
  nor (_09668_, _11209_, rst);
  nor (_11210_, _07230_, _06790_);
  and (_11211_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  and (_11212_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_11213_, _11212_, _11211_);
  and (_11215_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_11216_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  nor (_11217_, _11216_, _11215_);
  and (_11218_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  not (_11220_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  nor (_11221_, _07241_, _11220_);
  nor (_11223_, _11221_, _11218_);
  and (_11224_, _11223_, _11217_);
  and (_11225_, _11224_, _11213_);
  nor (_11226_, _11225_, _08374_);
  nor (_11227_, _11226_, _11210_);
  nor (_09673_, _11227_, rst);
  and (_11228_, _09939_, _08734_);
  and (_11229_, _08870_, _08623_);
  not (_11230_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_11231_, _10505_, _08874_);
  nor (_11232_, _11231_, _11230_);
  and (_11233_, _11231_, word_in[0]);
  or (_11234_, _11233_, _11232_);
  or (_11235_, _11234_, _11229_);
  not (_11236_, _11229_);
  or (_11237_, _11236_, word_in[8]);
  and (_11238_, _11237_, _11235_);
  or (_11240_, _11238_, _11228_);
  and (_11241_, _10500_, _08611_);
  not (_11242_, _11241_);
  not (_11243_, _11228_);
  or (_11244_, _11243_, _09837_);
  and (_11245_, _11244_, _11242_);
  and (_11246_, _11245_, _11240_);
  and (_11247_, _11241_, _09554_);
  or (_14563_, _11247_, _11246_);
  not (_11249_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_11250_, _11231_, _11249_);
  and (_11251_, _11231_, _09722_);
  or (_11253_, _11251_, _11250_);
  or (_11254_, _11253_, _11229_);
  or (_11255_, _11236_, word_in[9]);
  and (_11256_, _11255_, _11254_);
  or (_11257_, _11256_, _11228_);
  or (_11258_, _11243_, _09565_);
  and (_11259_, _11258_, _11242_);
  and (_11260_, _11259_, _11257_);
  and (_11261_, _08855_, word_in[25]);
  and (_11262_, _11241_, _11261_);
  or (_14564_, _11262_, _11260_);
  and (_11263_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  not (_11264_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  nor (_11265_, _07432_, _11264_);
  or (_11266_, _11265_, _11263_);
  and (_09708_, _11266_, _06444_);
  not (_11267_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_11268_, _11231_, _11267_);
  and (_11269_, _11231_, word_in[2]);
  or (_11270_, _11269_, _11268_);
  or (_11271_, _11270_, _11229_);
  or (_11272_, _11236_, word_in[10]);
  and (_11273_, _11272_, _11271_);
  or (_11274_, _11273_, _11228_);
  or (_11275_, _11243_, _10099_);
  and (_11276_, _11275_, _11242_);
  and (_11277_, _11276_, _11274_);
  and (_11278_, _11241_, _09582_);
  or (_14565_, _11278_, _11277_);
  not (_11279_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_11280_, _11231_, _11279_);
  and (_11281_, _11231_, word_in[3]);
  or (_11282_, _11281_, _11280_);
  or (_11283_, _11282_, _11229_);
  or (_11284_, _11236_, word_in[11]);
  and (_11285_, _11284_, _11283_);
  or (_11286_, _11285_, _11228_);
  or (_11287_, _11243_, _10116_);
  and (_11288_, _11287_, _11286_);
  or (_11289_, _11288_, _11241_);
  or (_11290_, _11242_, word_in[27]);
  and (_14566_, _11290_, _11289_);
  and (_11291_, _11228_, _10020_);
  not (_11292_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_11293_, _11231_, _11292_);
  and (_11294_, _11231_, word_in[4]);
  nor (_11295_, _11294_, _11293_);
  nor (_11296_, _11295_, _11229_);
  and (_11297_, _11229_, word_in[12]);
  or (_11299_, _11297_, _11296_);
  and (_11300_, _11299_, _11243_);
  or (_11301_, _11300_, _11291_);
  and (_11302_, _11301_, _11242_);
  and (_11303_, _11241_, word_in[28]);
  or (_14567_, _11303_, _11302_);
  not (_11305_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  nor (_11306_, _11231_, _11305_);
  and (_11307_, _11231_, _09777_);
  or (_11309_, _11307_, _11306_);
  or (_11310_, _11309_, _11229_);
  or (_11311_, _11236_, word_in[13]);
  and (_11312_, _11311_, _11310_);
  or (_11313_, _11312_, _11228_);
  or (_11314_, _11243_, _10149_);
  and (_11315_, _11314_, _11242_);
  and (_11316_, _11315_, _11313_);
  and (_11317_, _11241_, _09623_);
  or (_14568_, _11317_, _11316_);
  not (_11318_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  nor (_11319_, _11231_, _11318_);
  and (_11320_, _11231_, word_in[6]);
  or (_11321_, _11320_, _11319_);
  or (_11322_, _11321_, _11229_);
  or (_11323_, _11236_, word_in[14]);
  and (_11324_, _11323_, _11322_);
  or (_11325_, _11324_, _11228_);
  or (_11326_, _11243_, _10154_);
  and (_11327_, _11326_, _11242_);
  and (_11328_, _11327_, _11325_);
  and (_11329_, _11241_, _09626_);
  or (_14569_, _11329_, _11328_);
  nor (_11330_, _11231_, _08565_);
  and (_11331_, _11231_, word_in[7]);
  or (_11332_, _11331_, _11330_);
  or (_11333_, _11332_, _11229_);
  or (_11334_, _11236_, word_in[15]);
  and (_11335_, _11334_, _11333_);
  or (_11336_, _11335_, _11228_);
  or (_11337_, _11243_, _08886_);
  and (_11338_, _11337_, _11336_);
  or (_11339_, _11338_, _11241_);
  or (_11340_, _11242_, word_in[31]);
  and (_14570_, _11340_, _11339_);
  and (_11341_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_11342_, _07229_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_11343_, _11342_);
  or (_11344_, _08441_, _07232_);
  nor (_11345_, _07230_, \oc8051_top_1.oc8051_decoder1.op [4]);
  nor (_11346_, _11345_, _07265_);
  and (_11347_, _11346_, _11344_);
  not (_11348_, _09327_);
  or (_11349_, _08425_, _07232_);
  nor (_11350_, _07230_, \oc8051_top_1.oc8051_decoder1.op [3]);
  nor (_11351_, _11350_, _07265_);
  nand (_11352_, _11351_, _11349_);
  and (_11353_, _11352_, _11348_);
  and (_11354_, _11353_, _09477_);
  and (_11355_, _11354_, _07268_);
  and (_11356_, _11355_, _11347_);
  or (_11357_, _08457_, _07232_);
  nor (_11358_, _07230_, \oc8051_top_1.oc8051_decoder1.op [5]);
  nor (_11359_, _11358_, _07265_);
  nand (_11360_, _11359_, _11357_);
  or (_11361_, _08360_, _07232_);
  nor (_11362_, _07230_, \oc8051_top_1.oc8051_decoder1.op [7]);
  nor (_11363_, _11362_, _07265_);
  nand (_11364_, _11363_, _11361_);
  nand (_11365_, _08472_, _07231_);
  nor (_11366_, _07230_, \oc8051_top_1.oc8051_decoder1.op [6]);
  nor (_11367_, _11366_, _07265_);
  and (_11368_, _11367_, _11365_);
  nor (_11369_, _11368_, _11364_);
  and (_11370_, _11369_, _11360_);
  and (_11371_, _11370_, _11356_);
  and (_11372_, _11359_, _11357_);
  and (_11373_, _11368_, _11364_);
  and (_11374_, _11373_, _11372_);
  and (_11375_, _11356_, _11374_);
  not (_11376_, _11347_);
  and (_11377_, _11369_, _11372_);
  and (_11378_, _11377_, _11376_);
  and (_11379_, _11378_, _11355_);
  nor (_11380_, _11379_, _11375_);
  not (_11381_, _11380_);
  nor (_11382_, _11381_, _11371_);
  nor (_11383_, _11382_, _11343_);
  nor (_11384_, _09477_, _07268_);
  and (_11385_, _11384_, _11353_);
  not (_11386_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_11387_, \oc8051_top_1.oc8051_decoder1.state [1], _06308_);
  and (_11389_, _11387_, _11386_);
  and (_11390_, _11373_, _11389_);
  and (_11391_, _11390_, _11385_);
  not (_11392_, _11391_);
  and (_11393_, _11352_, _09327_);
  and (_11394_, _11384_, _11393_);
  and (_11395_, _11370_, _11376_);
  and (_11396_, _11395_, _11394_);
  and (_11398_, _11378_, _11394_);
  nor (_11399_, _11398_, _11396_);
  and (_11400_, _11399_, _11392_);
  not (_11401_, _11400_);
  nor (_11402_, _11401_, _11383_);
  nor (_11403_, _11402_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11404_, _11403_, _11341_);
  and (_11405_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11406_, _11393_, _09477_);
  and (_11407_, _11373_, _11360_);
  and (_11408_, _11407_, _11376_);
  and (_11409_, _11408_, _11406_);
  not (_11410_, _11364_);
  and (_11411_, _11360_, _11368_);
  and (_11412_, _11411_, _11410_);
  and (_11413_, _11385_, _11412_);
  and (_11414_, _11413_, _11347_);
  nor (_11415_, _11414_, _11409_);
  nand (_11416_, _11395_, _11406_);
  and (_11417_, _11372_, _11368_);
  and (_11418_, _11417_, _11410_);
  and (_11419_, _11418_, _11376_);
  nand (_11420_, _11419_, _11406_);
  and (_11421_, _11420_, _11416_);
  and (_11422_, _11421_, _11415_);
  and (_11423_, _11406_, _11347_);
  and (_11424_, _11423_, _11377_);
  not (_11425_, _11368_);
  and (_11426_, _11425_, _11364_);
  and (_11427_, _11426_, _11360_);
  and (_11428_, _11406_, _11427_);
  nor (_11429_, _11428_, _11424_);
  and (_11430_, _11354_, _07311_);
  and (_11431_, _11426_, _11372_);
  and (_11432_, _11431_, _11430_);
  and (_11433_, _11376_, _11374_);
  and (_11434_, _11433_, _11406_);
  nor (_11435_, _11434_, _11432_);
  and (_11436_, _11435_, _11429_);
  and (_11437_, _11407_, _11347_);
  and (_11438_, _11437_, _11406_);
  and (_11439_, _11406_, _11431_);
  or (_11440_, _11439_, _11438_);
  not (_11441_, _11440_);
  and (_11442_, _11406_, _11412_);
  and (_11443_, _11370_, _11347_);
  and (_11444_, _11443_, _11406_);
  nor (_11445_, _11444_, _11442_);
  and (_11446_, _11445_, _11441_);
  and (_11447_, _11446_, _11436_);
  and (_11448_, _11447_, _11422_);
  and (_11449_, _11448_, _11382_);
  nor (_11450_, _11449_, _11343_);
  and (_11451_, _11387_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_11452_, _11432_, _11451_);
  and (_11453_, _06308_, \oc8051_top_1.oc8051_decoder1.state [0]);
  and (_11454_, _11385_, _11431_);
  and (_11455_, _11454_, _11376_);
  and (_11456_, _11431_, _11347_);
  and (_11457_, _11456_, _11385_);
  and (_11458_, _11427_, _11347_);
  and (_11459_, _11385_, _11458_);
  or (_11460_, _11459_, _11457_);
  nor (_11461_, _11460_, _11455_);
  and (_11463_, _11391_, _11360_);
  not (_11464_, _11463_);
  and (_11465_, _11464_, _11461_);
  nor (_11466_, _11465_, _11453_);
  nor (_11467_, _11466_, _11392_);
  nor (_11468_, _11467_, _11452_);
  not (_11469_, _11468_);
  nor (_11470_, _11469_, _11450_);
  nor (_11471_, _11470_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11472_, _11471_, _11405_);
  not (_11473_, _11472_);
  and (_11474_, \oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_11475_, _11347_, _11374_);
  and (_11476_, _11475_, _11430_);
  and (_11477_, _11408_, _11354_);
  nor (_11478_, _11477_, _11476_);
  and (_11479_, _11378_, _11385_);
  not (_11480_, _09477_);
  and (_11481_, _11480_, _07268_);
  and (_11482_, _11393_, _11481_);
  and (_11483_, _11408_, _11482_);
  nor (_11484_, _11483_, _11479_);
  and (_11485_, _11484_, _11478_);
  and (_11486_, _11377_, _11347_);
  and (_11487_, _11385_, _11486_);
  not (_11488_, _11487_);
  and (_11489_, _11486_, _11430_);
  and (_11490_, _11412_, _11376_);
  and (_11491_, _11490_, _11430_);
  nor (_11492_, _11491_, _11489_);
  and (_11493_, _11412_, _11347_);
  and (_11494_, _11482_, _11493_);
  and (_11495_, _11482_, _11458_);
  nor (_11496_, _11495_, _11494_);
  and (_11497_, _11496_, _11492_);
  and (_11498_, _11497_, _11488_);
  and (_11499_, _11498_, _11485_);
  not (_11500_, _11482_);
  nor (_11501_, _11443_, _11486_);
  or (_11502_, _11501_, _11500_);
  and (_11503_, _11433_, _11482_);
  and (_11504_, _11490_, _11482_);
  nor (_11505_, _11504_, _11503_);
  not (_11507_, _11505_);
  or (_11508_, _11443_, _11493_);
  and (_11509_, _11508_, _11430_);
  nor (_11510_, _11509_, _11507_);
  and (_11511_, _11510_, _11502_);
  and (_11512_, _11395_, _11430_);
  and (_11513_, _11437_, _11354_);
  nor (_11514_, _11513_, _11512_);
  not (_11515_, _11514_);
  nor (_11516_, _11437_, _11431_);
  nor (_11517_, _11516_, _11500_);
  nor (_11518_, _11517_, _11515_);
  nor (_11519_, _11352_, _11347_);
  and (_11520_, _11519_, _11377_);
  or (_11521_, _11520_, _11413_);
  nor (_11522_, _11521_, _11432_);
  and (_11523_, _11427_, _11376_);
  and (_11524_, _11482_, _11523_);
  and (_11525_, _09477_, _09327_);
  not (_11526_, _11352_);
  nor (_11527_, _11526_, _11347_);
  and (_11528_, _11527_, _11525_);
  and (_11529_, _11528_, _11377_);
  nor (_11530_, _11529_, _11524_);
  and (_11531_, _11530_, _11522_);
  and (_11532_, _11531_, _11518_);
  and (_11533_, _11378_, _11430_);
  and (_11534_, _11395_, _11482_);
  nor (_11535_, _11534_, _11533_);
  and (_11536_, _11433_, _11354_);
  and (_11537_, _11419_, _11482_);
  nor (_11538_, _11537_, _11536_);
  and (_11539_, _11538_, _11535_);
  and (_11540_, _11539_, _11461_);
  and (_11541_, _11540_, _11532_);
  and (_11542_, _11541_, _11511_);
  and (_11543_, _11542_, _11499_);
  nor (_11544_, _11543_, _11343_);
  nor (_11545_, _11391_, _11452_);
  not (_11546_, _11545_);
  nor (_11547_, _11546_, _11544_);
  nor (_11548_, _11547_, \oc8051_top_1.oc8051_sfr1.wait_data );
  nor (_11549_, _11548_, _11474_);
  and (_11550_, _11549_, _11473_);
  and (_11551_, _11550_, _11404_);
  and (_11552_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_11553_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  nor (_11554_, _11553_, _11552_);
  and (_11555_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_11556_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  nor (_11557_, _11556_, _11555_);
  and (_11558_, _11557_, _11554_);
  and (_11559_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  and (_11560_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor (_11561_, _11560_, _11559_);
  and (_11562_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  and (_11563_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  nor (_11564_, _11563_, _11562_);
  and (_11565_, _11564_, _11561_);
  and (_11566_, _11565_, _11558_);
  nor (_11567_, _11566_, _07307_);
  not (_11568_, _06978_);
  and (_11569_, _07307_, _11568_);
  nor (_11570_, _11569_, _11567_);
  not (_11571_, _11570_);
  and (_11572_, _11571_, _11551_);
  not (_11573_, _11572_);
  not (_11574_, _11549_);
  not (_11575_, _11404_);
  nor (_11576_, _11472_, _11575_);
  and (_11577_, _11576_, _11574_);
  and (_11578_, _08978_, _06432_);
  and (_11579_, _11578_, _06978_);
  not (_11580_, _11578_);
  and (_11581_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3]);
  nor (_11582_, _11580_, _07300_);
  nor (_11583_, _11582_, _11581_);
  and (_11584_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2]);
  nor (_11585_, _06644_, _06604_);
  not (_11586_, _11585_);
  and (_11587_, _11586_, _09124_);
  and (_11588_, _11587_, _09121_);
  and (_11589_, _11588_, _09114_);
  nor (_11590_, _11589_, _11580_);
  nor (_11591_, _11590_, _11584_);
  and (_11592_, _11578_, _07070_);
  and (_11593_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1]);
  nor (_11594_, _11593_, _11592_);
  nor (_11595_, _11578_, _06401_);
  and (_11596_, _11578_, _09527_);
  nor (_11597_, _11596_, _11595_);
  and (_11598_, _11597_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  and (_11599_, _11598_, _11594_);
  and (_11600_, _11599_, _11591_);
  and (_11601_, _11600_, _11583_);
  nor (_11602_, _11580_, _07188_);
  and (_11603_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4]);
  nor (_11604_, _11603_, _11602_);
  and (_11605_, _11604_, _11601_);
  nor (_11606_, _11580_, _06666_);
  and (_11607_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5]);
  nor (_11608_, _11607_, _11606_);
  and (_11609_, _11608_, _11605_);
  nor (_11610_, _11580_, _10494_);
  and (_11611_, _11580_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6]);
  nor (_11612_, _11611_, _11610_);
  and (_11613_, _11612_, _11609_);
  nor (_11614_, _11578_, _06366_);
  nor (_11615_, _11614_, _11613_);
  and (_11616_, _11614_, _11613_);
  or (_11617_, _11616_, _11615_);
  nor (_11618_, _11617_, _06311_);
  nor (_11619_, _11578_, _06370_);
  not (_11620_, _11619_);
  nor (_11621_, _11620_, _11618_);
  nor (_11622_, _11621_, _11579_);
  and (_11623_, _11622_, _11577_);
  not (_11624_, _11623_);
  not (_11625_, _08376_);
  nor (_11626_, _11549_, _11473_);
  and (_11627_, _11626_, _11625_);
  nor (_11628_, _11627_, _11575_);
  and (_11629_, _11628_, _11624_);
  and (_11630_, _11629_, _11573_);
  nor (_11631_, _11630_, _08030_);
  and (_11632_, _11630_, _08030_);
  nor (_11633_, _11632_, _11631_);
  and (_11634_, _11472_, _11404_);
  and (_11635_, _11634_, _11574_);
  nor (_11636_, _07230_, _06747_);
  and (_11637_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  and (_11638_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  nor (_11639_, _11638_, _11637_);
  and (_11640_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_11641_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  nor (_11642_, _11641_, _11640_);
  and (_11643_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_11644_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  nor (_11645_, _11644_, _11643_);
  and (_11646_, _11645_, _11642_);
  and (_11647_, _11646_, _11639_);
  nor (_11648_, _11647_, _08374_);
  nor (_11649_, _11648_, _11636_);
  not (_11650_, _11649_);
  and (_11651_, _11650_, _11635_);
  and (_11652_, _11634_, _11549_);
  and (_11653_, _11652_, _07316_);
  nor (_11654_, _11653_, _11651_);
  not (_11655_, _07361_);
  and (_11656_, _11551_, _11655_);
  not (_11657_, _11656_);
  nor (_11658_, _11604_, _11601_);
  nor (_11659_, _11658_, _11605_);
  nor (_11660_, _11659_, _06311_);
  nor (_11661_, _11660_, _06315_);
  nor (_11662_, _11661_, _11578_);
  nor (_11663_, _11662_, _11602_);
  not (_11664_, _11663_);
  and (_11665_, _11664_, _11577_);
  and (_11666_, _11472_, _11575_);
  nor (_11667_, _11666_, _11665_);
  and (_11668_, _11667_, _11657_);
  and (_11669_, _11668_, _11654_);
  nor (_11670_, _11669_, _06337_);
  and (_11671_, _11669_, _06337_);
  nor (_11672_, _11671_, _11670_);
  not (_11673_, _07342_);
  and (_11674_, _11551_, _11673_);
  nor (_11675_, _07230_, _06770_);
  and (_11676_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  and (_11677_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_11678_, _11677_, _11676_);
  and (_11679_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_11680_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_11681_, _11680_, _11679_);
  and (_11682_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  and (_11683_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_11684_, _11683_, _11682_);
  and (_11685_, _11684_, _11681_);
  and (_11686_, _11685_, _11678_);
  nor (_11687_, _11686_, _08374_);
  nor (_11688_, _11687_, _11675_);
  not (_11689_, _11688_);
  and (_11690_, _11689_, _11635_);
  nor (_11691_, _11690_, _11674_);
  not (_11692_, _07302_);
  and (_11693_, _11652_, _11692_);
  nor (_11694_, _11600_, _11583_);
  nor (_11695_, _11694_, _11601_);
  nor (_11696_, _11695_, _06311_);
  nor (_11697_, _11696_, _06388_);
  nor (_11698_, _11697_, _11578_);
  nor (_11699_, _11698_, _11582_);
  not (_11700_, _11699_);
  and (_11701_, _11700_, _11577_);
  nor (_11702_, _11701_, _11693_);
  and (_11703_, _11702_, _11691_);
  nor (_11704_, _11703_, _06395_);
  and (_11705_, _11703_, _06395_);
  nor (_11706_, _11705_, _11704_);
  and (_11707_, _11706_, _11672_);
  not (_11708_, _07380_);
  and (_11709_, _11551_, _11708_);
  nor (_11710_, _07230_, _06474_);
  and (_11711_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  and (_11712_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_11713_, _11712_, _11711_);
  and (_11714_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_11715_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  nor (_11716_, _11715_, _11714_);
  and (_11717_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  not (_11718_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_11719_, _07241_, _11718_);
  nor (_11720_, _11719_, _11717_);
  and (_11721_, _11720_, _11716_);
  and (_11723_, _11721_, _11713_);
  nor (_11724_, _11723_, _08374_);
  nor (_11725_, _11724_, _11710_);
  not (_11726_, _11725_);
  and (_11727_, _11726_, _11635_);
  nor (_11728_, _11727_, _11709_);
  nor (_11729_, _11608_, _11605_);
  nor (_11730_, _11729_, _11609_);
  nor (_11731_, _11730_, _06311_);
  nor (_11732_, _11731_, _06342_);
  nor (_11733_, _11732_, _11578_);
  nor (_11734_, _11733_, _11606_);
  nor (_11735_, _11734_, _11472_);
  nor (_11736_, _11735_, _11575_);
  not (_11737_, _11736_);
  nor (_11738_, _11626_, _11550_);
  and (_11739_, _11738_, _11737_);
  not (_11740_, _11739_);
  and (_11741_, _11740_, _11728_);
  and (_11742_, _11741_, _06671_);
  nor (_11743_, _11741_, _06671_);
  nor (_11744_, _11743_, _11742_);
  and (_11745_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  and (_11746_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor (_11747_, _11746_, _11745_);
  and (_11749_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_11750_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  nor (_11751_, _11750_, _11749_);
  and (_11753_, _11751_, _11747_);
  and (_11754_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_11755_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  nor (_11756_, _11755_, _11754_);
  and (_11757_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [6]);
  and (_11758_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_11759_, _11758_, _11757_);
  and (_11760_, _11759_, _11756_);
  and (_11761_, _11760_, _11753_);
  nor (_11762_, _11761_, _07307_);
  not (_11763_, _10494_);
  and (_11764_, _11763_, _07307_);
  nor (_11765_, _11764_, _11762_);
  not (_11766_, _11765_);
  and (_11767_, _11766_, _11551_);
  nor (_11769_, _11612_, _11609_);
  nor (_11770_, _11769_, _11613_);
  nor (_11771_, _11770_, _06311_);
  nor (_11772_, _11771_, _06356_);
  nor (_11773_, _11772_, _11578_);
  nor (_11774_, _11773_, _11610_);
  not (_11775_, _11774_);
  and (_11776_, _11775_, _11577_);
  nor (_11777_, _11776_, _11767_);
  not (_11778_, _10734_);
  and (_11779_, _11635_, _11778_);
  nor (_11780_, _11550_, _11404_);
  nor (_11781_, _11780_, _11779_);
  and (_11782_, _11781_, _11777_);
  and (_11784_, _11782_, _06365_);
  nor (_11785_, _11782_, _06365_);
  nor (_11786_, _11785_, _11784_);
  and (_11787_, _11786_, _11744_);
  and (_11788_, _11787_, _11707_);
  and (_11789_, _11788_, _11633_);
  not (_11790_, _10995_);
  and (_11791_, _11551_, _11790_);
  not (_11792_, _11791_);
  and (_11793_, _11550_, _11575_);
  not (_11794_, _11227_);
  and (_11795_, _11635_, _11794_);
  nor (_11796_, _11795_, _11793_);
  nor (_11797_, _11598_, _11594_);
  nor (_11798_, _11797_, _11599_);
  nor (_11799_, _11798_, _06311_);
  nor (_11800_, _11799_, _06410_);
  nor (_11801_, _11800_, _11578_);
  nor (_11802_, _11801_, _11592_);
  not (_11803_, _11802_);
  and (_11804_, _11803_, _11577_);
  and (_11805_, _11652_, _09477_);
  nor (_11807_, _11805_, _11804_);
  and (_11808_, _11807_, _11796_);
  and (_11809_, _11808_, _11792_);
  nor (_11810_, _11809_, _06418_);
  and (_11811_, _11809_, _06418_);
  nor (_11812_, _11811_, _11810_);
  and (_11813_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_11814_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nor (_11815_, _11814_, _11813_);
  and (_11816_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_11817_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [0]);
  nor (_11818_, _11817_, _11816_);
  and (_11819_, _11818_, _11815_);
  and (_11820_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  and (_11821_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  nor (_11822_, _11821_, _11820_);
  and (_11823_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_11824_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  nor (_11825_, _11824_, _11823_);
  and (_11826_, _11825_, _11822_);
  and (_11827_, _11826_, _11819_);
  nor (_11828_, _11827_, _07307_);
  and (_11829_, _09527_, _07307_);
  nor (_11830_, _11829_, _11828_);
  not (_11831_, _11830_);
  and (_11832_, _11831_, _11551_);
  nor (_11833_, _07230_, _06801_);
  and (_11834_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  and (_11835_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [24]);
  nor (_11836_, _11835_, _11834_);
  and (_11837_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  not (_11838_, \oc8051_top_1.oc8051_memory_interface1.idat_old [16]);
  nor (_11839_, _07241_, _11838_);
  nor (_11840_, _11839_, _11837_);
  and (_11841_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  and (_11842_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nor (_11843_, _11842_, _11841_);
  and (_11844_, _11843_, _11840_);
  and (_11845_, _11844_, _11836_);
  nor (_11846_, _11845_, _08374_);
  nor (_11847_, _11846_, _11833_);
  not (_11848_, _11847_);
  and (_11849_, _11848_, _11635_);
  nor (_11850_, _11849_, _11832_);
  and (_11851_, _11652_, _07268_);
  nor (_11852_, _11597_, \oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop );
  nor (_11853_, _11852_, _11598_);
  nor (_11854_, _11853_, _06311_);
  nor (_11855_, _11854_, _06402_);
  nor (_11856_, _11855_, _11578_);
  nor (_11857_, _11856_, _11596_);
  not (_11858_, _11857_);
  and (_11859_, _11858_, _11577_);
  nor (_11860_, _11859_, _11851_);
  and (_11861_, _11860_, _11850_);
  and (_11862_, _11861_, _06407_);
  nor (_11863_, _11861_, _06407_);
  or (_11864_, _11863_, _11862_);
  nor (_11865_, _11864_, _11812_);
  and (_11866_, _07321_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  and (_11867_, _07327_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  nor (_11868_, _11867_, _11866_);
  and (_11869_, _07313_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_11870_, _07331_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_11871_, _11870_, _11869_);
  and (_11872_, _11871_, _11868_);
  and (_11873_, _07318_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  and (_11874_, _07333_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  nor (_11875_, _11874_, _11873_);
  and (_11876_, _07309_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  and (_11877_, _07325_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  nor (_11878_, _11877_, _11876_);
  and (_11879_, _11878_, _11875_);
  and (_11880_, _11879_, _11872_);
  nor (_11881_, _11880_, _07307_);
  not (_11882_, _11589_);
  and (_11883_, _11882_, _07307_);
  nor (_11884_, _11883_, _11881_);
  not (_11885_, _11884_);
  and (_11886_, _11885_, _11551_);
  not (_11887_, _11886_);
  and (_11888_, _11652_, _09327_);
  nor (_11889_, _07230_, _06780_);
  and (_11890_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  and (_11891_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_old [26]);
  nor (_11892_, _11891_, _11890_);
  and (_11893_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [18]);
  and (_11895_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  nor (_11896_, _11895_, _11893_);
  and (_11897_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  and (_11899_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [18]);
  nor (_11900_, _11899_, _11897_);
  and (_11901_, _11900_, _11896_);
  and (_11902_, _11901_, _11892_);
  nor (_11903_, _11902_, _08374_);
  nor (_11904_, _11903_, _11889_);
  not (_11905_, _11904_);
  and (_11906_, _11905_, _11635_);
  nor (_11907_, _11599_, _11591_);
  nor (_11908_, _11907_, _11600_);
  nor (_11909_, _11908_, _06311_);
  nor (_11910_, _11909_, _06421_);
  nor (_11911_, _11910_, _11578_);
  nor (_11912_, _11911_, _11590_);
  not (_11914_, _11912_);
  and (_11915_, _11914_, _11577_);
  or (_11917_, _11915_, _11906_);
  nor (_11918_, _11917_, _11888_);
  and (_11919_, _11918_, _11887_);
  nor (_11920_, _11919_, _06430_);
  and (_11921_, _11919_, _06430_);
  nor (_11922_, _11921_, _11920_);
  nor (_11923_, _11922_, _08925_);
  and (_11924_, _11923_, _11865_);
  and (_11925_, _11924_, _11789_);
  nor (_11926_, _06380_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_11927_, _11926_, _11925_);
  not (_11928_, _11927_);
  and (_11929_, _11466_, _11392_);
  nor (_11930_, _06933_, _06943_);
  and (_11931_, _11930_, _11789_);
  and (_11932_, _11931_, _11929_);
  and (_11933_, _11481_, _11353_);
  and (_11934_, _11427_, _11430_);
  nor (_11935_, _11934_, _11933_);
  nor (_11936_, _11935_, _11343_);
  not (_11937_, _11128_);
  not (_11938_, _11466_);
  nor (_11939_, _06822_, _06763_);
  and (_11940_, _11939_, _07991_);
  and (_11941_, _11940_, _09098_);
  and (_11942_, _11941_, _11392_);
  and (_11943_, _11942_, _08287_);
  not (_11944_, _11943_);
  nor (_11945_, _11944_, _08209_);
  and (_11946_, _11945_, _11938_);
  and (_11947_, _11946_, _08999_);
  and (_11948_, _11947_, _11937_);
  nor (_11949_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  nor (_11950_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_11951_, _11950_, _11949_);
  nor (_11952_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  nor (_11953_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_11954_, _11953_, _11952_);
  and (_11955_, _11954_, _11951_);
  and (_11957_, _11955_, _11467_);
  not (_11958_, _11957_);
  and (_11959_, _11929_, _06463_);
  and (_11960_, _11463_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_11961_, _11960_, _11959_);
  and (_11962_, _11961_, _11958_);
  not (_11963_, _11962_);
  nor (_11964_, _11963_, _11948_);
  and (_11965_, _11393_, _11480_);
  and (_11966_, _11965_, _11486_);
  nor (_11967_, _11966_, _11494_);
  and (_11968_, _11493_, _11526_);
  not (_11969_, _11968_);
  and (_11970_, _11969_, _11967_);
  not (_11971_, _11385_);
  nor (_11972_, _11437_, _11475_);
  nor (_11973_, _11972_, _11971_);
  not (_11974_, _11973_);
  not (_11975_, _11457_);
  and (_11976_, _11526_, _11347_);
  and (_11977_, _11976_, _11377_);
  nor (_11978_, _11977_, _11424_);
  and (_11979_, _11978_, _11975_);
  and (_11980_, _11979_, _11974_);
  and (_11981_, _11980_, _11970_);
  not (_11982_, _11981_);
  and (_11983_, _11982_, _11964_);
  not (_11984_, _11432_);
  and (_11986_, _11395_, _11385_);
  nor (_11987_, _11986_, _11375_);
  nand (_11989_, _11987_, _11984_);
  nor (_11990_, _11989_, _11983_);
  and (_11991_, _11431_, _11376_);
  and (_11993_, _11991_, _11385_);
  nor (_11994_, _11993_, _11459_);
  nand (_11995_, _11376_, _11373_);
  nor (_11996_, _11995_, _11971_);
  not (_11997_, _11996_);
  and (_11998_, _11997_, _11994_);
  nor (_11999_, _11998_, _11964_);
  not (_12001_, _11999_);
  and (_12002_, _12001_, _11990_);
  nor (_12003_, _11452_, _11389_);
  nor (_12004_, _12003_, _12002_);
  nor (_12005_, _12004_, _11936_);
  nor (_12006_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  not (_12008_, _12006_);
  nor (_12009_, _12008_, _07218_);
  nor (_12011_, _06395_, _06336_);
  and (_12012_, _12011_, _06677_);
  not (_12013_, _12012_);
  and (_12014_, _12013_, _12009_);
  nor (_12015_, _12014_, _11464_);
  not (_12016_, _08036_);
  and (_12017_, _11467_, _12016_);
  nor (_12018_, _12017_, _12015_);
  not (_12019_, _12018_);
  nor (_12020_, _12019_, _12005_);
  not (_12021_, _12020_);
  nor (_12022_, _12021_, _11932_);
  and (_12023_, _12022_, _11928_);
  not (_12024_, _09045_);
  and (_12025_, _11475_, _11355_);
  and (_12026_, _12025_, _11389_);
  nor (_12028_, _12026_, _11936_);
  and (_12029_, _11978_, _11461_);
  nand (_12030_, _12029_, _11967_);
  nand (_12031_, _12030_, _11389_);
  and (_12032_, _11934_, _11342_);
  not (_12033_, _12032_);
  and (_12034_, _11454_, _11342_);
  nor (_12035_, _12034_, _11452_);
  and (_12037_, _12035_, _12033_);
  nand (_12038_, _12037_, _12031_);
  not (_12039_, _11389_);
  and (_12040_, _11385_, _11373_);
  not (_12041_, _12040_);
  and (_12042_, _11970_, _12041_);
  and (_12043_, _12042_, _11987_);
  and (_12044_, _12043_, _12029_);
  nor (_12045_, _12044_, _12039_);
  nor (_12046_, _12045_, _12038_);
  and (_12047_, _12046_, _12028_);
  or (_12048_, _12047_, _12026_);
  and (_12050_, _12048_, _12024_);
  and (_12051_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  or (_12052_, _12038_, _12028_);
  nor (_12054_, _12052_, _12045_);
  and (_12055_, _12054_, _11778_);
  and (_12056_, _07429_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  or (_12058_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _07234_);
  and (_12059_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_12060_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [30]);
  or (_12061_, _12060_, _12059_);
  and (_12062_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [22]);
  and (_12063_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  and (_12064_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  or (_12065_, _12064_, _12063_);
  or (_12066_, _12065_, _12062_);
  or (_12067_, _12066_, _12061_);
  and (_12068_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [30]);
  or (_12069_, _12068_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_12070_, _12069_, _12067_);
  and (_12071_, _12070_, _07230_);
  and (_12072_, _12071_, _12058_);
  nor (_12073_, _12072_, _12056_);
  not (_12074_, _12073_);
  and (_12075_, _12074_, _12032_);
  or (_12076_, _12075_, _12055_);
  or (_12077_, _12076_, _12051_);
  not (_12078_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_12079_, _12037_, _12031_);
  and (_12080_, _12079_, _11778_);
  and (_12081_, _12074_, _12038_);
  nor (_12082_, _12081_, _12080_);
  nor (_12084_, _12082_, _12078_);
  and (_12085_, _12082_, _12078_);
  nor (_12086_, _12085_, _12084_);
  and (_12087_, _11725_, _12079_);
  and (_12088_, _07429_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  and (_12090_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12091_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  not (_12092_, \oc8051_top_1.oc8051_memory_interface1.idat_old [29]);
  nor (_12093_, _07241_, _12092_);
  nor (_12094_, _12093_, _12091_);
  and (_12095_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_12096_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [5]);
  nor (_12097_, _12096_, _12095_);
  and (_12098_, _12097_, _12094_);
  and (_12099_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_12100_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [21]);
  nor (_12101_, _12100_, _12099_);
  and (_12102_, _12101_, _12098_);
  nor (_12103_, _12102_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12104_, _12103_, _12090_);
  nor (_12105_, _12104_, _07429_);
  nor (_12106_, _12105_, _12088_);
  and (_12107_, _12106_, _12038_);
  nor (_12108_, _12107_, _12087_);
  nor (_12109_, _12108_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_12110_, _12108_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_12111_, _11649_, _12079_);
  and (_12112_, _07429_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  or (_12113_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _07234_);
  and (_12114_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_12115_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [28]);
  or (_12116_, _12115_, _12114_);
  and (_12117_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_12118_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_12119_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [4]);
  or (_12120_, _12119_, _12118_);
  or (_12121_, _12120_, _12117_);
  or (_12122_, _12121_, _12116_);
  and (_12123_, _07242_, \oc8051_top_1.oc8051_memory_interface1.idat_old [28]);
  or (_12124_, _12123_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  or (_12125_, _12124_, _12122_);
  and (_12126_, _12125_, _07230_);
  and (_12127_, _12126_, _12113_);
  nor (_12128_, _12127_, _12112_);
  and (_12129_, _12128_, _12038_);
  nor (_12130_, _12129_, _12111_);
  nand (_12131_, _12130_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_12132_, _11688_, _12079_);
  and (_12134_, _07429_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  and (_12135_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12136_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  not (_12137_, \oc8051_top_1.oc8051_memory_interface1.idat_old [27]);
  nor (_12138_, _07241_, _12137_);
  nor (_12139_, _12138_, _12136_);
  and (_12141_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [19]);
  and (_12142_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nor (_12144_, _12142_, _12141_);
  and (_12145_, _12144_, _12139_);
  and (_12146_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_12147_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [19]);
  nor (_12148_, _12147_, _12146_);
  and (_12149_, _12148_, _12145_);
  nor (_12150_, _12149_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12151_, _12150_, _12135_);
  nor (_12152_, _12151_, _07429_);
  nor (_12154_, _12152_, _12134_);
  and (_12155_, _12154_, _12038_);
  nor (_12156_, _12155_, _12132_);
  nor (_12157_, _12156_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_12158_, _12156_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  not (_12160_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  or (_12161_, _11905_, _12038_);
  not (_12162_, _11209_);
  or (_12163_, _12079_, _12162_);
  nand (_12164_, _12163_, _12161_);
  or (_12165_, _12164_, _12160_);
  not (_12166_, _12165_);
  or (_12167_, _12038_, _11794_);
  and (_12168_, _07429_, \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  and (_12169_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12170_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  not (_12171_, \oc8051_top_1.oc8051_memory_interface1.idat_old [25]);
  nor (_12172_, _07241_, _12171_);
  nor (_12173_, _12172_, _12170_);
  and (_12174_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_12175_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_12176_, _12175_, _12174_);
  and (_12177_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [17]);
  and (_12178_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_12179_, _12178_, _12177_);
  and (_12180_, _12179_, _12176_);
  and (_12181_, _12180_, _12173_);
  nor (_12182_, _12181_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12183_, _12182_, _12169_);
  nor (_12184_, _12183_, _07429_);
  nor (_12185_, _12184_, _12168_);
  not (_12186_, _12185_);
  or (_12187_, _12186_, _12079_);
  and (_12188_, _12187_, _12167_);
  nand (_12189_, _12188_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  or (_12190_, _11848_, _12038_);
  not (_12191_, _09672_);
  or (_12192_, _12079_, _12191_);
  and (_12193_, _12192_, _12190_);
  and (_12194_, _12193_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  or (_12195_, _12188_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_12196_, _12195_, _12189_);
  and (_12197_, _12196_, _12194_);
  not (_12198_, _12197_);
  nand (_12199_, _12198_, _12189_);
  nand (_12200_, _12164_, _12160_);
  and (_12201_, _12200_, _12165_);
  and (_12202_, _12201_, _12199_);
  or (_12203_, _12202_, _12166_);
  nor (_12204_, _12203_, _12158_);
  nor (_12205_, _12204_, _12157_);
  or (_12206_, _12130_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_12207_, _12206_, _12131_);
  nand (_12208_, _12207_, _12205_);
  nand (_12209_, _12208_, _12131_);
  nor (_12210_, _12209_, _12110_);
  nor (_12211_, _12210_, _12109_);
  and (_12212_, _12211_, _12086_);
  nor (_12213_, _12211_, _12086_);
  nor (_12214_, _12213_, _12212_);
  and (_12215_, _11385_, _11342_);
  and (_12216_, _12215_, _11431_);
  or (_12217_, _12216_, _12045_);
  and (_12218_, _12217_, _12052_);
  and (_12219_, _12218_, _12214_);
  or (_12220_, _12219_, _12077_);
  nor (_12221_, _12220_, _12050_);
  nand (_12222_, _12221_, _12023_);
  not (_12223_, _07432_);
  and (_12224_, _10949_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_12225_, _12224_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_12226_, _12225_, _12223_);
  and (_12227_, _12226_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_12228_, _12226_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_12229_, _12228_, _12227_);
  or (_12230_, _12229_, _12023_);
  and (_12231_, _12230_, _06444_);
  and (_09725_, _12231_, _12222_);
  nor (_09730_, _11884_, rst);
  or (_12232_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [5]);
  nand (_12233_, _07432_, _10716_);
  and (_12234_, _12233_, _06444_);
  and (_09742_, _12234_, _12232_);
  and (_12235_, _08866_, _08655_);
  not (_12236_, _12235_);
  and (_12237_, _08869_, _09400_);
  not (_12238_, _12237_);
  or (_12239_, _12238_, word_in[8]);
  not (_12240_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_12241_, _10069_, _08877_);
  nor (_12242_, _12241_, _12240_);
  and (_12243_, _12241_, word_in[0]);
  or (_12244_, _12243_, _12242_);
  or (_12245_, _12244_, _12237_);
  and (_12246_, _12245_, _12239_);
  and (_12247_, _12246_, _12236_);
  and (_12248_, _08855_, _09219_);
  and (_12249_, _12235_, _09837_);
  or (_12250_, _12249_, _12248_);
  or (_12251_, _12250_, _12247_);
  not (_12252_, _12248_);
  or (_12253_, _12252_, _09554_);
  and (_09784_, _12253_, _12251_);
  not (_12254_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_12255_, _12241_, _12254_);
  and (_12256_, _12241_, word_in[1]);
  or (_12257_, _12256_, _12255_);
  and (_12258_, _12257_, _12238_);
  and (_12260_, _12237_, word_in[9]);
  or (_12261_, _12260_, _12258_);
  and (_12262_, _12261_, _12236_);
  and (_12263_, _12235_, _09565_);
  or (_12264_, _12263_, _12248_);
  or (_12265_, _12264_, _12262_);
  or (_12266_, _12252_, _11261_);
  and (_09786_, _12266_, _12265_);
  not (_12267_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_12268_, _12241_, _12267_);
  and (_12269_, _12241_, word_in[2]);
  or (_12270_, _12269_, _12268_);
  and (_12271_, _12270_, _12238_);
  and (_12272_, _12237_, word_in[10]);
  or (_12273_, _12272_, _12271_);
  and (_12274_, _12273_, _12236_);
  and (_12275_, _12235_, _10099_);
  or (_12276_, _12275_, _12248_);
  or (_12277_, _12276_, _12274_);
  or (_12278_, _12252_, _09582_);
  and (_09789_, _12278_, _12277_);
  or (_12279_, _12238_, word_in[11]);
  not (_12280_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_12281_, _12241_, _12280_);
  and (_12282_, _12241_, word_in[3]);
  or (_12283_, _12282_, _12281_);
  or (_12284_, _12283_, _12237_);
  and (_12285_, _12284_, _12279_);
  and (_12286_, _12285_, _12236_);
  and (_12287_, _12235_, _10116_);
  or (_12288_, _12287_, _12248_);
  or (_12289_, _12288_, _12286_);
  or (_12290_, _12252_, _09596_);
  and (_09791_, _12290_, _12289_);
  or (_12291_, _12238_, word_in[12]);
  not (_12292_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_12293_, _12241_, _12292_);
  and (_12294_, _12241_, word_in[4]);
  or (_12295_, _12294_, _12293_);
  or (_12296_, _12295_, _12237_);
  and (_12297_, _12296_, _12291_);
  and (_12298_, _12297_, _12236_);
  and (_12299_, _12235_, _10020_);
  or (_12300_, _12299_, _12248_);
  or (_12301_, _12300_, _12298_);
  or (_12302_, _12252_, _09609_);
  and (_09793_, _12302_, _12301_);
  not (_12303_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_12305_, _12241_, _12303_);
  and (_12306_, _12241_, word_in[5]);
  or (_12307_, _12306_, _12305_);
  and (_12308_, _12307_, _12238_);
  and (_12309_, _12237_, word_in[13]);
  or (_12310_, _12309_, _12308_);
  and (_12311_, _12310_, _12236_);
  and (_12312_, _12235_, _10149_);
  or (_12313_, _12312_, _12248_);
  or (_12314_, _12313_, _12311_);
  or (_12315_, _12252_, _09623_);
  and (_09796_, _12315_, _12314_);
  or (_12316_, _12238_, word_in[14]);
  not (_12318_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_12319_, _12241_, _12318_);
  and (_12320_, _12241_, word_in[6]);
  or (_12321_, _12320_, _12319_);
  or (_12322_, _12321_, _12237_);
  and (_12323_, _12322_, _12316_);
  and (_12324_, _12323_, _12236_);
  and (_12325_, _12235_, _10154_);
  or (_12326_, _12325_, _12248_);
  or (_12327_, _12326_, _12324_);
  or (_12328_, _12252_, _09626_);
  and (_09799_, _12328_, _12327_);
  nor (_12329_, _12241_, _08685_);
  and (_12330_, _12241_, word_in[7]);
  or (_12331_, _12330_, _12329_);
  and (_12332_, _12331_, _12238_);
  and (_12333_, _12237_, word_in[15]);
  or (_12335_, _12333_, _12332_);
  and (_12336_, _12335_, _12236_);
  and (_12337_, _12235_, _08886_);
  or (_12338_, _12337_, _12248_);
  or (_12339_, _12338_, _12336_);
  or (_12340_, _12252_, _08856_);
  and (_09801_, _12340_, _12339_);
  nor (_09849_, _11765_, rst);
  nor (_09852_, _11847_, rst);
  nor (_09859_, _11649_, rst);
  nor (_09863_, _12185_, rst);
  and (_12342_, _08855_, _08655_);
  and (_12343_, _12342_, _08842_);
  not (_12344_, _12343_);
  and (_12345_, _08866_, _08613_);
  and (_12346_, _09695_, _08679_);
  not (_12347_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_12348_, _09699_, _08877_);
  nor (_12349_, _12348_, _12347_);
  and (_12350_, _12348_, word_in[0]);
  or (_12352_, _12350_, _12349_);
  or (_12353_, _12352_, _12346_);
  not (_12354_, _12346_);
  or (_12355_, _12354_, word_in[8]);
  and (_12357_, _12355_, _12353_);
  or (_12358_, _12357_, _12345_);
  not (_12359_, _12345_);
  or (_12360_, _12359_, _09837_);
  and (_12361_, _12360_, _12358_);
  and (_12362_, _12361_, _12344_);
  and (_12363_, _12343_, word_in[24]);
  or (_14571_, _12363_, _12362_);
  and (_12364_, _12348_, word_in[1]);
  not (_12365_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_12366_, _12348_, _12365_);
  nor (_12367_, _12366_, _12364_);
  nor (_12368_, _12367_, _12346_);
  and (_12369_, _12346_, word_in[9]);
  or (_12370_, _12369_, _12368_);
  and (_12371_, _12370_, _12359_);
  and (_12372_, _12345_, _09565_);
  or (_12373_, _12372_, _12371_);
  and (_12374_, _12373_, _12344_);
  and (_12376_, _12343_, word_in[25]);
  or (_09872_, _12376_, _12374_);
  and (_12377_, _12348_, word_in[2]);
  not (_12378_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_12379_, _12348_, _12378_);
  nor (_12381_, _12379_, _12377_);
  nor (_12382_, _12381_, _12346_);
  and (_12383_, _12346_, word_in[10]);
  or (_12384_, _12383_, _12382_);
  and (_12385_, _12384_, _12359_);
  and (_12386_, _12345_, _10099_);
  or (_12387_, _12386_, _12385_);
  and (_12388_, _12387_, _12344_);
  and (_12389_, _12343_, word_in[26]);
  or (_09877_, _12389_, _12388_);
  and (_12390_, _12348_, word_in[3]);
  not (_12391_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_12392_, _12348_, _12391_);
  nor (_12393_, _12392_, _12390_);
  nor (_12394_, _12393_, _12346_);
  and (_12395_, _12346_, word_in[11]);
  or (_12396_, _12395_, _12394_);
  and (_12397_, _12396_, _12359_);
  and (_12398_, _12345_, _10116_);
  or (_12399_, _12398_, _12397_);
  and (_12400_, _12399_, _12344_);
  and (_12401_, _12343_, word_in[27]);
  or (_09880_, _12401_, _12400_);
  and (_12402_, _12348_, word_in[4]);
  not (_12403_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_12404_, _12348_, _12403_);
  nor (_12405_, _12404_, _12402_);
  nor (_12406_, _12405_, _12346_);
  and (_12408_, _12346_, word_in[12]);
  or (_12410_, _12408_, _12406_);
  and (_12411_, _12410_, _12359_);
  and (_12412_, _12345_, _10020_);
  or (_12413_, _12412_, _12411_);
  and (_12414_, _12413_, _12344_);
  and (_12415_, _12343_, word_in[28]);
  or (_09884_, _12415_, _12414_);
  not (_12416_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_12417_, _12348_, _12416_);
  and (_12418_, _12348_, word_in[5]);
  nor (_12419_, _12418_, _12417_);
  nor (_12420_, _12419_, _12346_);
  and (_12421_, _12346_, word_in[13]);
  or (_12422_, _12421_, _12420_);
  and (_12423_, _12422_, _12359_);
  and (_12424_, _12345_, _10149_);
  or (_12425_, _12424_, _12423_);
  and (_12426_, _12425_, _12344_);
  and (_12427_, _12343_, word_in[29]);
  or (_09887_, _12427_, _12426_);
  and (_12428_, _12348_, word_in[6]);
  not (_12429_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_12430_, _12348_, _12429_);
  nor (_12431_, _12430_, _12428_);
  nor (_12432_, _12431_, _12346_);
  and (_12433_, _12346_, word_in[14]);
  or (_12434_, _12433_, _12432_);
  and (_12435_, _12434_, _12359_);
  and (_12436_, _12345_, _10154_);
  or (_12437_, _12436_, _12435_);
  and (_12438_, _12437_, _12344_);
  and (_12439_, _12343_, word_in[30]);
  or (_09890_, _12439_, _12438_);
  nor (_12440_, _12348_, _08571_);
  and (_12441_, _12348_, word_in[7]);
  nor (_12442_, _12441_, _12440_);
  nor (_12443_, _12442_, _12346_);
  and (_12444_, _12346_, word_in[15]);
  or (_12445_, _12444_, _12443_);
  and (_12446_, _12445_, _12359_);
  and (_12447_, _12345_, _08886_);
  or (_12448_, _12447_, _12446_);
  and (_12449_, _12448_, _12344_);
  and (_12450_, _12343_, word_in[31]);
  or (_09894_, _12450_, _12449_);
  or (_12451_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [3]);
  not (_12452_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [3]);
  nand (_12453_, _07432_, _12452_);
  and (_12454_, _12453_, _06444_);
  and (_09949_, _12454_, _12451_);
  and (_12455_, _09819_, _08679_);
  not (_12456_, _12455_);
  or (_12457_, _12456_, word_in[8]);
  and (_12458_, _08866_, _08611_);
  not (_12459_, _12458_);
  not (_12460_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_12461_, _09822_, _08819_);
  nor (_12462_, _12461_, _12460_);
  and (_12463_, _12461_, word_in[0]);
  or (_12464_, _12463_, _12462_);
  or (_12466_, _12464_, _12455_);
  and (_12467_, _12466_, _12459_);
  and (_12468_, _12467_, _12457_);
  and (_12469_, _09835_, _08842_);
  and (_12470_, _12458_, _09837_);
  or (_12471_, _12470_, _12469_);
  or (_12472_, _12471_, _12468_);
  not (_12473_, _12469_);
  or (_12474_, _12473_, word_in[24]);
  and (_09955_, _12474_, _12472_);
  and (_12475_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  and (_12476_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [12]);
  or (_12477_, _12476_, _12475_);
  and (_09958_, _12477_, _06444_);
  not (_12478_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  nor (_12479_, _12461_, _12478_);
  and (_12480_, _12461_, word_in[1]);
  nor (_12481_, _12480_, _12479_);
  nor (_12482_, _12481_, _12455_);
  and (_12483_, _12455_, word_in[9]);
  or (_12484_, _12483_, _12482_);
  and (_12485_, _12484_, _12459_);
  and (_12486_, _12458_, _09565_);
  or (_12488_, _12486_, _12469_);
  or (_12489_, _12488_, _12485_);
  or (_12490_, _12473_, word_in[25]);
  and (_09960_, _12490_, _12489_);
  or (_12491_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [8]);
  not (_12492_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [8]);
  nand (_12493_, _07432_, _12492_);
  and (_12494_, _12493_, _06444_);
  and (_09962_, _12494_, _12491_);
  not (_12495_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  nor (_12496_, _12461_, _12495_);
  and (_12497_, _12461_, word_in[2]);
  nor (_12498_, _12497_, _12496_);
  nor (_12499_, _12498_, _12455_);
  and (_12500_, _12455_, word_in[10]);
  or (_12501_, _12500_, _12499_);
  and (_12502_, _12501_, _12459_);
  and (_12503_, _12458_, _10099_);
  or (_12504_, _12503_, _12469_);
  or (_12505_, _12504_, _12502_);
  or (_12506_, _12473_, word_in[26]);
  and (_09964_, _12506_, _12505_);
  and (_12507_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  and (_12508_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [22]);
  or (_12509_, _12508_, _12507_);
  and (_09967_, _12509_, _06444_);
  not (_12510_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  nor (_12511_, _12461_, _12510_);
  and (_12512_, _12461_, word_in[3]);
  nor (_12513_, _12512_, _12511_);
  nor (_12514_, _12513_, _12455_);
  and (_12515_, _12455_, word_in[11]);
  or (_12516_, _12515_, _12514_);
  and (_12517_, _12516_, _12459_);
  and (_12518_, _12458_, _10116_);
  or (_12519_, _12518_, _12469_);
  or (_12520_, _12519_, _12517_);
  or (_12521_, _12473_, word_in[27]);
  and (_09969_, _12521_, _12520_);
  or (_12522_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [18]);
  nand (_12523_, _07432_, _10712_);
  and (_12524_, _12523_, _06444_);
  and (_09972_, _12524_, _12522_);
  and (_12525_, _12461_, word_in[4]);
  not (_12526_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  nor (_12527_, _12461_, _12526_);
  nor (_12528_, _12527_, _12525_);
  nor (_12529_, _12528_, _12455_);
  and (_12530_, _12455_, word_in[12]);
  or (_12531_, _12530_, _12529_);
  and (_12532_, _12531_, _12459_);
  and (_12533_, _12458_, _10020_);
  or (_12534_, _12533_, _12469_);
  or (_12535_, _12534_, _12532_);
  or (_12536_, _12473_, word_in[28]);
  and (_09974_, _12536_, _12535_);
  not (_12537_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  nor (_12538_, _12461_, _12537_);
  and (_12539_, _12461_, word_in[5]);
  nor (_12540_, _12539_, _12538_);
  nor (_12541_, _12540_, _12455_);
  and (_12542_, _12455_, word_in[13]);
  or (_12543_, _12542_, _12541_);
  and (_12544_, _12543_, _12459_);
  and (_12545_, _12458_, _10149_);
  or (_12546_, _12545_, _12469_);
  or (_12547_, _12546_, _12544_);
  or (_12548_, _12473_, word_in[29]);
  and (_09976_, _12548_, _12547_);
  or (_12549_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [28]);
  nand (_12550_, _07432_, _10708_);
  and (_12551_, _12550_, _06444_);
  and (_09979_, _12551_, _12549_);
  not (_12552_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  nor (_12553_, _12461_, _12552_);
  and (_12554_, _12461_, word_in[6]);
  nor (_12555_, _12554_, _12553_);
  nor (_12556_, _12555_, _12455_);
  and (_12557_, _12455_, word_in[14]);
  or (_12558_, _12557_, _12556_);
  and (_12559_, _12558_, _12459_);
  and (_12560_, _12458_, _10154_);
  or (_12561_, _12560_, _12469_);
  or (_12562_, _12561_, _12559_);
  or (_12563_, _12473_, word_in[30]);
  and (_09981_, _12563_, _12562_);
  nor (_12564_, _12461_, _08680_);
  and (_12565_, _12461_, word_in[7]);
  nor (_12566_, _12565_, _12564_);
  nor (_12567_, _12566_, _12455_);
  and (_12568_, _12455_, word_in[15]);
  or (_12569_, _12568_, _12567_);
  and (_12570_, _12569_, _12459_);
  and (_12571_, _12458_, _08886_);
  or (_12572_, _12571_, _12469_);
  or (_12573_, _12572_, _12570_);
  or (_12574_, _12473_, word_in[31]);
  and (_09983_, _12574_, _12573_);
  nor (_09996_, _11830_, rst);
  and (_12575_, _12048_, _08127_);
  and (_12576_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_12577_, _12106_, _12033_);
  and (_12578_, _12054_, _11726_);
  or (_12579_, _12578_, _12577_);
  or (_12580_, _12579_, _12576_);
  or (_12581_, _12110_, _12109_);
  and (_12582_, _12581_, _12209_);
  nor (_12583_, _12581_, _12209_);
  or (_12584_, _12583_, _12582_);
  and (_12585_, _12584_, _12218_);
  nor (_12586_, _12585_, _12580_);
  nand (_12587_, _12586_, _12023_);
  or (_12588_, _12587_, _12575_);
  and (_12589_, _10949_, _08483_);
  nor (_12590_, _12589_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  nor (_12591_, _12590_, _12226_);
  or (_12592_, _12591_, _12023_);
  and (_12593_, _12592_, _06444_);
  and (_10009_, _12593_, _12588_);
  or (_12594_, _12023_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_12595_, _12594_, _06444_);
  and (_12596_, _12048_, _08019_);
  and (_12597_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  and (_12598_, _12032_, _12191_);
  and (_12600_, _12054_, _11848_);
  or (_12601_, _12600_, _12598_);
  or (_12602_, _12601_, _12597_);
  or (_12603_, _12193_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  not (_12604_, _12194_);
  or (_12605_, _12045_, _12034_);
  and (_12606_, _12605_, _12052_);
  and (_12607_, _12606_, _12604_);
  and (_12608_, _12607_, _12603_);
  or (_12609_, _12608_, _12602_);
  nor (_12610_, _12609_, _12596_);
  nand (_12611_, _12610_, _12023_);
  and (_10012_, _12611_, _12595_);
  and (_12612_, _12227_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_12613_, _12612_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  and (_12614_, _12613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_12615_, _12614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_12616_, _12615_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_12617_, _12616_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nand (_12618_, _12616_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_12619_, _12618_, _12617_);
  or (_12620_, _12619_, _12023_);
  and (_12621_, _12620_, _06444_);
  and (_12622_, _11452_, _08230_);
  and (_12623_, _12026_, _08267_);
  and (_12624_, _11650_, _12032_);
  and (_12625_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  or (_12626_, _12625_, _12624_);
  or (_12627_, _12626_, _12623_);
  or (_12628_, _12627_, _12622_);
  and (_12629_, _12079_, _08376_);
  and (_12630_, _07429_, \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  and (_12631_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  and (_12632_, _07254_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  not (_12633_, \oc8051_top_1.oc8051_memory_interface1.idat_old [31]);
  nor (_12634_, _07241_, _12633_);
  nor (_12635_, _12634_, _12632_);
  and (_12636_, _07248_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [23]);
  and (_12637_, _07238_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_12638_, _12637_, _12636_);
  and (_12639_, _12638_, _12635_);
  and (_12640_, _07246_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_12641_, _07251_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_12643_, _12641_, _12640_);
  and (_12644_, _12643_, _12639_);
  nor (_12645_, _12644_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nor (_12646_, _12645_, _12631_);
  nor (_12647_, _12646_, _07429_);
  nor (_12648_, _12647_, _12630_);
  and (_12649_, _12648_, _12038_);
  nor (_12650_, _12649_, _12629_);
  and (_12651_, _12650_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_12652_, _12650_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_12653_, _12652_, _12651_);
  or (_12654_, _12212_, _12084_);
  and (_12655_, _12654_, _12653_);
  or (_12656_, _12655_, _12651_);
  or (_12657_, _12656_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_12658_, _12657_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  or (_12659_, _12658_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  or (_12660_, _12659_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand (_12661_, _12660_, _12650_);
  not (_12662_, _12650_);
  and (_12663_, \oc8051_top_1.oc8051_memory_interface1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_12664_, _12663_, _12656_);
  and (_12665_, _12664_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nand (_12666_, _12665_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nand (_12667_, _12666_, _12662_);
  nand (_12668_, _12667_, _12661_);
  nand (_12669_, _12668_, _08150_);
  or (_12670_, _12668_, _08150_);
  and (_12671_, _12670_, _12669_);
  and (_12672_, _12671_, _12218_);
  or (_12673_, _12672_, _12628_);
  and (_12674_, \oc8051_top_1.oc8051_memory_interface1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_12675_, \oc8051_top_1.oc8051_memory_interface1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  and (_12676_, _12675_, _12674_);
  and (_12677_, \oc8051_top_1.oc8051_memory_interface1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_12678_, \oc8051_top_1.oc8051_memory_interface1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_12679_, _12678_, _12663_);
  and (_12680_, _12679_, _12677_);
  and (_12681_, _12680_, _12676_);
  and (_12682_, _12681_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_12683_, _12682_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_12684_, _12682_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_12685_, _12684_, _12683_);
  nand (_12686_, _12685_, _12054_);
  nand (_12687_, _12686_, _12023_);
  or (_12688_, _12687_, _12673_);
  and (_10017_, _12688_, _12621_);
  or (_12689_, _10963_, _10957_);
  and (_12690_, _12689_, _10964_);
  or (_12691_, _12690_, _08374_);
  or (_12692_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  and (_12693_, _12692_, _10894_);
  and (_12694_, _12693_, _12691_);
  and (_12695_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_10025_, _12695_, _12694_);
  nor (_12696_, _10947_, _10933_);
  nor (_12697_, _12696_, _10948_);
  or (_12698_, _12697_, _08374_);
  or (_12699_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  and (_12700_, _12699_, _10894_);
  and (_12701_, _12700_, _12698_);
  and (_12702_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  or (_10029_, _12702_, _12701_);
  and (_12703_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _06444_);
  not (_12704_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  nor (_12705_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  nor (_12706_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_12707_, _12706_, _12705_);
  not (_12708_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  nor (_12709_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_12710_, _12709_, _12708_);
  and (_12711_, _12710_, _12707_);
  and (_12712_, _12711_, _12704_);
  and (_12713_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _06444_);
  and (_12714_, _12713_, _12712_);
  or (_10037_, _12714_, _12703_);
  and (_12715_, _09554_, _08859_);
  and (_12716_, _08878_, word_in[0]);
  not (_12717_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  nor (_12718_, _08878_, _12717_);
  nor (_12719_, _12718_, _12716_);
  nor (_12720_, _12719_, _08871_);
  and (_12721_, _08871_, word_in[8]);
  or (_12722_, _12721_, _12720_);
  and (_12723_, _12722_, _08868_);
  and (_12724_, _09837_, _08867_);
  or (_12725_, _12724_, _12723_);
  and (_12726_, _12725_, _08862_);
  or (_14572_, _12726_, _12715_);
  nor (_10040_, _11725_, rst);
  and (_12727_, _11261_, _08859_);
  and (_12728_, _08878_, word_in[1]);
  not (_12729_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  nor (_12730_, _08878_, _12729_);
  nor (_12731_, _12730_, _12728_);
  nor (_12732_, _12731_, _08871_);
  and (_12733_, _08871_, word_in[9]);
  or (_12734_, _12733_, _12732_);
  and (_12735_, _12734_, _08868_);
  and (_12736_, _09565_, _08867_);
  or (_12737_, _12736_, _12735_);
  and (_12738_, _12737_, _08862_);
  or (_14573_, _12738_, _12727_);
  and (_12739_, _09582_, _08859_);
  and (_12740_, _08878_, word_in[2]);
  not (_12741_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  nor (_12742_, _08878_, _12741_);
  nor (_12743_, _12742_, _12740_);
  nor (_12744_, _12743_, _08871_);
  and (_12745_, _08871_, word_in[10]);
  or (_12746_, _12745_, _12744_);
  and (_12747_, _12746_, _08868_);
  and (_12748_, _10099_, _08867_);
  or (_12750_, _12748_, _12747_);
  and (_12751_, _12750_, _08862_);
  or (_14574_, _12751_, _12739_);
  and (_12753_, _08878_, word_in[3]);
  not (_12754_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  nor (_12755_, _08878_, _12754_);
  nor (_12756_, _12755_, _12753_);
  nor (_12757_, _12756_, _08871_);
  and (_12758_, _08871_, word_in[11]);
  or (_12759_, _12758_, _12757_);
  and (_12760_, _12759_, _08868_);
  and (_12761_, _10116_, _08867_);
  or (_12762_, _12761_, _12760_);
  and (_12763_, _12762_, _08862_);
  and (_12764_, _08859_, word_in[27]);
  or (_14575_, _12764_, _12763_);
  and (_12765_, _08878_, word_in[4]);
  not (_12766_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  nor (_12767_, _08878_, _12766_);
  nor (_12768_, _12767_, _12765_);
  nor (_12770_, _12768_, _08871_);
  and (_12771_, _08871_, word_in[12]);
  or (_12772_, _12771_, _12770_);
  and (_12773_, _12772_, _08868_);
  and (_12774_, _10020_, _08867_);
  or (_12775_, _12774_, _12773_);
  and (_12776_, _12775_, _08862_);
  and (_12777_, _08859_, word_in[28]);
  or (_14576_, _12777_, _12776_);
  and (_12778_, _08878_, word_in[5]);
  not (_12779_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  nor (_12780_, _08878_, _12779_);
  nor (_12781_, _12780_, _12778_);
  nor (_12782_, _12781_, _08871_);
  and (_12783_, _08871_, word_in[13]);
  or (_12784_, _12783_, _12782_);
  and (_12785_, _12784_, _08868_);
  and (_12786_, _10149_, _08867_);
  or (_12787_, _12786_, _12785_);
  and (_12788_, _12787_, _08862_);
  and (_12789_, _08859_, word_in[29]);
  or (_14577_, _12789_, _12788_);
  and (_12790_, \oc8051_top_1.oc8051_memory_interface1.cdata [0], _08478_);
  and (_12791_, \oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_12792_, _12791_, _12790_);
  and (_10053_, _12792_, _06444_);
  and (_12793_, _08878_, word_in[6]);
  not (_12794_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  nor (_12795_, _08878_, _12794_);
  nor (_12796_, _12795_, _12793_);
  nor (_12797_, _12796_, _08871_);
  and (_12798_, _08871_, word_in[14]);
  or (_12799_, _12798_, _12797_);
  and (_12800_, _12799_, _08868_);
  and (_12801_, _10154_, _08867_);
  or (_12802_, _12801_, _12800_);
  and (_12803_, _12802_, _08862_);
  and (_12804_, _08859_, word_in[30]);
  or (_14578_, _12804_, _12803_);
  and (_12805_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [4]);
  nor (_12806_, _07432_, _11044_);
  or (_12807_, _12806_, _12805_);
  and (_10345_, _12807_, _06444_);
  or (_12808_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  nand (_12809_, _07432_, _11220_);
  and (_12810_, _12809_, _06444_);
  and (_10354_, _12810_, _12808_);
  and (_12811_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [9]);
  not (_12812_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [9]);
  nor (_12813_, _07432_, _12812_);
  or (_12814_, _12813_, _12811_);
  and (_10357_, _12814_, _06444_);
  or (_12815_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  nand (_12816_, _07432_, _12137_);
  and (_12817_, _12816_, _06444_);
  and (_10362_, _12817_, _12815_);
  or (_12818_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [22]);
  nand (_12819_, _07432_, _10728_);
  and (_12820_, _12819_, _06444_);
  and (_10364_, _12820_, _12818_);
  nor (_12821_, _06299_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1]);
  nor (_12822_, _12821_, _08473_);
  and (_10468_, _12822_, _06443_);
  and (_10560_, t2_i, _06444_);
  not (_12823_, _07159_);
  and (_12824_, _09331_, _12823_);
  or (_12825_, _12824_, _07158_);
  and (_12826_, _12825_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nand (_12827_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [2]);
  nor (_12828_, _12827_, _07415_);
  and (_12829_, _07416_, _06439_);
  not (_12830_, _12829_);
  nor (_12831_, _12830_, _11589_);
  or (_12832_, _12831_, _12828_);
  or (_12833_, _12832_, _12826_);
  and (_10727_, _12833_, _06444_);
  not (_12834_, _12824_);
  nor (_12835_, _07156_, _12834_);
  nand (_12836_, _07415_, _06439_);
  or (_12837_, _12836_, _12835_);
  and (_12838_, _12837_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nand (_12839_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [0]);
  nor (_12840_, _12839_, _07418_);
  nor (_12841_, _09526_, _07158_);
  and (_12842_, _12841_, _07044_);
  or (_12843_, _12842_, _12840_);
  or (_12844_, _12843_, _12838_);
  and (_10802_, _12844_, _06444_);
  and (_12845_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_12846_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_12847_, _08064_, _12846_);
  or (_12848_, _12847_, _12845_);
  and (_10809_, _12848_, _06444_);
  nor (_12849_, _11589_, _06449_);
  and (_12850_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [2]);
  or (_12851_, _12850_, _12849_);
  and (_10905_, _12851_, _06444_);
  or (_12852_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  nand (_12853_, _07432_, _12092_);
  and (_12854_, _12853_, _06444_);
  and (_10922_, _12854_, _12852_);
  and (_12855_, _08558_, word_in[0]);
  nand (_12856_, _08480_, _11230_);
  or (_12857_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_12858_, _12857_, _12856_);
  and (_12859_, _12858_, _08506_);
  nand (_12860_, _08480_, _12347_);
  or (_12861_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  and (_12862_, _12861_, _12860_);
  and (_12863_, _12862_, _08503_);
  nand (_12865_, _08480_, _10608_);
  or (_12866_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  and (_12867_, _12866_, _12865_);
  and (_12868_, _12867_, _08523_);
  or (_12869_, _12868_, _12863_);
  or (_12871_, _12869_, _12859_);
  nand (_12872_, _08480_, _12717_);
  or (_12873_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_12874_, _12873_, _12872_);
  and (_12875_, _12874_, _08513_);
  or (_12876_, _12875_, _08532_);
  or (_12877_, _12876_, _12871_);
  nand (_12878_, _08480_, _09941_);
  or (_12879_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_12880_, _12879_, _12878_);
  and (_12881_, _12880_, _08506_);
  nand (_12882_, _08480_, _09697_);
  or (_12883_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  and (_12884_, _12883_, _12882_);
  and (_12885_, _12884_, _08523_);
  nand (_12886_, _08480_, _10183_);
  or (_12887_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  and (_12888_, _12887_, _12886_);
  and (_12890_, _12888_, _08503_);
  or (_12891_, _12890_, _12885_);
  or (_12892_, _12891_, _12881_);
  nand (_12893_, _08480_, _10396_);
  or (_12894_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_12895_, _12894_, _12893_);
  and (_12896_, _12895_, _08513_);
  or (_12897_, _12896_, _08489_);
  or (_12898_, _12897_, _12892_);
  and (_12899_, _12898_, _12877_);
  and (_12900_, _12899_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [0], _12900_, _12855_);
  and (_12901_, _08558_, word_in[1]);
  nand (_12902_, _08480_, _10624_);
  or (_12903_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  and (_12904_, _12903_, _12902_);
  and (_12905_, _12904_, _08523_);
  nand (_12906_, _08480_, _11249_);
  or (_12907_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_12908_, _12907_, _12906_);
  and (_12909_, _12908_, _08506_);
  nand (_12910_, _08480_, _12365_);
  or (_12911_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  and (_12912_, _12911_, _12910_);
  and (_12913_, _12912_, _08503_);
  or (_12914_, _12913_, _12909_);
  or (_12915_, _12914_, _12905_);
  nand (_12916_, _08480_, _12729_);
  or (_12917_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_12918_, _12917_, _12916_);
  and (_12919_, _12918_, _08513_);
  or (_12920_, _12919_, _08532_);
  or (_12921_, _12920_, _12915_);
  nand (_12922_, _08480_, _09720_);
  or (_12923_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  and (_12924_, _12923_, _12922_);
  and (_12925_, _12924_, _08523_);
  nand (_12926_, _08480_, _09963_);
  or (_12927_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_12928_, _12927_, _12926_);
  and (_12929_, _12928_, _08506_);
  nand (_12930_, _08480_, _10197_);
  or (_12931_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  and (_12932_, _12931_, _12930_);
  and (_12933_, _12932_, _08503_);
  or (_12934_, _12933_, _12929_);
  or (_12935_, _12934_, _12925_);
  nand (_12936_, _08480_, _10406_);
  or (_12937_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_12938_, _12937_, _12936_);
  and (_12939_, _12938_, _08513_);
  or (_12940_, _12939_, _08489_);
  or (_12941_, _12940_, _12935_);
  and (_12942_, _12941_, _12921_);
  and (_12943_, _12942_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [1], _12943_, _12901_);
  and (_12944_, _08558_, word_in[2]);
  nand (_12945_, _08480_, _10636_);
  or (_12946_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  and (_12947_, _12946_, _12945_);
  and (_12948_, _12947_, _08523_);
  nand (_12949_, _08480_, _11267_);
  or (_12950_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_12951_, _12950_, _12949_);
  and (_12952_, _12951_, _08506_);
  nand (_12953_, _08480_, _12378_);
  or (_12954_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  and (_12955_, _12954_, _12953_);
  and (_12956_, _12955_, _08503_);
  or (_12957_, _12956_, _12952_);
  or (_12958_, _12957_, _12948_);
  nand (_12959_, _08480_, _12741_);
  or (_12960_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_12961_, _12960_, _12959_);
  and (_12962_, _12961_, _08513_);
  or (_12963_, _12962_, _08532_);
  or (_12964_, _12963_, _12958_);
  nand (_12965_, _08480_, _09734_);
  or (_12966_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  and (_12967_, _12966_, _12965_);
  and (_12968_, _12967_, _08523_);
  nand (_12969_, _08480_, _09985_);
  or (_12970_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_12971_, _12970_, _12969_);
  and (_12972_, _12971_, _08506_);
  nand (_12973_, _08480_, _10209_);
  or (_12974_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  and (_12975_, _12974_, _12973_);
  and (_12976_, _12975_, _08503_);
  or (_12977_, _12976_, _12972_);
  or (_12978_, _12977_, _12968_);
  nand (_12979_, _08480_, _10420_);
  or (_12980_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_12981_, _12980_, _12979_);
  and (_12982_, _12981_, _08513_);
  or (_12983_, _12982_, _08489_);
  or (_12984_, _12983_, _12978_);
  and (_12985_, _12984_, _12964_);
  and (_12986_, _12985_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [2], _12986_, _12944_);
  and (_12987_, _08558_, word_in[3]);
  nand (_12988_, _08480_, _10649_);
  or (_12989_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  and (_12990_, _12989_, _12988_);
  and (_12991_, _12990_, _08523_);
  nand (_12992_, _08480_, _11279_);
  or (_12993_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_12994_, _12993_, _12992_);
  and (_12995_, _12994_, _08506_);
  nand (_12996_, _08480_, _12391_);
  or (_12997_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  and (_12998_, _12997_, _12996_);
  and (_12999_, _12998_, _08503_);
  or (_13000_, _12999_, _12995_);
  or (_13001_, _13000_, _12991_);
  nand (_13002_, _08480_, _12754_);
  or (_13003_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_13004_, _13003_, _13002_);
  and (_13005_, _13004_, _08513_);
  or (_13006_, _13005_, _08532_);
  or (_13007_, _13006_, _13001_);
  nand (_13008_, _08480_, _09749_);
  or (_13009_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  and (_13010_, _13009_, _13008_);
  and (_13012_, _13010_, _08523_);
  nand (_13013_, _08480_, _09998_);
  or (_13014_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_13015_, _13014_, _13013_);
  and (_13016_, _13015_, _08506_);
  nand (_13017_, _08480_, _10221_);
  or (_13018_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  and (_13019_, _13018_, _13017_);
  and (_13020_, _13019_, _08503_);
  or (_13021_, _13020_, _13016_);
  or (_13022_, _13021_, _13012_);
  nand (_13024_, _08480_, _10431_);
  or (_13025_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_13026_, _13025_, _13024_);
  and (_13027_, _13026_, _08513_);
  or (_13028_, _13027_, _08489_);
  or (_13029_, _13028_, _13022_);
  and (_13030_, _13029_, _13007_);
  and (_13031_, _13030_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [3], _13031_, _12987_);
  and (_13032_, _08558_, word_in[4]);
  nand (_13033_, _08480_, _10660_);
  or (_13034_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  and (_13035_, _13034_, _13033_);
  and (_13036_, _13035_, _08523_);
  nand (_13037_, _08480_, _11292_);
  or (_13039_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_13040_, _13039_, _13037_);
  and (_13041_, _13040_, _08506_);
  nand (_13042_, _08480_, _12403_);
  or (_13043_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  and (_13044_, _13043_, _13042_);
  and (_13045_, _13044_, _08503_);
  or (_13047_, _13045_, _13041_);
  or (_13048_, _13047_, _13036_);
  nand (_13049_, _08480_, _12766_);
  or (_13051_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_13052_, _13051_, _13049_);
  and (_13053_, _13052_, _08513_);
  or (_13054_, _13053_, _08532_);
  or (_13055_, _13054_, _13048_);
  nand (_13056_, _08480_, _09761_);
  or (_13057_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  and (_13058_, _13057_, _13056_);
  and (_13059_, _13058_, _08523_);
  nand (_13060_, _08480_, _10011_);
  or (_13061_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_13062_, _13061_, _13060_);
  and (_13063_, _13062_, _08506_);
  nand (_13064_, _08480_, _10233_);
  or (_13065_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  and (_13066_, _13065_, _13064_);
  and (_13067_, _13066_, _08503_);
  or (_13068_, _13067_, _13063_);
  or (_13069_, _13068_, _13059_);
  nand (_13070_, _08480_, _10443_);
  or (_13071_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_13072_, _13071_, _13070_);
  and (_13073_, _13072_, _08513_);
  or (_13074_, _13073_, _08489_);
  or (_13075_, _13074_, _13069_);
  and (_13076_, _13075_, _13055_);
  and (_13077_, _13076_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [4], _13077_, _13032_);
  and (_13079_, _08558_, word_in[5]);
  nand (_13080_, _08480_, _10672_);
  or (_13081_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  and (_13082_, _13081_, _13080_);
  and (_13083_, _13082_, _08523_);
  nand (_13084_, _08480_, _11305_);
  or (_13085_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_13086_, _13085_, _13084_);
  and (_13087_, _13086_, _08506_);
  nand (_13088_, _08480_, _12416_);
  or (_13089_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  and (_13090_, _13089_, _13088_);
  and (_13091_, _13090_, _08503_);
  or (_13092_, _13091_, _13087_);
  or (_13093_, _13092_, _13083_);
  nand (_13094_, _08480_, _12779_);
  or (_13095_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_13096_, _13095_, _13094_);
  and (_13097_, _13096_, _08513_);
  or (_13098_, _13097_, _08532_);
  or (_13099_, _13098_, _13093_);
  nand (_13100_, _08480_, _09775_);
  or (_13101_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  and (_13102_, _13101_, _13100_);
  and (_13103_, _13102_, _08523_);
  nand (_13104_, _08480_, _10027_);
  or (_13105_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  and (_13106_, _13105_, _13104_);
  and (_13107_, _13106_, _08506_);
  nand (_13109_, _08480_, _10245_);
  or (_13110_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  and (_13111_, _13110_, _13109_);
  and (_13112_, _13111_, _08503_);
  or (_13113_, _13112_, _13107_);
  or (_13114_, _13113_, _13103_);
  nand (_13115_, _08480_, _10454_);
  or (_13116_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_13117_, _13116_, _13115_);
  and (_13118_, _13117_, _08513_);
  or (_13119_, _13118_, _08489_);
  or (_13120_, _13119_, _13114_);
  and (_13121_, _13120_, _13099_);
  and (_13122_, _13121_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [5], _13122_, _13079_);
  and (_13123_, _08558_, word_in[6]);
  nand (_13124_, _08480_, _11318_);
  or (_13125_, _08480_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_13126_, _13125_, _13124_);
  and (_13127_, _13126_, _08506_);
  nand (_13128_, _08480_, _12429_);
  or (_13129_, _08480_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  and (_13130_, _13129_, _13128_);
  and (_13131_, _13130_, _08503_);
  nand (_13132_, _08480_, _10685_);
  or (_13133_, _08480_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  and (_13134_, _13133_, _13132_);
  and (_13135_, _13134_, _08523_);
  or (_13136_, _13135_, _13131_);
  or (_13137_, _13136_, _13127_);
  nand (_13139_, _08480_, _12794_);
  or (_13140_, _08480_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_13141_, _13140_, _13139_);
  and (_13142_, _13141_, _08513_);
  or (_13143_, _13142_, _08532_);
  or (_13144_, _13143_, _13137_);
  nand (_13145_, _08480_, _10042_);
  or (_13146_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  and (_13147_, _13146_, _13145_);
  and (_13149_, _13147_, _08506_);
  nand (_13151_, _08480_, _09792_);
  or (_13152_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  and (_13153_, _13152_, _13151_);
  and (_13154_, _13153_, _08523_);
  nand (_13155_, _08480_, _10258_);
  or (_13156_, _08480_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  and (_13157_, _13156_, _13155_);
  and (_13158_, _13157_, _08503_);
  or (_13159_, _13158_, _13154_);
  or (_13160_, _13159_, _13149_);
  nand (_13162_, _08480_, _10469_);
  or (_13163_, _08480_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_13164_, _13163_, _13162_);
  and (_13165_, _13164_, _08513_);
  or (_13166_, _13165_, _08489_);
  or (_13167_, _13166_, _13160_);
  and (_13168_, _13167_, _13144_);
  and (_13169_, _13168_, _08557_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [6], _13169_, _13123_);
  and (_13170_, _08664_, word_in[8]);
  nand (_13171_, _08480_, _10998_);
  or (_13172_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_13173_, _13172_, _13171_);
  and (_13174_, _13173_, _08666_);
  nand (_13175_, _08480_, _10504_);
  or (_13176_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  and (_13177_, _13176_, _13175_);
  and (_13178_, _13177_, _08665_);
  or (_13179_, _13178_, _13174_);
  and (_13180_, _13179_, _08623_);
  nand (_13181_, _08480_, _12460_);
  or (_13182_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_13183_, _13182_, _13181_);
  and (_13184_, _13183_, _08666_);
  nand (_13185_, _08480_, _12240_);
  or (_13186_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  and (_13187_, _13186_, _13185_);
  and (_13188_, _13187_, _08665_);
  or (_13189_, _13188_, _13184_);
  and (_13190_, _13189_, _08679_);
  nand (_13191_, _08480_, _10290_);
  or (_13192_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_13193_, _13192_, _13191_);
  and (_13194_, _13193_, _08666_);
  nand (_13195_, _08480_, _10068_);
  or (_13196_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  and (_13197_, _13196_, _13195_);
  and (_13198_, _13197_, _08665_);
  or (_13199_, _13198_, _13194_);
  and (_13200_, _13199_, _08708_);
  nand (_13201_, _08480_, _09821_);
  or (_13202_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_13203_, _13202_, _13201_);
  and (_13204_, _13203_, _08666_);
  and (_13205_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_13206_, _08480_, _09697_);
  or (_13207_, _13206_, _13205_);
  and (_13208_, _13207_, _08665_);
  or (_13209_, _13208_, _13204_);
  and (_13210_, _13209_, _08626_);
  or (_13211_, _13210_, _13200_);
  or (_13212_, _13211_, _13190_);
  nor (_13213_, _13212_, _13180_);
  nor (_13214_, _13213_, _08664_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [8], _13214_, _13170_);
  and (_13215_, _08664_, word_in[9]);
  nand (_13216_, _08480_, _11019_);
  or (_13217_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  and (_13218_, _13217_, _13216_);
  and (_13219_, _13218_, _08666_);
  nand (_13220_, _08480_, _10522_);
  or (_13221_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_13222_, _13221_, _13220_);
  and (_13223_, _13222_, _08665_);
  or (_13224_, _13223_, _13219_);
  and (_13225_, _13224_, _08623_);
  nand (_13226_, _08480_, _12478_);
  or (_13227_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_13228_, _13227_, _13226_);
  and (_13229_, _13228_, _08666_);
  nand (_13230_, _08480_, _12254_);
  or (_13231_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  and (_13232_, _13231_, _13230_);
  and (_13233_, _13232_, _08665_);
  or (_13234_, _13233_, _13229_);
  and (_13235_, _13234_, _08679_);
  nand (_13236_, _08480_, _10301_);
  or (_13237_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_13238_, _13237_, _13236_);
  and (_13239_, _13238_, _08666_);
  nand (_13240_, _08480_, _10087_);
  or (_13241_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  and (_13242_, _13241_, _13240_);
  and (_13243_, _13242_, _08665_);
  or (_13244_, _13243_, _13239_);
  and (_13245_, _13244_, _08708_);
  nand (_13246_, _08480_, _09843_);
  or (_13247_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  and (_13248_, _13247_, _13246_);
  and (_13249_, _13248_, _08666_);
  nand (_13250_, _08480_, _09556_);
  or (_13251_, _08480_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_13252_, _13251_, _13250_);
  and (_13253_, _13252_, _08665_);
  or (_13254_, _13253_, _13249_);
  and (_13255_, _13254_, _08626_);
  or (_13256_, _13255_, _13245_);
  or (_13257_, _13256_, _13235_);
  nor (_13258_, _13257_, _13225_);
  nor (_13259_, _13258_, _08664_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [9], _13259_, _13215_);
  and (_13260_, _08664_, word_in[10]);
  nand (_13261_, _08480_, _11032_);
  or (_13262_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  and (_13263_, _13262_, _13261_);
  and (_13264_, _13263_, _08666_);
  nand (_13265_, _08480_, _10534_);
  or (_13266_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_13267_, _13266_, _13265_);
  and (_13268_, _13267_, _08665_);
  or (_13269_, _13268_, _13264_);
  and (_13270_, _13269_, _08623_);
  nand (_13271_, _08480_, _12495_);
  or (_13272_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_13273_, _13272_, _13271_);
  and (_13274_, _13273_, _08666_);
  nand (_13275_, _08480_, _12267_);
  or (_13276_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  and (_13277_, _13276_, _13275_);
  and (_13278_, _13277_, _08665_);
  or (_13279_, _13278_, _13274_);
  and (_13280_, _13279_, _08679_);
  nand (_13281_, _08480_, _10313_);
  or (_13282_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_13283_, _13282_, _13281_);
  and (_13284_, _13283_, _08666_);
  nand (_13285_, _08480_, _10101_);
  or (_13286_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  and (_13287_, _13286_, _13285_);
  and (_13288_, _13287_, _08665_);
  or (_13289_, _13288_, _13284_);
  and (_13290_, _13289_, _08708_);
  nand (_13291_, _08480_, _09857_);
  or (_13292_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_13293_, _13292_, _13291_);
  and (_13294_, _13293_, _08666_);
  and (_13295_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_13296_, _08480_, _09734_);
  or (_13297_, _13296_, _13295_);
  and (_13298_, _13297_, _08665_);
  or (_13299_, _13298_, _13294_);
  and (_13301_, _13299_, _08626_);
  or (_13302_, _13301_, _13290_);
  or (_13303_, _13302_, _13280_);
  nor (_13304_, _13303_, _13270_);
  nor (_13305_, _13304_, _08664_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [10], _13305_, _13260_);
  and (_13306_, _08664_, word_in[11]);
  nand (_13307_, _08480_, _11047_);
  or (_13308_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  and (_13309_, _13308_, _13307_);
  and (_13310_, _13309_, _08666_);
  nand (_13311_, _08480_, _10546_);
  or (_13312_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_13313_, _13312_, _13311_);
  and (_13314_, _13313_, _08665_);
  or (_13315_, _13314_, _13310_);
  and (_13316_, _13315_, _08623_);
  nand (_13317_, _08480_, _12510_);
  or (_13318_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_13319_, _13318_, _13317_);
  and (_13320_, _13319_, _08666_);
  nand (_13321_, _08480_, _12280_);
  or (_13322_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  and (_13323_, _13322_, _13321_);
  and (_13324_, _13323_, _08665_);
  or (_13325_, _13324_, _13320_);
  and (_13326_, _13325_, _08679_);
  nand (_13327_, _08480_, _10325_);
  or (_13328_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_13329_, _13328_, _13327_);
  and (_13330_, _13329_, _08666_);
  nand (_13331_, _08480_, _10118_);
  or (_13332_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  and (_13333_, _13332_, _13331_);
  and (_13334_, _13333_, _08665_);
  or (_13335_, _13334_, _13330_);
  and (_13336_, _13335_, _08708_);
  nand (_13337_, _08480_, _09871_);
  or (_13338_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_13340_, _13338_, _13337_);
  and (_13341_, _13340_, _08666_);
  and (_13342_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_13343_, _08480_, _09749_);
  or (_13344_, _13343_, _13342_);
  and (_13345_, _13344_, _08665_);
  or (_13346_, _13345_, _13341_);
  and (_13347_, _13346_, _08626_);
  or (_13348_, _13347_, _13336_);
  or (_13349_, _13348_, _13326_);
  nor (_13350_, _13349_, _13316_);
  nor (_13351_, _13350_, _08664_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [11], _13351_, _13306_);
  and (_13352_, _08664_, word_in[12]);
  nand (_13353_, _08480_, _11059_);
  or (_13354_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  and (_13355_, _13354_, _13353_);
  and (_13356_, _13355_, _08666_);
  nand (_13357_, _08480_, _10558_);
  or (_13358_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_13359_, _13358_, _13357_);
  and (_13360_, _13359_, _08665_);
  or (_13361_, _13360_, _13356_);
  and (_13362_, _13361_, _08623_);
  nand (_13363_, _08480_, _09889_);
  or (_13365_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_13366_, _13365_, _13363_);
  and (_13367_, _13366_, _08666_);
  and (_13368_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_13369_, _08480_, _09761_);
  or (_13370_, _13369_, _13368_);
  and (_13371_, _13370_, _08665_);
  or (_13372_, _13371_, _13367_);
  and (_13373_, _13372_, _08626_);
  nand (_13374_, _08480_, _10337_);
  or (_13375_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_13376_, _13375_, _13374_);
  and (_13377_, _13376_, _08666_);
  nand (_13378_, _08480_, _10129_);
  or (_13379_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  and (_13380_, _13379_, _13378_);
  and (_13381_, _13380_, _08665_);
  or (_13382_, _13381_, _13377_);
  and (_13383_, _13382_, _08708_);
  or (_13384_, _13383_, _13373_);
  nand (_13385_, _08480_, _12526_);
  or (_13386_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_13388_, _13386_, _13385_);
  and (_13389_, _13388_, _08666_);
  nand (_13390_, _08480_, _12292_);
  or (_13391_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  and (_13392_, _13391_, _13390_);
  and (_13393_, _13392_, _08665_);
  or (_13394_, _13393_, _13389_);
  and (_13395_, _13394_, _08679_);
  or (_13396_, _13395_, _13384_);
  nor (_13397_, _13396_, _13362_);
  nor (_13398_, _13397_, _08664_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [12], _13398_, _13352_);
  and (_13399_, _08664_, word_in[13]);
  nand (_13400_, _08480_, _11071_);
  or (_13401_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_13402_, _13401_, _13400_);
  and (_13403_, _13402_, _08666_);
  nand (_13404_, _08480_, _10571_);
  or (_13405_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  and (_13406_, _13405_, _13404_);
  and (_13407_, _13406_, _08665_);
  or (_13408_, _13407_, _13403_);
  and (_13409_, _13408_, _08623_);
  and (_13410_, _08480_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_13411_, _08480_, _10027_);
  or (_13412_, _13411_, _13410_);
  and (_13413_, _13412_, _08666_);
  and (_13414_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_13415_, _08480_, _09775_);
  or (_13416_, _13415_, _13414_);
  and (_13417_, _13416_, _08665_);
  or (_13418_, _13417_, _13413_);
  and (_13419_, _13418_, _08626_);
  nand (_13420_, _08480_, _10350_);
  or (_13421_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_13423_, _13421_, _13420_);
  and (_13424_, _13423_, _08666_);
  nand (_13425_, _08480_, _10141_);
  or (_13426_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  and (_13427_, _13426_, _13425_);
  and (_13428_, _13427_, _08665_);
  or (_13429_, _13428_, _13424_);
  and (_13430_, _13429_, _08708_);
  or (_13431_, _13430_, _13419_);
  nand (_13432_, _08480_, _12537_);
  or (_13433_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_13434_, _13433_, _13432_);
  and (_13435_, _13434_, _08666_);
  nand (_13436_, _08480_, _12303_);
  or (_13437_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  and (_13438_, _13437_, _13436_);
  and (_13439_, _13438_, _08665_);
  or (_13440_, _13439_, _13435_);
  and (_13441_, _13440_, _08679_);
  or (_13442_, _13441_, _13431_);
  nor (_13443_, _13442_, _13409_);
  nor (_13444_, _13443_, _08664_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [13], _13444_, _13399_);
  and (_13445_, _08664_, word_in[14]);
  nand (_13446_, _08480_, _11084_);
  or (_13447_, _08480_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_13448_, _13447_, _13446_);
  and (_13449_, _13448_, _08666_);
  nand (_13450_, _08480_, _10583_);
  or (_13451_, _08480_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  and (_13452_, _13451_, _13450_);
  and (_13453_, _13452_, _08665_);
  or (_13454_, _13453_, _13449_);
  and (_13455_, _13454_, _08623_);
  nand (_13456_, _08480_, _12552_);
  or (_13457_, _08480_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_13458_, _13457_, _13456_);
  and (_13459_, _13458_, _08666_);
  nand (_13460_, _08480_, _12318_);
  or (_13461_, _08480_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  and (_13462_, _13461_, _13460_);
  and (_13463_, _13462_, _08665_);
  or (_13464_, _13463_, _13459_);
  and (_13465_, _13464_, _08679_);
  nand (_13466_, _08480_, _10366_);
  or (_13467_, _08480_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_13468_, _13467_, _13466_);
  and (_13469_, _13468_, _08666_);
  nand (_13470_, _08480_, _10156_);
  or (_13471_, _08480_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  and (_13472_, _13471_, _13470_);
  and (_13473_, _13472_, _08665_);
  or (_13474_, _13473_, _13469_);
  and (_13475_, _13474_, _08708_);
  nand (_13476_, _08480_, _09915_);
  or (_13477_, _08480_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_13478_, _13477_, _13476_);
  and (_13479_, _13478_, _08666_);
  and (_13480_, _08480_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_13481_, _08480_, _09792_);
  or (_13482_, _13481_, _13480_);
  and (_13483_, _13482_, _08665_);
  or (_13484_, _13483_, _13479_);
  and (_13485_, _13484_, _08626_);
  or (_13486_, _13485_, _13475_);
  or (_13487_, _13486_, _13465_);
  nor (_13488_, _13487_, _13455_);
  nor (_13489_, _13488_, _08664_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [14], _13489_, _13445_);
  and (_13490_, _08769_, word_in[16]);
  and (_13491_, _12888_, _08506_);
  and (_13492_, _12884_, _08513_);
  or (_13493_, _13492_, _13491_);
  and (_13494_, _12895_, _08503_);
  and (_13495_, _12880_, _08523_);
  or (_13496_, _13495_, _13494_);
  or (_13497_, _13496_, _13493_);
  or (_13498_, _13497_, _08731_);
  and (_13499_, _12862_, _08506_);
  and (_13500_, _12867_, _08513_);
  or (_13501_, _13500_, _13499_);
  and (_13502_, _12874_, _08503_);
  and (_13503_, _12858_, _08523_);
  or (_13504_, _13503_, _13502_);
  or (_13505_, _13504_, _13501_);
  or (_13506_, _13505_, _08770_);
  nand (_13507_, _13506_, _13498_);
  nor (_13508_, _13507_, _08769_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [16], _13508_, _13490_);
  and (_13509_, _08769_, word_in[17]);
  and (_13510_, _12924_, _08513_);
  and (_13511_, _12938_, _08503_);
  or (_13512_, _13511_, _13510_);
  and (_13513_, _12932_, _08506_);
  and (_13514_, _12928_, _08523_);
  or (_13515_, _13514_, _13513_);
  or (_13516_, _13515_, _13512_);
  or (_13517_, _13516_, _08731_);
  and (_13518_, _12912_, _08506_);
  and (_13520_, _12904_, _08513_);
  or (_13521_, _13520_, _13518_);
  and (_13522_, _12918_, _08503_);
  and (_13523_, _12908_, _08523_);
  or (_13524_, _13523_, _13522_);
  or (_13526_, _13524_, _13521_);
  or (_13527_, _13526_, _08770_);
  nand (_13528_, _13527_, _13517_);
  nor (_13529_, _13528_, _08769_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [17], _13529_, _13509_);
  and (_13530_, _08769_, word_in[18]);
  and (_13531_, _12975_, _08506_);
  and (_13532_, _12967_, _08513_);
  or (_13533_, _13532_, _13531_);
  and (_13534_, _12981_, _08503_);
  and (_13535_, _12971_, _08523_);
  or (_13536_, _13535_, _13534_);
  or (_13537_, _13536_, _13533_);
  or (_13538_, _13537_, _08731_);
  and (_13539_, _12955_, _08506_);
  and (_13540_, _12947_, _08513_);
  or (_13541_, _13540_, _13539_);
  and (_13542_, _12961_, _08503_);
  and (_13543_, _12951_, _08523_);
  or (_13544_, _13543_, _13542_);
  or (_13545_, _13544_, _13541_);
  or (_13546_, _13545_, _08770_);
  nand (_13547_, _13546_, _13538_);
  nor (_13549_, _13547_, _08769_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [18], _13549_, _13530_);
  and (_13550_, _08769_, word_in[19]);
  and (_13552_, _13010_, _08513_);
  and (_13553_, _13026_, _08503_);
  or (_13554_, _13553_, _13552_);
  and (_13555_, _13019_, _08506_);
  and (_13556_, _13015_, _08523_);
  or (_13557_, _13556_, _13555_);
  or (_13558_, _13557_, _13554_);
  or (_13559_, _13558_, _08731_);
  and (_13560_, _12998_, _08506_);
  and (_13561_, _12990_, _08513_);
  or (_13562_, _13561_, _13560_);
  and (_13563_, _13004_, _08503_);
  and (_13564_, _12994_, _08523_);
  or (_13565_, _13564_, _13563_);
  or (_13566_, _13565_, _13562_);
  or (_13567_, _13566_, _08770_);
  nand (_13568_, _13567_, _13559_);
  nor (_13569_, _13568_, _08769_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [19], _13569_, _13550_);
  and (_13570_, _08769_, word_in[20]);
  and (_13571_, _13058_, _08513_);
  and (_13572_, _13072_, _08503_);
  or (_13573_, _13572_, _13571_);
  and (_13574_, _13066_, _08506_);
  and (_13575_, _13062_, _08523_);
  or (_13576_, _13575_, _13574_);
  or (_13577_, _13576_, _13573_);
  or (_13578_, _13577_, _08731_);
  and (_13579_, _13035_, _08513_);
  and (_13580_, _13052_, _08503_);
  or (_13581_, _13580_, _13579_);
  and (_13582_, _13044_, _08506_);
  and (_13583_, _13040_, _08523_);
  or (_13584_, _13583_, _13582_);
  or (_13585_, _13584_, _13581_);
  or (_13586_, _13585_, _08770_);
  nand (_13587_, _13586_, _13578_);
  nor (_13588_, _13587_, _08769_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [20], _13588_, _13570_);
  and (_13590_, _08769_, word_in[21]);
  and (_13591_, _13102_, _08513_);
  and (_13592_, _13117_, _08503_);
  or (_13593_, _13592_, _13591_);
  and (_13594_, _13111_, _08506_);
  and (_13595_, _13106_, _08523_);
  or (_13597_, _13595_, _13594_);
  or (_13598_, _13597_, _13593_);
  or (_13599_, _13598_, _08731_);
  and (_13600_, _13082_, _08513_);
  and (_13601_, _13096_, _08503_);
  or (_13602_, _13601_, _13600_);
  and (_13603_, _13090_, _08506_);
  and (_13604_, _13086_, _08523_);
  or (_13605_, _13604_, _13603_);
  or (_13606_, _13605_, _13602_);
  or (_13607_, _13606_, _08770_);
  nand (_13608_, _13607_, _13599_);
  nor (_13609_, _13608_, _08769_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [21], _13609_, _13590_);
  and (_13610_, _08769_, word_in[22]);
  and (_13611_, _13157_, _08506_);
  and (_13612_, _13153_, _08513_);
  or (_13613_, _13612_, _13611_);
  and (_13614_, _13164_, _08503_);
  and (_13615_, _13147_, _08523_);
  or (_13616_, _13615_, _13614_);
  or (_13617_, _13616_, _13613_);
  or (_13618_, _13617_, _08731_);
  and (_13619_, _13130_, _08506_);
  and (_13620_, _13134_, _08513_);
  or (_13621_, _13620_, _13619_);
  and (_13622_, _13141_, _08503_);
  and (_13623_, _13126_, _08523_);
  or (_13624_, _13623_, _13622_);
  or (_13625_, _13624_, _13621_);
  or (_13626_, _13625_, _08770_);
  nand (_13627_, _13626_, _13618_);
  nor (_13628_, _13627_, _08769_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [22], _13628_, _13610_);
  and (_13629_, _08828_, word_in[24]);
  and (_13630_, _13207_, _08666_);
  and (_13631_, _13203_, _08665_);
  or (_13632_, _13631_, _13630_);
  and (_13633_, _13632_, _08814_);
  and (_13635_, _13177_, _08666_);
  and (_13636_, _13173_, _08665_);
  or (_13638_, _13636_, _13635_);
  and (_13639_, _13638_, _08800_);
  and (_13640_, _13197_, _08666_);
  and (_13641_, _13193_, _08665_);
  or (_13642_, _13641_, _13640_);
  and (_13643_, _13642_, _08837_);
  and (_13644_, _13187_, _08666_);
  and (_13645_, _13183_, _08665_);
  or (_13646_, _13645_, _13644_);
  and (_13647_, _13646_, _08842_);
  or (_13648_, _13647_, _13643_);
  or (_13649_, _13648_, _13639_);
  nor (_13650_, _13649_, _13633_);
  nor (_13651_, _13650_, _08828_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [24], _13651_, _13629_);
  and (_13652_, _08828_, word_in[25]);
  and (_13653_, _13222_, _08666_);
  and (_13654_, _13218_, _08665_);
  or (_13655_, _13654_, _13653_);
  and (_13656_, _13655_, _08800_);
  and (_13657_, _13252_, _08666_);
  and (_13658_, _13248_, _08665_);
  or (_13659_, _13658_, _13657_);
  and (_13660_, _13659_, _08814_);
  and (_13662_, _13242_, _08666_);
  and (_13663_, _13238_, _08665_);
  or (_13664_, _13663_, _13662_);
  and (_13666_, _13664_, _08837_);
  and (_13667_, _13232_, _08666_);
  and (_13668_, _13228_, _08665_);
  or (_13669_, _13668_, _13667_);
  and (_13670_, _13669_, _08842_);
  or (_13671_, _13670_, _13666_);
  or (_13672_, _13671_, _13660_);
  nor (_13673_, _13672_, _13656_);
  nor (_13674_, _13673_, _08828_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [25], _13674_, _13652_);
  and (_13676_, _08828_, word_in[26]);
  and (_13677_, _13297_, _08666_);
  and (_13678_, _13293_, _08665_);
  or (_13679_, _13678_, _13677_);
  and (_13680_, _13679_, _08814_);
  and (_13681_, _13267_, _08666_);
  and (_13682_, _13263_, _08665_);
  or (_13683_, _13682_, _13681_);
  and (_13684_, _13683_, _08800_);
  and (_13685_, _13287_, _08666_);
  and (_13686_, _13283_, _08665_);
  or (_13687_, _13686_, _13685_);
  and (_13688_, _13687_, _08837_);
  and (_13689_, _13277_, _08666_);
  and (_13691_, _13273_, _08665_);
  or (_13692_, _13691_, _13689_);
  and (_13694_, _13692_, _08842_);
  or (_13695_, _13694_, _13688_);
  or (_13696_, _13695_, _13684_);
  nor (_13697_, _13696_, _13680_);
  nor (_13698_, _13697_, _08828_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [26], _13698_, _13676_);
  and (_13699_, _08828_, word_in[27]);
  and (_13700_, _13313_, _08666_);
  and (_13701_, _13309_, _08665_);
  or (_13702_, _13701_, _13700_);
  and (_13703_, _13702_, _08800_);
  and (_13704_, _13344_, _08666_);
  and (_13705_, _13340_, _08665_);
  or (_13706_, _13705_, _13704_);
  and (_13707_, _13706_, _08814_);
  and (_13708_, _13333_, _08666_);
  and (_13709_, _13329_, _08665_);
  or (_13710_, _13709_, _13708_);
  and (_13711_, _13710_, _08837_);
  and (_13712_, _13323_, _08666_);
  and (_13713_, _13319_, _08665_);
  or (_13715_, _13713_, _13712_);
  and (_13716_, _13715_, _08842_);
  or (_13717_, _13716_, _13711_);
  or (_13718_, _13717_, _13707_);
  nor (_13719_, _13718_, _13703_);
  nor (_13720_, _13719_, _08828_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [27], _13720_, _13699_);
  and (_13722_, _08828_, word_in[28]);
  and (_13723_, _13359_, _08666_);
  and (_13724_, _13355_, _08665_);
  or (_13725_, _13724_, _13723_);
  and (_13726_, _13725_, _08800_);
  and (_13728_, _13370_, _08666_);
  and (_13729_, _13366_, _08665_);
  or (_13730_, _13729_, _13728_);
  and (_13731_, _13730_, _08814_);
  and (_13732_, _13380_, _08666_);
  and (_13733_, _13376_, _08665_);
  or (_13734_, _13733_, _13732_);
  and (_13735_, _13734_, _08837_);
  and (_13736_, _13392_, _08666_);
  and (_13737_, _13388_, _08665_);
  or (_13738_, _13737_, _13736_);
  and (_13740_, _13738_, _08842_);
  or (_13741_, _13740_, _13735_);
  or (_13743_, _13741_, _13731_);
  nor (_13744_, _13743_, _13726_);
  nor (_13746_, _13744_, _08828_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [28], _13746_, _13722_);
  and (_13748_, _08828_, word_in[29]);
  and (_13749_, _13406_, _08666_);
  and (_13750_, _13402_, _08665_);
  or (_13751_, _13750_, _13749_);
  and (_13752_, _13751_, _08800_);
  and (_13753_, _13416_, _08666_);
  and (_13755_, _13412_, _08665_);
  or (_13756_, _13755_, _13753_);
  and (_13757_, _13756_, _08814_);
  and (_13758_, _13427_, _08666_);
  and (_13759_, _13423_, _08665_);
  or (_13760_, _13759_, _13758_);
  and (_13761_, _13760_, _08837_);
  and (_13762_, _13438_, _08666_);
  and (_13763_, _13434_, _08665_);
  or (_13764_, _13763_, _13762_);
  and (_13765_, _13764_, _08842_);
  or (_13766_, _13765_, _13761_);
  or (_13767_, _13766_, _13757_);
  nor (_13768_, _13767_, _13752_);
  nor (_13769_, _13768_, _08828_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [29], _13769_, _13748_);
  and (_13770_, _08828_, word_in[30]);
  and (_13771_, _13482_, _08666_);
  and (_13772_, _13478_, _08665_);
  or (_13773_, _13772_, _13771_);
  and (_13774_, _13773_, _08814_);
  and (_13775_, _13452_, _08666_);
  and (_13776_, _13448_, _08665_);
  or (_13777_, _13776_, _13775_);
  and (_13778_, _13777_, _08800_);
  and (_13779_, _13472_, _08666_);
  and (_13780_, _13468_, _08665_);
  or (_13781_, _13780_, _13779_);
  and (_13782_, _13781_, _08837_);
  and (_13784_, _13462_, _08666_);
  and (_13785_, _13458_, _08665_);
  or (_13786_, _13785_, _13784_);
  and (_13787_, _13786_, _08842_);
  or (_13788_, _13787_, _13782_);
  or (_13789_, _13788_, _13778_);
  nor (_13790_, _13789_, _13774_);
  nor (_13791_, _13790_, _08828_);
  or (\oc8051_symbolic_cxrom1.cxrom_data_out [30], _13791_, _13770_);
  and (_11141_, _07987_, _06444_);
  and (_11154_, _09095_, _06444_);
  and (_11159_, _07927_, _06444_);
  nor (_13792_, _07602_, _07606_);
  and (_13793_, _07602_, _07606_);
  or (_13794_, _13793_, _13792_);
  and (_11176_, _13794_, _06444_);
  and (_11198_, _08097_, _06444_);
  and (_11214_, _08205_, _06444_);
  and (_11219_, _09196_, _06444_);
  and (_11222_, _09275_, _06444_);
  and (_11239_, _08284_, _06444_);
  and (_11248_, _07635_, _06444_);
  and (_11252_, _07628_, _06444_);
  and (_11298_, _08163_, _06444_);
  and (_11304_, _08246_, _06444_);
  and (_11308_, _08332_, _06444_);
  and (_13795_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  not (_13796_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_13797_, _08064_, _13796_);
  or (_13798_, _13797_, _13795_);
  and (_11397_, _13798_, _06444_);
  or (_13799_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  nand (_13800_, _07432_, _11718_);
  and (_13801_, _13800_, _06444_);
  and (_11462_, _13801_, _13799_);
  and (_13802_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [20]);
  and (_13803_, _12223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  or (_13804_, _13803_, _13802_);
  and (_11506_, _13804_, _06444_);
  and (_13806_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [23]);
  nor (_13807_, _07432_, _11016_);
  or (_13808_, _13807_, _13806_);
  and (_11748_, _13808_, _06444_);
  or (_13809_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  nand (_13810_, _07432_, _11194_);
  and (_13811_, _13810_, _06444_);
  and (_11752_, _13811_, _13809_);
  or (_13812_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  nand (_13813_, _07432_, _12171_);
  and (_13814_, _13813_, _06444_);
  and (_11768_, _13814_, _13812_);
  or (_13815_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  nand (_13816_, _07432_, _09662_);
  and (_13817_, _13816_, _06444_);
  and (_11783_, _13817_, _13815_);
  nand (_13818_, _11589_, _10112_);
  or (_13819_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [2]);
  and (_13820_, _13819_, _06444_);
  and (_11806_, _13820_, _13818_);
  or (_13821_, _09339_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  or (_13822_, _09467_, _09373_);
  and (_11894_, _13822_, _13821_);
  and (_11898_, _07765_, _06444_);
  and (_11913_, _08278_, _06444_);
  nor (_11916_, _09092_, rst);
  nor (_13823_, _07190_, _06666_);
  and (_13824_, _07190_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [5]);
  or (_13825_, _13824_, _13823_);
  and (_11956_, _13825_, _06444_);
  nand (_13826_, _08474_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  or (_13827_, _08474_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3]);
  and (_13828_, _13827_, _13826_);
  and (_11985_, _13828_, _06443_);
  and (_13830_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [8]);
  nor (_13832_, _07432_, _12492_);
  or (_13833_, _13832_, _13830_);
  and (_11988_, _13833_, _06444_);
  and (_13835_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , \oc8051_top_1.oc8051_sfr1.pres_ow );
  and (_13836_, _13835_, _06295_);
  nor (_13837_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nor (_13838_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  and (_13840_, _13838_, _13837_);
  nor (_13841_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  nor (_13842_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  nor (_13843_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  and (_13845_, _13843_, _13842_);
  and (_13846_, _13845_, _13841_);
  and (_13847_, _13846_, _13840_);
  and (_13848_, _13847_, _13836_);
  not (_13849_, _13836_);
  nand (_13850_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_13851_, _13850_, _06298_);
  nor (_13852_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2]);
  nor (_13853_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0]);
  and (_13854_, _13853_, _13852_);
  not (_13855_, _13854_);
  nor (_13856_, _13855_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand (_13857_, _13856_, _13847_);
  nand (_13858_, _13855_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done );
  nand (_13859_, _13858_, _13857_);
  and (_13860_, _13859_, _06298_);
  or (_13861_, _13860_, _13851_);
  and (_13862_, _13861_, _13849_);
  or (_13863_, _13862_, _13848_);
  and (_11992_, _13863_, _06443_);
  and (_13864_, _06440_, _06382_);
  and (_13865_, _13864_, _06434_);
  not (_13866_, _06297_);
  or (_13867_, _13857_, _13866_);
  nand (_13868_, _13867_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans );
  nor (_13869_, _13868_, _13848_);
  or (_13870_, _13869_, _13865_);
  and (_12000_, _13870_, _06444_);
  not (_13871_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  and (_13872_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  not (_13873_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_13874_, _07382_, _13873_);
  not (_13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  nor (_13876_, _13875_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_13877_, _13876_, _13874_);
  nor (_13878_, _13877_, _13872_);
  nand (_13879_, _13878_, _13871_);
  nor (_13880_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nor (_13881_, _13880_, _13878_);
  nand (_13882_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr );
  nand (_13883_, _13882_, _13881_);
  and (_13884_, _13883_, _06444_);
  and (_12007_, _13884_, _13879_);
  and (_12010_, _13881_, _06444_);
  and (_13885_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [7]);
  not (_13886_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [7]);
  nor (_13887_, _07432_, _13886_);
  or (_13888_, _13887_, _13885_);
  and (_12027_, _13888_, _06444_);
  and (_13889_, _07214_, _06933_);
  and (_13890_, _13889_, _07402_);
  or (_13891_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  and (_13892_, _13891_, _06444_);
  and (_13893_, _08978_, _06933_);
  nand (_13894_, _13893_, _06978_);
  and (_12036_, _13894_, _13892_);
  and (_13895_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [6]);
  not (_13896_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [6]);
  nor (_13898_, _07432_, _13896_);
  or (_13899_, _13898_, _13895_);
  and (_12049_, _13899_, _06444_);
  nor (_13900_, _06394_, _06336_);
  and (_13901_, _07401_, _06676_);
  and (_13902_, _13901_, _13900_);
  and (_13903_, _13902_, _06933_);
  nand (_13904_, _13903_, _06930_);
  or (_13905_, _13903_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_13906_, _06945_, _06382_);
  not (_13907_, _13906_);
  and (_13908_, _13907_, _13905_);
  and (_13909_, _13908_, _13904_);
  nor (_13910_, _13907_, _06978_);
  or (_13911_, _13910_, _13909_);
  and (_12053_, _13911_, _06444_);
  and (_12057_, _08078_, _06444_);
  and (_13912_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  not (_13913_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_13914_, _07382_, _13913_);
  or (_13915_, _13914_, _13876_);
  nor (_13916_, _13915_, _13912_);
  or (_13917_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  nand (_13918_, _13917_, _06444_);
  nor (_12083_, _13918_, _13916_);
  nor (_12089_, _07381_, rst);
  not (_13919_, rxd_i);
  nand (_13920_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _13919_);
  nand (_13921_, _13920_, _09353_);
  or (_13922_, _09354_, _09343_);
  and (_13923_, _13922_, _13921_);
  not (_13924_, _09340_);
  nand (_13926_, _09427_, _13924_);
  or (_13927_, _13926_, _13923_);
  and (_12133_, _13927_, _09373_);
  and (_13929_, _09678_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_13930_, _13929_, _09345_);
  and (_13931_, _09677_, _13930_);
  not (_13932_, _09344_);
  nor (_13933_, _13929_, _13932_);
  or (_13934_, _13933_, _09675_);
  and (_13935_, _13934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3]);
  or (_13936_, _13935_, _13931_);
  and (_12140_, _13936_, _06444_);
  and (_13937_, _09679_, _09346_);
  and (_13938_, _09677_, _13937_);
  nand (_13939_, _13938_, _13919_);
  or (_13940_, _13938_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  and (_13941_, _13940_, _06444_);
  and (_12143_, _13941_, _13939_);
  not (_13942_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r );
  nor (_13943_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _09355_);
  not (_13944_, _13943_);
  nor (_13945_, _06295_, _09339_);
  and (_13946_, _13945_, _13944_);
  and (_13947_, _13946_, _13932_);
  nor (_13948_, _13947_, _13942_);
  and (_13949_, _13947_, rxd_i);
  or (_13950_, _13949_, rst);
  or (_12153_, _13950_, _13948_);
  or (_13951_, _09351_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0]);
  or (_13952_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_13953_, _13952_, _06295_);
  or (_13954_, _13953_, _09344_);
  nand (_13955_, _13954_, _13951_);
  nand (_12159_, _13955_, _09373_);
  and (_13956_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_13957_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [4]);
  and (_13958_, _13957_, _09332_);
  and (_13959_, _07425_, _07359_);
  or (_13960_, _13959_, _13958_);
  or (_13961_, _13960_, _13956_);
  and (_12259_, _13961_, _06444_);
  nand (_13962_, _07613_, _07602_);
  or (_13963_, _07602_, \oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1]);
  and (_13964_, _13963_, _06444_);
  and (_12304_, _13964_, _13962_);
  and (_12317_, _08990_, _06444_);
  and (_13967_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [11]);
  not (_13968_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [11]);
  nor (_13969_, _07432_, _13968_);
  or (_13970_, _13969_, _13967_);
  and (_12334_, _13970_, _06444_);
  or (_13971_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  nand (_13972_, _07432_, _11838_);
  and (_13973_, _13972_, _06444_);
  and (_12341_, _13973_, _13971_);
  nand (_13975_, _12829_, _10494_);
  or (_13976_, _12829_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [6]);
  and (_13977_, _13976_, _06444_);
  and (_12351_, _13977_, _13975_);
  and (_13979_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [15]);
  not (_13980_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [15]);
  nor (_13982_, _07432_, _13980_);
  or (_13983_, _13982_, _13979_);
  and (_12356_, _13983_, _06444_);
  and (_13984_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [14]);
  not (_13985_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [14]);
  nor (_13986_, _07432_, _13985_);
  or (_13987_, _13986_, _13984_);
  and (_12375_, _13987_, _06444_);
  and (_13989_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [13]);
  not (_13990_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [13]);
  nor (_13992_, _07432_, _13990_);
  or (_13993_, _13992_, _13989_);
  and (_12380_, _13993_, _06444_);
  and (_13994_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [12]);
  and (_13995_, _12223_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [12]);
  or (_13997_, _13995_, _13994_);
  and (_12407_, _13997_, _06444_);
  and (_13998_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [10]);
  not (_13999_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [10]);
  nor (_14001_, _07432_, _13999_);
  or (_14002_, _14001_, _13998_);
  and (_12409_, _14002_, _06444_);
  and (_14003_, _07425_, _07378_);
  and (_14004_, _07153_, _07271_);
  or (_14005_, _14004_, _07420_);
  and (_14006_, _14005_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [5]);
  or (_14007_, _14006_, _14003_);
  and (_12465_, _14007_, _06444_);
  and (_14008_, _07190_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [7]);
  nor (_14010_, _07190_, _06978_);
  or (_14011_, _14010_, _14008_);
  and (_12599_, _14011_, _06444_);
  nor (_14013_, _12830_, _06666_);
  not (_14014_, _07415_);
  or (_14015_, _12825_, _14014_);
  and (_14016_, _14015_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [5]);
  or (_14017_, _14016_, _14013_);
  and (_12642_, _14017_, _06444_);
  and (_14018_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [3]);
  nor (_14019_, _07300_, _07046_);
  or (_14020_, _14019_, _14018_);
  and (_12752_, _14020_, _06444_);
  and (_14022_, _07070_, _06448_);
  and (_14024_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [1]);
  or (_14025_, _14024_, _14022_);
  and (_12864_, _14025_, _06444_);
  and (_14027_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_12870_, _14027_, _09425_);
  and (_12889_, _06444_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  and (_14028_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_13011_, _14028_, _09418_);
  or (_14029_, _09431_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1]);
  or (_14030_, _14029_, _13932_);
  and (_14031_, _14030_, _09430_);
  or (_14033_, _14031_, rxd_i);
  and (_14034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], rxd_i);
  nor (_14035_, _14034_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  and (_14036_, _14035_, _09349_);
  and (_14038_, _14036_, _09344_);
  nor (_14039_, _14038_, _09360_);
  and (_14041_, _14039_, _14033_);
  or (_14042_, _14041_, _09339_);
  nor (_14043_, _09351_, _09339_);
  or (_14044_, _14043_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  and (_14045_, _14044_, _06444_);
  and (_13023_, _14045_, _14042_);
  and (_14046_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [3]);
  nor (_14048_, _07432_, _12452_);
  or (_14049_, _14048_, _14046_);
  and (_13038_, _14049_, _06444_);
  and (_13046_, _06444_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  and (_13050_, _07586_, _06444_);
  and (_14050_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [2]);
  not (_14051_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [2]);
  nor (_14052_, _07432_, _14051_);
  or (_14053_, _14052_, _14050_);
  and (_13078_, _14053_, _06444_);
  and (_14054_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [1]);
  not (_14056_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [1]);
  nor (_14057_, _07432_, _14056_);
  or (_14058_, _14057_, _14054_);
  and (_13108_, _14058_, _06444_);
  and (_14059_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_old [0]);
  not (_14060_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [0]);
  nor (_14061_, _07432_, _14060_);
  or (_14062_, _14061_, _14059_);
  and (_13138_, _14062_, _06444_);
  nor (_14063_, _11589_, _09146_);
  and (_14064_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  or (_14065_, _14064_, _14063_);
  or (_14066_, _14065_, _07158_);
  or (_14067_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [2]);
  and (_14068_, _14067_, _06444_);
  and (_13148_, _14068_, _14066_);
  and (_14069_, _07154_, _06439_);
  not (_14070_, _14069_);
  and (_14071_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [2]);
  nor (_14072_, _14070_, _11589_);
  or (_14074_, _14072_, _14071_);
  and (_13161_, _14074_, _06444_);
  nand (_14075_, _10112_, _07188_);
  or (_14076_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [4]);
  and (_14077_, _14076_, _06444_);
  and (_13300_, _14077_, _14075_);
  nor (_14078_, _11919_, _11703_);
  and (_14079_, _11861_, _11809_);
  and (_14080_, _14079_, _14078_);
  and (_14081_, _11669_, _11741_);
  nor (_14082_, _11630_, _11782_);
  and (_14083_, _14082_, _14081_);
  and (_14084_, _14083_, _14080_);
  not (_14085_, _11703_);
  and (_14086_, _11919_, _14085_);
  and (_14087_, _14079_, _14086_);
  and (_14088_, _14083_, _14087_);
  nor (_14089_, _14088_, _14084_);
  not (_14090_, _11861_);
  nor (_14091_, _14090_, _11809_);
  and (_14092_, _14091_, _14086_);
  and (_14093_, _14083_, _14092_);
  and (_14094_, _14090_, _11809_);
  and (_14095_, _14094_, _14078_);
  and (_14096_, _14083_, _14095_);
  nor (_14097_, _14096_, _14093_);
  and (_14098_, _14097_, _14089_);
  not (_14099_, _11782_);
  nor (_14100_, _11630_, _14099_);
  and (_14101_, _14081_, _14100_);
  and (_14102_, _14087_, _14101_);
  nor (_14103_, _11861_, _11809_);
  and (_14104_, _14086_, _14103_);
  and (_14105_, _14083_, _14104_);
  nor (_14106_, _14105_, _14102_);
  not (_14107_, _11741_);
  and (_14108_, _14100_, _14107_);
  and (_14109_, _14108_, _11669_);
  and (_14110_, _14109_, _14087_);
  not (_14111_, _11669_);
  and (_14112_, _14108_, _14111_);
  not (_14113_, _11919_);
  and (_14114_, _14103_, _14113_);
  and (_14115_, _14114_, _11703_);
  and (_14116_, _14115_, _14112_);
  nor (_14117_, _14116_, _14110_);
  and (_14118_, _14117_, _14106_);
  and (_14119_, _14118_, _14098_);
  and (_14120_, _14104_, _14101_);
  and (_14121_, _14094_, _14086_);
  and (_14122_, _14121_, _14101_);
  nor (_14123_, _14122_, _14120_);
  and (_14124_, _14095_, _14101_);
  and (_14125_, _14092_, _14101_);
  nor (_14126_, _14125_, _14124_);
  and (_14127_, _14126_, _14123_);
  and (_14128_, _14100_, _11741_);
  and (_14129_, _14128_, _14111_);
  and (_14130_, _14129_, _14121_);
  and (_14131_, _14129_, _14087_);
  nor (_14132_, _14131_, _14130_);
  and (_14133_, _14080_, _14101_);
  and (_14134_, _14115_, _14101_);
  nor (_14135_, _14134_, _14133_);
  and (_14136_, _14135_, _14132_);
  and (_14137_, _14136_, _14127_);
  and (_14138_, _14137_, _14119_);
  and (_14139_, _11919_, _11703_);
  and (_14140_, _14139_, _14079_);
  and (_14141_, _14140_, _14111_);
  and (_14142_, _14082_, _11741_);
  and (_14143_, _14142_, _14141_);
  and (_14144_, _14082_, _14107_);
  and (_14145_, _14140_, _11669_);
  and (_14146_, _14145_, _14144_);
  nor (_14147_, _14146_, _14143_);
  nand (_14148_, _14140_, _14100_);
  and (_14149_, _14139_, _14101_);
  and (_14150_, _14149_, _14091_);
  and (_14151_, _14139_, _14103_);
  and (_14152_, _14151_, _14101_);
  nor (_14153_, _14152_, _14150_);
  and (_14154_, _14144_, _14141_);
  and (_14155_, _14139_, _14094_);
  and (_14156_, _14155_, _14101_);
  nor (_14157_, _14156_, _14154_);
  and (_14158_, _14157_, _14153_);
  and (_14159_, _14158_, _14148_);
  and (_14160_, _14159_, _14147_);
  nand (_14161_, _14160_, _14138_);
  and (_14162_, _14143_, _12008_);
  and (_14163_, _14149_, _14103_);
  and (_14164_, _14163_, _08975_);
  nor (_14165_, _14164_, _14162_);
  nor (_14166_, _14165_, \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_14167_, _14166_);
  not (_14168_, _06676_);
  nor (_14169_, _14114_, _14168_);
  nand (_14170_, _14169_, _11789_);
  nand (_14171_, _14146_, _08025_);
  and (_14172_, _14171_, _14170_);
  and (_14173_, _14172_, _11928_);
  and (_14174_, _14173_, _14167_);
  nand (_14175_, _14174_, _14161_);
  and (_14176_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  and (_14178_, _14150_, _08975_);
  and (_14179_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  and (_14181_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_14183_, _14181_, _14179_);
  and (_14184_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_14185_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_14186_, _14185_, _14184_);
  or (_14187_, _14186_, _14183_);
  and (_14188_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_14189_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_14190_, _14189_, _14188_);
  and (_14191_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_14192_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  or (_14193_, _14192_, _14191_);
  or (_14194_, _14193_, _14190_);
  or (_14195_, _14194_, _14187_);
  and (_14196_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_14198_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  or (_14199_, _14198_, _14196_);
  and (_14200_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_14201_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  or (_14202_, _14201_, _14200_);
  or (_14203_, _14202_, _14199_);
  and (_14204_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  and (_14205_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  or (_14206_, _14205_, _14204_);
  and (_14208_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_14209_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  or (_14210_, _14209_, _14208_);
  or (_14211_, _14210_, _14206_);
  or (_14212_, _14211_, _14203_);
  or (_14213_, _14212_, _14195_);
  and (_14214_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  and (_14215_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_14216_, _14215_, _14214_);
  and (_14217_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_14218_, _14156_, _11775_);
  or (_14219_, _14218_, _14217_);
  and (_14220_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  and (_14221_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  or (_14222_, _14221_, _14220_);
  or (_14223_, _14222_, _14219_);
  and (_14224_, _14140_, _14101_);
  and (_14225_, _11437_, _11965_);
  or (_14226_, _14225_, _11513_);
  nor (_14227_, _14226_, _11512_);
  and (_14228_, _11528_, _11374_);
  not (_14229_, _14228_);
  nor (_14230_, _11536_, _11428_);
  and (_14231_, _14230_, _14229_);
  and (_14232_, _11493_, _11430_);
  nor (_14233_, _14232_, _11524_);
  and (_14234_, _11519_, _11374_);
  nor (_14235_, _14234_, _11503_);
  and (_14236_, _14235_, _14233_);
  nor (_14237_, _11352_, _11372_);
  and (_14238_, _14237_, _11364_);
  and (_14239_, _11976_, _11412_);
  and (_14240_, _11407_, _11406_);
  or (_14241_, _14240_, _14239_);
  nor (_14242_, _14241_, _14238_);
  and (_14243_, _14242_, _14236_);
  and (_14244_, _14243_, _14231_);
  and (_14245_, _14244_, _11499_);
  and (_14246_, _14245_, _14227_);
  nor (_14247_, _14246_, _11343_);
  or (_14248_, _14247_, p0_in[6]);
  not (_14249_, _14247_);
  or (_14250_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_14251_, _14250_, _14248_);
  and (_14252_, _14251_, _14224_);
  and (_14253_, _14129_, _14140_);
  or (_14254_, _14247_, p1_in[6]);
  or (_14255_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_14256_, _14255_, _14254_);
  and (_14258_, _14256_, _14253_);
  or (_14259_, _14258_, _14252_);
  and (_14260_, _14112_, _14140_);
  or (_14261_, _14247_, p3_in[6]);
  or (_14262_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_14263_, _14262_, _14261_);
  and (_14264_, _14263_, _14260_);
  and (_14265_, _14109_, _14140_);
  or (_14266_, _14247_, p2_in[6]);
  or (_14267_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_14268_, _14267_, _14266_);
  and (_14269_, _14268_, _14265_);
  or (_14270_, _14269_, _14264_);
  or (_14271_, _14270_, _14259_);
  or (_14272_, _14271_, _14223_);
  or (_14273_, _14272_, _14216_);
  or (_14274_, _14273_, _14213_);
  and (_14275_, _14274_, _14174_);
  or (_14276_, _14275_, _14178_);
  or (_14277_, _14276_, _14176_);
  nand (_14278_, _14178_, _09045_);
  and (_14279_, _14278_, _06444_);
  and (_13364_, _14279_, _14277_);
  and (_14280_, _07189_, _07070_);
  and (_14281_, _10497_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [1]);
  or (_14282_, _14281_, _14280_);
  and (_13387_, _14282_, _06444_);
  and (_13422_, _07757_, _06444_);
  and (_14283_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  and (_14284_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_14285_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_14286_, _14285_, _14284_);
  and (_14287_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  and (_14288_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_14289_, _14288_, _14287_);
  or (_14290_, _14289_, _14286_);
  and (_14291_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_14292_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or (_14293_, _14292_, _14291_);
  and (_14294_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_14296_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  or (_14297_, _14296_, _14294_);
  or (_14298_, _14297_, _14293_);
  or (_14299_, _14298_, _14290_);
  and (_14300_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_14301_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  or (_14302_, _14301_, _14300_);
  and (_14303_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_14304_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_14305_, _14304_, _14303_);
  or (_14306_, _14305_, _14302_);
  and (_14307_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_14308_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_14309_, _14308_, _14307_);
  and (_14310_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  and (_14311_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  or (_14312_, _14311_, _14310_);
  or (_14313_, _14312_, _14309_);
  or (_14314_, _14313_, _14306_);
  or (_14315_, _14314_, _14299_);
  and (_14316_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_14317_, _14156_, _11700_);
  or (_14318_, _14317_, _14316_);
  and (_14319_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  and (_14320_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  or (_14321_, _14320_, _14319_);
  or (_14322_, _14321_, _14318_);
  or (_14323_, _14247_, p0_in[3]);
  or (_14324_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_14325_, _14324_, _14323_);
  and (_14326_, _14325_, _14224_);
  or (_14327_, _14247_, p1_in[3]);
  or (_14328_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_14329_, _14328_, _14327_);
  and (_14330_, _14329_, _14253_);
  or (_14331_, _14330_, _14326_);
  or (_14332_, _14247_, p2_in[3]);
  or (_14333_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_14334_, _14333_, _14332_);
  and (_14335_, _14334_, _14265_);
  or (_14336_, _14247_, p3_in[3]);
  or (_14337_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_14338_, _14337_, _14336_);
  and (_14339_, _14338_, _14260_);
  or (_14340_, _14339_, _14335_);
  or (_14341_, _14340_, _14331_);
  or (_14342_, _14341_, _14322_);
  and (_14343_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  and (_14344_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  or (_14345_, _14344_, _14343_);
  or (_14347_, _14345_, _14342_);
  or (_14349_, _14347_, _14315_);
  and (_14350_, _14349_, _14174_);
  or (_14351_, _14350_, _14178_);
  or (_14352_, _14351_, _14283_);
  not (_14353_, _14178_);
  or (_14354_, _14353_, _08308_);
  and (_14355_, _14354_, _06444_);
  and (_13519_, _14355_, _14352_);
  and (_14357_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  and (_14358_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_14359_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_14360_, _14359_, _14358_);
  and (_14361_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_14362_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  or (_14363_, _14362_, _14361_);
  or (_14364_, _14363_, _14360_);
  and (_14366_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_14367_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_14368_, _14367_, _14366_);
  and (_14369_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  and (_14370_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_14371_, _14370_, _14369_);
  or (_14372_, _14371_, _14368_);
  or (_14373_, _14372_, _14364_);
  and (_14374_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_14375_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_14376_, _14375_, _14374_);
  and (_14377_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_14378_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  or (_14379_, _14378_, _14377_);
  or (_14380_, _14379_, _14376_);
  and (_14381_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  and (_14382_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_14383_, _14382_, _14381_);
  and (_14384_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_14385_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  or (_14386_, _14385_, _14384_);
  or (_14387_, _14386_, _14383_);
  or (_14388_, _14387_, _14380_);
  or (_14389_, _14388_, _14373_);
  and (_14390_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  and (_14391_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_14393_, _14391_, _14390_);
  and (_14394_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  and (_14395_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  or (_14396_, _14395_, _14394_);
  and (_14397_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_14398_, _14156_, _11914_);
  or (_14399_, _14398_, _14397_);
  or (_14400_, _14399_, _14396_);
  or (_14401_, _14247_, p2_in[2]);
  or (_14402_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_14403_, _14402_, _14401_);
  and (_14404_, _14403_, _14265_);
  or (_14405_, _14247_, p3_in[2]);
  or (_14406_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_14407_, _14406_, _14405_);
  and (_14408_, _14407_, _14260_);
  or (_14409_, _14408_, _14404_);
  or (_14410_, _14247_, p0_in[2]);
  or (_14411_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_14412_, _14411_, _14410_);
  and (_14413_, _14412_, _14224_);
  or (_14414_, _14247_, p1_in[2]);
  or (_14415_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_14417_, _14415_, _14414_);
  and (_14418_, _14417_, _14253_);
  or (_14419_, _14418_, _14413_);
  or (_14420_, _14419_, _14409_);
  or (_14421_, _14420_, _14400_);
  or (_14422_, _14421_, _14393_);
  or (_14423_, _14422_, _14389_);
  and (_14424_, _14423_, _14174_);
  or (_14425_, _14424_, _14178_);
  or (_14426_, _14425_, _14357_);
  nand (_14427_, _14178_, _09138_);
  and (_14428_, _14427_, _06444_);
  and (_13525_, _14428_, _14426_);
  and (_14429_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  and (_14430_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_14431_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_14432_, _14431_, _14430_);
  and (_14433_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_14434_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_14435_, _14434_, _14433_);
  or (_14436_, _14435_, _14432_);
  and (_14437_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  and (_14438_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_14439_, _14438_, _14437_);
  and (_14440_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_14441_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_14442_, _14441_, _14440_);
  or (_14443_, _14442_, _14439_);
  or (_14444_, _14443_, _14436_);
  and (_14445_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_14446_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_14447_, _14446_, _14445_);
  and (_14448_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_14449_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  or (_14450_, _14449_, _14448_);
  or (_14451_, _14450_, _14447_);
  and (_14452_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  and (_14453_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_14454_, _14453_, _14452_);
  and (_14455_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_14456_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  or (_14457_, _14456_, _14455_);
  or (_14458_, _14457_, _14454_);
  or (_14459_, _14458_, _14451_);
  or (_14460_, _14459_, _14444_);
  and (_14461_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_14462_, _14156_, _11803_);
  or (_14463_, _14462_, _14461_);
  and (_14464_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  and (_14465_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  or (_14466_, _14465_, _14464_);
  or (_14467_, _14466_, _14463_);
  or (_14468_, _14247_, p3_in[1]);
  or (_14469_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_14470_, _14469_, _14468_);
  and (_14471_, _14470_, _14260_);
  or (_14472_, _14247_, p2_in[1]);
  or (_14473_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_14474_, _14473_, _14472_);
  and (_14475_, _14474_, _14265_);
  or (_14476_, _14475_, _14471_);
  or (_14477_, _14247_, p0_in[1]);
  or (_14478_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_14479_, _14478_, _14477_);
  and (_14480_, _14479_, _14224_);
  or (_14481_, _14247_, p1_in[1]);
  or (_14482_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_14483_, _14482_, _14481_);
  and (_14484_, _14483_, _14253_);
  or (_14485_, _14484_, _14480_);
  or (_14486_, _14485_, _14476_);
  or (_14487_, _14486_, _14467_);
  and (_14488_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_14489_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_14490_, _14489_, _14488_);
  or (_14491_, _14490_, _14487_);
  or (_14492_, _14491_, _14460_);
  and (_14493_, _14492_, _14174_);
  or (_14494_, _14493_, _14178_);
  or (_14495_, _14494_, _14429_);
  nor (_14496_, _14178_, rst);
  and (_14497_, _07959_, _06444_);
  or (_14498_, _14497_, _14496_);
  and (_13548_, _14498_, _14495_);
  nor (_14499_, _07300_, _06449_);
  and (_14500_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [3]);
  or (_14501_, _14500_, _14499_);
  and (_13551_, _14501_, _06444_);
  or (_14502_, _11137_, _08980_);
  or (_14503_, _08982_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_14504_, _14503_, _06444_);
  and (_13589_, _14504_, _14502_);
  and (_14505_, _11137_, _09157_);
  and (_14506_, _09158_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_14507_, _14506_, _08975_);
  or (_14508_, _14507_, _14505_);
  or (_14509_, _11177_, _09208_);
  and (_14510_, _14509_, _06444_);
  and (_13596_, _14510_, _14508_);
  and (_14511_, _07402_, _06434_);
  and (_14512_, _14511_, _06440_);
  nand (_14513_, _14512_, _11589_);
  or (_14514_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_14516_, _14514_, _06444_);
  and (_13634_, _14516_, _14513_);
  nand (_14517_, _14512_, _07069_);
  or (_14518_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_14519_, _14518_, _06444_);
  and (_13637_, _14519_, _14517_);
  or (_14520_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  and (_14521_, _14520_, _06444_);
  nand (_14523_, _14512_, _07300_);
  and (_13661_, _14523_, _14521_);
  or (_14525_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  and (_14526_, _14525_, _06444_);
  nand (_14527_, _14512_, _07188_);
  and (_13665_, _14527_, _14526_);
  not (_14528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nor (_14529_, _14512_, _14528_);
  and (_14530_, _14512_, _09527_);
  or (_14531_, _14530_, _14529_);
  and (_13675_, _14531_, _06444_);
  and (_14532_, _07402_, _06984_);
  nand (_14533_, _14532_, _06666_);
  and (_14534_, _14528_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_14535_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_14536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _14535_);
  or (_14537_, _14536_, _14534_);
  not (_14538_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_14539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_14540_, _14539_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_14541_, _14540_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_14542_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_14543_, _14542_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_14545_, t0_i);
  and (_14546_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  and (_14547_, _14546_, _14545_);
  or (_14548_, _14547_, _14543_);
  and (_14549_, _14548_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_14550_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_14551_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_14552_, _14551_, _14550_);
  and (_14553_, _14552_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_14554_, _14553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  and (_00001_, _14554_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00002_, _00001_, _14549_);
  and (_00003_, _00002_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_00004_, _00003_, _14541_);
  and (_00005_, _00004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_00006_, _00005_, _14535_);
  nor (_00007_, _00006_, _14538_);
  and (_00008_, _00006_, _14538_);
  or (_00009_, _00008_, _00007_);
  and (_00010_, _00009_, _14537_);
  and (_00011_, \oc8051_top_1.oc8051_sfr1.pres_ow , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_00012_, _00011_, _14541_);
  and (_00013_, _00012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_00014_, _00013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00015_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00016_, _00013_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  not (_00017_, _00016_);
  and (_00018_, _00017_, _00015_);
  and (_00019_, _00018_, _00014_);
  and (_00020_, _14549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  and (_00021_, _00020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  and (_00022_, _00021_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  and (_00023_, _00022_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  and (_00024_, _00023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_00025_, _00024_, _14541_);
  and (_00026_, _00025_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_00027_, _00026_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_00028_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  not (_00029_, _00028_);
  and (_00030_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_00031_, _00030_, _14541_);
  and (_00032_, _00031_, _00024_);
  nor (_00033_, _00032_, _00029_);
  and (_00034_, _00033_, _00027_);
  or (_00035_, _00034_, _00019_);
  or (_00036_, _00035_, _00010_);
  or (_00037_, _00036_, _14532_);
  and (_00039_, _09483_, _07402_);
  not (_00040_, _00039_);
  and (_00041_, _00040_, _00037_);
  and (_00042_, _00041_, _14533_);
  and (_00043_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  or (_00044_, _00043_, _00042_);
  and (_13690_, _00044_, _06444_);
  nand (_00045_, _14532_, _10494_);
  and (_00046_, _00032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_00047_, _00032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_00048_, _00047_, _00028_);
  nor (_00049_, _00048_, _00046_);
  and (_00050_, _00031_, _00003_);
  or (_00051_, _00050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00052_, _00050_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  not (_00053_, _00052_);
  and (_00054_, _00053_, _14536_);
  and (_00055_, _00054_, _00051_);
  and (_00057_, _00016_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  or (_00058_, _00057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  nand (_00059_, _00057_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00060_, _00059_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00062_, _00060_, _00058_);
  or (_00063_, _00062_, _00055_);
  or (_00065_, _00063_, _00049_);
  or (_00067_, _00065_, _14532_);
  and (_00068_, _00067_, _00040_);
  and (_00069_, _00068_, _00045_);
  and (_00070_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  or (_00071_, _00070_, _00069_);
  and (_13693_, _00071_, _06444_);
  nand (_00072_, _14532_, _09526_);
  or (_00073_, _00024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_00074_, _00024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_00075_, _00074_, _00029_);
  and (_00076_, _00075_, _00073_);
  not (_00077_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_00078_, _00003_, _14535_);
  and (_00079_, _00078_, _00077_);
  nor (_00080_, _00078_, _00077_);
  or (_00081_, _00080_, _00079_);
  and (_00083_, _00081_, _14537_);
  and (_00084_, _00011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  or (_00086_, _00011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nand (_00087_, _00086_, _00015_);
  nor (_00089_, _00087_, _00084_);
  or (_00090_, _00089_, _00083_);
  or (_00091_, _00090_, _00076_);
  or (_00092_, _00091_, _14532_);
  and (_00093_, _00092_, _00072_);
  or (_00094_, _00093_, _00039_);
  nand (_00095_, _00039_, _00077_);
  and (_00096_, _00095_, _06444_);
  and (_13714_, _00096_, _00094_);
  nand (_00097_, _00039_, _10494_);
  or (_00098_, _00028_, _14532_);
  and (_00099_, _00098_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00100_, _00024_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_00101_, _00100_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  nor (_00102_, _00028_, _00002_);
  and (_00103_, _00102_, _00101_);
  and (_00104_, _14534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_00105_, _00104_, _00003_);
  nor (_00106_, _00105_, _00103_);
  nor (_00107_, _00106_, _14532_);
  or (_00108_, _00107_, _00099_);
  or (_00109_, _00108_, _00039_);
  and (_00110_, _00109_, _06444_);
  and (_13721_, _00110_, _00097_);
  nand (_00111_, _00039_, _06666_);
  and (_00112_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  and (_00113_, _00112_, _14549_);
  and (_00114_, _00113_, _14553_);
  and (_00115_, _14534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_00116_, _00115_, _00114_);
  nand (_00117_, _00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  nor (_00118_, _00028_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  nand (_00119_, _00118_, _00024_);
  and (_00120_, _00119_, _00117_);
  nor (_00121_, _00120_, _14532_);
  not (_00122_, _00024_);
  or (_00123_, _00098_, _00122_);
  and (_00124_, _00123_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_00125_, _00124_, _00121_);
  or (_00126_, _00125_, _00039_);
  and (_00127_, _00126_, _06444_);
  and (_13727_, _00127_, _00111_);
  nand (_00128_, _14532_, _11589_);
  and (_00129_, _00003_, _14539_);
  or (_00130_, _00129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nand (_00131_, _00129_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00132_, _00131_, _14536_);
  and (_00133_, _00132_, _00130_);
  not (_00134_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00135_, _14553_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_00136_, _14549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00137_, _00136_, _00135_);
  and (_00138_, _00137_, _00134_);
  nor (_00139_, _00137_, _00134_);
  or (_00140_, _00139_, _00138_);
  and (_00141_, _00140_, _00028_);
  and (_00142_, _00011_, _14539_);
  and (_00144_, _00142_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  nand (_00146_, _00144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_00148_, _00144_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  and (_00150_, _00148_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  and (_00152_, _00150_, _00146_);
  or (_00154_, _00152_, _00141_);
  or (_00155_, _00154_, _00133_);
  or (_00156_, _00155_, _14532_);
  and (_00157_, _00156_, _00040_);
  and (_00158_, _00157_, _00128_);
  and (_00159_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  or (_00160_, _00159_, _00158_);
  and (_13739_, _00160_, _06444_);
  nand (_00161_, _14532_, _07188_);
  nor (_00163_, _00025_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_00165_, _00163_, _00026_);
  and (_00167_, _00165_, _00028_);
  or (_00168_, _00004_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  not (_00170_, _00005_);
  and (_00171_, _00170_, _14536_);
  and (_00173_, _00171_, _00168_);
  and (_00174_, _14534_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_00175_, _00012_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  nor (_00176_, _00175_, _00013_);
  and (_00178_, _00176_, _00015_);
  or (_00179_, _00178_, _00174_);
  or (_00180_, _00179_, _00173_);
  or (_00181_, _00180_, _00167_);
  or (_00182_, _00181_, _14532_);
  and (_00183_, _00182_, _00040_);
  and (_00184_, _00183_, _00161_);
  and (_00185_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  or (_00186_, _00185_, _00184_);
  and (_13742_, _00186_, _06444_);
  nand (_00187_, _14532_, _07300_);
  and (_00188_, _00024_, _14540_);
  or (_00190_, _00188_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_00192_, _00025_, _00029_);
  and (_00193_, _00192_, _00190_);
  and (_00194_, _00078_, _14540_);
  or (_00195_, _00194_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_00196_, _00004_);
  or (_00197_, _00196_, _14534_);
  and (_00198_, _00197_, _14537_);
  and (_00199_, _00198_, _00195_);
  and (_00200_, _00011_, _14540_);
  or (_00201_, _00200_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  not (_00202_, _00012_);
  and (_00203_, _00015_, _00202_);
  and (_00204_, _00203_, _00201_);
  or (_00206_, _00204_, _00199_);
  or (_00207_, _00206_, _00193_);
  or (_00208_, _00207_, _14532_);
  and (_00209_, _00208_, _00040_);
  and (_00210_, _00209_, _00187_);
  and (_00212_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  or (_00213_, _00212_, _00210_);
  and (_13745_, _00213_, _06444_);
  not (_00214_, _00074_);
  nor (_00215_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  and (_00216_, _00214_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_00217_, _00216_, _00215_);
  and (_00218_, _00217_, _00028_);
  or (_00219_, _00084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_00220_, _00142_);
  and (_00221_, _00015_, _00220_);
  and (_00222_, _00221_, _00219_);
  and (_00223_, _00003_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_00224_, _00223_, _14535_);
  or (_00225_, _00224_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  not (_00226_, _00129_);
  and (_00227_, _00226_, _14536_);
  or (_00228_, _00227_, _14534_);
  and (_00229_, _00228_, _00225_);
  or (_00230_, _00229_, _00222_);
  or (_00231_, _00230_, _00218_);
  or (_00232_, _00231_, _14532_);
  nand (_00233_, _14532_, _07069_);
  and (_00234_, _00233_, _00040_);
  and (_00235_, _00234_, _00232_);
  and (_00236_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  or (_00237_, _00236_, _00235_);
  and (_13747_, _00237_, _06444_);
  nor (_00238_, _06430_, _06418_);
  and (_00240_, _00238_, _06406_);
  and (_00241_, _13902_, _00240_);
  nand (_00242_, _00241_, _06930_);
  or (_00243_, _00241_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  and (_00244_, _00243_, _13907_);
  and (_00245_, _00244_, _00242_);
  nor (_00246_, _13907_, _10494_);
  or (_00248_, _00246_, _00245_);
  and (_13754_, _00248_, _06444_);
  and (_00249_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [25]);
  and (_00250_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [25]);
  or (_00251_, _00250_, _00249_);
  and (_13783_, _00251_, _06444_);
  and (_00253_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [27]);
  and (_00254_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [27]);
  or (_00255_, _00254_, _00253_);
  and (_13805_, _00255_, _06444_);
  nor (_00257_, _00022_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  nor (_00258_, _00257_, _00023_);
  and (_00259_, _00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  nor (_00260_, _00259_, _00258_);
  nor (_00261_, _00260_, _14532_);
  and (_00262_, _14532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  or (_00263_, _00262_, _00261_);
  and (_00264_, _00263_, _00040_);
  nor (_00265_, _00040_, _07300_);
  or (_00266_, _00265_, _00264_);
  and (_13829_, _00266_, _06444_);
  nand (_00267_, _00039_, _07188_);
  nor (_00268_, _00023_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  nor (_00269_, _00268_, _00024_);
  and (_00270_, _00174_, _00003_);
  nor (_00271_, _00270_, _00269_);
  nor (_00273_, _00271_, _14532_);
  and (_00275_, _14532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  or (_00277_, _00275_, _00273_);
  or (_00279_, _00277_, _00039_);
  and (_00281_, _00279_, _06444_);
  and (_13831_, _00281_, _00267_);
  nor (_00283_, _00021_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  nor (_00284_, _00283_, _00022_);
  and (_00285_, _00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  nor (_00286_, _00285_, _00284_);
  nor (_00288_, _00286_, _14532_);
  and (_00289_, _14532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  or (_00290_, _00289_, _00288_);
  and (_00291_, _00290_, _00040_);
  nor (_00292_, _00040_, _11589_);
  or (_00293_, _00292_, _00291_);
  and (_13834_, _00293_, _06444_);
  or (_00294_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00296_, _00294_, _06444_);
  nand (_00297_, _14512_, _10494_);
  and (_13839_, _00297_, _00296_);
  or (_00298_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00300_, _00298_, _06444_);
  nand (_00301_, _14512_, _06666_);
  and (_13844_, _00301_, _00300_);
  and (_00302_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [26]);
  and (_00303_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [26]);
  or (_00304_, _00303_, _00302_);
  and (_13897_, _00304_, _06444_);
  nor (_00305_, _14549_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  nor (_00306_, _00305_, _00020_);
  and (_00307_, _00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  nor (_00308_, _00307_, _00306_);
  nor (_00309_, _00308_, _14532_);
  and (_00310_, _14532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or (_00311_, _00310_, _00309_);
  and (_00312_, _00311_, _00040_);
  and (_00313_, _00039_, _09527_);
  or (_00314_, _00313_, _00312_);
  and (_13925_, _00314_, _06444_);
  nor (_00315_, _00020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  nor (_00316_, _00315_, _00021_);
  and (_00317_, _00116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  nor (_00318_, _00317_, _00316_);
  nor (_00319_, _00318_, _14532_);
  and (_00320_, _14532_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  or (_00321_, _00320_, _00319_);
  and (_00322_, _00321_, _00040_);
  nor (_00323_, _00040_, _07069_);
  or (_00324_, _00323_, _00322_);
  and (_13928_, _00324_, _06444_);
  and (_00325_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  and (_00327_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [31]);
  or (_00328_, _00327_, _00325_);
  and (_13965_, _00328_, _06444_);
  nor (_00329_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , rst);
  and (_13966_, _00329_, \oc8051_top_1.oc8051_memory_interface1.int_ack_buff );
  and (_00330_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [24]);
  and (_00332_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [24]);
  or (_00333_, _00332_, _00330_);
  and (_13974_, _00333_, _06444_);
  and (_00334_, _07402_, _06988_);
  nand (_00335_, _00334_, _10494_);
  not (_00336_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_00337_, _00336_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  not (_00338_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00340_, _00338_, \oc8051_top_1.oc8051_sfr1.pres_ow );
  not (_00341_, t1_i);
  and (_00343_, _00341_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  and (_00344_, _00343_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff );
  or (_00346_, _00344_, _00340_);
  and (_00347_, _00346_, _00337_);
  and (_00348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00349_, _00348_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_00351_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00352_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_00353_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  and (_00354_, _00353_, _00352_);
  and (_00355_, _00354_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00356_, _00355_, _00351_);
  and (_00357_, _00356_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00358_, _00357_, _00349_);
  and (_00359_, _00358_, _00347_);
  or (_00360_, _00359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00361_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_00362_, _00361_);
  and (_00363_, _00359_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00364_, _00363_, _00362_);
  not (_00365_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00366_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _00365_);
  and (_00367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  and (_00369_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_00370_, _00369_, _00367_);
  and (_00372_, _00370_, _00354_);
  and (_00373_, _00372_, _00351_);
  and (_00374_, _00373_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00375_, _00374_, _00347_);
  and (_00376_, _00375_, _00349_);
  nand (_00377_, _00376_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_00378_, _00377_, _00366_);
  or (_00379_, _00378_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  and (_00380_, _00367_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_00381_, _00366_, _00380_);
  or (_00382_, _00381_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  and (_00383_, _00382_, _00379_);
  or (_00384_, _00383_, _00364_);
  and (_00385_, _00384_, _00360_);
  or (_00386_, _00385_, _00334_);
  and (_00387_, _09478_, _07402_);
  not (_00388_, _00387_);
  and (_00389_, _00388_, _00386_);
  and (_00390_, _00389_, _00335_);
  and (_00391_, _00387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_00392_, _00391_, _00390_);
  and (_13978_, _00392_, _06444_);
  nand (_00393_, _00334_, _06666_);
  not (_00394_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  not (_00395_, _00366_);
  nor (_00396_, _00375_, _00395_);
  not (_00397_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00398_, _00361_, _00397_);
  and (_00399_, _00355_, _00347_);
  and (_00400_, _00399_, _00351_);
  nor (_00401_, _00362_, _00400_);
  nor (_00402_, _00401_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  not (_00403_, _00402_);
  nor (_00404_, _00403_, _00398_);
  not (_00405_, _00404_);
  or (_00406_, _00405_, _00396_);
  not (_00407_, _00406_);
  and (_00408_, _00407_, _00348_);
  nor (_00409_, _00408_, _00394_);
  and (_00410_, _00408_, _00394_);
  or (_00411_, _00410_, _00409_);
  or (_00412_, _00411_, _00334_);
  and (_00413_, _00412_, _00388_);
  and (_00414_, _00413_, _00393_);
  and (_00415_, _00387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  or (_00416_, _00415_, _00414_);
  and (_13981_, _00416_, _06444_);
  nand (_00417_, _00334_, _07300_);
  nor (_00418_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  and (_00419_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_00420_, _00419_, _00418_);
  or (_00421_, _00420_, _00334_);
  and (_00422_, _00421_, _00388_);
  and (_00423_, _00422_, _00417_);
  and (_00424_, _00387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  or (_00425_, _00424_, _00423_);
  and (_13988_, _00425_, _06444_);
  nand (_00426_, _00334_, _07188_);
  not (_00427_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  and (_00428_, _00407_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_00429_, _00428_, _00427_);
  and (_00430_, _00428_, _00427_);
  or (_00431_, _00430_, _00429_);
  or (_00432_, _00431_, _00334_);
  and (_00433_, _00432_, _00426_);
  or (_00435_, _00433_, _00387_);
  nand (_00436_, _00387_, _00427_);
  and (_00437_, _00436_, _06444_);
  and (_13991_, _00437_, _00435_);
  nand (_00438_, _00334_, _07069_);
  and (_00439_, _00399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00440_, _00439_, _00380_);
  nor (_00441_, _00440_, _00395_);
  or (_00442_, _00441_, _00403_);
  and (_00443_, _00442_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00444_, _00439_, _00401_);
  nor (_00445_, _00395_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00446_, _00445_, _00440_);
  or (_00448_, _00446_, _00444_);
  or (_00449_, _00448_, _00443_);
  or (_00450_, _00449_, _00334_);
  and (_00451_, _00450_, _00438_);
  or (_00452_, _00451_, _00387_);
  or (_00453_, _00388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  and (_00454_, _00453_, _06444_);
  and (_13996_, _00454_, _00452_);
  nand (_00455_, _00334_, _11589_);
  and (_00456_, _00406_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  and (_00457_, _00366_, _00397_);
  and (_00458_, _00457_, _00380_);
  or (_00459_, _00458_, _00398_);
  and (_00460_, _00459_, _00400_);
  or (_00461_, _00460_, _00456_);
  or (_00462_, _00461_, _00334_);
  and (_00463_, _00462_, _00455_);
  or (_00464_, _00463_, _00387_);
  nand (_00465_, _00387_, _00397_);
  and (_00466_, _00465_, _06444_);
  and (_14000_, _00466_, _00464_);
  not (_00467_, \oc8051_top_1.oc8051_sfr1.prescaler [2]);
  and (_00468_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  and (_00469_, _00468_, _00467_);
  and (_00470_, _00469_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nor (_00472_, _00468_, _00467_);
  or (_00473_, _00472_, _00469_);
  nand (_00474_, _00473_, _06444_);
  nor (_14009_, _00474_, _00470_);
  or (_00476_, \oc8051_top_1.oc8051_sfr1.prescaler [0], \oc8051_top_1.oc8051_sfr1.prescaler [1]);
  nor (_00477_, _00468_, rst);
  and (_14012_, _00477_, _00476_);
  and (_00478_, _00399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_00479_, _00399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  nor (_00480_, _00479_, _00478_);
  nor (_00481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _00365_);
  nor (_00482_, _00481_, _00366_);
  nor (_00483_, _00482_, _00334_);
  and (_00484_, _00483_, _00480_);
  not (_00485_, _00483_);
  and (_00486_, _00485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_00487_, _00380_, _00399_);
  and (_00488_, _00481_, _00487_);
  nand (_00489_, _00488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  nor (_00490_, _00489_, _00334_);
  or (_00491_, _00490_, _00486_);
  or (_00492_, _00491_, _00484_);
  and (_00493_, _00492_, _00388_);
  nor (_00494_, _00388_, _06666_);
  or (_00495_, _00494_, _00493_);
  and (_14021_, _00495_, _06444_);
  nand (_00496_, _00387_, _10494_);
  and (_00497_, _00478_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_00498_, _00478_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nor (_00499_, _00498_, _00497_);
  and (_00500_, _00499_, _00483_);
  and (_00502_, _00485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  nand (_00503_, _00488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  nor (_00505_, _00503_, _00334_);
  or (_00506_, _00505_, _00502_);
  or (_00507_, _00506_, _00500_);
  or (_00508_, _00507_, _00387_);
  and (_00510_, _00508_, _06444_);
  and (_14023_, _00510_, _00496_);
  and (_00511_, _00347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  and (_00512_, _00511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_00513_, _00512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_00514_, _00513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_00515_, _00514_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  nor (_00516_, _00515_, _00399_);
  and (_00517_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  nor (_00518_, _00517_, _00334_);
  and (_00519_, _00518_, _00516_);
  not (_00520_, _00518_);
  and (_00521_, _00520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_00522_, _00481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  nand (_00523_, _00522_, _00487_);
  nor (_00524_, _00523_, _00334_);
  or (_00525_, _00524_, _00521_);
  or (_00526_, _00525_, _00519_);
  and (_00527_, _00526_, _00388_);
  nor (_00528_, _00388_, _07188_);
  or (_00529_, _00528_, _00527_);
  and (_14026_, _00529_, _06444_);
  nor (_00530_, _00512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  or (_00531_, _00530_, _00513_);
  nand (_00532_, _00531_, _00518_);
  or (_00533_, _00518_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  and (_00534_, _00533_, _00532_);
  and (_00535_, _00497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_00536_, _00481_, _00535_);
  nand (_00537_, _00536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  nor (_00538_, _00537_, _00334_);
  or (_00539_, _00538_, _00387_);
  or (_00540_, _00539_, _00534_);
  nand (_00541_, _00387_, _11589_);
  and (_00542_, _00541_, _06444_);
  and (_14032_, _00542_, _00540_);
  and (_00543_, _00520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nand (_00545_, _00536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  nor (_00546_, _00545_, _00334_);
  or (_00547_, _00546_, _00543_);
  nor (_00548_, _00513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  nor (_00549_, _00548_, _00514_);
  and (_00551_, _00549_, _00518_);
  or (_00552_, _00551_, _00387_);
  or (_00553_, _00552_, _00547_);
  nand (_00554_, _00387_, _07300_);
  and (_00555_, _00554_, _06444_);
  and (_14037_, _00555_, _00553_);
  nor (_00556_, _00511_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  or (_00557_, _00556_, _00512_);
  nand (_00558_, _00557_, _00518_);
  or (_00559_, _00518_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  and (_00560_, _00559_, _00558_);
  nand (_00561_, _00536_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  nor (_00562_, _00561_, _00334_);
  or (_00563_, _00562_, _00387_);
  or (_00564_, _00563_, _00560_);
  nand (_00565_, _00387_, _07069_);
  and (_00566_, _00565_, _06444_);
  and (_14040_, _00566_, _00564_);
  or (_00567_, _00388_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00568_, _00567_, _06444_);
  or (_00570_, _00399_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  nor (_00571_, _00439_, _00362_);
  and (_00573_, _00571_, _00570_);
  or (_00574_, _00487_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_00575_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  or (_00576_, _00575_, _00441_);
  and (_00577_, _00576_, _00574_);
  nor (_00578_, _00577_, _00573_);
  nor (_00579_, _00578_, _00334_);
  and (_00580_, _00334_, _09527_);
  or (_00581_, _00580_, _00579_);
  or (_00582_, _00581_, _00387_);
  and (_14047_, _00582_, _00568_);
  and (_00583_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  not (_00584_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  nor (_00585_, _08064_, _00584_);
  or (_00586_, _00585_, _00583_);
  and (_14073_, _00586_, _06444_);
  nor (_14177_, _11630_, rst);
  and (_00587_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  and (_00588_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_00589_, _00588_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_00590_, _00588_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2]);
  nor (_00591_, _00590_, _00589_);
  or (_00592_, _00591_, _00587_);
  and (_14180_, _00592_, _06444_);
  not (_00593_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0]);
  nor (_00594_, _00587_, _00593_);
  nor (_00595_, _00594_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  and (_00596_, _00594_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1]);
  or (_00597_, _00596_, _00595_);
  nor (_14182_, _00597_, rst);
  and (_00598_, _00587_, _00593_);
  nor (_00599_, _00598_, _00594_);
  and (_14197_, _00599_, _06444_);
  and (_00600_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  not (_00601_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_00602_, _08064_, _00601_);
  or (_00603_, _00602_, _00600_);
  and (_14207_, _00603_, _06444_);
  and (_00604_, _12011_, _08030_);
  and (_00605_, _00604_, _07401_);
  and (_00606_, _00605_, _06933_);
  nand (_00607_, _00606_, _06930_);
  or (_00609_, _00606_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_00610_, _00609_, _06674_);
  and (_00611_, _00610_, _00607_);
  and (_00612_, _07150_, _06382_);
  nand (_00613_, _00612_, _06978_);
  or (_00614_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_00615_, _00614_, _06440_);
  and (_00616_, _00615_, _00613_);
  and (_00617_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  or (_00618_, _00617_, rst);
  or (_00619_, _00618_, _00616_);
  or (_14346_, _00619_, _00611_);
  and (_00620_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  not (_00621_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_00622_, _08064_, _00621_);
  or (_00623_, _00622_, _00620_);
  and (_14348_, _00623_, _06444_);
  nand (_00624_, _10112_, _06978_);
  or (_00625_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [7]);
  and (_00626_, _00625_, _06444_);
  and (_14356_, _00626_, _00624_);
  and (_00627_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  or (_14365_, _00627_, _09368_);
  and (_00628_, _00520_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or (_00630_, _00347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  nor (_00631_, _00511_, _00517_);
  and (_00632_, _00631_, _00630_);
  and (_00633_, _00481_, _00440_);
  nor (_00634_, _00633_, _00632_);
  nor (_00635_, _00634_, _00334_);
  or (_00636_, _00635_, _00387_);
  or (_00637_, _00636_, _00628_);
  nand (_00638_, _00387_, _09526_);
  and (_00639_, _00638_, _06444_);
  and (_14392_, _00639_, _00637_);
  and (_00640_, _07402_, _06394_);
  and (_00641_, _00640_, _06933_);
  nand (_00642_, _00641_, _06930_);
  or (_00643_, _00641_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_00644_, _00643_, _06674_);
  and (_00645_, _00644_, _00642_);
  and (_00646_, _07402_, _07150_);
  nand (_00647_, _00646_, _06978_);
  or (_00648_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_00649_, _00648_, _06440_);
  and (_00651_, _00649_, _00647_);
  and (_00652_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  or (_00653_, _00652_, rst);
  or (_00654_, _00653_, _00651_);
  or (_14416_, _00654_, _00645_);
  nand (_00656_, _10112_, _07069_);
  or (_00657_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [1]);
  and (_00658_, _00657_, _06444_);
  and (_14515_, _00658_, _00656_);
  and (_00659_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  not (_00660_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_00661_, _08064_, _00660_);
  or (_00662_, _00661_, _00659_);
  and (_14522_, _00662_, _06444_);
  or (_00663_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  not (_00664_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  nand (_00665_, _08064_, _00664_);
  and (_00666_, _00665_, _06444_);
  and (_14524_, _00666_, _00663_);
  and (_00667_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  or (_14544_, _00667_, _09376_);
  and (_00668_, _08912_, _06676_);
  and (_00669_, _00668_, _13900_);
  and (_00670_, _00669_, _00240_);
  nand (_00672_, _00670_, _06930_);
  or (_00673_, _00670_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nor (_00674_, _06350_, _06336_);
  and (_00675_, _00674_, _06381_);
  and (_00677_, _00675_, _13889_);
  not (_00678_, _00677_);
  and (_00679_, _00678_, _00673_);
  and (_00680_, _00679_, _00672_);
  nor (_00681_, _00678_, _10494_);
  or (_00682_, _00681_, _00680_);
  and (_00038_, _00682_, _06444_);
  and (_00683_, _00669_, _06987_);
  nand (_00684_, _00683_, _06930_);
  or (_00685_, _00683_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  and (_00686_, _00685_, _00678_);
  and (_00687_, _00686_, _00684_);
  nor (_00689_, _00678_, _06666_);
  or (_00690_, _00689_, _00687_);
  and (_00056_, _00690_, _06444_);
  and (_00692_, _06430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_00693_, _00692_, _08233_);
  and (_00694_, _00693_, _00669_);
  not (_00696_, _00669_);
  nor (_00697_, _06982_, _06430_);
  or (_00698_, _00697_, _00696_);
  and (_00699_, _00698_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_00700_, _00699_, _00677_);
  or (_00702_, _00700_, _00694_);
  nand (_00703_, _00677_, _07188_);
  and (_00704_, _00703_, _06444_);
  and (_00061_, _00704_, _00702_);
  and (_00705_, _00669_, _08310_);
  nand (_00706_, _00705_, _06930_);
  or (_00707_, _00705_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  and (_00708_, _00707_, _00678_);
  and (_00709_, _00708_, _00706_);
  nor (_00710_, _00678_, _07300_);
  or (_00711_, _00710_, _00709_);
  and (_00064_, _00711_, _06444_);
  not (_00712_, _08977_);
  nor (_00713_, _00712_, _06930_);
  and (_00714_, _06431_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_00715_, _00714_, _00713_);
  and (_00716_, _00715_, _00669_);
  or (_00717_, _06932_, _06931_);
  or (_00718_, _00696_, _00717_);
  and (_00719_, _00718_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  or (_00720_, _00719_, _00677_);
  or (_00721_, _00720_, _00716_);
  nand (_00722_, _00677_, _11589_);
  and (_00723_, _00722_, _06444_);
  and (_00066_, _00723_, _00721_);
  and (_00725_, _00669_, _06432_);
  nand (_00726_, _00725_, _06930_);
  or (_00727_, _00725_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  and (_00728_, _00727_, _00678_);
  and (_00729_, _00728_, _00726_);
  nor (_00730_, _00678_, _07069_);
  or (_00731_, _00730_, _00729_);
  and (_00082_, _00731_, _06444_);
  and (_00732_, _00669_, _06942_);
  nand (_00733_, _00732_, _06930_);
  or (_00734_, _00732_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  and (_00735_, _00734_, _00678_);
  and (_00736_, _00735_, _00733_);
  and (_00737_, _00677_, _09527_);
  or (_00738_, _00737_, _00736_);
  and (_00085_, _00738_, _06444_);
  or (_00739_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [30]);
  nand (_00740_, _07432_, _07434_);
  and (_00741_, _00740_, _06444_);
  and (_00088_, _00741_, _00739_);
  and (_00742_, _00668_, _06670_);
  and (_00743_, _00742_, _08310_);
  nand (_00744_, _00743_, _06930_);
  or (_00745_, _00743_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_00746_, _08912_, _06945_);
  and (_00747_, _00746_, _06940_);
  not (_00748_, _00747_);
  and (_00749_, _00748_, _00745_);
  and (_00750_, _00749_, _00744_);
  nor (_00751_, _00748_, _07300_);
  or (_00752_, _00751_, _00750_);
  and (_00143_, _00752_, _06444_);
  and (_00753_, _00742_, _00240_);
  nand (_00754_, _00753_, _06930_);
  or (_00755_, _00753_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_00756_, _00755_, _00748_);
  and (_00757_, _00756_, _00754_);
  nor (_00758_, _00748_, _10494_);
  or (_00759_, _00758_, _00757_);
  and (_00145_, _00759_, _06444_);
  and (_00760_, _00742_, _06987_);
  nand (_00761_, _00760_, _06930_);
  or (_00762_, _00760_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_00763_, _00762_, _00748_);
  and (_00764_, _00763_, _00761_);
  nor (_00765_, _00748_, _06666_);
  or (_00766_, _00765_, _00764_);
  and (_00147_, _00766_, _06444_);
  and (_00767_, _06430_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_00768_, _00767_, _08233_);
  and (_00769_, _00768_, _00742_);
  not (_00770_, _00742_);
  or (_00771_, _00770_, _00697_);
  and (_00772_, _00771_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  or (_00773_, _00772_, _00747_);
  or (_00774_, _00773_, _00769_);
  nand (_00775_, _00747_, _07188_);
  and (_00776_, _00775_, _06444_);
  and (_00149_, _00776_, _00774_);
  and (_00777_, \oc8051_top_1.oc8051_memory_interface1.cdata [2], _08478_);
  and (_00778_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [2]);
  or (_00779_, _00778_, _00777_);
  and (_00151_, _00779_, _06444_);
  and (_00780_, _06431_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_00781_, _00780_, _00713_);
  and (_00782_, _00781_, _00742_);
  or (_00783_, _00770_, _00717_);
  and (_00784_, _00783_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_00785_, _00784_, _00747_);
  or (_00786_, _00785_, _00782_);
  nand (_00787_, _00747_, _11589_);
  and (_00788_, _00787_, _06444_);
  and (_00153_, _00788_, _00786_);
  and (_00789_, \oc8051_top_1.oc8051_memory_interface1.cdata [6], _08478_);
  and (_00790_, \oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00791_, _00790_, _00789_);
  and (_00162_, _00791_, _06444_);
  and (_00792_, _08478_, \oc8051_top_1.oc8051_memory_interface1.cdata [5]);
  and (_00793_, \oc8051_top_1.oc8051_memory_interface1.istb_t , \oc8051_top_1.oc8051_rom1.data_o [5]);
  or (_00794_, _00793_, _00792_);
  and (_00164_, _00794_, _06444_);
  and (_00795_, \oc8051_top_1.oc8051_memory_interface1.cdata [4], _08478_);
  and (_00796_, \oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00797_, _00796_, _00795_);
  and (_00166_, _00797_, _06444_);
  and (_00798_, _00742_, _06432_);
  nand (_00799_, _00798_, _06930_);
  or (_00800_, _00798_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  and (_00801_, _00800_, _00748_);
  and (_00802_, _00801_, _00799_);
  nor (_00803_, _00748_, _07069_);
  or (_00804_, _00803_, _00802_);
  and (_00169_, _00804_, _06444_);
  and (_00805_, _00742_, _06942_);
  nand (_00806_, _00805_, _06930_);
  or (_00807_, _00805_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_00808_, _00807_, _00748_);
  and (_00809_, _00808_, _00806_);
  and (_00810_, _00747_, _09527_);
  or (_00811_, _00810_, _00809_);
  and (_00172_, _00811_, _06444_);
  and (_00812_, \oc8051_top_1.oc8051_memory_interface1.cdata [3], _08478_);
  and (_00813_, \oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00814_, _00813_, _00812_);
  and (_00177_, _00814_, _06444_);
  and (_00815_, \oc8051_top_1.oc8051_memory_interface1.cdata [1], _08478_);
  and (_00816_, \oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_00817_, _00816_, _00815_);
  and (_00189_, _00817_, _06444_);
  and (_00818_, _13901_, _06670_);
  and (_00819_, _00818_, _06983_);
  nand (_00820_, _00819_, _06930_);
  or (_00821_, _00819_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_00822_, _00821_, _07408_);
  and (_00823_, _00822_, _00820_);
  nor (_00824_, _07408_, _07188_);
  or (_00825_, _00824_, _00823_);
  and (_00191_, _00825_, _06444_);
  and (_00826_, _00818_, _08977_);
  nand (_00827_, _00826_, _06930_);
  or (_00828_, _00826_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  and (_00829_, _00828_, _07408_);
  and (_00830_, _00829_, _00827_);
  nor (_00831_, _11589_, _07408_);
  or (_00832_, _00831_, _00830_);
  and (_00205_, _00832_, _06444_);
  and (_00833_, _00818_, _06942_);
  or (_00834_, _00833_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_00835_, _00834_, _07408_);
  nand (_00836_, _00833_, _06930_);
  and (_00837_, _00836_, _00835_);
  and (_00838_, _09527_, _07407_);
  or (_00839_, _00838_, _00837_);
  and (_00211_, _00839_, _06444_);
  and (_00840_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  or (_00841_, _00840_, _09452_);
  and (_00239_, _00841_, _06444_);
  nor (_00842_, _13916_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_00843_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  nand (_00844_, _00842_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re );
  and (_00845_, _00844_, _06444_);
  and (_00247_, _00845_, _00843_);
  nand (_00846_, _07199_, _07195_);
  and (_00847_, _07199_, _07108_);
  or (_00848_, _00847_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0]);
  and (_00849_, _00848_, _06444_);
  and (_00252_, _00849_, _00846_);
  nor (_00850_, _07073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nand (_00851_, _00850_, _07195_);
  and (_00852_, _00850_, _07108_);
  or (_00853_, _00852_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0]);
  and (_00854_, _00853_, _06444_);
  and (_00256_, _00854_, _00851_);
  not (_00855_, _11452_);
  and (_00856_, _12023_, _00855_);
  and (_00272_, _00856_, _06444_);
  or (_00857_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00858_, _00857_, _07120_);
  or (_00859_, _00858_, _07126_);
  and (_00860_, _07111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_00861_, _00860_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00862_, _07113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_00863_, _00862_, _07116_);
  and (_00864_, _00863_, _00861_);
  nand (_00865_, _07394_, _07116_);
  nand (_00866_, _00865_, _07125_);
  or (_00867_, _00866_, _00864_);
  and (_00868_, _00867_, _00859_);
  and (_00869_, _07394_, _07119_);
  or (_00870_, _00869_, _07130_);
  or (_00871_, _00870_, _00868_);
  or (_00872_, _07131_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00873_, _00872_, _00871_);
  and (_00874_, _00873_, _07134_);
  and (_00875_, _00857_, _07085_);
  or (_00876_, _00875_, _07091_);
  and (_00877_, _07095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  or (_00878_, _00877_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  nor (_00879_, _07101_, _07077_);
  nor (_00880_, _00879_, _07104_);
  and (_00881_, _00880_, _00878_);
  nand (_00882_, _07394_, _07104_);
  nand (_00883_, _00882_, _07090_);
  or (_00884_, _00883_, _00881_);
  and (_00885_, _00884_, _00876_);
  and (_00886_, _07394_, _07084_);
  or (_00887_, _00886_, _00885_);
  and (_00888_, _00887_, _07108_);
  or (_00889_, _00888_, _07073_);
  or (_00890_, _00889_, _00874_);
  or (_00891_, _07075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1]);
  and (_00892_, _00891_, _06444_);
  and (_00274_, _00892_, _00890_);
  or (_00893_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_00894_, _00893_, _07085_);
  not (_00895_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  or (_00896_, _00877_, _00895_);
  nand (_00897_, _00896_, _00880_);
  or (_00898_, _07385_, _07105_);
  and (_00899_, _00898_, _00897_);
  or (_00900_, _00899_, _07089_);
  not (_00901_, _07087_);
  not (_00902_, _07089_);
  or (_00903_, _00893_, _00902_);
  and (_00904_, _00903_, _00901_);
  and (_00905_, _00904_, _00900_);
  and (_00906_, _07385_, _07087_);
  or (_00907_, _00906_, _07084_);
  or (_00908_, _00907_, _00905_);
  and (_00909_, _00908_, _00894_);
  or (_00910_, _00909_, _07134_);
  or (_00911_, _00893_, _07120_);
  or (_00912_, _00860_, _00895_);
  nand (_00913_, _00912_, _00863_);
  or (_00914_, _07385_, _07117_);
  and (_00915_, _00914_, _00913_);
  or (_00916_, _00915_, _07124_);
  not (_00917_, _07122_);
  not (_00918_, _07124_);
  or (_00919_, _00893_, _00918_);
  and (_00920_, _00919_, _00917_);
  and (_00921_, _00920_, _00916_);
  and (_00922_, _07385_, _07122_);
  or (_00923_, _00922_, _07119_);
  or (_00924_, _00923_, _00921_);
  and (_00925_, _00924_, _00911_);
  or (_00926_, _00925_, _07196_);
  and (_00927_, _00926_, _00910_);
  or (_00928_, _00927_, _07073_);
  nor (_00929_, _07132_, _07073_);
  or (_00930_, _00929_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0]);
  and (_00931_, _00930_, _06444_);
  and (_00276_, _00931_, _00928_);
  or (_00932_, _00589_, \oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3]);
  and (_00278_, _00932_, _06444_);
  and (_00933_, _06442_, _06444_);
  and (_00934_, _00933_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_00935_, _13854_, _06298_);
  nor (_00936_, _00935_, _13836_);
  and (_00937_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_00938_, _00937_, _06443_);
  or (_00280_, _00938_, _00934_);
  nor (_00282_, _12648_, rst);
  and (_00287_, _11576_, _06444_);
  or (_00939_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_00940_, _00939_, _07120_);
  or (_00941_, _00940_, _07126_);
  and (_00942_, _07111_, _07077_);
  or (_00943_, _00942_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_00944_, _07113_, _07077_);
  nor (_00945_, _00944_, _07116_);
  and (_00946_, _00945_, _00943_);
  nand (_00947_, _07393_, _07116_);
  nand (_00948_, _00947_, _07125_);
  or (_00949_, _00948_, _00946_);
  and (_00950_, _00949_, _00941_);
  and (_00951_, _07393_, _07119_);
  or (_00952_, _00951_, _07130_);
  or (_00953_, _00952_, _00950_);
  or (_00954_, _07131_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_00955_, _00954_, _00953_);
  and (_00956_, _00955_, _07134_);
  and (_00957_, _00939_, _07085_);
  or (_00958_, _00957_, _07091_);
  and (_00959_, _07393_, _07104_);
  nor (_00960_, _07101_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0]);
  nor (_00961_, _00960_, _07104_);
  and (_00962_, _07095_, _07077_);
  or (_00963_, _00962_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  nand (_00964_, _00963_, _00961_);
  nand (_00965_, _00964_, _07090_);
  or (_00966_, _00965_, _00959_);
  and (_00967_, _00966_, _00958_);
  and (_00968_, _07393_, _07084_);
  or (_00969_, _00968_, _00967_);
  and (_00970_, _00969_, _07108_);
  or (_00971_, _00970_, _00956_);
  or (_00972_, _00971_, _07073_);
  or (_00973_, _07075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1]);
  and (_00974_, _00973_, _06444_);
  and (_00295_, _00974_, _00972_);
  or (_00975_, _07077_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_00977_, _00975_, _07120_);
  or (_00978_, _07384_, _00917_);
  not (_00979_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  or (_00980_, _00942_, _00979_);
  nand (_00981_, _00980_, _00945_);
  or (_00982_, _07384_, _07117_);
  and (_00983_, _00982_, _00918_);
  and (_00984_, _00983_, _00981_);
  and (_00985_, _00975_, _07124_);
  or (_00986_, _00985_, _07122_);
  or (_00987_, _00986_, _00984_);
  and (_00988_, _00987_, _00978_);
  or (_00989_, _00988_, _07119_);
  and (_00990_, _00989_, _00977_);
  or (_00991_, _00990_, _07196_);
  or (_00992_, _00975_, _07085_);
  or (_00993_, _00962_, _00979_);
  nand (_00994_, _00993_, _00961_);
  or (_00995_, _07384_, _07105_);
  and (_00996_, _00995_, _00994_);
  or (_00997_, _00996_, _07089_);
  or (_00998_, _00975_, _00902_);
  and (_01000_, _00998_, _00901_);
  and (_01001_, _01000_, _00997_);
  and (_01002_, _07384_, _07087_);
  or (_01003_, _01002_, _07084_);
  or (_01004_, _01003_, _01001_);
  and (_01005_, _01004_, _00992_);
  or (_01006_, _01005_, _07134_);
  and (_01007_, _01006_, _00991_);
  or (_01008_, _01007_, _07073_);
  or (_01009_, _00929_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0]);
  and (_01010_, _01009_, _06444_);
  and (_00299_, _01010_, _01008_);
  nor (_01011_, _07108_, _07073_);
  or (_01012_, _01011_, _07077_);
  nand (_01013_, _00850_, _07132_);
  and (_01014_, _01013_, _06444_);
  and (_00326_, _01014_, _01012_);
  and (_01015_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _06444_);
  and (_00331_, _01015_, _07073_);
  nand (_01016_, _07127_, _07203_);
  nor (_01017_, _01016_, _07108_);
  and (_01018_, _07073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  or (_01019_, _07104_, _07073_);
  nor (_01020_, _01019_, _07082_);
  not (_01021_, _07091_);
  nor (_01022_, _07102_, _01021_);
  and (_01023_, _01022_, _01020_);
  or (_01024_, _01023_, _01018_);
  or (_01025_, _01024_, _01017_);
  and (_00339_, _01025_, _06444_);
  or (_01026_, _07124_, _07116_);
  and (_01027_, _07114_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_01028_, _01027_, _01026_);
  and (_01029_, _01028_, _00917_);
  and (_01030_, _07195_, _07120_);
  and (_01031_, _01030_, _01029_);
  or (_01032_, _07104_, _07089_);
  and (_01033_, _07102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  or (_01034_, _01033_, _01032_);
  and (_01035_, _01034_, _00901_);
  and (_01036_, _07108_, _07085_);
  and (_01037_, _01036_, _01035_);
  or (_01038_, _01037_, _07073_);
  or (_01039_, _01038_, _01031_);
  or (_01040_, _07075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_01041_, _01040_, _06444_);
  and (_00342_, _01041_, _01039_);
  nor (_01042_, _07111_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  nor (_01043_, _01042_, _07113_);
  or (_01044_, _01043_, _07116_);
  and (_01045_, _01044_, _00918_);
  or (_01046_, _01045_, _07122_);
  and (_01047_, _01046_, _01030_);
  or (_01048_, _07095_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01049_, _01048_, _07101_);
  or (_01050_, _01049_, _07104_);
  and (_01051_, _01050_, _00902_);
  or (_01052_, _01051_, _07087_);
  and (_01053_, _01052_, _01036_);
  or (_01054_, _01053_, _07073_);
  or (_01055_, _01054_, _01047_);
  or (_01056_, _07075_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01057_, _01056_, _06444_);
  and (_00345_, _01057_, _01055_);
  and (_00350_, _12703_, _07073_);
  and (_01058_, _07073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  or (_01059_, _01058_, _00929_);
  and (_00368_, _01059_, _06444_);
  and (_01060_, _07073_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  or (_01061_, _01060_, _00929_);
  and (_00371_, _01061_, _06444_);
  and (_01062_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [29]);
  and (_01063_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [29]);
  or (_01064_, _01063_, _01062_);
  and (_00434_, _01064_, _06444_);
  and (_01065_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  not (_01066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_01067_, _08064_, _01066_);
  or (_01068_, _01067_, _01065_);
  and (_00447_, _01068_, _06444_);
  and (_01069_, _12825_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nand (_01070_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [1]);
  nor (_01071_, _01070_, _07415_);
  and (_01072_, _12829_, _07070_);
  or (_01073_, _01072_, _01071_);
  or (_01074_, _01073_, _01069_);
  and (_00471_, _01074_, _06444_);
  or (_01075_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  not (_01076_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nand (_01077_, _08064_, _01076_);
  and (_01078_, _01077_, _06444_);
  and (_00475_, _01078_, _01075_);
  and (_01079_, _00604_, _08912_);
  and (_01080_, _01079_, _06933_);
  nand (_01081_, _01080_, _06930_);
  or (_01082_, _01080_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_01083_, _01082_, _06674_);
  and (_01084_, _01083_, _01081_);
  and (_01085_, _00674_, _07150_);
  and (_01086_, _01085_, _06381_);
  not (_01087_, _01086_);
  nor (_01088_, _01087_, _06978_);
  and (_01089_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_01090_, _01089_, _01088_);
  and (_01091_, _01090_, _06440_);
  and (_01092_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  or (_01093_, _01092_, rst);
  or (_01094_, _01093_, _01091_);
  or (_00501_, _01094_, _01084_);
  and (_01095_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [4]);
  nor (_01096_, _14070_, _07188_);
  or (_01097_, _01096_, _01095_);
  and (_00504_, _01097_, _06444_);
  nor (_01098_, _12830_, _07300_);
  nor (_01099_, _07415_, _07158_);
  or (_01100_, _01099_, _12825_);
  and (_01101_, _01100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [3]);
  or (_01102_, _01101_, _01098_);
  and (_00509_, _01102_, _06444_);
  and (_01103_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  or (_00544_, _01103_, _09383_);
  and (_01104_, _09373_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_00550_, _01104_, _09390_);
  or (_01105_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  not (_01106_, \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  nand (_01107_, _08064_, _01106_);
  and (_01108_, _01107_, _06444_);
  and (_00569_, _01108_, _01105_);
  and (_01109_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  not (_01110_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_01111_, _08064_, _01110_);
  or (_01112_, _01111_, _01109_);
  and (_00572_, _01112_, _06444_);
  nor (_00608_, _11688_, rst);
  nor (_01113_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_01114_, _01113_, _06296_);
  and (_01115_, _01114_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11]);
  not (_01116_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  nor (_01117_, _01114_, _01116_);
  or (_01118_, _01117_, _01115_);
  or (_01119_, _01118_, _13902_);
  or (_01120_, _08977_, _01116_);
  nand (_01121_, _01120_, _13902_);
  or (_01122_, _01121_, _00713_);
  and (_01123_, _01122_, _01119_);
  or (_01124_, _01123_, _13906_);
  nand (_01125_, _13906_, _11589_);
  and (_01126_, _01125_, _06444_);
  and (_00629_, _01126_, _01124_);
  and (_01127_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  not (_01128_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nor (_01129_, _08064_, _01128_);
  or (_01130_, _01129_, _01127_);
  and (_00650_, _01130_, _06444_);
  and (_01131_, _10891_, \oc8051_top_1.oc8051_memory_interface1.op_pos [0]);
  or (_01132_, _10882_, _07236_);
  nand (_01133_, _10882_, _07236_);
  and (_01134_, _01133_, _01132_);
  nand (_01135_, _01134_, _01131_);
  or (_01136_, _01134_, _01131_);
  and (_01137_, _01136_, _01135_);
  or (_01138_, _01137_, _07429_);
  or (_01139_, _07230_, \oc8051_top_1.oc8051_memory_interface1.op_pos [1]);
  and (_01140_, _01139_, _10894_);
  and (_00655_, _01140_, _01138_);
  or (_01141_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  not (_01142_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_01143_, _08064_, _01142_);
  and (_01144_, _01143_, _06444_);
  and (_00671_, _01144_, _01141_);
  and (_01146_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  nor (_01147_, _08064_, _01142_);
  or (_01148_, _01147_, _01146_);
  and (_00676_, _01148_, _06444_);
  or (_01149_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  not (_01150_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_01151_, _08064_, _01150_);
  and (_01152_, _01151_, _06444_);
  and (_00688_, _01152_, _01149_);
  and (_01153_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  not (_01154_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_01155_, _08064_, _01154_);
  or (_01156_, _01155_, _01153_);
  and (_00691_, _01156_, _06444_);
  and (_01158_, _13902_, _06987_);
  nand (_01160_, _01158_, _06930_);
  or (_01161_, _01158_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_01162_, _01161_, _13907_);
  and (_01163_, _01162_, _01160_);
  nor (_01165_, _13907_, _06666_);
  or (_01166_, _01165_, _01163_);
  and (_00695_, _01166_, _06444_);
  and (_01167_, _13902_, _06983_);
  nand (_01168_, _01167_, _06930_);
  or (_01169_, _01167_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_01170_, _01169_, _13907_);
  and (_01171_, _01170_, _01168_);
  nor (_01172_, _13907_, _07188_);
  or (_01173_, _01172_, _01171_);
  and (_00701_, _01173_, _06444_);
  or (_01174_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [14]);
  nand (_01175_, _07432_, _13985_);
  and (_01176_, _01175_, _06444_);
  and (_00724_, _01176_, _01174_);
  and (_01177_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1]);
  or (_01178_, _01177_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  and (_00976_, _01178_, _06444_);
  and (_01179_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0]);
  or (_01180_, _01179_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  and (_00999_, _01180_, _06444_);
  nor (_01181_, _06978_, _06449_);
  and (_01182_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [7]);
  or (_01184_, _01182_, _01181_);
  and (_01157_, _01184_, _06444_);
  and (_01185_, _13902_, _08310_);
  nand (_01186_, _01185_, _06930_);
  or (_01187_, _01185_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_01188_, _01187_, _13907_);
  and (_01189_, _01188_, _01186_);
  nor (_01190_, _13907_, _07300_);
  or (_01191_, _01190_, _01189_);
  and (_01159_, _01191_, _06444_);
  and (_01192_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  and (_01193_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_01194_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  or (_01195_, _01194_, _01193_);
  and (_01196_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_01197_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_01198_, _01197_, _01196_);
  or (_01199_, _01198_, _01195_);
  and (_01200_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_01201_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  or (_01202_, _01201_, _01200_);
  and (_01203_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_01204_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  or (_01205_, _01204_, _01203_);
  or (_01206_, _01205_, _01202_);
  or (_01207_, _01206_, _01199_);
  and (_01208_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  and (_01209_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  or (_01210_, _01209_, _01208_);
  and (_01211_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  and (_01212_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  or (_01213_, _01212_, _01211_);
  or (_01214_, _01213_, _01210_);
  and (_01215_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  and (_01216_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  or (_01217_, _01216_, _01215_);
  and (_01219_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  and (_01220_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  or (_01221_, _01220_, _01219_);
  or (_01222_, _01221_, _01217_);
  or (_01223_, _01222_, _01214_);
  or (_01224_, _01223_, _01207_);
  and (_01225_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  not (_01226_, _11734_);
  and (_01227_, _14156_, _01226_);
  or (_01228_, _01227_, _01225_);
  and (_01229_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  and (_01230_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  or (_01231_, _01230_, _01229_);
  or (_01232_, _01231_, _01228_);
  or (_01233_, _14247_, p3_in[5]);
  or (_01234_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_01235_, _01234_, _01233_);
  and (_01236_, _01235_, _14260_);
  or (_01237_, _14247_, p2_in[5]);
  or (_01238_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_01239_, _01238_, _01237_);
  and (_01240_, _01239_, _14265_);
  or (_01241_, _01240_, _01236_);
  or (_01242_, _14247_, p0_in[5]);
  or (_01243_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01244_, _01243_, _01242_);
  and (_01245_, _01244_, _14224_);
  or (_01246_, _14247_, p1_in[5]);
  or (_01248_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_01249_, _01248_, _01246_);
  and (_01250_, _01249_, _14253_);
  or (_01251_, _01250_, _01245_);
  or (_01252_, _01251_, _01241_);
  or (_01253_, _01252_, _01232_);
  and (_01254_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_01255_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  or (_01256_, _01255_, _01254_);
  or (_01257_, _01256_, _01253_);
  or (_01258_, _01257_, _01224_);
  and (_01259_, _01258_, _14174_);
  or (_01260_, _01259_, _14178_);
  or (_01261_, _01260_, _01192_);
  or (_01262_, _14353_, _08127_);
  and (_01263_, _01262_, _06444_);
  and (_01164_, _01263_, _01261_);
  nor (_01264_, _11589_, _07190_);
  and (_01265_, _10497_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [2]);
  or (_01266_, _01265_, _01264_);
  and (_01183_, _01266_, _06444_);
  and (_01267_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [0]);
  and (_01268_, _12841_, _06447_);
  or (_01269_, _01268_, _01267_);
  and (_01218_, _01269_, _06444_);
  and (_01270_, _07414_, _06439_);
  or (_01271_, _01270_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [0]);
  nand (_01272_, _01270_, _09526_);
  and (_01273_, _01272_, _06444_);
  and (_01247_, _01273_, _01271_);
  or (_01274_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  not (_01275_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  nand (_01276_, _08064_, _01275_);
  and (_01277_, _01276_, _06444_);
  and (_01378_, _01277_, _01274_);
  and (_01278_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  not (_01279_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_01280_, _08064_, _01279_);
  or (_01281_, _01280_, _01278_);
  and (_01394_, _01281_, _06444_);
  nor (_01282_, _14070_, _07300_);
  and (_01283_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [3]);
  or (_01284_, _01283_, _01282_);
  and (_01641_, _01284_, _06444_);
  nor (_01285_, \oc8051_top_1.oc8051_decoder1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  and (_01286_, _01285_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  not (_01287_, _01286_);
  or (_01288_, _01287_, _08308_);
  or (_01289_, _01286_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [3]);
  and (_01290_, _01289_, _06444_);
  and (_01650_, _01290_, _01288_);
  and (_01291_, _12711_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6]);
  or (_01292_, _01291_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  and (_01676_, _01292_, _06444_);
  and (_01293_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5]);
  or (_01294_, _01293_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  and (_01679_, _01294_, _06444_);
  and (_01295_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4]);
  or (_01296_, _01295_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  and (_01684_, _01296_, _06444_);
  nand (_01297_, _01286_, _09138_);
  or (_01298_, _01286_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [2]);
  and (_01299_, _01298_, _06444_);
  and (_01697_, _01299_, _01297_);
  not (_01300_, _06432_);
  nor (_01301_, _06930_, _01300_);
  nand (_01302_, _01300_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  nand (_01303_, _01302_, _13902_);
  or (_01304_, _01303_, _01301_);
  or (_01305_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_01306_, _01305_, _13902_);
  and (_01307_, _01306_, _01304_);
  or (_01308_, _01307_, _13906_);
  nand (_01309_, _13906_, _07069_);
  and (_01310_, _01309_, _06444_);
  and (_01700_, _01310_, _01308_);
  not (_01311_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  or (_01312_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _01311_);
  or (_01313_, _01312_, _06295_);
  and (_01314_, _01313_, _01113_);
  or (_01315_, _01314_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_01316_, _01315_, _13902_);
  nand (_01317_, _08021_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  nand (_01318_, _01317_, _13902_);
  or (_01319_, _01318_, _08022_);
  and (_01320_, _01319_, _01316_);
  or (_01321_, _01320_, _13906_);
  nand (_01322_, _13906_, _09526_);
  and (_01323_, _01322_, _06444_);
  and (_01702_, _01323_, _01321_);
  and (_01324_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [17]);
  and (_01325_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [17]);
  or (_01326_, _01325_, _01324_);
  and (_01708_, _01326_, _06444_);
  and (_01327_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3]);
  or (_01328_, _01327_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  and (_01716_, _01328_, _06444_);
  and (_01329_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [6]);
  nor (_01330_, _14070_, _10494_);
  or (_01331_, _01330_, _01329_);
  and (_01734_, _01331_, _06444_);
  or (_01332_, _01287_, _07959_);
  or (_01333_, _01286_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [1]);
  and (_01334_, _01333_, _06444_);
  and (_01752_, _01334_, _01332_);
  or (_01335_, _01287_, _08019_);
  or (_01336_, _01286_, \oc8051_top_1.oc8051_memory_interface1.iadr_t [0]);
  and (_01337_, _01336_, _06444_);
  and (_01786_, _01337_, _01335_);
  and (_01338_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  nor (_01339_, _08064_, _00664_);
  or (_01340_, _01339_, _01338_);
  and (_01790_, _01340_, _06444_);
  and (_01341_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [16]);
  and (_01343_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [16]);
  or (_01344_, _01343_, _01341_);
  and (_01803_, _01344_, _06444_);
  nor (_01806_, \oc8051_top_1.oc8051_sfr1.prescaler [0], rst);
  and (_01345_, _08230_, _06444_);
  or (_01346_, _01345_, _14496_);
  and (_01347_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  and (_01348_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  and (_01349_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  or (_01350_, _01349_, _01348_);
  and (_01351_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_01352_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  or (_01353_, _01352_, _01351_);
  or (_01354_, _01353_, _01350_);
  and (_01355_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_01356_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_01357_, _01356_, _01355_);
  and (_01358_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  and (_01359_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  or (_01360_, _01359_, _01358_);
  or (_01361_, _01360_, _01357_);
  or (_01362_, _01361_, _01354_);
  and (_01363_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  and (_01364_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  or (_01365_, _01364_, _01363_);
  and (_01366_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  and (_01367_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  or (_01368_, _01367_, _01366_);
  or (_01369_, _01368_, _01365_);
  and (_01370_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  and (_01371_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  or (_01372_, _01371_, _01370_);
  and (_01373_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  and (_01374_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  or (_01375_, _01374_, _01373_);
  or (_01376_, _01375_, _01372_);
  or (_01377_, _01376_, _01369_);
  or (_01379_, _01377_, _01362_);
  and (_01380_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  and (_01381_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  or (_01382_, _01381_, _01380_);
  and (_01383_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_01384_, _14156_, _11664_);
  or (_01385_, _01384_, _01383_);
  or (_01386_, _01385_, _01382_);
  or (_01387_, _14247_, p0_in[4]);
  or (_01388_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_01389_, _01388_, _01387_);
  and (_01390_, _01389_, _14224_);
  or (_01391_, _14247_, p1_in[4]);
  or (_01392_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_01393_, _01392_, _01391_);
  and (_01395_, _01393_, _14253_);
  or (_01396_, _01395_, _01390_);
  or (_01397_, _14247_, p3_in[4]);
  or (_01398_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_01399_, _01398_, _01397_);
  and (_01400_, _01399_, _14260_);
  or (_01401_, _14247_, p2_in[4]);
  or (_01402_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_01403_, _01402_, _01401_);
  and (_01404_, _01403_, _14265_);
  or (_01405_, _01404_, _01400_);
  or (_01406_, _01405_, _01396_);
  or (_01407_, _01406_, _01386_);
  and (_01408_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_01409_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_01410_, _01409_, _01408_);
  or (_01411_, _01410_, _01407_);
  or (_01412_, _01411_, _01379_);
  and (_01413_, _01412_, _14174_);
  or (_01414_, _01413_, _14178_);
  or (_01415_, _01414_, _01347_);
  and (_01808_, _01415_, _01346_);
  and (_01416_, _08019_, _06444_);
  or (_01417_, _01416_, _14496_);
  and (_01418_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_01419_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_01420_, _01419_, _01418_);
  and (_01421_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_01422_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_01423_, _01422_, _01421_);
  or (_01424_, _01423_, _01420_);
  and (_01425_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_01426_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or (_01427_, _01426_, _01425_);
  and (_01428_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  and (_01429_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  or (_01430_, _01429_, _01428_);
  or (_01431_, _01430_, _01427_);
  or (_01432_, _01431_, _01424_);
  and (_01433_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  and (_01434_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  or (_01435_, _01434_, _01433_);
  and (_01436_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  and (_01437_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  or (_01438_, _01437_, _01436_);
  or (_01439_, _01438_, _01435_);
  and (_01440_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  and (_01441_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  or (_01442_, _01441_, _01440_);
  and (_01443_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  and (_01444_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  or (_01445_, _01444_, _01443_);
  or (_01446_, _01445_, _01442_);
  or (_01447_, _01446_, _01439_);
  or (_01448_, _01447_, _01432_);
  and (_01449_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  and (_01450_, _14156_, _11858_);
  or (_01451_, _01450_, _01449_);
  and (_01452_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  and (_01453_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  or (_01454_, _01453_, _01452_);
  or (_01455_, _01454_, _01451_);
  or (_01456_, _14247_, p3_in[0]);
  or (_01457_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_01458_, _01457_, _01456_);
  and (_01459_, _01458_, _14260_);
  or (_01460_, _14247_, p2_in[0]);
  or (_01461_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_01462_, _01461_, _01460_);
  and (_01463_, _01462_, _14265_);
  or (_01464_, _01463_, _01459_);
  or (_01465_, _14247_, p0_in[0]);
  or (_01466_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_01467_, _01466_, _01465_);
  and (_01468_, _01467_, _14224_);
  or (_01469_, _14247_, p1_in[0]);
  or (_01470_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_01471_, _01470_, _01469_);
  and (_01472_, _01471_, _14253_);
  or (_01473_, _01472_, _01468_);
  or (_01474_, _01473_, _01464_);
  or (_01475_, _01474_, _01455_);
  or (_01476_, _08269_, _08196_);
  nand (_01477_, _08269_, _08196_);
  nand (_01478_, _01477_, _01476_);
  or (_01479_, _09045_, _07652_);
  not (_01480_, _00240_);
  nor (_01481_, _01480_, _06930_);
  nor (_01482_, _00240_, _06736_);
  nor (_01483_, _01482_, _01481_);
  nor (_01484_, _01483_, _08028_);
  and (_01485_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_01486_, _01485_, _07439_);
  nor (_01487_, _01486_, _01484_);
  nand (_01488_, _01487_, _01479_);
  and (_01489_, _09201_, _07439_);
  not (_01490_, _01489_);
  and (_01491_, _01490_, _01488_);
  or (_01492_, _01491_, _11179_);
  nand (_01493_, _01491_, _11179_);
  and (_01494_, _01493_, _01492_);
  nand (_01495_, _01494_, _01478_);
  or (_01496_, _01494_, _01478_);
  and (_01497_, _01496_, _01495_);
  or (_01498_, _08063_, _07976_);
  nand (_01499_, _08063_, _07976_);
  nand (_01500_, _01499_, _01498_);
  or (_01501_, _09138_, _07652_);
  nor (_01502_, _08977_, _06782_);
  nor (_01503_, _01502_, _00713_);
  nor (_01504_, _01503_, _08028_);
  and (_01505_, _08036_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_01506_, _01505_, _07439_);
  nor (_01507_, _01506_, _01504_);
  and (_01508_, _01507_, _01501_);
  and (_01509_, _09280_, _07439_);
  or (_01510_, _01509_, _01508_);
  nand (_01511_, _01510_, _08344_);
  or (_01512_, _01510_, _08344_);
  and (_01513_, _01512_, _01511_);
  nand (_01514_, _01513_, _01500_);
  or (_01515_, _01513_, _01500_);
  and (_01516_, _01515_, _01514_);
  nor (_01517_, _01516_, _01497_);
  and (_01518_, _01516_, _01497_);
  or (_01519_, _01518_, _01517_);
  and (_01520_, _01519_, _14143_);
  and (_01521_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_01522_, _01521_, _01520_);
  or (_01523_, _01522_, _01475_);
  or (_01524_, _01523_, _01448_);
  and (_01525_, _01524_, _14174_);
  and (_01526_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  or (_01527_, _01526_, _14178_);
  or (_01528_, _01527_, _01525_);
  and (_01810_, _01528_, _01417_);
  not (_01529_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  not (_01530_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  and (_01531_, _10967_, _01530_);
  and (_01532_, _01531_, _01529_);
  nor (_01533_, _01531_, _01529_);
  nor (_01534_, _01533_, _01532_);
  not (_01535_, _01534_);
  nor (_01536_, _10967_, _01530_);
  or (_01537_, _01536_, _01531_);
  and (_01538_, _01537_, _10970_);
  and (_01539_, _01538_, _01535_);
  nor (_01540_, _01538_, _01535_);
  nor (_01541_, _01540_, _01539_);
  or (_01542_, _01541_, _08374_);
  or (_01543_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_01544_, _01543_, _10894_);
  and (_01545_, _01544_, _01542_);
  and (_01546_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_01846_, _01546_, _01545_);
  not (_01547_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  not (_01548_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  not (_01549_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  and (_01550_, _01532_, _01549_);
  and (_01551_, _01550_, _01548_);
  nor (_01552_, _01551_, _01547_);
  and (_01553_, _01551_, _01547_);
  nor (_01554_, _01553_, _01552_);
  not (_01555_, _01554_);
  nor (_01556_, _01550_, _01548_);
  or (_01557_, _01556_, _01551_);
  nor (_01558_, _01532_, _01549_);
  nor (_01559_, _01558_, _01550_);
  not (_01561_, _01559_);
  and (_01562_, _01561_, _01539_);
  and (_01563_, _01562_, _01557_);
  and (_01564_, _01563_, _01555_);
  nor (_01565_, _01563_, _01555_);
  nor (_01566_, _01565_, _01564_);
  or (_01567_, _01566_, _08374_);
  or (_01568_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  and (_01569_, _01568_, _10894_);
  and (_01570_, _01569_, _01567_);
  and (_01571_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_01849_, _01571_, _01570_);
  nor (_01572_, _01562_, _01557_);
  nor (_01573_, _01572_, _01563_);
  or (_01574_, _01573_, _08374_);
  or (_01575_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_01576_, _01575_, _10894_);
  and (_01577_, _01576_, _01574_);
  and (_01578_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_01854_, _01578_, _01577_);
  and (_01579_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  not (_01580_, \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  nor (_01581_, _08064_, _01580_);
  or (_01582_, _01581_, _01579_);
  and (_01974_, _01582_, _06444_);
  and (_01583_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nor (_01584_, _01561_, _01539_);
  nor (_01585_, _01584_, _01562_);
  or (_01586_, _01585_, _08374_);
  or (_01587_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  and (_01588_, _01587_, _10894_);
  and (_01589_, _01588_, _01586_);
  or (_02013_, _01589_, _01583_);
  and (_01590_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_01591_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nor (_01592_, _08064_, _01591_);
  or (_01593_, _01592_, _01590_);
  and (_02042_, _01593_, _06444_);
  nor (_01594_, _01537_, _10970_);
  nor (_01595_, _01594_, _01538_);
  or (_01596_, _01595_, _08374_);
  or (_01597_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  and (_01598_, _01597_, _10894_);
  and (_01599_, _01598_, _01596_);
  and (_01600_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_02046_, _01600_, _01599_);
  and (_01601_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  not (_01602_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_01603_, _08064_, _01602_);
  or (_01604_, _01603_, _01601_);
  and (_02090_, _01604_, _06444_);
  and (_01605_, _07425_, _11568_);
  and (_01606_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_01607_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [7]);
  and (_01608_, _01607_, _09332_);
  or (_01609_, _01608_, _01606_);
  or (_01610_, _01609_, _01605_);
  and (_02146_, _01610_, _06444_);
  or (_01611_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  and (_01612_, _01611_, _06444_);
  nand (_01613_, _13893_, _06666_);
  and (_02191_, _01613_, _01612_);
  or (_01614_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  and (_01615_, _01614_, _06444_);
  nand (_01616_, _13893_, _10494_);
  and (_02204_, _01616_, _01615_);
  or (_01617_, _09675_, _09347_);
  or (_01618_, _09677_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0]);
  and (_01619_, _01618_, _06444_);
  and (_02236_, _01619_, _01617_);
  or (_01620_, _13931_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0]);
  nand (_01621_, _13931_, _13919_);
  and (_01622_, _01621_, _06444_);
  and (_02250_, _01622_, _01620_);
  and (_01623_, _06449_, \oc8051_top_1.oc8051_indi_addr1.buff[7] [6]);
  nor (_01624_, _10494_, _06449_);
  or (_01625_, _01624_, _01623_);
  and (_02266_, _01625_, _06444_);
  nor (_01626_, _07188_, _09146_);
  and (_01627_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  or (_01628_, _01627_, _07158_);
  or (_01629_, _01628_, _01626_);
  or (_01630_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [4]);
  and (_01631_, _01630_, _06444_);
  and (_02269_, _01631_, _01629_);
  or (_01632_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  and (_01633_, _01632_, _06444_);
  nand (_01634_, _13893_, _07188_);
  and (_02313_, _01634_, _01633_);
  and (_02560_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _06444_);
  or (_01635_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [15]);
  nand (_01636_, _07432_, _13980_);
  and (_01637_, _01636_, _06444_);
  and (_02566_, _01637_, _01635_);
  or (_01638_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [31]);
  nand (_01639_, _07432_, _12633_);
  and (_01640_, _01639_, _06444_);
  and (_02583_, _01640_, _01638_);
  or (_01642_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  and (_01643_, _01642_, _06444_);
  nand (_01644_, _13893_, _07300_);
  and (_02632_, _01644_, _01643_);
  and (_01645_, _09527_, _07148_);
  and (_01646_, _07190_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  or (_01647_, _01646_, _01645_);
  or (_01648_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[6] [0]);
  and (_01649_, _01648_, _06444_);
  and (_02645_, _01649_, _01647_);
  or (_01651_, _14512_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  and (_01652_, _01651_, _06444_);
  nand (_01653_, _14512_, _06978_);
  and (_02649_, _01653_, _01652_);
  nand (_01654_, _14532_, _06978_);
  or (_01655_, _00046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_01656_, _01655_, _00028_);
  and (_01657_, _00046_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_01658_, _01657_, _01656_);
  and (_01659_, _00016_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  and (_01660_, _01659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01661_, _01659_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_01662_, _01661_, _00015_);
  nor (_01663_, _01662_, _01660_);
  and (_01664_, _00052_, _14535_);
  or (_01665_, _01664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nand (_01666_, _01664_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_01667_, _01666_, _01665_);
  and (_01668_, _01667_, _14537_);
  or (_01669_, _01668_, _01663_);
  or (_01670_, _01669_, _01658_);
  or (_01671_, _01670_, _14532_);
  and (_01672_, _01671_, _00040_);
  and (_01673_, _01672_, _01654_);
  and (_01674_, _00039_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01675_, _01674_, _01673_);
  and (_02652_, _01675_, _06444_);
  not (_01677_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 );
  nor (_01678_, _00011_, _01677_);
  or (_01680_, _01678_, _01660_);
  and (_01681_, _01680_, _00015_);
  not (_01682_, _14532_);
  nor (_01683_, _00039_, rst);
  and (_01685_, _01683_, _01682_);
  and (_02658_, _01685_, _01681_);
  nand (_01686_, _00039_, _06978_);
  not (_01687_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  and (_01688_, _00029_, _00002_);
  and (_01689_, _01688_, _01682_);
  nor (_01690_, _01689_, _01687_);
  and (_01691_, _01689_, _01687_);
  or (_01692_, _01691_, _01690_);
  and (_01693_, _00115_, _00002_);
  nand (_01694_, _01693_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  nor (_01695_, _01694_, _14532_);
  or (_01696_, _01695_, _01692_);
  or (_01698_, _01696_, _00039_);
  and (_01699_, _01698_, _06444_);
  and (_02661_, _01699_, _01686_);
  not (_01701_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  nor (_01703_, _14549_, _01701_);
  or (_01704_, _01703_, _01657_);
  and (_01705_, _01704_, _00028_);
  and (_01706_, _00052_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  or (_01707_, _01706_, _01703_);
  and (_01709_, _01707_, _14536_);
  or (_01710_, _01703_, _00003_);
  and (_01711_, _01710_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  or (_01712_, _01711_, _01709_);
  or (_01713_, _01712_, _01705_);
  and (_02664_, _01713_, _01685_);
  and (_01714_, _00517_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  not (_01715_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 );
  nor (_01717_, _00347_, _01715_);
  and (_01718_, _01717_, _00481_);
  or (_01719_, _01718_, _01714_);
  and (_01720_, _00347_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_01721_, _01720_, _00349_);
  and (_01722_, _01721_, _00374_);
  and (_01723_, _01722_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  or (_01724_, _01723_, _01717_);
  and (_01725_, _01724_, _00366_);
  or (_01726_, _01725_, _01719_);
  and (_01727_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_01728_, _01727_, _01717_);
  and (_01729_, _01728_, _00361_);
  or (_01730_, _01729_, _00536_);
  or (_01731_, _01730_, _01726_);
  and (_01732_, _01731_, _06444_);
  nand (_01733_, _01732_, _00388_);
  nor (_02666_, _01733_, _00334_);
  and (_02670_, t0_i, _06444_);
  nand (_01735_, _00334_, _06978_);
  or (_01736_, _00363_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_01737_, _01727_, _00362_);
  and (_01738_, _01737_, _01736_);
  and (_01739_, _00379_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_01740_, _00377_, _00395_);
  nor (_01741_, _01740_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_01742_, _01741_, _01739_);
  or (_01743_, _01742_, _01738_);
  or (_01744_, _01743_, _00334_);
  and (_01745_, _01744_, _00388_);
  and (_01746_, _01745_, _01735_);
  and (_01747_, _00387_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  or (_01748_, _01747_, _01746_);
  and (_02673_, _01748_, _06444_);
  nand (_01749_, _00387_, _06978_);
  nor (_01750_, _00497_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nor (_01751_, _01750_, _00487_);
  and (_01753_, _01751_, _00483_);
  and (_01754_, _00485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  nand (_01755_, _00488_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  nor (_01756_, _01755_, _00334_);
  or (_01757_, _01756_, _01754_);
  or (_01758_, _01757_, _01753_);
  or (_01759_, _01758_, _00387_);
  and (_01760_, _01759_, _06444_);
  and (_02676_, _01760_, _01749_);
  and (_02679_, t1_i, _06444_);
  nand (_01761_, _12829_, _06978_);
  or (_01762_, _12829_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [7]);
  and (_01763_, _01762_, _06444_);
  and (_02763_, _01763_, _01761_);
  and (_01764_, _01079_, _06432_);
  nand (_01765_, _01764_, _06930_);
  or (_01766_, _01764_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  and (_01767_, _01766_, _06674_);
  and (_01768_, _01767_, _01765_);
  nor (_01769_, _01087_, _07069_);
  and (_01770_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_01771_, _01770_, _01769_);
  and (_01772_, _01771_, _06440_);
  and (_01773_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  or (_01774_, _01773_, rst);
  or (_01775_, _01774_, _01772_);
  or (_02879_, _01775_, _01768_);
  and (_01776_, _01079_, _06987_);
  nand (_01777_, _01776_, _06930_);
  or (_01778_, _01776_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  and (_01779_, _01778_, _06674_);
  and (_01780_, _01779_, _01777_);
  nor (_01781_, _01087_, _06666_);
  and (_01782_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_01783_, _01782_, _01781_);
  and (_01784_, _01783_, _06440_);
  and (_01785_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  or (_01787_, _01785_, rst);
  or (_01788_, _01787_, _01784_);
  or (_02881_, _01788_, _01780_);
  and (_01789_, _08913_, _06432_);
  nand (_01791_, _01789_, _06930_);
  or (_01792_, _01789_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  and (_01793_, _01792_, _06674_);
  and (_01794_, _01793_, _01791_);
  and (_01795_, _08919_, _07070_);
  and (_01796_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_01797_, _01796_, _01795_);
  and (_01798_, _01797_, _06440_);
  and (_01799_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  or (_01800_, _01799_, rst);
  or (_01801_, _01800_, _01798_);
  or (_02883_, _01801_, _01794_);
  and (_01802_, _08913_, _06987_);
  nand (_01804_, _01802_, _06930_);
  or (_01805_, _01802_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  and (_01807_, _01805_, _06674_);
  and (_01809_, _01807_, _01804_);
  nor (_01811_, _08920_, _06666_);
  and (_01812_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_01813_, _01812_, _01811_);
  and (_01814_, _01813_, _06440_);
  and (_01815_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  or (_01816_, _01815_, rst);
  or (_01817_, _01816_, _01814_);
  or (_02886_, _01817_, _01809_);
  and (_01818_, _00605_, _08977_);
  nand (_01819_, _01818_, _06930_);
  or (_01820_, _01818_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_01821_, _01820_, _06674_);
  and (_01822_, _01821_, _01819_);
  nand (_01823_, _11589_, _00612_);
  or (_01824_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  and (_01825_, _01824_, _06440_);
  and (_01826_, _01825_, _01823_);
  and (_01827_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  or (_01828_, _01827_, rst);
  or (_01829_, _01828_, _01826_);
  or (_02888_, _01829_, _01822_);
  and (_01830_, _00640_, _06987_);
  nand (_01831_, _01830_, _06930_);
  or (_01832_, _01830_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01833_, _01832_, _06674_);
  and (_01834_, _01833_, _01831_);
  nand (_01835_, _00646_, _06666_);
  or (_01836_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  and (_01837_, _01836_, _06440_);
  and (_01838_, _01837_, _01835_);
  and (_01839_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  or (_01840_, _01839_, rst);
  or (_01841_, _01840_, _01838_);
  or (_02890_, _01841_, _01834_);
  and (_01842_, _07402_, _07043_);
  nand (_01843_, _01842_, _06930_);
  or (_01844_, _01842_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_01845_, _01844_, _06674_);
  and (_01847_, _01845_, _01843_);
  nand (_01848_, _00646_, _07069_);
  or (_01850_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  and (_01851_, _01850_, _06440_);
  and (_01852_, _01851_, _01848_);
  and (_01853_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  or (_01855_, _01853_, rst);
  or (_01856_, _01855_, _01852_);
  or (_02893_, _01856_, _01847_);
  and (_01857_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nor (_01858_, _08064_, _01150_);
  or (_01859_, _01858_, _01857_);
  and (_02898_, _01859_, _06444_);
  and (_01860_, _06934_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  or (_01861_, _01860_, _06935_);
  and (_01862_, _01861_, _12012_);
  nand (_01863_, _12008_, _06930_);
  nor (_01864_, _12008_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  nor (_01865_, _01864_, _12012_);
  and (_01866_, _01865_, _01863_);
  or (_01867_, _01866_, _07218_);
  or (_01868_, _01867_, _01862_);
  nand (_01869_, _07218_, _06978_);
  and (_01870_, _01869_, _06444_);
  and (_02905_, _01870_, _01868_);
  and (_01871_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  not (_01872_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nor (_01873_, _08064_, _01872_);
  or (_01874_, _01873_, _01871_);
  and (_02908_, _01874_, _06444_);
  and (_01875_, _01079_, _06942_);
  nand (_01876_, _01875_, _06930_);
  or (_01877_, _01875_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  and (_01878_, _01877_, _06674_);
  and (_01879_, _01878_, _01876_);
  and (_01880_, _01086_, _09527_);
  and (_01881_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_01882_, _01881_, _01880_);
  and (_01883_, _01882_, _06440_);
  and (_01884_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  or (_01885_, _01884_, rst);
  or (_01886_, _01885_, _01883_);
  or (_02914_, _01886_, _01879_);
  and (_01887_, _01079_, _08310_);
  nand (_01888_, _01887_, _06930_);
  or (_01889_, _01887_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  and (_01890_, _01889_, _06674_);
  and (_01891_, _01890_, _01888_);
  nor (_01892_, _01087_, _07300_);
  and (_01893_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_01894_, _01893_, _01892_);
  and (_01895_, _01894_, _06440_);
  and (_01896_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  or (_01897_, _01896_, rst);
  or (_01898_, _01897_, _01895_);
  or (_02916_, _01898_, _01891_);
  and (_01899_, _00605_, _00240_);
  nand (_01900_, _01899_, _06930_);
  or (_01901_, _01899_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_01902_, _01901_, _06674_);
  and (_01903_, _01902_, _01900_);
  nand (_01904_, _10494_, _00612_);
  or (_01905_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  and (_01906_, _01905_, _06440_);
  and (_01907_, _01906_, _01904_);
  and (_01908_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  or (_01909_, _01908_, rst);
  or (_01910_, _01909_, _01907_);
  or (_02919_, _01910_, _01903_);
  nand (_01911_, _00612_, _06930_);
  or (_01912_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  and (_01913_, _01912_, _06674_);
  and (_01914_, _01913_, _01911_);
  nand (_01915_, _09526_, _00612_);
  and (_01916_, _01915_, _06440_);
  and (_01917_, _01916_, _01912_);
  and (_01918_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  or (_01919_, _01918_, rst);
  or (_01920_, _01919_, _01917_);
  or (_02921_, _01920_, _01914_);
  nand (_01921_, _00646_, _06930_);
  or (_01922_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  and (_01923_, _01922_, _06674_);
  and (_01924_, _01923_, _01921_);
  nand (_01925_, _09526_, _00646_);
  and (_01926_, _01922_, _06440_);
  and (_01927_, _01926_, _01925_);
  and (_01928_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  or (_01929_, _01928_, rst);
  or (_01930_, _01929_, _01927_);
  or (_02924_, _01930_, _01924_);
  and (_01931_, _00640_, _08310_);
  nand (_01932_, _01931_, _06930_);
  or (_01933_, _01931_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_01934_, _01933_, _06674_);
  and (_01935_, _01934_, _01932_);
  nand (_01937_, _00646_, _07300_);
  or (_01938_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  and (_01939_, _01938_, _06440_);
  and (_01940_, _01939_, _01937_);
  and (_01941_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  or (_01942_, _01941_, rst);
  or (_01943_, _01942_, _01940_);
  or (_02926_, _01943_, _01935_);
  and (_01944_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  nor (_01945_, _08064_, _01076_);
  or (_01946_, _01945_, _01944_);
  and (_02945_, _01946_, _06444_);
  nand (_01947_, _12829_, _09526_);
  or (_01948_, _12829_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [0]);
  and (_01949_, _01948_, _01947_);
  and (_03036_, _01949_, _06444_);
  and (_01950_, _00605_, _06987_);
  nand (_01951_, _01950_, _06930_);
  or (_01952_, _01950_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_01953_, _01952_, _06674_);
  and (_01954_, _01953_, _01951_);
  nand (_01955_, _00612_, _06666_);
  or (_01956_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  and (_01957_, _01956_, _06440_);
  and (_01958_, _01957_, _01955_);
  and (_01959_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  or (_01960_, _01959_, rst);
  or (_01961_, _01960_, _01958_);
  or (_03040_, _01961_, _01954_);
  and (_01962_, _00605_, _06983_);
  nand (_01963_, _01962_, _06930_);
  or (_01964_, _01962_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_01965_, _01964_, _06674_);
  and (_01966_, _01965_, _01963_);
  nand (_01967_, _00612_, _07188_);
  or (_01968_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  and (_01969_, _01968_, _06440_);
  and (_01970_, _01969_, _01967_);
  and (_01971_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  or (_01972_, _01971_, rst);
  or (_01973_, _01972_, _01970_);
  or (_03042_, _01973_, _01966_);
  and (_01975_, _08913_, _06983_);
  nand (_01976_, _01975_, _06930_);
  or (_01977_, _01975_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  and (_01978_, _01977_, _06674_);
  and (_01979_, _01978_, _01976_);
  nor (_01980_, _08920_, _07188_);
  and (_01981_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_01982_, _01981_, _01980_);
  and (_01983_, _01982_, _06440_);
  and (_01984_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  or (_01985_, _01984_, rst);
  or (_01986_, _01985_, _01983_);
  or (_03044_, _01986_, _01979_);
  and (_01987_, _08913_, _08310_);
  nand (_01988_, _01987_, _06930_);
  or (_01989_, _01987_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  and (_01990_, _01989_, _06674_);
  and (_01991_, _01990_, _01988_);
  nor (_01992_, _08920_, _07300_);
  and (_01993_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_01994_, _01993_, _01992_);
  and (_01995_, _01994_, _06440_);
  and (_01996_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  or (_01997_, _01996_, rst);
  or (_01998_, _01997_, _01995_);
  or (_03046_, _01998_, _01991_);
  nand (_01999_, _13890_, _11589_);
  or (_02000_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  and (_02001_, _02000_, _06444_);
  and (_03049_, _02001_, _01999_);
  nand (_02002_, _13890_, _07069_);
  or (_02003_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  and (_02004_, _02003_, _06444_);
  and (_03061_, _02004_, _02002_);
  and (_02005_, _00640_, _00240_);
  nand (_02006_, _02005_, _06930_);
  or (_02007_, _02005_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02008_, _02007_, _06674_);
  and (_02009_, _02008_, _02006_);
  nand (_02010_, _10494_, _00646_);
  or (_02011_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  and (_02012_, _02011_, _06440_);
  and (_02014_, _02012_, _02010_);
  and (_02015_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  or (_02016_, _02015_, rst);
  or (_02017_, _02016_, _02014_);
  or (_03070_, _02017_, _02009_);
  and (_02018_, _00640_, _06983_);
  nand (_02019_, _02018_, _06930_);
  or (_02020_, _02018_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02021_, _02020_, _06674_);
  and (_02022_, _02021_, _02019_);
  nand (_02023_, _00646_, _07188_);
  or (_02024_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  and (_02025_, _02024_, _06440_);
  and (_02026_, _02025_, _02023_);
  and (_02027_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  or (_02028_, _02027_, rst);
  or (_02029_, _02028_, _02026_);
  or (_03072_, _02029_, _02022_);
  not (_02030_, _00640_);
  or (_02031_, _02030_, _00717_);
  and (_02032_, _02031_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02033_, _06431_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_02034_, _02033_, _00713_);
  and (_02035_, _02034_, _00640_);
  or (_02036_, _02035_, _02032_);
  and (_02037_, _02036_, _06674_);
  nand (_02038_, _11589_, _00646_);
  or (_02039_, _00646_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  and (_02040_, _02039_, _06440_);
  and (_02041_, _02040_, _02038_);
  and (_02043_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  or (_02044_, _02043_, rst);
  or (_02045_, _02044_, _02041_);
  or (_03074_, _02045_, _02037_);
  and (_02047_, _00605_, _08310_);
  nand (_02048_, _02047_, _06930_);
  or (_02049_, _02047_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02050_, _02049_, _06674_);
  and (_02051_, _02050_, _02048_);
  nand (_02052_, _00612_, _07300_);
  or (_02053_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  and (_02054_, _02053_, _06440_);
  and (_02055_, _02054_, _02052_);
  and (_02056_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  or (_02057_, _02056_, rst);
  or (_02058_, _02057_, _02055_);
  or (_03076_, _02058_, _02051_);
  and (_02059_, _08913_, _00240_);
  nand (_02060_, _02059_, _06930_);
  or (_02061_, _02059_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  and (_02062_, _02061_, _06674_);
  and (_02063_, _02062_, _02060_);
  nor (_02064_, _10494_, _08920_);
  and (_02065_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02066_, _02065_, _02064_);
  and (_02067_, _02066_, _06440_);
  and (_02068_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  or (_02069_, _02068_, rst);
  or (_02070_, _02069_, _02067_);
  or (_03078_, _02070_, _02063_);
  and (_02071_, _00605_, _06432_);
  nand (_02072_, _02071_, _06930_);
  or (_02073_, _02071_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  and (_02074_, _02073_, _06674_);
  and (_02075_, _02074_, _02072_);
  or (_02076_, _00612_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  nand (_02077_, _00612_, _07069_);
  and (_02078_, _02077_, _06440_);
  and (_02079_, _02078_, _02076_);
  and (_02080_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  or (_02081_, _02080_, rst);
  or (_02082_, _02081_, _02079_);
  or (_03080_, _02082_, _02075_);
  and (_02083_, _08913_, _08977_);
  nand (_02084_, _02083_, _06930_);
  or (_02085_, _02083_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  and (_02086_, _02085_, _06674_);
  and (_02087_, _02086_, _02084_);
  nor (_02088_, _11589_, _08920_);
  and (_02089_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02091_, _02089_, _02088_);
  and (_02092_, _02091_, _06440_);
  and (_02093_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  or (_02094_, _02093_, rst);
  or (_02095_, _02094_, _02092_);
  or (_03081_, _02095_, _02087_);
  nand (_02096_, _08919_, _06930_);
  or (_02097_, _08919_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  and (_02098_, _02097_, _06674_);
  and (_02099_, _02098_, _02096_);
  and (_02100_, _09527_, _08919_);
  and (_02101_, _08920_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_02102_, _02101_, _02100_);
  and (_02103_, _02102_, _06440_);
  and (_02104_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  or (_02105_, _02104_, rst);
  or (_02106_, _02105_, _02103_);
  or (_03084_, _02106_, _02099_);
  and (_02107_, _01079_, _00240_);
  nand (_02108_, _02107_, _06930_);
  or (_02109_, _02107_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  and (_02110_, _02109_, _06674_);
  and (_02111_, _02110_, _02108_);
  nor (_02112_, _01087_, _10494_);
  and (_02113_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_02114_, _02113_, _02112_);
  and (_02115_, _02114_, _06440_);
  and (_02116_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  or (_02117_, _02116_, rst);
  or (_02118_, _02117_, _02115_);
  or (_03086_, _02118_, _02111_);
  and (_02119_, _01079_, _06983_);
  nand (_02120_, _02119_, _06930_);
  or (_02121_, _02119_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  and (_02122_, _02121_, _06674_);
  and (_02123_, _02122_, _02120_);
  nor (_02124_, _01087_, _07188_);
  and (_02125_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_02126_, _02125_, _02124_);
  and (_02127_, _02126_, _06440_);
  and (_02128_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  or (_02129_, _02128_, rst);
  or (_02130_, _02129_, _02127_);
  or (_03088_, _02130_, _02123_);
  and (_02131_, _01079_, _08977_);
  nand (_02132_, _02131_, _06930_);
  or (_02133_, _02131_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  and (_02134_, _02133_, _06674_);
  and (_02135_, _02134_, _02132_);
  nor (_02136_, _01087_, _11589_);
  and (_02137_, _01087_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_02138_, _02137_, _02136_);
  and (_02139_, _02138_, _06440_);
  and (_02140_, _08925_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  or (_02141_, _02140_, rst);
  or (_02142_, _02141_, _02139_);
  or (_03091_, _02142_, _02135_);
  nand (_02143_, _13890_, _09526_);
  or (_02144_, _13890_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  and (_02145_, _02144_, _06444_);
  and (_03118_, _02145_, _02143_);
  and (_03132_, _01286_, _06444_);
  and (_03406_, \oc8051_top_1.oc8051_memory_interface1.istb_t , _06444_);
  and (_02147_, _03406_, \oc8051_top_1.oc8051_memory_interface1.imem_wait );
  or (_03144_, _02147_, _03132_);
  or (_02148_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [13]);
  nand (_02149_, _07432_, _13990_);
  and (_02150_, _02149_, _06444_);
  and (_03147_, _02150_, _02148_);
  nand (_02151_, _07226_, \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  and (_03150_, _02151_, _06444_);
  and (_03196_, _00287_, _11574_);
  and (_03293_, _07982_, _06444_);
  nor (_02152_, _07432_, _07429_);
  nand (_02153_, _01135_, _01132_);
  and (_02154_, _02153_, _07230_);
  and (_02155_, _02154_, _07235_);
  nor (_02156_, _02154_, _07235_);
  nor (_02157_, _02156_, _02155_);
  nor (_02158_, _02157_, _02152_);
  and (_02159_, _07240_, \oc8051_top_1.oc8051_memory_interface1.op_pos [2]);
  and (_02160_, _02159_, _02152_);
  and (_02161_, _02160_, _10890_);
  or (_02162_, _02161_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02163_, _02162_, _02158_);
  and (_03295_, _02163_, _06444_);
  and (_03300_, _11622_, _06444_);
  and (_02164_, _12712_, \oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7]);
  or (_02165_, _02164_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  and (_03304_, _02165_, _06444_);
  and (_03307_, _01491_, _06444_);
  not (_02166_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  nand (_02167_, _07230_, _02166_);
  nand (_02168_, _02167_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t );
  nand (_02169_, _02168_, _12712_);
  and (_03309_, _02169_, _06444_);
  and (_02170_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [0]);
  and (_02171_, _12841_, _07154_);
  or (_02172_, _02171_, _02170_);
  and (_03321_, _02172_, _06444_);
  nor (_02173_, _12830_, _07188_);
  and (_02174_, _01100_, \oc8051_top_1.oc8051_indi_addr1.buff[2] [4]);
  or (_02175_, _02174_, _02173_);
  and (_03325_, _02175_, _06444_);
  and (_03331_, \oc8051_top_1.oc8051_memory_interface1.int_ack_t , _06444_);
  and (_02176_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [4]);
  nor (_02177_, _07188_, _07046_);
  or (_02178_, _02177_, _02176_);
  and (_03344_, _02178_, _06444_);
  nor (_03350_, _01510_, rst);
  nor (_02179_, _10946_, _10944_);
  nor (_02180_, _02179_, _10947_);
  or (_02181_, _02180_, _08374_);
  or (_02182_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  and (_02183_, _02182_, _10894_);
  and (_02184_, _02183_, _02181_);
  and (_02185_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  or (_03355_, _02185_, _02184_);
  and (_02186_, _14069_, _07070_);
  and (_02187_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [1]);
  or (_02188_, _02187_, _02186_);
  and (_03357_, _02188_, _06444_);
  or (_02189_, _10942_, _10940_);
  and (_02190_, _02189_, _10943_);
  or (_02192_, _02190_, _08374_);
  or (_02193_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  and (_02194_, _02193_, _10894_);
  and (_02195_, _02194_, _02192_);
  and (_02196_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  or (_03360_, _02196_, _02195_);
  nor (_02197_, _10939_, _10891_);
  nor (_02198_, _02197_, _10940_);
  or (_02199_, _02198_, _08374_);
  or (_02200_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  and (_02201_, _02200_, _10894_);
  and (_02202_, _02201_, _02199_);
  and (_02203_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  or (_03385_, _02203_, _02202_);
  not (_02205_, _00599_);
  and (_02206_, _02205_, _00597_);
  and (_02207_, _00278_, _00592_);
  and (_03398_, _02207_, _02206_);
  and (_02208_, \oc8051_top_1.oc8051_memory_interface1.cdata [7], _08478_);
  and (_02209_, \oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_top_1.oc8051_memory_interface1.istb_t );
  or (_02210_, _02209_, _02208_);
  and (_03414_, _02210_, _06444_);
  and (_02211_, _11763_, _07425_);
  and (_02212_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_02213_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [6]);
  and (_02214_, _02213_, _09332_);
  or (_02215_, _02214_, _02212_);
  or (_02216_, _02215_, _02211_);
  and (_03425_, _02216_, _06444_);
  and (_02217_, _08421_, _08356_);
  and (_02218_, _02217_, _08453_);
  and (_02219_, _08437_, _08405_);
  and (_02220_, _02219_, _08468_);
  and (_02221_, _07231_, _06444_);
  and (_02222_, _02221_, _08388_);
  and (_02223_, _02222_, _07259_);
  and (_02224_, _02223_, _02220_);
  and (_03428_, _02224_, _02218_);
  nor (_02225_, _14070_, _06666_);
  and (_02226_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [5]);
  or (_02227_, _02226_, _02225_);
  and (_03429_, _02227_, _06444_);
  or (_02228_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [19]);
  nand (_02229_, _07432_, _11264_);
  and (_02230_, _02229_, _06444_);
  and (_03460_, _02230_, _02228_);
  and (_02231_, _13934_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2]);
  and (_02232_, _09678_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done );
  and (_02233_, _02232_, _13933_);
  or (_02234_, _02233_, _02231_);
  and (_03483_, _02234_, _06444_);
  and (_02235_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [21]);
  and (_02237_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [21]);
  or (_02238_, _02237_, _02235_);
  and (_03495_, _02238_, _06444_);
  and (_02239_, _07432_, \oc8051_top_1.oc8051_memory_interface1.idat_cur [20]);
  and (_02240_, _12223_, \oc8051_top_1.oc8051_rom1.data_o [20]);
  or (_02241_, _02240_, _02239_);
  and (_03502_, _02241_, _06444_);
  not (_02242_, _00850_);
  or (_02243_, _02242_, _07198_);
  and (_02244_, _00850_, _07208_);
  and (_02245_, _02244_, _07206_);
  or (_02246_, _02245_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2]);
  and (_02247_, _02246_, _06444_);
  and (_03515_, _02247_, _02243_);
  nor (_03523_, _11570_, rst);
  nor (_03532_, _07222_, rst);
  and (_02248_, _11443_, _11385_);
  and (_02249_, _11408_, _11394_);
  or (_02251_, _02249_, _11483_);
  or (_02252_, _02251_, _02248_);
  and (_02253_, _11394_, _11523_);
  and (_02254_, _11394_, _11493_);
  and (_02255_, _11394_, _11458_);
  or (_02256_, _02255_, _02254_);
  or (_02257_, _02256_, _02253_);
  or (_02258_, _11519_, _11394_);
  and (_02259_, _02258_, _11418_);
  and (_02260_, _11426_, _11355_);
  or (_02261_, _02260_, _02259_);
  or (_02262_, _02261_, _02257_);
  and (_02263_, _11433_, _11965_);
  and (_02264_, _11443_, _11965_);
  or (_02265_, _02264_, _02263_);
  or (_02267_, _02265_, _11379_);
  and (_02268_, _11370_, _11423_);
  and (_02270_, _11528_, _11418_);
  or (_02271_, _14240_, _02270_);
  or (_02272_, _02271_, _02268_);
  or (_02273_, _02272_, _02267_);
  or (_02274_, _02273_, _02262_);
  and (_02275_, _11431_, _11965_);
  and (_02276_, _11407_, _11976_);
  and (_02277_, _11431_, _11526_);
  or (_02278_, _02277_, _02276_);
  and (_02279_, _11370_, _11976_);
  or (_02280_, _02279_, _11439_);
  or (_02281_, _02280_, _02278_);
  or (_02282_, _02281_, _02275_);
  and (_02283_, _11394_, _11475_);
  or (_02284_, _02283_, _14234_);
  and (_02285_, _11519_, _11407_);
  or (_02286_, _02285_, _11537_);
  or (_02287_, _02286_, _02284_);
  or (_02288_, _14225_, _14228_);
  or (_02289_, _02288_, _02287_);
  or (_02290_, _02289_, _02282_);
  or (_02291_, _02290_, _02274_);
  or (_02292_, _02291_, _02252_);
  and (_02293_, _02292_, _07230_);
  and (_02294_, \oc8051_top_1.oc8051_decoder1.wr_sfr [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  not (_02295_, \oc8051_top_1.oc8051_decoder1.state [1]);
  and (_02296_, _11453_, _02295_);
  and (_02297_, _11370_, _11355_);
  nor (_02298_, _11385_, _11354_);
  not (_02299_, _02298_);
  and (_02300_, _02299_, _11419_);
  nor (_02301_, _02300_, _02297_);
  not (_02302_, _02301_);
  and (_02303_, _02302_, _02296_);
  or (_02304_, _02303_, _02294_);
  or (_02305_, _02304_, _02293_);
  and (_03537_, _02305_, _06444_);
  and (_02306_, _06444_, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_02307_, _02306_, \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  or (_02308_, _11394_, _11526_);
  and (_02309_, _02308_, _11486_);
  and (_02310_, _11528_, _11373_);
  or (_02311_, _02310_, _11442_);
  or (_02312_, _02311_, _11424_);
  or (_02314_, _02312_, _02309_);
  not (_02315_, _11430_);
  or (_02316_, _11995_, _02315_);
  nand (_02317_, _02316_, _11505_);
  or (_02318_, _02317_, _02314_);
  or (_02319_, _02318_, _02252_);
  or (_02320_, _02264_, _14225_);
  or (_02321_, _02320_, _02263_);
  and (_02322_, _02321_, _07311_);
  and (_02323_, _11519_, _11411_);
  or (_02324_, _14234_, _02323_);
  and (_02325_, _11395_, _11355_);
  or (_02326_, _11419_, _11431_);
  and (_02327_, _02326_, _11394_);
  or (_02328_, _02327_, _02325_);
  or (_02329_, _02328_, _02324_);
  or (_02330_, _02329_, _02322_);
  or (_02331_, _02330_, _02319_);
  and (_02332_, _07230_, _06444_);
  and (_02333_, _02332_, _02331_);
  or (_03545_, _02333_, _02307_);
  and (_02334_, \oc8051_top_1.oc8051_decoder1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_02335_, _02334_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  and (_02336_, _06870_, _06847_);
  and (_02337_, _06838_, _06680_);
  nand (_02338_, _06640_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  nand (_02339_, _02338_, _02334_);
  or (_02340_, _02339_, _02337_);
  or (_02341_, _02340_, _02336_);
  and (_02342_, _02341_, _02335_);
  or (_02343_, _02342_, _12012_);
  or (_02344_, _00240_, _08294_);
  nand (_02345_, _02344_, _12012_);
  or (_02346_, _02345_, _01481_);
  and (_02347_, _02346_, _02343_);
  or (_02348_, _02347_, _07218_);
  nand (_02349_, _10494_, _07218_);
  and (_02350_, _02349_, _06444_);
  and (_03547_, _02350_, _02348_);
  and (_02351_, _11459_, _11389_);
  not (_02352_, _11399_);
  and (_02353_, _02352_, _02296_);
  and (_02354_, _11934_, _11347_);
  and (_02355_, _11933_, _11347_);
  or (_02356_, _02355_, _02354_);
  and (_02357_, _02356_, _11389_);
  or (_02358_, _02357_, _02353_);
  or (_02359_, _02358_, _02351_);
  and (_02360_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02361_, _11524_, _11494_);
  or (_02362_, _02361_, _11509_);
  not (_02363_, _11354_);
  nor (_02364_, _11995_, _02363_);
  or (_02365_, _02364_, _02354_);
  or (_02366_, _02365_, _02362_);
  and (_02367_, _11482_, _11347_);
  and (_02368_, _02367_, _11417_);
  or (_02369_, _11534_, _11504_);
  or (_02370_, _02369_, _02368_);
  nor (_02371_, _11495_, _11413_);
  nand (_02372_, _02371_, _11492_);
  or (_02373_, _02372_, _02370_);
  or (_02374_, _02373_, _02366_);
  not (_02375_, _11513_);
  nand (_02376_, _02375_, _11416_);
  and (_02377_, _11519_, _11370_);
  or (_02378_, _02377_, _02355_);
  or (_02379_, _02378_, _02376_);
  or (_02380_, _02379_, _02374_);
  and (_02381_, _02380_, _07230_);
  or (_02382_, _02381_, _02360_);
  or (_02383_, _02382_, _02359_);
  and (_03554_, _02383_, _06444_);
  and (_02384_, _11423_, _11417_);
  or (_02385_, _11529_, _11428_);
  or (_02386_, _02385_, _02384_);
  and (_02387_, _11413_, _11376_);
  or (_02388_, _02387_, _11442_);
  or (_02389_, _02388_, _02356_);
  or (_02390_, _02389_, _02386_);
  and (_02391_, _02390_, _07230_);
  and (_02392_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02393_, _02392_, _02358_);
  or (_02394_, _02393_, _02391_);
  and (_03573_, _02394_, _06444_);
  nand (_02395_, _01480_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  nand (_02396_, _02395_, _06678_);
  or (_02397_, _02396_, _01481_);
  and (_02398_, _07015_, _06981_);
  or (_02399_, _02398_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_02400_, _02399_, _06678_);
  and (_02401_, _02400_, _02397_);
  or (_02402_, _02401_, _06946_);
  nand (_02403_, _10494_, _06946_);
  and (_02404_, _02403_, _06444_);
  and (_03597_, _02404_, _02402_);
  and (_02405_, _07147_, _06440_);
  and (_02406_, _02405_, _06941_);
  and (_02407_, _06987_, _06678_);
  nand (_02408_, _02407_, _06930_);
  or (_02409_, _02407_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  and (_02410_, _02409_, _02408_);
  or (_02411_, _02410_, _02406_);
  nand (_02412_, _06946_, _06666_);
  and (_02413_, _02412_, _06444_);
  and (_03599_, _02413_, _02411_);
  and (_02414_, _06983_, _06678_);
  nand (_02415_, _02414_, _06930_);
  not (_02416_, _06946_);
  or (_02417_, _02414_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_02418_, _02417_, _02416_);
  and (_02419_, _02418_, _02415_);
  nor (_02420_, _07188_, _02416_);
  or (_02421_, _02420_, _02419_);
  and (_03606_, _02421_, _06444_);
  and (_02422_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_02423_, _10956_, _10920_);
  nor (_02424_, _02423_, _10957_);
  or (_02425_, _02424_, _08374_);
  or (_02426_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  and (_02427_, _02426_, _10894_);
  and (_02428_, _02427_, _02425_);
  or (_03621_, _02428_, _02422_);
  nor (_03623_, _11402_, rst);
  nand (_02429_, _02332_, _11418_);
  or (_03625_, _02429_, _02298_);
  and (_02430_, _10839_, _10751_);
  and (_02431_, _02430_, _10836_);
  and (_02432_, _10850_, _10746_);
  and (_02433_, _10874_, _10836_);
  or (_02434_, _02433_, _02432_);
  or (_02435_, _02434_, _02431_);
  nor (_02436_, _10884_, _10848_);
  nand (_02437_, _02436_, _10786_);
  or (_02438_, _02437_, _02435_);
  nand (_02439_, _10822_, _10776_);
  or (_02440_, _02439_, _02438_);
  and (_02441_, _10820_, _10753_);
  and (_02442_, _10743_, _08425_);
  and (_02443_, _10739_, _08457_);
  and (_02444_, _10770_, _02443_);
  or (_02445_, _02444_, _02442_);
  or (_02446_, _02445_, _02441_);
  or (_02447_, _10831_, _10826_);
  and (_02448_, _10799_, _10753_);
  and (_02449_, _02448_, _10812_);
  and (_02450_, _10736_, _10812_);
  and (_02451_, _10782_, _02450_);
  and (_02452_, _10736_, _10741_);
  and (_02453_, _10850_, _02452_);
  or (_02454_, _02453_, _02451_);
  or (_02455_, _02454_, _02449_);
  or (_02456_, _02455_, _02447_);
  or (_02457_, _02456_, _02446_);
  or (_02458_, _02457_, _02440_);
  and (_02459_, _02458_, _07231_);
  and (_02460_, _07228_, _06308_);
  and (_02461_, _02460_, _11386_);
  nor (_02462_, _02461_, _02295_);
  or (_02463_, _02462_, rst);
  or (_03627_, _02463_, _02459_);
  not (_02464_, _07229_);
  or (_02465_, _08360_, _02464_);
  or (_02466_, _07229_, \oc8051_top_1.oc8051_decoder1.op [7]);
  and (_02467_, _02466_, _06444_);
  and (_03630_, _02467_, _02465_);
  and (_02468_, _02306_, \oc8051_top_1.oc8051_decoder1.src_sel3 );
  and (_02469_, _11490_, _11355_);
  or (_02470_, _02469_, _11986_);
  and (_02471_, _11419_, _11394_);
  and (_02472_, _11493_, _11354_);
  or (_02473_, _02472_, _02471_);
  or (_02474_, _02473_, _02470_);
  or (_02475_, _11491_, _12040_);
  or (_02476_, _02475_, _02325_);
  nor (_02477_, _02476_, _02474_);
  nand (_02478_, _02477_, _11461_);
  and (_02479_, _02478_, _02332_);
  or (_03632_, _02479_, _02468_);
  or (_02480_, _02248_, _11379_);
  and (_02481_, _11519_, _11412_);
  or (_02482_, _02481_, _11442_);
  and (_02483_, _11490_, _11965_);
  or (_02484_, _02483_, _02482_);
  or (_02485_, _02484_, _02480_);
  and (_02486_, _02485_, _07230_);
  and (_02487_, \oc8051_top_1.oc8051_decoder1.wr_sfr [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02488_, _02487_, _02353_);
  or (_02489_, _02488_, _02486_);
  and (_03634_, _02489_, _06444_);
  and (_02490_, _02306_, \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  and (_02491_, _11443_, _11394_);
  not (_02492_, _11429_);
  and (_02493_, _11427_, _11526_);
  or (_02494_, _02493_, _14239_);
  or (_02495_, _02494_, _02492_);
  or (_02496_, _02495_, _02491_);
  and (_02497_, _11965_, _11458_);
  or (_02498_, _02361_, _02253_);
  or (_02499_, _02498_, _02497_);
  or (_02500_, _02480_, _02309_);
  or (_02501_, _02500_, _02499_);
  or (_02502_, _02501_, _02496_);
  and (_02503_, _02502_, _02332_);
  or (_03637_, _02503_, _02490_);
  and (_02504_, _12012_, _06987_);
  nand (_02505_, _02504_, _06930_);
  or (_02506_, _02504_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_02507_, _02506_, _07219_);
  and (_02508_, _02507_, _02505_);
  nor (_02509_, _07219_, _06666_);
  or (_02510_, _02509_, _02508_);
  and (_03640_, _02510_, _06444_);
  and (_02511_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_02512_, _02511_, _07026_);
  and (_02513_, _07011_, _06994_);
  or (_02514_, _02513_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  nand (_02515_, _07011_, _06995_);
  and (_02516_, _02515_, _02514_);
  or (_02517_, _02516_, _02512_);
  and (_02518_, _02517_, _07035_);
  and (_02519_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_02520_, _02519_, _06985_);
  or (_02521_, _02520_, _02518_);
  nand (_02522_, _07188_, _06985_);
  and (_02523_, _02522_, _09503_);
  and (_02524_, _02523_, _02521_);
  and (_02525_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_02526_, _02525_, _02524_);
  and (_03644_, _02526_, _06444_);
  and (_02527_, \oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_02528_, _11534_, _07230_);
  or (_02529_, _02528_, _02527_);
  or (_02530_, _02529_, _02353_);
  and (_03646_, _02530_, _06444_);
  or (_02531_, _02356_, _02325_);
  and (_02532_, _02531_, _11342_);
  or (_02533_, _02303_, \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02534_, _02533_, _02357_);
  or (_02535_, _02534_, _02532_);
  or (_02536_, \oc8051_top_1.oc8051_decoder1.src_sel1 [2], _06308_);
  and (_02537_, _02536_, _06444_);
  and (_03648_, _02537_, _02535_);
  not (_02538_, _06985_);
  and (_02539_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_02540_, _07011_, _06993_);
  nor (_02541_, _02540_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  nor (_02542_, _02541_, _02513_);
  and (_02543_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_02544_, _02543_, _07026_);
  or (_02545_, _02544_, _02542_);
  and (_02546_, _02545_, _07035_);
  or (_02547_, _02546_, _02539_);
  and (_02548_, _02547_, _02538_);
  nor (_02549_, _07300_, _02538_);
  or (_02550_, _02549_, _06989_);
  or (_02551_, _02550_, _02548_);
  or (_02552_, _09503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  and (_02553_, _02552_, _06444_);
  and (_03651_, _02553_, _02551_);
  and (_02554_, _02306_, \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  or (_02555_, _11412_, _11427_);
  and (_02556_, _02555_, _11976_);
  or (_02557_, _11379_, _11494_);
  or (_02558_, _02557_, _02556_);
  or (_02559_, _02481_, _11504_);
  or (_02561_, _11533_, _11489_);
  or (_02562_, _02561_, _02559_);
  or (_02563_, _02472_, _02497_);
  and (_02564_, _11490_, _11406_);
  and (_02565_, _11406_, _11458_);
  or (_02567_, _02565_, _02564_);
  or (_02568_, _02567_, _02563_);
  or (_02569_, _02568_, _02562_);
  or (_02570_, _02569_, _02558_);
  and (_02571_, _02570_, _02332_);
  or (_03653_, _02571_, _02554_);
  and (_02572_, _02306_, \oc8051_top_1.oc8051_decoder1.alu_op [3]);
  not (_02573_, _11478_);
  or (_02574_, _02249_, _02573_);
  or (_02575_, _02311_, _02260_);
  or (_02576_, _02575_, _02494_);
  nor (_02577_, _02576_, _02574_);
  and (_02578_, _02577_, _11488_);
  or (_02579_, _02483_, _02263_);
  nor (_02580_, _02579_, _02324_);
  nand (_02581_, _02580_, _11484_);
  nor (_02582_, _02581_, _02499_);
  and (_02584_, _02582_, _14230_);
  nand (_02585_, _02584_, _02578_);
  and (_02586_, _02585_, _02332_);
  or (_03656_, _02586_, _02572_);
  or (_02587_, _02275_, _02268_);
  or (_02588_, _02280_, _02277_);
  or (_02589_, _02588_, _02587_);
  or (_02590_, _02264_, _02352_);
  or (_02591_, _02590_, _02589_);
  and (_02592_, _02591_, _02332_);
  nor (_02593_, _11399_, _11342_);
  and (_02594_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02595_, _02594_, _02593_);
  and (_02596_, _02595_, _06444_);
  or (_03658_, _02596_, _02592_);
  and (_02597_, _11976_, _11417_);
  or (_02598_, _02597_, _02355_);
  and (_02599_, _11519_, _11369_);
  or (_02600_, _02599_, _02482_);
  or (_02601_, _02600_, _02598_);
  or (_02602_, _02601_, _02376_);
  or (_02603_, _02494_, _02386_);
  or (_02604_, _02603_, _02602_);
  or (_02605_, _02604_, _02374_);
  and (_02606_, _02605_, _07230_);
  and (_02607_, \oc8051_top_1.oc8051_decoder1.wr , \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02608_, _02607_, _02359_);
  or (_02609_, _02608_, _02606_);
  and (_03660_, _02609_, _06444_);
  and (_02610_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_02611_, _07011_, _06992_);
  nor (_02612_, _02611_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_02613_, _02612_, _02540_);
  and (_02614_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_02615_, _02614_, _07026_);
  or (_02616_, _02615_, _02613_);
  and (_02617_, _02616_, _07035_);
  or (_02618_, _02617_, _02610_);
  and (_02619_, _02618_, _02538_);
  nor (_02620_, _11589_, _02538_);
  or (_02621_, _02620_, _06989_);
  or (_02622_, _02621_, _02619_);
  or (_02623_, _09503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  and (_02624_, _02623_, _06444_);
  and (_03663_, _02624_, _02622_);
  and (_02625_, _07011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  nor (_02626_, _02625_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  nor (_02627_, _02626_, _02611_);
  and (_02628_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_02629_, _02628_, _07026_);
  or (_02630_, _02629_, _02627_);
  and (_02631_, _02630_, _07035_);
  and (_02633_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_02634_, _02633_, _06985_);
  or (_02635_, _02634_, _02631_);
  nand (_02636_, _07069_, _06985_);
  and (_02637_, _02636_, _09503_);
  and (_02638_, _02637_, _02635_);
  and (_02639_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  or (_02640_, _02639_, _02638_);
  and (_03667_, _02640_, _06444_);
  and (_02641_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  nor (_02642_, _10955_, _10925_);
  nor (_02643_, _02642_, _10956_);
  or (_02644_, _02643_, _08374_);
  or (_02646_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  and (_02647_, _02646_, _10894_);
  and (_02648_, _02647_, _02644_);
  or (_03669_, _02648_, _02641_);
  nand (_02650_, _01085_, _07216_);
  or (_02651_, _02650_, _08230_);
  not (_02653_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  nand (_02654_, _02650_, _02653_);
  and (_02655_, _02654_, _06440_);
  and (_02656_, _02655_, _02651_);
  nor (_02657_, _06673_, _02653_);
  and (_02659_, _00604_, _07963_);
  and (_02660_, _02659_, _06983_);
  nand (_02662_, _02660_, _06930_);
  or (_02663_, _02660_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  and (_02665_, _02663_, _06674_);
  and (_02667_, _02665_, _02662_);
  or (_02668_, _02667_, _02657_);
  or (_02669_, _02668_, _02656_);
  and (_03678_, _02669_, _06444_);
  and (_02671_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  nand (_02672_, _02671_, _07006_);
  nand (_02674_, _02672_, _02625_);
  or (_02675_, _07011_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_02677_, _02675_, _07035_);
  and (_02678_, _02677_, _02674_);
  and (_02680_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_02681_, _02680_, _06985_);
  or (_02682_, _02681_, _02678_);
  nand (_02683_, _09526_, _06985_);
  and (_02684_, _02683_, _09503_);
  and (_02685_, _02684_, _02682_);
  and (_02686_, _06989_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  or (_02687_, _02686_, _02685_);
  and (_03685_, _02687_, _06444_);
  not (_02688_, _02332_);
  or (_03688_, _02688_, _02301_);
  or (_02689_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [7]);
  nand (_02690_, _07432_, _13886_);
  and (_02691_, _02690_, _06444_);
  and (_03692_, _02691_, _02689_);
  or (_02692_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [6]);
  nand (_02693_, _07432_, _13896_);
  and (_02694_, _02693_, _06444_);
  and (_03700_, _02694_, _02692_);
  or (_02695_, _02650_, _08019_);
  not (_02696_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  nand (_02697_, _02650_, _02696_);
  and (_02698_, _02697_, _06440_);
  and (_02699_, _02698_, _02695_);
  nor (_02700_, _06673_, _02696_);
  or (_02701_, _02650_, _08232_);
  and (_02702_, _02697_, _06674_);
  and (_02703_, _02702_, _02701_);
  or (_02704_, _02703_, _02700_);
  or (_02705_, _02704_, _02699_);
  and (_03705_, _02705_, _06444_);
  or (_02706_, _02650_, _08127_);
  not (_02707_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  nand (_02708_, _02650_, _02707_);
  and (_02709_, _02708_, _06440_);
  and (_02710_, _02709_, _02706_);
  nor (_02711_, _06673_, _02707_);
  and (_02712_, _02659_, _06987_);
  nand (_02713_, _02712_, _06930_);
  or (_02714_, _02712_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_02715_, _02714_, _06674_);
  and (_02716_, _02715_, _02713_);
  or (_02717_, _02716_, _02711_);
  or (_02718_, _02717_, _02710_);
  and (_03708_, _02718_, _06444_);
  and (_02719_, _11418_, _11347_);
  and (_02720_, _02719_, _11394_);
  or (_02721_, _02720_, _02257_);
  or (_02722_, _02471_, _11966_);
  or (_02723_, _02722_, _11396_);
  or (_02724_, _02723_, _02721_);
  or (_02725_, _02249_, _02283_);
  or (_02726_, _02598_, _02384_);
  or (_02727_, _02726_, _02725_);
  and (_02728_, _02263_, _07311_);
  or (_02729_, _02728_, _02354_);
  or (_02730_, _02729_, _02727_);
  or (_02731_, _14225_, _11398_);
  and (_02732_, _11456_, _11965_);
  or (_02733_, _02297_, _02732_);
  or (_02734_, _02733_, _02731_);
  and (_02735_, _02367_, _11418_);
  and (_02736_, _11437_, _11430_);
  and (_02737_, _02275_, _11376_);
  or (_02738_, _02737_, _02736_);
  or (_02739_, _02738_, _02735_);
  or (_02740_, _02739_, _02734_);
  or (_02741_, _02740_, _02730_);
  or (_02742_, _02279_, _02260_);
  or (_02743_, _02742_, _11440_);
  or (_02744_, _02743_, _02278_);
  and (_02745_, _02483_, _07311_);
  or (_02746_, _02264_, _11444_);
  or (_02747_, _02746_, _11375_);
  or (_02748_, _02747_, _02745_);
  or (_02749_, _02748_, _02744_);
  or (_02750_, _02749_, _02741_);
  or (_02751_, _02750_, _02724_);
  and (_02752_, _02751_, _07230_);
  and (_02753_, \oc8051_top_1.oc8051_sfr1.wait_data , \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  or (_02754_, _02593_, _02303_);
  or (_02755_, _02754_, _02753_);
  or (_02756_, _02755_, _02752_);
  and (_03710_, _02756_, _06444_);
  or (_02757_, _10954_, _10929_);
  nor (_02758_, _10955_, _08374_);
  and (_02759_, _02758_, _02757_);
  and (_02760_, _08374_, \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  or (_02761_, _02760_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 );
  or (_02762_, _02761_, _02759_);
  or (_02764_, _02166_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [5]);
  and (_02765_, _02764_, _06444_);
  and (_03712_, _02765_, _02762_);
  and (_02766_, _11418_, _11385_);
  nor (_02767_, _02766_, _02297_);
  or (_03715_, _02767_, _02688_);
  or (_02768_, _02448_, \oc8051_top_1.oc8051_decoder1.state [1]);
  or (_02769_, _02768_, _02454_);
  and (_02770_, _02769_, _02461_);
  nor (_02771_, _02460_, _11386_);
  or (_02772_, _02771_, rst);
  or (_03718_, _02772_, _02770_);
  and (_02773_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_02774_, _01553_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_02775_, _01553_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  nor (_02776_, _02775_, _02774_);
  not (_02777_, _02776_);
  nor (_02778_, _02777_, _01564_);
  and (_02779_, _02777_, _01564_);
  or (_02780_, _02779_, _02778_);
  or (_02781_, _02780_, _08374_);
  or (_02782_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  and (_02783_, _02782_, _10894_);
  and (_02784_, _02783_, _02781_);
  or (_03720_, _02784_, _02773_);
  and (_02785_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8], \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  and (_02786_, _12225_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [6]);
  and (_02787_, _02786_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  and (_02788_, _02787_, _02785_);
  and (_02789_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11], \oc8051_top_1.oc8051_memory_interface1.pc_buf [12]);
  nand (_02790_, _02789_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_02791_, _02790_, _07432_);
  and (_02792_, _02791_, _02788_);
  and (_02793_, _02792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  and (_02794_, _02793_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nand (_02795_, _02794_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_02796_, _02794_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  and (_02797_, _02796_, _02795_);
  or (_02798_, _02797_, _12023_);
  and (_02799_, _02798_, _06444_);
  and (_02800_, _11452_, _11137_);
  and (_02801_, _12026_, _11177_);
  and (_02802_, _12032_, _11625_);
  and (_02803_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [15]);
  or (_02804_, _02803_, _02802_);
  or (_02805_, _02804_, _02801_);
  or (_02806_, _02805_, _02800_);
  or (_02807_, \oc8051_top_1.oc8051_memory_interface1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  or (_02808_, _02807_, _12660_);
  or (_02809_, _02808_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nand (_02810_, _02809_, _12650_);
  or (_02811_, _12666_, _08150_);
  or (_02812_, _02811_, _08155_);
  or (_02813_, _02812_, _09186_);
  nand (_02814_, _02813_, _12662_);
  nand (_02815_, _02814_, _02810_);
  nand (_02816_, _02815_, _11165_);
  or (_02817_, _02815_, _11165_);
  and (_02818_, _02817_, _12218_);
  and (_02819_, _02818_, _02816_);
  or (_02820_, _02819_, _02806_);
  and (_02821_, _12683_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  and (_02822_, _02821_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_02823_, _02822_, _11165_);
  and (_02824_, _02822_, _11165_);
  or (_02825_, _02824_, _02823_);
  nand (_02826_, _02825_, _12054_);
  nand (_02827_, _02826_, _12023_);
  or (_02828_, _02827_, _02820_);
  and (_03733_, _02828_, _02799_);
  or (_02829_, _02650_, _12024_);
  not (_02830_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  nand (_02831_, _02650_, _02830_);
  and (_02832_, _02831_, _06440_);
  and (_02833_, _02832_, _02829_);
  nor (_02834_, _06673_, _02830_);
  and (_02835_, _02659_, _00240_);
  nand (_02836_, _02835_, _06930_);
  or (_02837_, _02835_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  and (_02838_, _02837_, _06674_);
  and (_02839_, _02838_, _02836_);
  or (_02840_, _02839_, _02834_);
  or (_02841_, _02840_, _02833_);
  and (_03737_, _02841_, _06444_);
  and (_02842_, _11418_, _11976_);
  or (_02843_, _02842_, _11513_);
  or (_02844_, _02843_, _11517_);
  and (_02845_, _02384_, _11410_);
  or (_02846_, _02845_, _11371_);
  or (_02847_, _02846_, _02844_);
  and (_02848_, _02364_, _07268_);
  or (_02849_, _02248_, _11398_);
  or (_02850_, _02849_, _02368_);
  or (_02851_, _02850_, _02848_);
  or (_02852_, _02851_, _02847_);
  or (_02853_, _02852_, _02749_);
  or (_02854_, _02853_, _02724_);
  and (_02855_, _02854_, _07230_);
  and (_02856_, \oc8051_top_1.oc8051_decoder1.src_sel1 [1], \oc8051_top_1.oc8051_sfr1.wait_data );
  or (_02857_, _02856_, _02754_);
  or (_02858_, _02857_, _02855_);
  and (_03743_, _02858_, _06444_);
  nor (_03747_, _12073_, rst);
  and (_03752_, \oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _06444_);
  nand (_02859_, _10494_, _09479_);
  not (_02860_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  nor (_02861_, _09485_, _02860_);
  and (_02862_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_02863_, _02862_, _02861_);
  or (_02864_, _02863_, _09479_);
  and (_02865_, _02864_, _06444_);
  and (_03756_, _02865_, _02859_);
  nor (_03758_, _11547_, rst);
  nand (_02866_, _10112_, _09526_);
  or (_02867_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [0]);
  and (_02868_, _02867_, _02866_);
  and (_03765_, _02868_, _06444_);
  and (_02869_, _12012_, _06983_);
  nand (_02870_, _02869_, _06930_);
  or (_02871_, _02869_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_02872_, _02871_, _07219_);
  and (_02873_, _02872_, _02870_);
  or (_02874_, _02873_, _07221_);
  and (_03784_, _02874_, _06444_);
  or (_02875_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  or (_02876_, _09486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  and (_02877_, _02876_, _02875_);
  or (_02878_, _02877_, _09479_);
  nand (_02880_, _09479_, _07069_);
  and (_02882_, _02880_, _06444_);
  and (_03787_, _02882_, _02878_);
  nand (_02884_, _09479_, _06666_);
  or (_02885_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  not (_02887_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  nand (_02889_, _09485_, _02887_);
  and (_02891_, _02889_, _02885_);
  or (_02892_, _02891_, _09479_);
  and (_02894_, _02892_, _06444_);
  and (_03791_, _02894_, _02884_);
  nor (_03794_, _11470_, rst);
  nand (_02895_, _09479_, _07188_);
  and (_02896_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_02897_, _09486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_02899_, _02897_, _02896_);
  or (_02900_, _02899_, _09479_);
  and (_02901_, _02900_, _06444_);
  and (_03797_, _02901_, _02895_);
  and (_02902_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  not (_02903_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  nor (_02904_, _09485_, _02903_);
  or (_02906_, _02904_, _02902_);
  or (_02907_, _02906_, _09479_);
  nand (_02909_, _09479_, _07300_);
  and (_02910_, _02909_, _06444_);
  and (_03800_, _02910_, _02907_);
  nor (_03802_, _12106_, rst);
  or (_02911_, _02650_, _07959_);
  not (_02912_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  nand (_02913_, _02650_, _02912_);
  and (_02915_, _02913_, _06440_);
  and (_02917_, _02915_, _02911_);
  nor (_02918_, _06673_, _02912_);
  and (_02920_, _02659_, _06432_);
  nand (_02922_, _02920_, _06930_);
  or (_02923_, _02920_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_02925_, _02923_, _06674_);
  and (_02927_, _02925_, _02922_);
  or (_02928_, _02927_, _02918_);
  or (_02929_, _02928_, _02917_);
  and (_03804_, _02929_, _06444_);
  or (_02930_, _02650_, _08308_);
  not (_02931_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  nand (_02932_, _02650_, _02931_);
  and (_02933_, _02932_, _06440_);
  and (_02934_, _02933_, _02930_);
  nor (_02935_, _06673_, _02931_);
  and (_02936_, _02659_, _08310_);
  nand (_02937_, _02936_, _06930_);
  or (_02938_, _02936_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  and (_02939_, _02938_, _06674_);
  and (_02940_, _02939_, _02937_);
  or (_02941_, _02940_, _02935_);
  or (_02942_, _02941_, _02934_);
  and (_03807_, _02942_, _06444_);
  nor (_03812_, _12128_, rst);
  and (_02943_, _02306_, \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  or (_02944_, _11479_, _11476_);
  or (_02946_, _11512_, _11487_);
  or (_02947_, _02946_, _02944_);
  or (_02948_, _02947_, _02558_);
  and (_02949_, _02555_, _11356_);
  or (_02950_, _11456_, _11486_);
  and (_02951_, _02950_, _11355_);
  or (_02952_, _02951_, _02949_);
  or (_02953_, _02481_, _02264_);
  or (_02954_, _02953_, _02279_);
  or (_02955_, _02954_, _02952_);
  or (_02956_, _02955_, _02948_);
  and (_02957_, _02497_, _07311_);
  or (_02958_, _02957_, _02254_);
  or (_02959_, _02958_, _11495_);
  or (_02960_, _02564_, _02732_);
  and (_02961_, _11456_, _11526_);
  and (_02962_, _11423_, _11426_);
  or (_02963_, _02962_, _02961_);
  or (_02964_, _02963_, _02960_);
  or (_02965_, _11504_, _11444_);
  or (_02966_, _02965_, _11509_);
  or (_02967_, _02966_, _02964_);
  or (_02968_, _02967_, _02959_);
  or (_02969_, _02968_, _02956_);
  and (_02970_, _02969_, _02332_);
  or (_03816_, _02970_, _02943_);
  and (_02971_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_02972_, _09486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  or (_02973_, _02972_, _02971_);
  or (_02974_, _02973_, _09479_);
  nand (_02975_, _11589_, _09479_);
  and (_02976_, _02975_, _06444_);
  and (_03821_, _02976_, _02974_);
  not (_02977_, _09138_);
  or (_02978_, _02650_, _02977_);
  not (_02979_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  nand (_02980_, _02650_, _02979_);
  and (_02981_, _02980_, _06440_);
  and (_02982_, _02981_, _02978_);
  nor (_02983_, _06673_, _02979_);
  not (_02984_, _02659_);
  or (_02985_, _02984_, _00717_);
  and (_02986_, _02985_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  and (_02987_, _06431_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_02988_, _02987_, _00713_);
  and (_02989_, _02988_, _02659_);
  or (_02990_, _02989_, _02986_);
  and (_02991_, _02990_, _06674_);
  or (_02992_, _02991_, _02983_);
  or (_02993_, _02992_, _02982_);
  and (_03824_, _02993_, _06444_);
  and (_02994_, _12012_, _08310_);
  or (_02995_, _02994_, _07278_);
  nand (_02996_, _02994_, _06930_);
  and (_02997_, _02996_, _02995_);
  or (_02998_, _02997_, _07301_);
  and (_03828_, _02998_, _06444_);
  or (_02999_, _07263_, _02464_);
  or (_03000_, _07229_, \oc8051_top_1.oc8051_decoder1.op [0]);
  and (_03001_, _03000_, _06444_);
  and (_03831_, _03001_, _02999_);
  or (_03002_, _08392_, _02464_);
  or (_03003_, _07229_, \oc8051_top_1.oc8051_decoder1.op [1]);
  and (_03004_, _03003_, _06444_);
  and (_03833_, _03004_, _03002_);
  nand (_03005_, _08408_, _07229_);
  or (_03006_, _07229_, \oc8051_top_1.oc8051_decoder1.op [2]);
  and (_03007_, _03006_, _06444_);
  and (_03835_, _03007_, _03005_);
  or (_03008_, _08425_, _02464_);
  or (_03009_, _07229_, \oc8051_top_1.oc8051_decoder1.op [3]);
  and (_03010_, _03009_, _06444_);
  and (_03837_, _03010_, _03008_);
  or (_03011_, _08441_, _02464_);
  or (_03012_, _07229_, \oc8051_top_1.oc8051_decoder1.op [4]);
  and (_03013_, _03012_, _06444_);
  and (_03839_, _03013_, _03011_);
  or (_03014_, _08457_, _02464_);
  or (_03015_, _07229_, \oc8051_top_1.oc8051_decoder1.op [5]);
  and (_03016_, _03015_, _06444_);
  and (_03840_, _03016_, _03014_);
  nor (_03017_, _10953_, _10948_);
  nor (_03018_, _03017_, _10954_);
  or (_03019_, _03018_, _08374_);
  or (_03020_, _08373_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  and (_03021_, _03020_, _10894_);
  and (_03022_, _03021_, _03019_);
  and (_03023_, _10976_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  or (_03842_, _03023_, _03022_);
  nand (_03024_, _08472_, _07229_);
  or (_03025_, _07229_, \oc8051_top_1.oc8051_decoder1.op [6]);
  and (_03026_, _03025_, _06444_);
  and (_03851_, _03026_, _03024_);
  or (_03027_, \oc8051_top_1.oc8051_decoder1.psw_set [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03028_, _07987_, _07927_);
  or (_03029_, _03028_, _09095_);
  or (_03030_, _03029_, _08284_);
  or (_03031_, _03030_, _08097_);
  or (_03032_, _03031_, _08996_);
  and (_03033_, _03032_, _07602_);
  or (_03034_, _06844_, _06842_);
  not (_03035_, _06706_);
  nand (_03037_, _06842_, _03035_);
  and (_03038_, _03037_, _06680_);
  and (_03039_, _03038_, _03034_);
  not (_03041_, _06707_);
  nand (_03043_, _06877_, _03041_);
  nor (_03045_, _06878_, _06848_);
  and (_03047_, _03045_, _03043_);
  and (_03048_, _06752_, _06482_);
  and (_03050_, _03048_, _07578_);
  and (_03051_, _03050_, _08167_);
  nand (_03052_, _03051_, _07459_);
  nand (_03053_, _03052_, \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  or (_03054_, _03053_, _03047_);
  or (_03055_, _03054_, _03039_);
  nor (_03056_, _03055_, _08206_);
  nand (_03057_, _03056_, _11108_);
  or (_03058_, _03057_, _03033_);
  and (_03059_, _03058_, _03027_);
  or (_03060_, _03059_, _12012_);
  and (_03062_, _00712_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  or (_03063_, _03062_, _00713_);
  or (_03064_, _03063_, _12013_);
  and (_03065_, _03064_, _03060_);
  or (_03066_, _03065_, _07218_);
  nand (_03067_, _11589_, _07218_);
  and (_03068_, _03067_, _06444_);
  and (_03860_, _03068_, _03066_);
  or (_03069_, _09485_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  or (_03071_, _09486_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  and (_03073_, _03071_, _03069_);
  or (_03075_, _03073_, _09479_);
  nand (_03077_, _09526_, _09479_);
  and (_03079_, _03077_, _06444_);
  and (_03864_, _03079_, _03075_);
  and (_03082_, _12012_, _06432_);
  nand (_03083_, _03082_, _06930_);
  or (_03085_, _03082_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  and (_03087_, _03085_, _07219_);
  and (_03089_, _03087_, _03083_);
  nor (_03090_, _07219_, _07069_);
  or (_03092_, _03090_, _03089_);
  and (_03869_, _03092_, _06444_);
  nand (_03093_, _09484_, _07300_);
  and (_03094_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  and (_03095_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  or (_03096_, _03095_, _03094_);
  or (_03097_, _03096_, _09484_);
  and (_03098_, _03097_, _09684_);
  and (_03099_, _03098_, _03093_);
  and (_03100_, _09479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  or (_03101_, _03100_, _03099_);
  and (_03911_, _03101_, _06444_);
  nand (_03102_, _10494_, _09484_);
  and (_03103_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_03104_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  or (_03105_, _03104_, _03103_);
  or (_03106_, _03105_, _09484_);
  and (_03107_, _03106_, _09684_);
  and (_03108_, _03107_, _03102_);
  and (_03109_, _09479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  or (_03110_, _03109_, _03108_);
  and (_03914_, _03110_, _06444_);
  and (_03111_, _06430_, _06395_);
  and (_03112_, _08976_, _03111_);
  and (_03113_, _03112_, _06941_);
  and (_03114_, _03113_, _06440_);
  or (_03115_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  not (_03116_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  nand (_03117_, _09481_, _03116_);
  nand (_03119_, _03117_, _03115_);
  nor (_03120_, _03119_, _03114_);
  not (_03121_, _03114_);
  nor (_03122_, _03121_, _06666_);
  or (_03123_, _03122_, _03120_);
  or (_03124_, _03123_, _09479_);
  or (_03125_, _09684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_03126_, _03125_, _06444_);
  and (_03917_, _03126_, _03124_);
  nand (_03127_, _09484_, _07188_);
  and (_03128_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  and (_03129_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  or (_03130_, _03129_, _03128_);
  or (_03131_, _03130_, _09484_);
  and (_03133_, _03131_, _09684_);
  and (_03134_, _03133_, _03127_);
  and (_03135_, _09479_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  or (_03136_, _03135_, _03134_);
  and (_03923_, _03136_, _06444_);
  and (_03137_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_03138_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  nor (_03139_, _03138_, _03137_);
  nor (_03140_, _03139_, _03114_);
  nor (_03141_, _11589_, _03121_);
  or (_03142_, _03141_, _03140_);
  or (_03143_, _03142_, _09479_);
  or (_03145_, _09684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  and (_03146_, _03145_, _06444_);
  and (_03935_, _03146_, _03143_);
  and (_03148_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [2]);
  nor (_03149_, _11589_, _07046_);
  or (_03151_, _03149_, _03148_);
  and (_03944_, _03151_, _06444_);
  or (_03152_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  or (_03153_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  and (_03154_, _03153_, _03152_);
  or (_03155_, _03154_, _09484_);
  nand (_03156_, _09484_, _07069_);
  and (_03157_, _03156_, _03155_);
  or (_03158_, _03157_, _09479_);
  or (_03159_, _09684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  and (_03160_, _03159_, _06444_);
  and (_03958_, _03160_, _03158_);
  nand (_03161_, _09526_, _09484_);
  or (_03162_, _09481_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  or (_03163_, _09482_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  and (_03164_, _03163_, _03162_);
  or (_03165_, _03164_, _09484_);
  and (_03166_, _03165_, _03161_);
  or (_03167_, _03166_, _09479_);
  or (_03168_, _09684_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  and (_03169_, _03168_, _06444_);
  and (_03962_, _03169_, _03167_);
  and (_03170_, _02306_, \oc8051_top_1.oc8051_decoder1.alu_op [0]);
  or (_03171_, _02574_, _11381_);
  or (_03172_, _03171_, _02734_);
  and (_03173_, _02260_, _11347_);
  or (_03174_, _02278_, _11440_);
  or (_03175_, _03174_, _03173_);
  or (_03176_, _02254_, _11409_);
  or (_03177_, _02737_, _02483_);
  or (_03178_, _03177_, _03176_);
  or (_03179_, _02323_, _11343_);
  or (_03180_, _03179_, _11442_);
  nor (_03181_, _03180_, _11483_);
  nand (_03182_, _03181_, _11514_);
  or (_03183_, _03182_, _03178_);
  or (_03184_, _03183_, _03175_);
  or (_03185_, _03184_, _03172_);
  or (_03186_, _11398_, _11342_);
  nor (_03187_, rst, \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_03188_, _03187_, _03186_);
  and (_03189_, _03188_, _03185_);
  or (_03981_, _03189_, _03170_);
  nor (_03190_, _14070_, _06978_);
  and (_03191_, _14070_, \oc8051_top_1.oc8051_indi_addr1.buff[3] [7]);
  or (_03192_, _03191_, _03190_);
  and (_03986_, _03192_, _06444_);
  and (_03193_, _02306_, \oc8051_top_1.oc8051_decoder1.alu_op [1]);
  or (_03194_, _02276_, _11977_);
  or (_03195_, _02483_, _11438_);
  nor (_03197_, _03195_, _03194_);
  nand (_03198_, _03197_, _14227_);
  and (_03199_, _11486_, _11355_);
  or (_03200_, _02720_, _11489_);
  or (_03201_, _03200_, _03199_);
  or (_03202_, _03201_, _02954_);
  or (_03203_, _03202_, _03198_);
  nor (_03204_, _11479_, _11398_);
  nand (_03205_, _03204_, _11445_);
  and (_03206_, _11431_, _11355_);
  or (_03207_, _02722_, _03206_);
  or (_03208_, _03207_, _03205_);
  or (_03209_, _03208_, _02495_);
  or (_03210_, _03209_, _02499_);
  or (_03211_, _03210_, _03203_);
  and (_03212_, _03211_, _03188_);
  or (_03989_, _03212_, _03193_);
  or (_03213_, _11442_, _11428_);
  or (_03214_, _03213_, _02276_);
  or (_03215_, _03214_, _11438_);
  or (_03216_, _03215_, _02494_);
  or (_03217_, _03201_, _02498_);
  or (_03218_, _03217_, _03216_);
  or (_03219_, _02559_, _14226_);
  and (_03220_, _02260_, _11360_);
  or (_03221_, _03220_, _02946_);
  or (_03222_, _03221_, _03219_);
  or (_03223_, _03222_, _02959_);
  or (_03224_, _03223_, _03218_);
  and (_03225_, _03224_, _07230_);
  and (_03226_, \oc8051_top_1.oc8051_decoder1.alu_op [2], \oc8051_top_1.oc8051_sfr1.wait_data );
  and (_03227_, _11396_, _06308_);
  or (_03228_, _03227_, _03226_);
  or (_03229_, _03228_, _03225_);
  and (_03994_, _03229_, _06444_);
  and (_03230_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [5]);
  nor (_03231_, _07046_, _06666_);
  or (_03232_, _03231_, _03230_);
  and (_03996_, _03232_, _06444_);
  nor (_04000_, _12154_, rst);
  and (_03233_, _02306_, \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  or (_03234_, _02254_, _02264_);
  or (_03235_, _03234_, _02469_);
  nor (_03236_, _11533_, _11966_);
  nand (_03237_, _03236_, _11978_);
  or (_03238_, _03237_, _03235_);
  or (_03239_, _02952_, _02947_);
  or (_03240_, _03239_, _03238_);
  or (_03241_, _03240_, _02589_);
  and (_03242_, _03241_, _02332_);
  or (_04011_, _03242_, _03233_);
  nor (_03243_, _06978_, _09146_);
  and (_03244_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  or (_03245_, _03244_, _07158_);
  or (_03246_, _03245_, _03243_);
  or (_03247_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [7]);
  and (_03248_, _03247_, _06444_);
  and (_04025_, _03248_, _03246_);
  or (_03249_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [11]);
  nand (_03250_, _07432_, _13968_);
  and (_03251_, _03250_, _06444_);
  and (_04050_, _03251_, _03249_);
  or (_03252_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [10]);
  nand (_03253_, _07432_, _13999_);
  and (_03254_, _03253_, _06444_);
  and (_04052_, _03254_, _03252_);
  or (_03255_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [9]);
  nand (_03256_, _07432_, _12812_);
  and (_03257_, _03256_, _06444_);
  and (_04057_, _03257_, _03255_);
  and (_04074_, _06444_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  and (_03258_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  or (_03259_, _07459_, \oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0]);
  nand (_03260_, _03259_, _06444_);
  nor (_04088_, _03260_, _03258_);
  and (_04094_, _08201_, _06444_);
  and (_03261_, _09328_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  and (_03262_, _11882_, _07151_);
  and (_03263_, _09332_, \oc8051_top_1.oc8051_indi_addr1.buff[4] [2]);
  or (_03264_, _03263_, _03262_);
  and (_03265_, _03264_, _06439_);
  or (_03266_, _03265_, _03261_);
  and (_04095_, _03266_, _06444_);
  nand (_03267_, _10494_, _10112_);
  or (_03268_, _10112_, \oc8051_top_1.oc8051_indi_addr1.buff[0] [6]);
  and (_03269_, _03268_, _06444_);
  and (_04105_, _03269_, _03267_);
  nor (_03270_, _12615_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  nor (_03271_, _03270_, _12616_);
  or (_03272_, _03271_, _12023_);
  and (_03273_, _03272_, _06444_);
  not (_03274_, _12023_);
  and (_03275_, _12659_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  or (_03276_, _03275_, _12661_);
  or (_03277_, _12665_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  and (_03278_, _03277_, _12666_);
  or (_03279_, _03278_, _12650_);
  and (_03280_, _03279_, _12218_);
  and (_03281_, _03280_, _03276_);
  nor (_03282_, _12681_, \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  nor (_03283_, _03282_, _12682_);
  and (_03284_, _03283_, _12054_);
  and (_03285_, _11452_, _08308_);
  and (_03286_, _12026_, _08342_);
  and (_03287_, _11689_, _12032_);
  and (_03288_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [11]);
  or (_03289_, _03288_, _03287_);
  or (_03290_, _03289_, _03286_);
  or (_03291_, _03290_, _03285_);
  or (_03292_, _03291_, _03284_);
  or (_03294_, _03292_, _03281_);
  or (_03296_, _03294_, _03274_);
  and (_04109_, _03296_, _03273_);
  nor (_03297_, _00855_, _09138_);
  not (_03298_, _12026_);
  nor (_03299_, _03298_, _09280_);
  and (_03301_, _11905_, _12032_);
  and (_03302_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  or (_03303_, _03302_, _03301_);
  or (_03305_, _03303_, _03299_);
  or (_03306_, _03305_, _03297_);
  and (_03308_, _12658_, _12650_);
  nor (_03310_, _12664_, _12650_);
  or (_03311_, _03310_, _03308_);
  nand (_03312_, _03311_, _08143_);
  or (_03313_, _03311_, _08143_);
  and (_03314_, _03313_, _03312_);
  and (_03315_, _03314_, _12218_);
  or (_03316_, _03315_, _03306_);
  nand (_03317_, _12054_, _08360_);
  nand (_03318_, _03317_, _12023_);
  or (_03319_, _03318_, _03316_);
  nor (_03320_, _12614_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [10]);
  nor (_03322_, _03320_, _12615_);
  or (_03323_, _03322_, _12023_);
  and (_03324_, _03323_, _06444_);
  and (_04113_, _03324_, _03319_);
  and (_03326_, _12656_, \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  or (_03327_, _03326_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  and (_03328_, _03327_, _03310_);
  nand (_03329_, _12657_, \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  nand (_03330_, _03329_, _12658_);
  and (_03332_, _03330_, _12650_);
  or (_03333_, _03332_, _03328_);
  and (_03334_, _03333_, _12218_);
  nor (_03335_, _03298_, _07640_);
  and (_03336_, _11452_, _07959_);
  and (_03337_, _12032_, _11794_);
  and (_03338_, _12054_, _10739_);
  and (_03339_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  or (_03340_, _03339_, _03338_);
  or (_03341_, _03340_, _03337_);
  or (_03342_, _03341_, _03336_);
  or (_03343_, _03342_, _03335_);
  or (_03345_, _03343_, _03334_);
  or (_03346_, _03345_, _03274_);
  nor (_03347_, _12613_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [9]);
  nor (_03348_, _03347_, _12614_);
  or (_03349_, _03348_, _12023_);
  and (_03351_, _03349_, _06444_);
  and (_04123_, _03351_, _03346_);
  and (_03352_, _11452_, _08019_);
  and (_03353_, _12054_, _08457_);
  nor (_03354_, _03298_, _08060_);
  and (_03356_, _11848_, _12032_);
  and (_03358_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  or (_03359_, _03358_, _03356_);
  or (_03361_, _03359_, _03354_);
  or (_03362_, _03361_, _03353_);
  nor (_03363_, _03362_, _03352_);
  nand (_03364_, _03363_, _12023_);
  nand (_03365_, _12656_, _07589_);
  or (_03366_, _12656_, _07589_);
  and (_03367_, _03366_, _03365_);
  nor (_03368_, _03367_, _12650_);
  and (_03369_, _03367_, _12650_);
  or (_03370_, _03369_, _03368_);
  and (_03371_, _03370_, _12606_);
  or (_03372_, _03371_, _03364_);
  nor (_03373_, _12612_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [8]);
  nor (_03374_, _03373_, _12613_);
  or (_03375_, _03374_, _12023_);
  and (_03376_, _03375_, _06444_);
  and (_04126_, _03376_, _03372_);
  nor (_03377_, _12227_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_03378_, _03377_, _12612_);
  or (_03379_, _03378_, _12023_);
  and (_03380_, _03379_, _06444_);
  nor (_03381_, _12654_, _12653_);
  nor (_03382_, _03381_, _12655_);
  and (_03383_, _03382_, _12218_);
  and (_03384_, _12048_, _11137_);
  and (_03386_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [7]);
  nor (_03387_, _12648_, _12033_);
  and (_03388_, _12054_, _11625_);
  or (_03389_, _03388_, _03387_);
  or (_03390_, _03389_, _03386_);
  or (_03391_, _03390_, _03384_);
  nor (_03392_, _03391_, _03383_);
  nand (_03393_, _03392_, _12023_);
  and (_04131_, _03393_, _03380_);
  nor (_03394_, _03258_, _07471_);
  and (_03395_, _03258_, _07471_);
  or (_03396_, _03395_, _03394_);
  and (_04192_, _03396_, _06444_);
  and (_04195_, _11102_, _06444_);
  and (_04203_, _06444_, \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  or (_03397_, _07414_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  nand (_03399_, _07069_, _07414_);
  and (_03400_, _03399_, _03397_);
  or (_03401_, _03400_, _07158_);
  or (_03402_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [1]);
  and (_03403_, _03402_, _06444_);
  and (_04204_, _03403_, _03401_);
  not (_03404_, _00936_);
  or (_03405_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_03407_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10]);
  and (_03408_, _03407_, _03405_);
  and (_03409_, _03408_, _06443_);
  and (_03410_, _06442_, _06296_);
  or (_03411_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _13875_);
  and (_03412_, _03411_, _06444_);
  and (_03413_, _03412_, _03410_);
  or (_04206_, _03413_, _03409_);
  nor (_03415_, _07300_, _09146_);
  and (_03416_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  or (_03417_, _03416_, _07158_);
  or (_03418_, _03417_, _03415_);
  or (_03419_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [3]);
  and (_03420_, _03419_, _06444_);
  and (_04208_, _03420_, _03418_);
  nor (_03421_, _10494_, _09146_);
  and (_03422_, _09146_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  or (_03423_, _03422_, _07158_);
  or (_03424_, _03423_, _03421_);
  or (_03426_, _06439_, \oc8051_top_1.oc8051_indi_addr1.buff[1] [6]);
  and (_03427_, _03426_, _06444_);
  and (_04210_, _03427_, _03424_);
  nor (_03430_, _14085_, _11669_);
  and (_03431_, _03430_, _14142_);
  or (_03432_, _01519_, _14113_);
  or (_03433_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  and (_03434_, _03433_, _14079_);
  and (_03435_, _03434_, _03432_);
  and (_03436_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  and (_03437_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  or (_03438_, _03437_, _03436_);
  and (_03439_, _03438_, _14094_);
  or (_03440_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  or (_03441_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_03442_, _03441_, _14103_);
  and (_03443_, _03442_, _03440_);
  or (_03444_, _03443_, _03439_);
  or (_03445_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  or (_03446_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  and (_03447_, _03446_, _14091_);
  and (_03448_, _03447_, _03445_);
  or (_03449_, _03448_, _03444_);
  or (_03450_, _03449_, _03435_);
  and (_03451_, _03450_, _03431_);
  nor (_03452_, _11919_, _07098_);
  and (_03453_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  or (_03454_, _03453_, _03452_);
  and (_03455_, _03454_, _14079_);
  or (_03456_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  or (_03457_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  and (_03458_, _03457_, _14094_);
  and (_03459_, _03458_, _03456_);
  or (_03461_, _03459_, _03455_);
  and (_03462_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  and (_03463_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  or (_03464_, _03463_, _03462_);
  and (_03465_, _03464_, _14091_);
  or (_03466_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  or (_03467_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  and (_03468_, _03467_, _14103_);
  and (_03469_, _03468_, _03466_);
  or (_03470_, _03469_, _03465_);
  or (_03471_, _03470_, _03461_);
  and (_03472_, _03471_, _14109_);
  or (_03473_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  or (_03474_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  and (_03475_, _03474_, _14079_);
  and (_03476_, _03475_, _03473_);
  or (_03477_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  or (_03478_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  and (_03479_, _03478_, _14094_);
  and (_03480_, _03479_, _03477_);
  or (_03481_, _03480_, _03476_);
  and (_03482_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  and (_03484_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  or (_03485_, _03484_, _03482_);
  and (_03486_, _03485_, _14091_);
  or (_03487_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  or (_03488_, _14113_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  and (_03489_, _03488_, _14103_);
  and (_03490_, _03489_, _03487_);
  or (_03491_, _03490_, _03486_);
  or (_03492_, _03491_, _03481_);
  and (_03493_, _03492_, _14101_);
  nor (_03494_, _11919_, _07110_);
  and (_03496_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  or (_03497_, _03496_, _03494_);
  and (_03498_, _03497_, _14094_);
  nand (_03499_, _11919_, _07118_);
  or (_03500_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  and (_03501_, _03500_, _14079_);
  and (_03503_, _03501_, _03499_);
  or (_03504_, _03503_, _03498_);
  or (_03505_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  nand (_03506_, _11919_, _07115_);
  and (_03507_, _03506_, _14103_);
  and (_03508_, _03507_, _03505_);
  or (_03509_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  nand (_03510_, _11919_, _07123_);
  and (_03511_, _03510_, _14091_);
  and (_03512_, _03511_, _03509_);
  or (_03513_, _03512_, _03508_);
  or (_03514_, _03513_, _03504_);
  and (_03516_, _03514_, _14112_);
  or (_03517_, _03516_, _03493_);
  or (_03518_, _03517_, _03472_);
  and (_03519_, _03518_, _14085_);
  and (_03520_, _14108_, _11703_);
  nor (_03521_, _03431_, _03520_);
  nand (_03522_, _14144_, _11703_);
  and (_03524_, _03522_, _03521_);
  nand (_03525_, _14129_, _11703_);
  and (_03526_, _14083_, _14085_);
  and (_03527_, _14101_, _11703_);
  nand (_03528_, _14100_, _14085_);
  nand (_03529_, _03528_, \oc8051_top_1.oc8051_sfr1.bit_out );
  or (_03530_, _03529_, _03527_);
  nor (_03531_, _03530_, _03526_);
  and (_03533_, _03531_, _03525_);
  and (_03534_, _03533_, _03524_);
  and (_03535_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  and (_03536_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  or (_03538_, _03536_, _11919_);
  or (_03539_, _03538_, _03535_);
  and (_03540_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  and (_03541_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  or (_03542_, _03541_, _14113_);
  or (_03543_, _03542_, _03540_);
  and (_03544_, _03543_, _03539_);
  or (_03546_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  nand (_03548_, _11919_, _01116_);
  and (_03549_, _03548_, _14091_);
  and (_03550_, _03549_, _03546_);
  nor (_03551_, _11919_, _01311_);
  and (_03552_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  or (_03553_, _03552_, _03551_);
  and (_03555_, _03553_, _14094_);
  or (_03556_, _03555_, _11703_);
  or (_03557_, _03556_, _03550_);
  or (_03558_, _03557_, _03544_);
  or (_03559_, _14247_, p1_in[7]);
  or (_03560_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  and (_03561_, _03560_, _03559_);
  and (_03562_, _03561_, _14103_);
  and (_03563_, _14256_, _14091_);
  or (_03564_, _03563_, _11919_);
  or (_03565_, _03564_, _03562_);
  and (_03566_, _14329_, _14103_);
  and (_03567_, _14417_, _14091_);
  or (_03568_, _03567_, _14113_);
  or (_03569_, _03568_, _03566_);
  and (_03570_, _03569_, _03565_);
  or (_03571_, _01471_, _14113_);
  or (_03572_, _01393_, _11919_);
  and (_03574_, _03572_, _14079_);
  and (_03575_, _03574_, _03571_);
  or (_03576_, _14483_, _14113_);
  or (_03577_, _01249_, _11919_);
  and (_03578_, _03577_, _14094_);
  and (_03579_, _03578_, _03576_);
  or (_03580_, _03579_, _14085_);
  or (_03581_, _03580_, _03575_);
  or (_03582_, _03581_, _03570_);
  and (_03583_, _03582_, _14129_);
  and (_03584_, _03583_, _03558_);
  and (_03585_, _11925_, \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  and (_03586_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  and (_03587_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  or (_03588_, _03587_, _03586_);
  and (_03589_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_03590_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  or (_03591_, _03590_, _03589_);
  or (_03592_, _03591_, _03588_);
  and (_03593_, _03592_, _14113_);
  and (_03594_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_03595_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_03596_, _03595_, _03594_);
  and (_03598_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_03600_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  or (_03601_, _03600_, _03598_);
  or (_03602_, _03601_, _03596_);
  and (_03603_, _03602_, _11919_);
  or (_03604_, _03603_, _03593_);
  and (_03605_, _03604_, _03526_);
  or (_03607_, _03605_, _03585_);
  or (_03608_, _03607_, _03584_);
  or (_03609_, _03608_, _03534_);
  or (_03610_, _14474_, _14113_);
  or (_03611_, _01239_, _11919_);
  and (_03612_, _03611_, _14094_);
  and (_03613_, _03612_, _03610_);
  or (_03614_, _14268_, _11919_);
  or (_03615_, _14403_, _14113_);
  and (_03616_, _03615_, _14091_);
  and (_03617_, _03616_, _03614_);
  or (_03618_, _03617_, _03613_);
  or (_03619_, _01462_, _14113_);
  or (_03620_, _01403_, _11919_);
  and (_03622_, _03620_, _14079_);
  and (_03624_, _03622_, _03619_);
  or (_03626_, _14334_, _14113_);
  or (_03628_, _14247_, p2_in[7]);
  or (_03629_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  and (_03631_, _03629_, _03628_);
  or (_03633_, _03631_, _11919_);
  and (_03635_, _03633_, _14103_);
  and (_03636_, _03635_, _03626_);
  or (_03638_, _03636_, _03624_);
  or (_03639_, _03638_, _03618_);
  and (_03641_, _03639_, _11669_);
  and (_03642_, _01399_, _14079_);
  or (_03643_, _03642_, _11919_);
  and (_03645_, _14263_, _14091_);
  and (_03647_, _01235_, _14094_);
  or (_03649_, _14247_, p3_in[7]);
  or (_03650_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  and (_03652_, _03650_, _03649_);
  and (_03654_, _03652_, _14103_);
  or (_03655_, _03654_, _03647_);
  or (_03657_, _03655_, _03645_);
  or (_03659_, _03657_, _03643_);
  and (_03661_, _14470_, _14094_);
  or (_03662_, _03661_, _14113_);
  and (_03664_, _01458_, _14079_);
  and (_03665_, _14338_, _14103_);
  and (_03666_, _14407_, _14091_);
  or (_03668_, _03666_, _03665_);
  or (_03670_, _03668_, _03664_);
  or (_03671_, _03670_, _03662_);
  and (_03672_, _03671_, _14111_);
  and (_03673_, _03672_, _03659_);
  or (_03674_, _03673_, _03641_);
  and (_03675_, _03674_, _03520_);
  and (_03676_, _01389_, _14113_);
  and (_03677_, _01467_, _11919_);
  or (_03679_, _03677_, _03676_);
  and (_03680_, _03679_, _14079_);
  or (_03681_, _14479_, _14113_);
  or (_03682_, _01244_, _11919_);
  and (_03683_, _03682_, _14094_);
  and (_03684_, _03683_, _03681_);
  or (_03686_, _14412_, _14113_);
  or (_03687_, _14251_, _11919_);
  and (_03689_, _03687_, _14091_);
  and (_03690_, _03689_, _03686_);
  or (_03691_, _14325_, _14113_);
  or (_03693_, _14247_, p0_in[7]);
  or (_03694_, _14249_, \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  and (_03695_, _03694_, _03693_);
  or (_03696_, _03695_, _11919_);
  and (_03697_, _03696_, _14103_);
  and (_03698_, _03697_, _03691_);
  or (_03699_, _03698_, _03690_);
  or (_03701_, _03699_, _03684_);
  or (_03702_, _03701_, _03680_);
  and (_03703_, _03702_, _03527_);
  and (_03704_, _03430_, _14144_);
  and (_03706_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  and (_03707_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  or (_03709_, _03707_, _03706_);
  and (_03711_, _03709_, _14113_);
  and (_03713_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  and (_03714_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  or (_03716_, _03714_, _03713_);
  and (_03717_, _03716_, _11919_);
  not (_03719_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  nor (_03721_, _11919_, _03719_);
  and (_03722_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  or (_03723_, _03722_, _03721_);
  and (_03724_, _03723_, _14103_);
  nor (_03725_, _11919_, _02653_);
  and (_03726_, _11919_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  or (_03727_, _03726_, _03725_);
  and (_03728_, _03727_, _14079_);
  or (_03729_, _03728_, _03724_);
  or (_03730_, _03729_, _03717_);
  or (_03731_, _03730_, _03711_);
  and (_03732_, _03731_, _03704_);
  and (_03734_, _11703_, _11669_);
  and (_03735_, _03734_, _14144_);
  and (_03736_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  and (_03738_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  or (_03739_, _03738_, _03736_);
  and (_03740_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  and (_03741_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  or (_03742_, _03741_, _03740_);
  or (_03744_, _03742_, _03739_);
  and (_03745_, _03744_, _11919_);
  and (_03746_, _14094_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  and (_03748_, _14091_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  or (_03749_, _03748_, _03746_);
  and (_03750_, _14103_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  and (_03751_, _14079_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  or (_03753_, _03751_, _03750_);
  or (_03754_, _03753_, _03749_);
  and (_03755_, _03754_, _14113_);
  or (_03757_, _03755_, _03745_);
  and (_03759_, _03757_, _03735_);
  or (_03760_, _03759_, _03732_);
  or (_03761_, _03760_, _03703_);
  or (_03762_, _03761_, _03675_);
  or (_03763_, _03762_, _03609_);
  or (_03764_, _03763_, _03519_);
  or (_03766_, _03764_, _03451_);
  and (_03767_, _03735_, _07646_);
  nor (_03768_, _03767_, _11931_);
  nand (_03769_, _03585_, _06930_);
  and (_03770_, _03769_, _03768_);
  and (_03771_, _03770_, _03766_);
  and (_03772_, _14103_, _11568_);
  and (_03773_, _14091_, _11763_);
  or (_03774_, _03773_, _03772_);
  and (_03775_, _03774_, _14113_);
  and (_03776_, _14103_, _07340_);
  and (_03777_, _14091_, _11882_);
  or (_03778_, _03777_, _03776_);
  and (_03779_, _03778_, _11919_);
  nor (_03780_, _11919_, _06666_);
  and (_03781_, _11919_, _07070_);
  or (_03782_, _03781_, _03780_);
  and (_03783_, _03782_, _14094_);
  nor (_03785_, _11919_, _07188_);
  and (_03786_, _11919_, _09527_);
  or (_03788_, _03786_, _03785_);
  and (_03789_, _03788_, _14079_);
  or (_03790_, _03789_, _03783_);
  or (_03792_, _03790_, _03779_);
  nor (_03793_, _03792_, _03775_);
  nor (_03795_, _03793_, _03768_);
  or (_03796_, _03795_, _03771_);
  and (_04214_, _03796_, _06444_);
  nor (_03798_, _00469_, rst);
  or (_03799_, _00468_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  nand (_03801_, _00468_, \oc8051_top_1.oc8051_sfr1.prescaler [3]);
  and (_03803_, _03801_, _03799_);
  and (_04218_, _03803_, _03798_);
  and (_04220_, _00470_, _06444_);
  nor (_03805_, _02821_, \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  nor (_03806_, _03805_, _02822_);
  and (_03808_, _03806_, _12054_);
  nor (_03809_, _00855_, _09045_);
  nor (_03810_, _03298_, _09201_);
  and (_03811_, _12032_, _11778_);
  and (_03813_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  or (_03814_, _03813_, _03811_);
  or (_03815_, _03814_, _03810_);
  or (_03817_, _03815_, _03809_);
  or (_03818_, _03817_, _03808_);
  and (_03819_, _02812_, _12662_);
  and (_03820_, _02808_, _12650_);
  or (_03822_, _03820_, _03819_);
  nand (_03823_, _03822_, _09186_);
  or (_03825_, _03822_, _09186_);
  and (_03826_, _03825_, _03823_);
  and (_03827_, _03826_, _12218_);
  or (_03829_, _03827_, _03818_);
  or (_03830_, _03829_, _03274_);
  nor (_03832_, _02793_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [14]);
  nor (_03834_, _03832_, _02794_);
  or (_03836_, _03834_, _12023_);
  and (_03838_, _03836_, _06444_);
  and (_04222_, _03838_, _03830_);
  or (_03841_, _12683_, \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  not (_03843_, _02821_);
  and (_03844_, _03843_, _12054_);
  and (_03845_, _03844_, _03841_);
  and (_03846_, _11452_, _08127_);
  and (_03847_, _12026_, _08194_);
  and (_03848_, _11726_, _12032_);
  and (_03849_, _12047_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  or (_03850_, _03849_, _03848_);
  or (_03852_, _03850_, _03847_);
  or (_03853_, _03852_, _03846_);
  nand (_03854_, _12650_, _08150_);
  nor (_03855_, _03854_, _12660_);
  nor (_03856_, _02811_, _12650_);
  nor (_03857_, _03856_, _03855_);
  nand (_03858_, _03857_, _08155_);
  or (_03859_, _03857_, _08155_);
  and (_03861_, _03859_, _03858_);
  and (_03862_, _03861_, _12218_);
  or (_03863_, _03862_, _03853_);
  or (_03865_, _03863_, _03845_);
  or (_03866_, _03865_, _03274_);
  nor (_03867_, _02792_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [13]);
  nor (_03868_, _03867_, _02793_);
  or (_03870_, _03868_, _12023_);
  and (_03871_, _03870_, _06444_);
  and (_04226_, _03871_, _03866_);
  or (_03872_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [0]);
  nand (_03873_, _07432_, _14060_);
  and (_03874_, _03873_, _06444_);
  and (_04313_, _03874_, _03872_);
  or (_03875_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [2]);
  nand (_03876_, _07432_, _14051_);
  and (_03877_, _03876_, _06444_);
  and (_04362_, _03877_, _03875_);
  not (_03878_, _11453_);
  and (_03879_, _11460_, _03878_);
  nor (_03880_, _11533_, _11455_);
  nand (_03881_, _03880_, _11492_);
  or (_03882_, _03881_, _11509_);
  or (_03883_, _03882_, _02947_);
  and (_03884_, _03883_, _11342_);
  or (_03885_, _03884_, _03879_);
  and (_04364_, _03885_, _06444_);
  and (_03886_, _14088_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  and (_03887_, _14084_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  or (_03888_, _03887_, _03886_);
  and (_03889_, _14096_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  and (_03890_, _14093_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  or (_03891_, _03890_, _03889_);
  or (_03892_, _03891_, _03888_);
  and (_03893_, _14102_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  and (_03894_, _14105_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  or (_03895_, _03894_, _03893_);
  and (_03896_, _14110_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_03897_, _14116_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  or (_03898_, _03897_, _03896_);
  or (_03899_, _03898_, _03895_);
  or (_03900_, _03899_, _03892_);
  and (_03901_, _14120_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  and (_03902_, _14122_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  or (_03903_, _03902_, _03901_);
  and (_03904_, _14124_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  and (_03905_, _14125_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  or (_03906_, _03905_, _03904_);
  or (_03907_, _03906_, _03903_);
  and (_03908_, _14130_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  and (_03909_, _14131_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  or (_03910_, _03909_, _03908_);
  and (_03912_, _14133_, \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  and (_03913_, _14134_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  or (_03915_, _03913_, _03912_);
  or (_03916_, _03915_, _03910_);
  or (_03918_, _03916_, _03907_);
  or (_03919_, _03918_, _03900_);
  and (_03920_, _14154_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03921_, _14156_, _11622_);
  or (_03922_, _03921_, _03920_);
  and (_03924_, _14150_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  and (_03925_, _14152_, \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  or (_03926_, _03925_, _03924_);
  or (_03927_, _03926_, _03922_);
  and (_03928_, _03631_, _14265_);
  and (_03929_, _03652_, _14260_);
  or (_03930_, _03929_, _03928_);
  and (_03931_, _03695_, _14224_);
  and (_03932_, _03561_, _14253_);
  or (_03933_, _03932_, _03931_);
  or (_03934_, _03933_, _03930_);
  or (_03936_, _03934_, _03927_);
  and (_03937_, _14143_, \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  and (_03938_, _14146_, \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  or (_03939_, _03938_, _03937_);
  or (_03940_, _03939_, _03936_);
  or (_03941_, _03940_, _03919_);
  and (_03942_, _03941_, _14174_);
  and (_03943_, _14175_, \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  or (_03945_, _03943_, _03942_);
  or (_03946_, _03945_, _14178_);
  or (_03947_, _14353_, _11137_);
  and (_03948_, _03947_, _06444_);
  and (_04366_, _03948_, _03946_);
  or (_03949_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9]);
  or (_03950_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_03951_, _03950_, _03949_);
  or (_03952_, _03951_, _06442_);
  and (_03953_, _03952_, _06444_);
  nand (_03954_, _03410_, _06978_);
  and (_04369_, _03954_, _03953_);
  or (_03955_, _02650_, _11137_);
  nand (_03956_, _02650_, _03719_);
  and (_03957_, _03956_, _06440_);
  and (_03959_, _03957_, _03955_);
  nor (_03960_, _06673_, _03719_);
  and (_03961_, _02659_, _06933_);
  nand (_03963_, _03961_, _06930_);
  or (_03964_, _03961_, \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  and (_03965_, _03964_, _06674_);
  and (_03966_, _03965_, _03963_);
  or (_03967_, _03966_, _03960_);
  or (_03968_, _03967_, _03959_);
  and (_04377_, _03968_, _06444_);
  or (_03969_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_03970_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8]);
  and (_03971_, _03970_, _03969_);
  and (_03972_, _03971_, _06443_);
  nand (_03973_, _06978_, _06295_);
  nand (_03974_, _10494_, _06296_);
  and (_03975_, _03974_, _00933_);
  and (_03976_, _03975_, _03973_);
  or (_04379_, _03976_, _03972_);
  and (_03977_, _06442_, _06295_);
  and (_03978_, _03977_, _11763_);
  or (_03979_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7]);
  or (_03980_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nand (_03982_, _03980_, _03979_);
  nor (_03983_, _03982_, _06442_);
  and (_03984_, _03410_, _07378_);
  or (_03985_, _03984_, _03983_);
  or (_03987_, _03985_, _03978_);
  and (_04383_, _03987_, _06444_);
  nor (_04491_, _11904_, rst);
  nand (_03988_, _06406_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  nor (_03990_, _03988_, _00238_);
  or (_03991_, _03990_, _01481_);
  and (_03992_, _03991_, _00818_);
  nand (_03993_, _00818_, _06406_);
  and (_03995_, _03993_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  or (_03997_, _03995_, _07407_);
  or (_03998_, _03997_, _03992_);
  nand (_03999_, _10494_, _07407_);
  and (_04001_, _03999_, _06444_);
  and (_04530_, _04001_, _03998_);
  or (_04002_, _07432_, \oc8051_top_1.oc8051_rom1.data_o [1]);
  nand (_04003_, _07432_, _14056_);
  and (_04004_, _04003_, _06444_);
  and (_04533_, _04004_, _04002_);
  and (_04005_, _00742_, _06933_);
  nand (_04006_, _04005_, _06930_);
  or (_04007_, _04005_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  and (_04008_, _04007_, _00748_);
  and (_04009_, _04008_, _04006_);
  nor (_04010_, _00748_, _06978_);
  or (_04012_, _04010_, _04009_);
  and (_04535_, _04012_, _06444_);
  and (_04013_, _00669_, _06933_);
  nand (_04014_, _04013_, _06930_);
  or (_04015_, _04013_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  and (_04016_, _04015_, _00678_);
  and (_04017_, _04016_, _04014_);
  nor (_04018_, _00678_, _06978_);
  or (_04019_, _04018_, _04017_);
  and (_04538_, _04019_, _06444_);
  and (_04020_, _08310_, _06678_);
  nand (_04021_, _04020_, _06930_);
  or (_04022_, _04020_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  and (_04023_, _04022_, _02416_);
  and (_04024_, _04023_, _04021_);
  nor (_04026_, _07300_, _02416_);
  or (_04027_, _04026_, _04024_);
  and (_04545_, _04027_, _06444_);
  and (_04028_, _06431_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_04029_, _04028_, _00713_);
  and (_04030_, _04029_, _06678_);
  not (_04031_, _06678_);
  or (_04032_, _00717_, _04031_);
  and (_04033_, _04032_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  or (_04034_, _04033_, _06946_);
  or (_04035_, _04034_, _04030_);
  nand (_04036_, _11589_, _06946_);
  and (_04037_, _04036_, _06444_);
  and (_04548_, _04037_, _04035_);
  and (_04038_, _06678_, _06432_);
  nand (_04039_, _04038_, _06930_);
  or (_04040_, _04038_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  and (_04041_, _04040_, _04039_);
  or (_04042_, _04041_, _02406_);
  nand (_04043_, _07069_, _06946_);
  and (_04044_, _04043_, _06444_);
  and (_04551_, _04044_, _04042_);
  and (_04045_, _06678_, _06942_);
  nand (_04046_, _04045_, _06930_);
  or (_04047_, _04045_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  and (_04048_, _04047_, _04046_);
  or (_04049_, _04048_, _02406_);
  nand (_04051_, _09526_, _06946_);
  and (_04053_, _04051_, _06444_);
  and (_04555_, _04053_, _04049_);
  not (_04054_, _14174_);
  and (_04557_, _14496_, _04054_);
  nor (_04055_, _08484_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_04056_, _04055_, _12589_);
  or (_04058_, _04056_, _12023_);
  and (_04059_, _12048_, _08230_);
  and (_04060_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [4]);
  nor (_04061_, _12128_, _12033_);
  and (_04062_, _12054_, _11650_);
  or (_04063_, _04062_, _04061_);
  or (_04064_, _04063_, _04060_);
  or (_04065_, _12207_, _12205_);
  and (_04066_, _04065_, _12208_);
  and (_04067_, _04066_, _12218_);
  or (_04068_, _04067_, _04064_);
  nor (_04069_, _04068_, _04059_);
  nand (_04070_, _04069_, _12023_);
  and (_04071_, _04070_, _06444_);
  and (_04562_, _04071_, _04058_);
  or (_04072_, _12023_, _08486_);
  and (_04073_, _12048_, _08308_);
  and (_04075_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [3]);
  nor (_04076_, _12154_, _12033_);
  and (_04077_, _12054_, _11689_);
  or (_04078_, _04077_, _04076_);
  or (_04079_, _04078_, _04075_);
  or (_04080_, _12157_, _12158_);
  not (_04081_, _04080_);
  nand (_04082_, _04081_, _12203_);
  or (_04083_, _04081_, _12203_);
  and (_04084_, _04083_, _12606_);
  and (_04085_, _04084_, _04082_);
  or (_04086_, _04085_, _04079_);
  nor (_04087_, _04086_, _04073_);
  nand (_04089_, _04087_, _12023_);
  and (_04090_, _04089_, _06444_);
  and (_04564_, _04090_, _04072_);
  and (_04091_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  nor (_04092_, _08064_, _01106_);
  or (_04093_, _04092_, _04091_);
  and (_04566_, _04093_, _06444_);
  and (_04096_, _03977_, _07378_);
  or (_04097_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or (_04098_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6]);
  nand (_04099_, _04098_, _04097_);
  nor (_04100_, _04099_, _06442_);
  and (_04101_, _03410_, _07359_);
  or (_04102_, _04101_, _04100_);
  or (_04103_, _04102_, _04096_);
  and (_04573_, _04103_, _06444_);
  and (_04104_, _12048_, _02977_);
  and (_04106_, _11452_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [2]);
  and (_04107_, _12032_, _12162_);
  and (_04108_, _12054_, _11905_);
  or (_04110_, _04108_, _04107_);
  or (_04111_, _04110_, _04106_);
  nor (_04112_, _12201_, _12199_);
  nor (_04114_, _04112_, _12202_);
  and (_04115_, _04114_, _12218_);
  or (_04116_, _04115_, _04111_);
  or (_04117_, _04116_, _04104_);
  and (_04118_, _04117_, _12023_);
  and (_04119_, _03274_, _08499_);
  or (_04120_, _04119_, _04118_);
  and (_04576_, _04120_, _06444_);
  and (_04121_, _03977_, _07359_);
  or (_04122_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5]);
  or (_04124_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nand (_04125_, _04124_, _04122_);
  nor (_04127_, _04125_, _06442_);
  and (_04128_, _03410_, _07340_);
  or (_04129_, _04128_, _04127_);
  or (_04130_, _04129_, _04121_);
  and (_04580_, _04130_, _06444_);
  not (_04132_, \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  nor (_04133_, _00856_, _04132_);
  and (_04134_, _12054_, _11794_);
  and (_04135_, _12186_, _12032_);
  or (_04136_, _04135_, _04134_);
  or (_04137_, _12196_, _12194_);
  and (_04138_, _12606_, _12198_);
  and (_04139_, _04138_, _04137_);
  or (_04140_, _04139_, _04136_);
  and (_04141_, _12048_, _07959_);
  or (_04142_, _04141_, _04140_);
  and (_04143_, _04142_, _12023_);
  or (_04144_, _04143_, _04133_);
  and (_04582_, _04144_, _06444_);
  and (_04145_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [7]);
  nor (_04146_, _07046_, _06978_);
  or (_04147_, _04146_, _04145_);
  and (_04587_, _04147_, _06444_);
  or (_04148_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or (_04149_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4]);
  nand (_04150_, _04149_, _04148_);
  nor (_04151_, _04150_, _06442_);
  and (_04152_, _03410_, _11882_);
  or (_04153_, _04152_, _04151_);
  and (_04154_, _13865_, _06295_);
  and (_04155_, _04154_, _07340_);
  or (_04156_, _04155_, _04153_);
  and (_04590_, _04156_, _06444_);
  and (_04157_, _07403_, _07402_);
  nand (_04158_, _04157_, _08310_);
  nor (_04159_, _04158_, _06930_);
  and (_04160_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  nand (_04161_, _07387_, \oc8051_top_1.oc8051_memory_interface1.int_ack );
  nor (_04162_, _07396_, _07076_);
  not (_04163_, _04162_);
  or (_04164_, _04163_, _07392_);
  or (_04165_, _04164_, _04161_);
  and (_04166_, _04165_, _04160_);
  and (_04167_, _04166_, _04158_);
  or (_04168_, _04167_, _07407_);
  or (_04169_, _04168_, _04159_);
  nand (_04170_, _07407_, _07300_);
  and (_04171_, _04170_, _06444_);
  and (_04592_, _04171_, _04169_);
  and (_04172_, _07011_, _07004_);
  nor (_04173_, _04172_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  or (_04174_, _04173_, _07024_);
  nor (_04175_, _07028_, _02860_);
  nand (_04176_, _04175_, _07026_);
  and (_04177_, _04176_, _04174_);
  nor (_04178_, _04177_, _07017_);
  and (_04179_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  or (_04180_, _04179_, _06985_);
  or (_04181_, _04180_, _04178_);
  or (_04182_, _02538_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  and (_04183_, _04182_, _09503_);
  and (_04184_, _04183_, _04181_);
  nor (_04185_, _10494_, _09503_);
  or (_04186_, _04185_, _04184_);
  and (_04595_, _04186_, _06444_);
  and (_04187_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_04188_, _04187_, _07026_);
  nand (_04189_, _07011_, _07003_);
  and (_04190_, _04189_, _02887_);
  nor (_04191_, _04190_, _04172_);
  or (_04193_, _04191_, _07017_);
  or (_04194_, _04193_, _04188_);
  or (_04196_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  and (_04197_, _04196_, _06990_);
  and (_04198_, _04197_, _04194_);
  nor (_04199_, _09503_, _06666_);
  and (_04200_, _06985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  or (_04201_, _04200_, _04199_);
  or (_04202_, _04201_, _04198_);
  and (_04597_, _04202_, _06444_);
  or (_04205_, _04162_, _07392_);
  or (_04207_, _04205_, _04161_);
  nand (_04209_, _04207_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  nand (_04211_, _04209_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  and (_04212_, _14511_, _06674_);
  or (_04213_, _04212_, _04211_);
  and (_04215_, _04213_, _07408_);
  nand (_04216_, _04212_, _06930_);
  and (_04217_, _04216_, _04215_);
  nor (_04219_, _07408_, _07069_);
  or (_04221_, _04219_, _04217_);
  and (_04803_, _04221_, _06444_);
  nand (_04806_, _11857_, _06444_);
  nand (_04808_, _11802_, _06444_);
  nand (_04810_, _11912_, _06444_);
  nor (_04812_, _11699_, rst);
  nor (_04814_, _11663_, rst);
  nor (_04822_, _11734_, rst);
  nor (_04824_, _11774_, rst);
  nor (_04223_, _01701_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff );
  or (_04224_, _04164_, _07388_);
  and (_04225_, _04224_, \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  or (_04227_, _04225_, _04223_);
  and (_04228_, _04157_, _06987_);
  or (_04229_, _04228_, _04227_);
  and (_04230_, _04229_, _07408_);
  nand (_04231_, _04228_, _06930_);
  and (_04232_, _04231_, _04230_);
  nor (_04233_, _07408_, _06666_);
  or (_04234_, _04233_, _04232_);
  and (_04826_, _04234_, _06444_);
  and (_04235_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04236_, _04235_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  and (_04237_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  and (_04238_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_04239_, _04238_, _04237_);
  and (_04240_, _04239_, _04236_);
  and (_04241_, _04240_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_04242_, _04241_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_04243_, _04242_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_04244_, _04243_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  and (_04245_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  and (_04246_, _04245_, _04244_);
  and (_04247_, _04246_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04248_, _04246_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_04249_, _04248_, _04247_);
  nor (_04250_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not (_04251_, _04250_);
  and (_04252_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  and (_04253_, _04252_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04254_, _04252_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  nor (_04255_, _04254_, _04253_);
  not (_04256_, _04255_);
  and (_04257_, _04253_, _01279_);
  nor (_04258_, _04253_, _01279_);
  nor (_04259_, _04258_, _04257_);
  nor (_04260_, _04259_, _08481_);
  and (_04261_, _04259_, \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_04262_, _04261_, _04260_);
  nor (_04263_, _04262_, _04256_);
  and (_04264_, _04259_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nor (_04265_, _04259_, _08521_);
  nor (_04266_, _04265_, _04264_);
  nor (_04267_, _04266_, _04255_);
  nor (_04268_, _04267_, _04263_);
  nor (_04269_, _04268_, _04251_);
  and (_04270_, _13796_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not (_04271_, _04270_);
  nor (_04272_, _04259_, _08515_);
  and (_04273_, _04259_, \oc8051_symbolic_cxrom1.regvalid [7]);
  nor (_04274_, _04273_, _04272_);
  nor (_04275_, _04274_, _04256_);
  and (_04276_, _04259_, \oc8051_symbolic_cxrom1.regvalid [3]);
  not (_04277_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_04278_, _04259_, _04277_);
  nor (_04279_, _04278_, _04276_);
  nor (_04280_, _04279_, _04255_);
  nor (_04281_, _04280_, _04275_);
  nor (_04282_, _04281_, _04271_);
  nor (_04283_, _04282_, _04269_);
  and (_04284_, _04259_, \oc8051_symbolic_cxrom1.regvalid [4]);
  not (_04285_, \oc8051_symbolic_cxrom1.regvalid [12]);
  nor (_04286_, _04259_, _04285_);
  nor (_04287_, _04286_, _04284_);
  nor (_04288_, _04287_, _04256_);
  and (_04289_, _04259_, \oc8051_symbolic_cxrom1.regvalid [0]);
  not (_04290_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_04291_, _04259_, _04290_);
  nor (_04292_, _04291_, _04289_);
  nor (_04293_, _04292_, _01154_);
  or (_04294_, _04293_, _04288_);
  and (_04295_, _04294_, _04252_);
  and (_04296_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _12846_);
  not (_04297_, _04296_);
  nor (_04298_, _04259_, _08546_);
  and (_04299_, _04259_, \oc8051_symbolic_cxrom1.regvalid [6]);
  nor (_04300_, _04299_, _04298_);
  nor (_04301_, _04300_, _04256_);
  and (_04302_, _04259_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_04303_, _04259_, _09302_);
  nor (_04304_, _04303_, _04302_);
  nor (_04305_, _04304_, _04255_);
  nor (_04306_, _04305_, _04301_);
  nor (_04307_, _04306_, _04297_);
  nor (_04308_, _04307_, _04295_);
  and (_04309_, _04308_, _04283_);
  and (_04310_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_04311_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [7]);
  nor (_04312_, _04311_, _04310_);
  and (_04314_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [7]);
  and (_04315_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [7]);
  nor (_04316_, _04315_, _04314_);
  and (_04317_, _04316_, _04312_);
  and (_04318_, _04317_, _04256_);
  not (_04319_, _04259_);
  and (_04320_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [7]);
  and (_04321_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [7]);
  nor (_04322_, _04321_, _04320_);
  and (_04323_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_04324_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [7]);
  nor (_04325_, _04324_, _04323_);
  and (_04326_, _04325_, _04322_);
  and (_04327_, _04326_, _04255_);
  or (_04328_, _04327_, _04319_);
  nor (_04329_, _04328_, _04318_);
  and (_04330_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_04331_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [7]);
  nor (_04332_, _04331_, _04330_);
  and (_04333_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [7]);
  and (_04334_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [7]);
  nor (_04335_, _04334_, _04333_);
  and (_04336_, _04335_, _04332_);
  and (_04337_, _04336_, _04256_);
  and (_04338_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_04339_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [7]);
  nor (_04340_, _04339_, _04338_);
  and (_04341_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [7]);
  and (_04342_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [7]);
  nor (_04343_, _04342_, _04341_);
  and (_04344_, _04343_, _04340_);
  and (_04345_, _04344_, _04255_);
  or (_04346_, _04345_, _04259_);
  nor (_04347_, _04346_, _04337_);
  nor (_04348_, _04347_, _04329_);
  nor (_04349_, _04348_, _04309_);
  and (_04350_, _04349_, _04249_);
  nor (_04351_, _04349_, _04249_);
  nor (_04352_, _04351_, _04350_);
  and (_04353_, _04244_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_04354_, _04353_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_04355_, _04354_, _04246_);
  and (_04356_, _04355_, _04349_);
  nor (_04357_, _04355_, _04349_);
  nor (_04358_, _04244_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_04359_, _04358_, _04353_);
  and (_04360_, _04359_, _04349_);
  nor (_04361_, _04243_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_04363_, _04361_, _04244_);
  and (_04365_, _04363_, _04349_);
  nor (_04367_, _04242_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_04368_, _04367_, _04243_);
  and (_04370_, _04368_, _04349_);
  nor (_04371_, _04363_, _04349_);
  nor (_04372_, _04371_, _04365_);
  nor (_04373_, _04368_, _04349_);
  nor (_04374_, _04373_, _04370_);
  not (_04375_, _04374_);
  nor (_04376_, _04241_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nor (_04378_, _04376_, _04242_);
  and (_04380_, _04378_, _04349_);
  nor (_04381_, _04378_, _04349_);
  nor (_04382_, _04240_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_04384_, _04382_, _04241_);
  and (_04385_, _04384_, _04349_);
  and (_04386_, _04237_, _04236_);
  and (_04387_, _04386_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_04388_, _04387_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_04389_, _04388_, _04240_);
  and (_04390_, _04389_, _04349_);
  nor (_04391_, _04389_, _04349_);
  nor (_04392_, _04386_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_04393_, _04392_, _04387_);
  and (_04394_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [6]);
  and (_04395_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [6]);
  nor (_04396_, _04395_, _04394_);
  and (_04397_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [6]);
  and (_04398_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [6]);
  nor (_04399_, _04398_, _04397_);
  and (_04400_, _04399_, _04396_);
  and (_04401_, _04400_, _04256_);
  and (_04402_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [6]);
  and (_04403_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [6]);
  nor (_04404_, _04403_, _04402_);
  and (_04405_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [6]);
  and (_04406_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [6]);
  nor (_04407_, _04406_, _04405_);
  and (_04408_, _04407_, _04404_);
  and (_04409_, _04408_, _04255_);
  or (_04410_, _04409_, _04259_);
  nor (_04411_, _04410_, _04401_);
  and (_04412_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [6]);
  and (_04413_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [6]);
  nor (_04414_, _04413_, _04412_);
  and (_04415_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [6]);
  and (_04416_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [6]);
  nor (_04417_, _04416_, _04415_);
  and (_04418_, _04417_, _04414_);
  nor (_04419_, _04418_, _04255_);
  and (_04420_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [6]);
  and (_04421_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [6]);
  nor (_04422_, _04421_, _04420_);
  and (_04423_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [6]);
  and (_04424_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [6]);
  nor (_04425_, _04424_, _04423_);
  and (_04426_, _04425_, _04422_);
  nor (_04427_, _04426_, _04256_);
  or (_04428_, _04427_, _04419_);
  and (_04429_, _04428_, _04259_);
  nor (_04430_, _04429_, _04411_);
  nor (_04431_, _04430_, _04309_);
  and (_04432_, _04431_, _04393_);
  nor (_04433_, _04431_, _04393_);
  nor (_04434_, _04433_, _04432_);
  not (_04435_, _04434_);
  and (_04436_, _04236_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_04437_, _04436_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  nor (_04438_, _04437_, _04386_);
  and (_04439_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [5]);
  and (_04440_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [5]);
  nor (_04441_, _04440_, _04439_);
  and (_04442_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [5]);
  and (_04443_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [5]);
  nor (_04444_, _04443_, _04442_);
  and (_04445_, _04444_, _04441_);
  and (_04446_, _04445_, _04256_);
  and (_04447_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [5]);
  and (_04448_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [5]);
  nor (_04449_, _04448_, _04447_);
  and (_04450_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [5]);
  and (_04451_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [5]);
  nor (_04452_, _04451_, _04450_);
  and (_04453_, _04452_, _04449_);
  and (_04454_, _04453_, _04255_);
  or (_04455_, _04454_, _04259_);
  nor (_04456_, _04455_, _04446_);
  and (_04457_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [5]);
  and (_04458_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [5]);
  nor (_04459_, _04458_, _04457_);
  and (_04460_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [5]);
  and (_04461_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [5]);
  nor (_04462_, _04461_, _04460_);
  and (_04463_, _04462_, _04459_);
  nor (_04464_, _04463_, _04255_);
  and (_04465_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [5]);
  and (_04466_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [5]);
  nor (_04467_, _04466_, _04465_);
  and (_04468_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [5]);
  and (_04469_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [5]);
  nor (_04470_, _04469_, _04468_);
  and (_04471_, _04470_, _04467_);
  nor (_04472_, _04471_, _04256_);
  or (_04473_, _04472_, _04464_);
  and (_04474_, _04473_, _04259_);
  nor (_04475_, _04474_, _04456_);
  nor (_04476_, _04475_, _04309_);
  and (_04477_, _04476_, _04438_);
  nor (_04478_, _04476_, _04438_);
  nor (_04479_, _04478_, _04477_);
  not (_04480_, _04479_);
  nor (_04481_, _04236_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_04482_, _04481_, _04436_);
  and (_04483_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [4]);
  and (_04484_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [4]);
  nor (_04485_, _04484_, _04483_);
  and (_04486_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [4]);
  and (_04487_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [4]);
  nor (_04488_, _04487_, _04486_);
  and (_04489_, _04488_, _04485_);
  and (_04490_, _04489_, _04256_);
  and (_04492_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [4]);
  and (_04493_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [4]);
  nor (_04494_, _04493_, _04492_);
  and (_04495_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [4]);
  and (_04496_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [4]);
  nor (_04497_, _04496_, _04495_);
  and (_04498_, _04497_, _04494_);
  and (_04499_, _04498_, _04255_);
  or (_04500_, _04499_, _04319_);
  nor (_04501_, _04500_, _04490_);
  and (_04502_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [4]);
  and (_04503_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [4]);
  nor (_04504_, _04503_, _04502_);
  and (_04505_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [4]);
  and (_04506_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [4]);
  nor (_04507_, _04506_, _04505_);
  and (_04508_, _04507_, _04504_);
  and (_04509_, _04508_, _04256_);
  and (_04510_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [4]);
  and (_04511_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [4]);
  nor (_04512_, _04511_, _04510_);
  and (_04513_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [4]);
  and (_04514_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [4]);
  nor (_04515_, _04514_, _04513_);
  and (_04516_, _04515_, _04512_);
  and (_04517_, _04516_, _04255_);
  or (_04518_, _04517_, _04259_);
  nor (_04519_, _04518_, _04509_);
  nor (_04520_, _04519_, _04501_);
  nor (_04521_, _04520_, _04309_);
  and (_04522_, _04521_, _04482_);
  and (_04523_, _04235_, _01279_);
  nor (_04524_, _04235_, _01279_);
  nor (_04525_, _04524_, _04523_);
  not (_04526_, _04525_);
  and (_04527_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [3]);
  and (_04528_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [3]);
  nor (_04529_, _04528_, _04527_);
  and (_04531_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [3]);
  and (_04532_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [3]);
  nor (_04534_, _04532_, _04531_);
  and (_04536_, _04534_, _04529_);
  and (_04537_, _04536_, _04256_);
  and (_04539_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [3]);
  and (_04540_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [3]);
  nor (_04541_, _04540_, _04539_);
  and (_04542_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [3]);
  and (_04543_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [3]);
  nor (_04544_, _04543_, _04542_);
  and (_04546_, _04544_, _04541_);
  and (_04547_, _04546_, _04255_);
  or (_04549_, _04547_, _04319_);
  nor (_04550_, _04549_, _04537_);
  and (_04552_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [3]);
  and (_04553_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [3]);
  nor (_04554_, _04553_, _04552_);
  and (_04556_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [3]);
  and (_04558_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [3]);
  nor (_04559_, _04558_, _04556_);
  and (_04560_, _04559_, _04554_);
  and (_04561_, _04560_, _04256_);
  and (_04563_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [3]);
  and (_04565_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [3]);
  nor (_04567_, _04565_, _04563_);
  and (_04568_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [3]);
  and (_04569_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [3]);
  nor (_04570_, _04569_, _04568_);
  and (_04571_, _04570_, _04567_);
  and (_04572_, _04571_, _04255_);
  or (_04574_, _04572_, _04259_);
  nor (_04575_, _04574_, _04561_);
  nor (_04577_, _04575_, _04550_);
  nor (_04578_, _04577_, _04309_);
  and (_04579_, _04578_, _04526_);
  nor (_04581_, _04578_, _04526_);
  nor (_04583_, _04581_, _04579_);
  not (_04584_, _04583_);
  and (_04585_, _12846_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_04586_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _01154_);
  nor (_04588_, _04586_, _04585_);
  not (_04589_, _04588_);
  and (_04591_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [2]);
  and (_04593_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [2]);
  nor (_04594_, _04593_, _04591_);
  and (_04596_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [2]);
  and (_04598_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [2]);
  nor (_04599_, _04598_, _04596_);
  and (_04600_, _04599_, _04594_);
  and (_04601_, _04600_, _04256_);
  and (_04602_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [2]);
  and (_04603_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [2]);
  nor (_04604_, _04603_, _04602_);
  and (_04605_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [2]);
  and (_04606_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [2]);
  nor (_04607_, _04606_, _04605_);
  and (_04608_, _04607_, _04604_);
  and (_04609_, _04608_, _04255_);
  or (_04610_, _04609_, _04319_);
  nor (_04611_, _04610_, _04601_);
  and (_04612_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [2]);
  and (_04613_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [2]);
  nor (_04614_, _04613_, _04612_);
  and (_04615_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [2]);
  and (_04616_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [2]);
  nor (_04617_, _04616_, _04615_);
  and (_04618_, _04617_, _04614_);
  and (_04619_, _04618_, _04256_);
  and (_04620_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [2]);
  and (_04621_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [2]);
  nor (_04622_, _04621_, _04620_);
  and (_04623_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [2]);
  and (_04624_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [2]);
  nor (_04625_, _04624_, _04623_);
  and (_04626_, _04625_, _04622_);
  and (_04627_, _04626_, _04255_);
  or (_04628_, _04627_, _04259_);
  nor (_04629_, _04628_, _04619_);
  nor (_04630_, _04629_, _04611_);
  nor (_04631_, _04630_, _04309_);
  and (_04632_, _04631_, _04589_);
  and (_04633_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [1]);
  and (_04634_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [1]);
  nor (_04635_, _04634_, _04633_);
  and (_04636_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [1]);
  and (_04637_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [1]);
  nor (_04638_, _04637_, _04636_);
  and (_04639_, _04638_, _04635_);
  and (_04640_, _04639_, _04256_);
  and (_04641_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [1]);
  and (_04642_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [1]);
  nor (_04643_, _04642_, _04641_);
  and (_04644_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [1]);
  and (_04645_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [1]);
  nor (_04646_, _04645_, _04644_);
  and (_04647_, _04646_, _04643_);
  and (_04648_, _04647_, _04255_);
  or (_04649_, _04648_, _04319_);
  nor (_04650_, _04649_, _04640_);
  and (_04651_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [1]);
  and (_04652_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [1]);
  nor (_04653_, _04652_, _04651_);
  and (_04654_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [1]);
  and (_04655_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [1]);
  nor (_04656_, _04655_, _04654_);
  and (_04657_, _04656_, _04653_);
  and (_04658_, _04657_, _04256_);
  and (_04659_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [1]);
  and (_04660_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [1]);
  nor (_04661_, _04660_, _04659_);
  and (_04662_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [1]);
  and (_04663_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [1]);
  nor (_04664_, _04663_, _04662_);
  and (_04665_, _04664_, _04661_);
  and (_04666_, _04665_, _04255_);
  or (_04667_, _04666_, _04259_);
  nor (_04668_, _04667_, _04658_);
  nor (_04669_, _04668_, _04650_);
  nor (_04670_, _04669_, _04309_);
  and (_04671_, _04670_, _12846_);
  and (_04672_, _04296_, \oc8051_symbolic_cxrom1.regarray[2] [0]);
  and (_04673_, _04252_, \oc8051_symbolic_cxrom1.regarray[0] [0]);
  nor (_04674_, _04673_, _04672_);
  and (_04675_, _04270_, \oc8051_symbolic_cxrom1.regarray[3] [0]);
  and (_04676_, _04250_, \oc8051_symbolic_cxrom1.regarray[1] [0]);
  nor (_04677_, _04676_, _04675_);
  and (_04678_, _04677_, _04674_);
  and (_04679_, _04678_, _04256_);
  and (_04680_, _04270_, \oc8051_symbolic_cxrom1.regarray[7] [0]);
  and (_04681_, _04250_, \oc8051_symbolic_cxrom1.regarray[5] [0]);
  nor (_04682_, _04681_, _04680_);
  and (_04683_, _04296_, \oc8051_symbolic_cxrom1.regarray[6] [0]);
  and (_04684_, _04252_, \oc8051_symbolic_cxrom1.regarray[4] [0]);
  nor (_04685_, _04684_, _04683_);
  and (_04686_, _04685_, _04682_);
  and (_04687_, _04686_, _04255_);
  or (_04688_, _04687_, _04319_);
  nor (_04689_, _04688_, _04679_);
  and (_04690_, _04296_, \oc8051_symbolic_cxrom1.regarray[10] [0]);
  and (_04691_, _04252_, \oc8051_symbolic_cxrom1.regarray[8] [0]);
  nor (_04692_, _04691_, _04690_);
  and (_04693_, _04270_, \oc8051_symbolic_cxrom1.regarray[11] [0]);
  and (_04694_, _04250_, \oc8051_symbolic_cxrom1.regarray[9] [0]);
  nor (_04695_, _04694_, _04693_);
  and (_04696_, _04695_, _04692_);
  nor (_04697_, _04696_, _04255_);
  and (_04698_, _04270_, \oc8051_symbolic_cxrom1.regarray[15] [0]);
  and (_04699_, _04250_, \oc8051_symbolic_cxrom1.regarray[13] [0]);
  nor (_04700_, _04699_, _04698_);
  and (_04701_, _04296_, \oc8051_symbolic_cxrom1.regarray[14] [0]);
  and (_04702_, _04252_, \oc8051_symbolic_cxrom1.regarray[12] [0]);
  nor (_04703_, _04702_, _04701_);
  and (_04704_, _04703_, _04700_);
  nor (_04705_, _04704_, _04256_);
  or (_04706_, _04705_, _04697_);
  and (_04707_, _04706_, _04319_);
  nor (_04708_, _04707_, _04689_);
  nor (_04709_, _04708_, _04309_);
  and (_04710_, _04709_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04711_, _04670_, _12846_);
  nor (_04712_, _04711_, _04671_);
  and (_04713_, _04712_, _04710_);
  nor (_04714_, _04713_, _04671_);
  nor (_04715_, _04631_, _04589_);
  nor (_04716_, _04715_, _04632_);
  not (_04717_, _04716_);
  nor (_04718_, _04717_, _04714_);
  nor (_04719_, _04718_, _04632_);
  nor (_04720_, _04719_, _04584_);
  nor (_04721_, _04720_, _04579_);
  nor (_04722_, _04521_, _04482_);
  nor (_04723_, _04722_, _04522_);
  not (_04724_, _04723_);
  nor (_04725_, _04724_, _04721_);
  nor (_04726_, _04725_, _04522_);
  nor (_04727_, _04726_, _04480_);
  nor (_04728_, _04727_, _04477_);
  nor (_04729_, _04728_, _04435_);
  nor (_04730_, _04729_, _04432_);
  nor (_04731_, _04730_, _04391_);
  or (_04732_, _04731_, _04390_);
  nor (_04733_, _04384_, _04349_);
  nor (_04734_, _04733_, _04385_);
  and (_04735_, _04734_, _04732_);
  nor (_04736_, _04735_, _04385_);
  nor (_04737_, _04736_, _04381_);
  nor (_04738_, _04737_, _04380_);
  nor (_04739_, _04738_, _04375_);
  and (_04740_, _04739_, _04372_);
  or (_04741_, _04740_, _04370_);
  nor (_04742_, _04741_, _04365_);
  nor (_04743_, _04359_, _04349_);
  nor (_04744_, _04743_, _04360_);
  not (_04745_, _04744_);
  nor (_04746_, _04745_, _04742_);
  nor (_04747_, _04746_, _04360_);
  nor (_04748_, _04747_, _04357_);
  or (_04749_, _04748_, _04356_);
  and (_04750_, _04749_, _04352_);
  nor (_04751_, _04750_, _04350_);
  nor (_04752_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_04753_, \oc8051_top_1.oc8051_memory_interface1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_04754_, _04753_, _04752_);
  nor (_04755_, _04754_, _04247_);
  and (_04756_, _04754_, _04247_);
  nor (_04757_, _04756_, _04755_);
  nor (_04758_, _04757_, _04349_);
  and (_04759_, _04757_, _04349_);
  nor (_04760_, _04759_, _04758_);
  nor (_04761_, _04760_, _04751_);
  and (_04762_, _04745_, _04742_);
  nor (_04763_, _04762_, _04746_);
  nor (_04764_, _04763_, _00664_);
  nor (_04765_, _04739_, _04370_);
  nand (_04766_, _04372_, _01602_);
  or (_04767_, _04372_, _01602_);
  and (_04768_, _04767_, _04766_);
  not (_04769_, _04768_);
  nor (_04770_, _04769_, _04765_);
  not (_04771_, _04349_);
  nor (_04772_, _04378_, _01150_);
  and (_04773_, _04378_, _01150_);
  or (_04774_, _04773_, _04772_);
  nand (_04775_, _04774_, _04771_);
  or (_04776_, _04774_, _04771_);
  and (_04777_, _04776_, _04775_);
  or (_04778_, _04777_, _04736_);
  nand (_04779_, _04777_, _04736_);
  and (_04780_, _04779_, _04778_);
  nor (_04781_, _04734_, _04732_);
  nor (_04782_, _04781_, _04735_);
  nor (_04783_, _04782_, _01872_);
  and (_04784_, _04782_, _01872_);
  nor (_04785_, _04390_, _04391_);
  nor (_04786_, _04785_, _04730_);
  and (_04787_, _04785_, _04730_);
  nor (_04788_, _04787_, _04786_);
  and (_04789_, _04788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  nor (_04790_, _04788_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_04791_, _04728_, _04435_);
  nor (_04792_, _04791_, _04729_);
  and (_04793_, _04792_, _01106_);
  nor (_04794_, _04792_, _01106_);
  and (_04795_, _04726_, _04480_);
  nor (_04796_, _04795_, _04727_);
  nor (_04797_, _04796_, _01128_);
  and (_04798_, _04796_, _01128_);
  and (_04799_, _04724_, _04721_);
  nor (_04800_, _04799_, _04725_);
  nor (_04801_, _04800_, _01275_);
  not (_04802_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04804_, _04719_, _04584_);
  nor (_04805_, _04804_, _04720_);
  nor (_04807_, _04805_, _04802_);
  and (_04809_, _04805_, _04802_);
  not (_04811_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04813_, _04717_, _04714_);
  nor (_04815_, _04813_, _04718_);
  and (_04816_, _04815_, _04811_);
  and (_04817_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_04818_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_04819_, _04818_, _04817_);
  not (_04820_, _04819_);
  nand (_04821_, _04820_, _04709_);
  or (_04823_, _04820_, _04709_);
  and (_04825_, _04823_, _04821_);
  not (_04827_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nor (_04828_, _04712_, _04710_);
  nor (_04829_, _04828_, _04713_);
  nor (_04830_, _04829_, _04827_);
  and (_04831_, _04829_, _04827_);
  or (_04832_, _04831_, _04830_);
  or (_04833_, _04832_, _04825_);
  nor (_04834_, _04815_, _04811_);
  or (_04835_, _04834_, _04833_);
  or (_04836_, _04835_, _04816_);
  or (_04837_, _04836_, _04809_);
  or (_04838_, _04837_, _04807_);
  and (_04839_, _04800_, _01275_);
  or (_04840_, _04839_, _04838_);
  or (_04841_, _04840_, _04801_);
  or (_04842_, _04841_, _04798_);
  or (_04843_, _04842_, _04797_);
  or (_04844_, _04843_, _04794_);
  or (_04845_, _04844_, _04793_);
  or (_04846_, _04845_, _04790_);
  or (_04847_, _04846_, _04789_);
  or (_04848_, _04847_, _04784_);
  or (_04849_, _04848_, _04783_);
  or (_04850_, _04849_, _04780_);
  or (_04851_, _04850_, _04770_);
  and (_04852_, _04738_, _04375_);
  nor (_04853_, _04852_, _04739_);
  nor (_04854_, _04853_, _01142_);
  and (_04855_, _04769_, _04765_);
  and (_04856_, _04853_, _01142_);
  or (_04857_, _04856_, _04855_);
  or (_04858_, _04857_, _04854_);
  or (_04859_, _04858_, _04851_);
  or (_04860_, _04859_, _04764_);
  nor (_04861_, _04355_, _01591_);
  and (_04862_, _04355_, _01591_);
  or (_04863_, _04862_, _04861_);
  nand (_04864_, _04863_, _04349_);
  or (_04865_, _04863_, _04349_);
  and (_04866_, _04865_, _04864_);
  and (_04867_, _04866_, _04747_);
  and (_04868_, _04763_, _00664_);
  nor (_04869_, _04866_, _04747_);
  or (_04870_, _04869_, _04868_);
  or (_04871_, _04870_, _04867_);
  or (_04872_, _04871_, _04860_);
  or (_04873_, _04872_, _04761_);
  nor (_04874_, _04749_, _04352_);
  nor (_04875_, _04874_, _04750_);
  nor (_04876_, _04875_, _01580_);
  and (_04877_, _04760_, _04751_);
  and (_04878_, _04875_, _01580_);
  or (_04879_, _04878_, _04877_);
  or (_04880_, _04879_, _04876_);
  or (_04881_, _04880_, _04873_);
  or (_04882_, _04802_, \oc8051_symbolic_cxrom1.regvalid [13]);
  or (_04883_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_04884_, _04883_, _04882_);
  and (_04885_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], _04811_);
  and (_04886_, _04885_, _04884_);
  or (_04887_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_04888_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_04889_, _04802_, \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_04890_, _04889_, _04888_);
  and (_04891_, _04890_, _04887_);
  or (_04892_, _04891_, _04886_);
  nor (_04893_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_04895_, _04893_, _04811_);
  nor (_04896_, _04895_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04897_, _04895_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_04898_, _04897_, _04896_);
  and (_04899_, _04898_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_04900_, _04893_, _04811_);
  nor (_04901_, _04900_, _04895_);
  or (_04902_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], _09063_);
  nand (_04903_, _04902_, _04901_);
  or (_04904_, _04903_, _04899_);
  and (_04905_, _04904_, _04827_);
  nand (_04906_, _04898_, _04277_);
  or (_04907_, _04898_, \oc8051_symbolic_cxrom1.regvalid [3]);
  and (_04908_, _04907_, _04906_);
  or (_04909_, _04901_, _04908_);
  and (_04911_, _04909_, _04905_);
  or (_04912_, _04911_, _04892_);
  and (_04913_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  and (_04914_, _04802_, \oc8051_symbolic_cxrom1.regvalid [0]);
  or (_04915_, _04914_, _04913_);
  and (_04917_, _04915_, _04811_);
  and (_04918_, _04802_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_04919_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_04920_, _04919_, _04918_);
  and (_04921_, _04920_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_04922_, _04921_, _04917_);
  and (_04923_, _04922_, _04827_);
  and (_04924_, _04888_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_04925_, _04924_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_04927_, _04924_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_04928_, _04927_, _04925_);
  or (_04929_, _04928_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_04930_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  nor (_04931_, _04930_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_04932_, _04931_, _04924_);
  and (_04933_, _04932_, _04882_);
  and (_04934_, _04933_, _04929_);
  or (_04936_, _04928_, \oc8051_symbolic_cxrom1.regvalid [1]);
  not (_04938_, _04932_);
  nand (_04939_, _04928_, _08521_);
  and (_04940_, _04939_, _04938_);
  and (_04941_, _04940_, _04936_);
  or (_04942_, _04941_, _04934_);
  and (_04944_, _04942_, _04923_);
  or (_04946_, _04928_, \oc8051_symbolic_cxrom1.regvalid [7]);
  or (_04947_, _04802_, \oc8051_symbolic_cxrom1.regvalid [15]);
  and (_04948_, _04947_, _04932_);
  and (_04949_, _04948_, _04946_);
  or (_04951_, _04928_, \oc8051_symbolic_cxrom1.regvalid [3]);
  nand (_04952_, _04928_, _04277_);
  and (_04953_, _04952_, _04938_);
  and (_04954_, _04953_, _04951_);
  or (_04955_, _04954_, _04949_);
  and (_04956_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_04957_, _04802_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_04958_, _04957_, _04811_);
  or (_04959_, _04958_, _04956_);
  or (_04961_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_04962_, _04802_, \oc8051_symbolic_cxrom1.regvalid [10]);
  and (_04963_, _04962_, _04961_);
  or (_04964_, _04963_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_04965_, _04964_, _04959_);
  and (_04967_, _04965_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_04968_, _04920_, _04885_);
  or (_04969_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_04970_, _04802_, \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_04971_, _04970_, _04888_);
  and (_04972_, _04971_, _04969_);
  or (_04973_, _04972_, _04968_);
  and (_04974_, _04973_, _04967_);
  and (_04975_, _04974_, _04955_);
  or (_04976_, _04975_, _04944_);
  not (_04977_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_04978_, _04973_, _04965_);
  and (_04979_, _04978_, _04977_);
  and (_04980_, _04979_, _04976_);
  and (_04981_, _04980_, _04912_);
  or (_04982_, _04827_, \oc8051_symbolic_cxrom1.regvalid [2]);
  or (_04983_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [0]);
  and (_04985_, _04983_, _04982_);
  or (_04987_, _04985_, _04898_);
  or (_04988_, _04827_, \oc8051_symbolic_cxrom1.regvalid [10]);
  or (_04989_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_symbolic_cxrom1.regvalid [8]);
  nand (_04991_, _04989_, _04988_);
  and (_04992_, _04991_, _04898_);
  nor (_04993_, _04992_, _04901_);
  and (_04994_, _04993_, _04987_);
  and (_04995_, _04898_, \oc8051_symbolic_cxrom1.regvalid [12]);
  or (_04996_, _04918_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  or (_04997_, _04996_, _04995_);
  and (_04998_, _04898_, \oc8051_symbolic_cxrom1.regvalid [14]);
  or (_04999_, _04957_, _04827_);
  or (_05000_, _04999_, _04998_);
  and (_05001_, _05000_, _04901_);
  and (_05002_, _05001_, _04997_);
  or (_05003_, _05002_, _04994_);
  or (_05004_, _04928_, \oc8051_symbolic_cxrom1.regvalid [6]);
  or (_05005_, _04802_, \oc8051_symbolic_cxrom1.regvalid [14]);
  and (_05006_, _05005_, _05004_);
  or (_05007_, _05006_, _04938_);
  nand (_05008_, _04928_, _09302_);
  or (_05009_, _04928_, \oc8051_symbolic_cxrom1.regvalid [2]);
  and (_05010_, _05009_, _05008_);
  or (_05011_, _05010_, _04932_);
  and (_05012_, _05011_, _05007_);
  or (_05013_, _05012_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  not (_05014_, \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_05015_, _04928_, _05014_);
  and (_05016_, _04928_, \oc8051_symbolic_cxrom1.regvalid [8]);
  or (_05017_, _05016_, _05015_);
  and (_05018_, _05017_, _04938_);
  or (_05019_, _04928_, \oc8051_symbolic_cxrom1.regvalid [4]);
  or (_05021_, _04802_, \oc8051_symbolic_cxrom1.regvalid [12]);
  and (_05022_, _05021_, _04932_);
  and (_05023_, _05022_, _05019_);
  or (_05024_, _05023_, _04827_);
  or (_05025_, _05024_, _05018_);
  or (_05026_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  and (_05027_, _05026_, _04947_);
  or (_05028_, _05027_, _04811_);
  or (_05029_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  or (_05030_, _04802_, \oc8051_symbolic_cxrom1.regvalid [11]);
  and (_05032_, _05030_, _05029_);
  or (_05033_, _05032_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05034_, _05033_, _05028_);
  and (_05035_, _05034_, _04930_);
  and (_05036_, _04827_, \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  or (_05037_, _04884_, _04811_);
  or (_05038_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  or (_05039_, _04802_, \oc8051_symbolic_cxrom1.regvalid [9]);
  and (_05040_, _05039_, _05038_);
  or (_05041_, _05040_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05042_, _05041_, _05037_);
  and (_05043_, _05042_, _05036_);
  or (_05044_, _05043_, _05035_);
  and (_05045_, _05034_, _04827_);
  or (_05046_, _05045_, _04892_);
  and (_05047_, _05046_, _05044_);
  and (_05048_, _05047_, _05025_);
  and (_05049_, _05048_, _05013_);
  and (_05050_, _05049_, _05003_);
  or (_05051_, _05050_, _04981_);
  nor (_05052_, _04250_, _01154_);
  and (_05053_, _05052_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_05054_, _05052_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_05055_, _05054_, _05053_);
  nand (_05056_, _05055_, _08515_);
  nor (_05057_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05058_, _05057_, _13796_);
  nor (_05059_, _05058_, _05052_);
  nor (_05060_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [7]);
  not (_05061_, _05060_);
  and (_05062_, _05061_, _05059_);
  and (_05063_, _05062_, _05056_);
  not (_05064_, _05059_);
  and (_05065_, _05055_, \oc8051_symbolic_cxrom1.regvalid [11]);
  nor (_05066_, _05055_, _08508_);
  or (_05067_, _05066_, _05065_);
  and (_05068_, _05067_, _05064_);
  or (_05069_, _05068_, _05063_);
  and (_05070_, _05069_, _04250_);
  or (_05071_, _05055_, \oc8051_symbolic_cxrom1.regvalid [4]);
  and (_05072_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04285_);
  nor (_05073_, _05072_, _05064_);
  and (_05074_, _05073_, _05071_);
  and (_05075_, _05055_, \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_05076_, _05055_, _05014_);
  or (_05077_, _05076_, _05075_);
  and (_05078_, _05077_, _05064_);
  or (_05079_, _05078_, _05074_);
  and (_05080_, _05079_, _04296_);
  or (_05081_, _05080_, _05070_);
  nand (_05082_, _05055_, _08546_);
  nor (_05083_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [6]);
  not (_05084_, _05083_);
  and (_05085_, _05084_, _05059_);
  and (_05086_, _05085_, _05082_);
  or (_05087_, _05055_, \oc8051_symbolic_cxrom1.regvalid [2]);
  nand (_05088_, _05055_, _09302_);
  and (_05089_, _05088_, _05087_);
  and (_05090_, _05089_, _05064_);
  or (_05091_, _05090_, _05086_);
  and (_05092_, _05091_, _04252_);
  or (_05093_, _05055_, \oc8051_symbolic_cxrom1.regvalid [5]);
  and (_05094_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08481_);
  nor (_05095_, _05094_, _05064_);
  and (_05096_, _05095_, _05093_);
  or (_05097_, _05055_, \oc8051_symbolic_cxrom1.regvalid [1]);
  nand (_05098_, _05055_, _08521_);
  and (_05099_, _05098_, _05064_);
  and (_05100_, _05099_, _05097_);
  or (_05101_, _05100_, _05096_);
  and (_05102_, _05101_, _04270_);
  or (_05103_, _05102_, _05092_);
  or (_05104_, _05103_, _05081_);
  and (_05105_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08515_);
  nor (_05106_, _05105_, _01154_);
  and (_05107_, _05106_, _05061_);
  and (_05108_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04277_);
  nor (_05109_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [3]);
  nor (_05110_, _05109_, _05108_);
  and (_05111_, _05110_, _01154_);
  nor (_05112_, _05111_, _05107_);
  nor (_05113_, _05112_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  not (_05114_, _04235_);
  and (_05115_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_05116_, _01279_, \oc8051_symbolic_cxrom1.regvalid [9]);
  nor (_05117_, _05116_, _05115_);
  nor (_05118_, _05117_, _05114_);
  nor (_05119_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [5]);
  nor (_05120_, _05119_, _05094_);
  and (_05121_, _05120_, _04586_);
  nor (_05122_, _05121_, _05118_);
  not (_05123_, _05122_);
  nor (_05124_, _05123_, _05113_);
  nor (_05125_, _05124_, _13796_);
  not (_05126_, _05125_);
  and (_05127_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08546_);
  nor (_05128_, _05127_, _01154_);
  and (_05129_, _05128_, _05084_);
  and (_05130_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _09302_);
  nor (_05131_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [2]);
  nor (_05132_, _05131_, _05130_);
  and (_05133_, _05132_, _01154_);
  nor (_05134_, _05133_, _05129_);
  nor (_05135_, _05134_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_05136_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [4]);
  nor (_05137_, _05136_, _05072_);
  and (_05138_, _05137_, _04586_);
  nor (_05139_, _05138_, _05135_);
  nor (_05140_, _05139_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05141_, _04270_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  and (_05142_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _05014_);
  nor (_05143_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [8]);
  nor (_05144_, _05143_, _05142_);
  and (_05145_, _05144_, _05141_);
  nor (_05146_, _05145_, _05140_);
  and (_05147_, _05146_, _05126_);
  and (_05148_, _05137_, _04585_);
  nor (_05149_, _05148_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05150_, _05134_, _12846_);
  and (_05151_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _04290_);
  nor (_05152_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [0]);
  nor (_05153_, _05152_, _05151_);
  and (_05154_, _05153_, _05057_);
  nor (_05155_, _05154_, _05150_);
  and (_05156_, _05155_, _05149_);
  nor (_05157_, _05112_, _12846_);
  nor (_05158_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], \oc8051_symbolic_cxrom1.regvalid [1]);
  and (_05159_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _08521_);
  nor (_05160_, _05159_, _05158_);
  and (_05161_, _05160_, _05057_);
  and (_05162_, _05120_, _04585_);
  or (_05163_, _05162_, _13796_);
  or (_05164_, _05163_, _05161_);
  nor (_05165_, _05164_, _05157_);
  nor (_05166_, _05165_, _05156_);
  not (_05167_, _08064_);
  nor (_05168_, _05167_, first_instr);
  nand (_05169_, _05168_, _05166_);
  or (_05170_, _05169_, _05147_);
  nor (_05171_, _05170_, _04309_);
  and (_05172_, _05171_, _05104_);
  and (_05173_, _05172_, _05051_);
  nor (_05174_, \oc8051_symbolic_cxrom1.regarray[0] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05175_, _09720_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05176_, _05175_, _05174_);
  and (_05177_, _05176_, _05057_);
  nor (_05178_, _05177_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_05179_, \oc8051_symbolic_cxrom1.regarray[4] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05180_, _10197_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05181_, _05180_, _05179_);
  and (_05182_, _05181_, _04585_);
  not (_05183_, _05182_);
  nor (_05184_, \oc8051_symbolic_cxrom1.regarray[2] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05185_, _09963_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05186_, _05185_, _05184_);
  and (_05187_, _05186_, _04586_);
  nor (_05188_, \oc8051_symbolic_cxrom1.regarray[6] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05189_, _10406_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05190_, _05189_, _05188_);
  and (_05191_, _05190_, _04235_);
  nor (_05192_, _05191_, _05187_);
  and (_05193_, _05192_, _05183_);
  and (_05194_, _05193_, _05178_);
  nor (_05195_, \oc8051_symbolic_cxrom1.regarray[8] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05196_, _10624_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05197_, _05196_, _05195_);
  and (_05198_, _05197_, _05057_);
  nor (_05199_, _05198_, _01279_);
  nor (_05200_, \oc8051_symbolic_cxrom1.regarray[12] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05201_, _12365_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05202_, _05201_, _05200_);
  and (_05203_, _05202_, _04585_);
  not (_05204_, _05203_);
  nor (_05205_, \oc8051_symbolic_cxrom1.regarray[10] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05206_, _11249_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05207_, _05206_, _05205_);
  and (_05208_, _05207_, _04586_);
  nor (_05209_, \oc8051_symbolic_cxrom1.regarray[14] [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05210_, _12729_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05211_, _05210_, _05209_);
  and (_05212_, _05211_, _04235_);
  nor (_05213_, _05212_, _05208_);
  and (_05214_, _05213_, _05204_);
  and (_05215_, _05214_, _05199_);
  nor (_05216_, _05215_, _05194_);
  and (_05217_, _05216_, _05166_);
  nor (_05218_, \oc8051_symbolic_cxrom1.regarray[0] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05219_, _09697_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05220_, _05219_, _05218_);
  and (_05221_, _05220_, _05057_);
  nor (_05222_, _05221_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_05223_, \oc8051_symbolic_cxrom1.regarray[4] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05224_, _10183_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05225_, _05224_, _05223_);
  and (_05226_, _05225_, _04585_);
  not (_05227_, _05226_);
  nor (_05228_, \oc8051_symbolic_cxrom1.regarray[2] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05229_, _09941_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05230_, _05229_, _05228_);
  and (_05231_, _05230_, _04586_);
  nor (_05232_, \oc8051_symbolic_cxrom1.regarray[6] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05233_, _10396_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05234_, _05233_, _05232_);
  and (_05235_, _05234_, _04235_);
  nor (_05236_, _05235_, _05231_);
  and (_05237_, _05236_, _05227_);
  and (_05238_, _05237_, _05222_);
  nor (_05239_, \oc8051_symbolic_cxrom1.regarray[8] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05240_, _10608_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05241_, _05240_, _05239_);
  and (_05242_, _05241_, _05057_);
  nor (_05243_, _05242_, _01279_);
  nor (_05244_, \oc8051_symbolic_cxrom1.regarray[12] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05245_, _12347_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05246_, _05245_, _05244_);
  and (_05247_, _05246_, _04585_);
  not (_05248_, _05247_);
  nor (_05249_, \oc8051_symbolic_cxrom1.regarray[10] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05250_, _11230_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05251_, _05250_, _05249_);
  and (_05252_, _05251_, _04586_);
  nor (_05253_, \oc8051_symbolic_cxrom1.regarray[14] [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05254_, _12717_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05255_, _05254_, _05253_);
  and (_05256_, _05255_, _04235_);
  nor (_05257_, _05256_, _05252_);
  and (_05258_, _05257_, _05248_);
  and (_05259_, _05258_, _05243_);
  nor (_05260_, _05259_, _05238_);
  and (_05261_, _05260_, _05166_);
  nor (_05262_, _05261_, _05217_);
  nor (_05263_, \oc8051_symbolic_cxrom1.regarray[0] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05264_, _09775_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05265_, _05264_, _05263_);
  and (_05266_, _05265_, _05057_);
  nor (_05267_, _05266_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_05268_, \oc8051_symbolic_cxrom1.regarray[4] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05269_, _10245_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05270_, _05269_, _05268_);
  and (_05271_, _05270_, _04585_);
  not (_05272_, _05271_);
  nor (_05273_, \oc8051_symbolic_cxrom1.regarray[2] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05274_, _10027_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05275_, _05274_, _05273_);
  and (_05276_, _05275_, _04586_);
  nor (_05277_, \oc8051_symbolic_cxrom1.regarray[6] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05278_, _10454_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05279_, _05278_, _05277_);
  and (_05280_, _05279_, _04235_);
  nor (_05281_, _05280_, _05276_);
  and (_05282_, _05281_, _05272_);
  and (_05283_, _05282_, _05267_);
  nor (_05284_, \oc8051_symbolic_cxrom1.regarray[8] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05285_, _10672_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05286_, _05285_, _05284_);
  and (_05287_, _05286_, _05057_);
  nor (_05288_, _05287_, _01279_);
  nor (_05289_, \oc8051_symbolic_cxrom1.regarray[12] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05290_, _12416_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05291_, _05290_, _05289_);
  and (_05292_, _05291_, _04585_);
  not (_05293_, _05292_);
  nor (_05294_, \oc8051_symbolic_cxrom1.regarray[10] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05295_, _11305_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05296_, _05295_, _05294_);
  and (_05297_, _05296_, _04586_);
  nor (_05298_, \oc8051_symbolic_cxrom1.regarray[14] [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05299_, _12779_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05300_, _05299_, _05298_);
  and (_05301_, _05300_, _04235_);
  nor (_05302_, _05301_, _05297_);
  and (_05303_, _05302_, _05293_);
  and (_05304_, _05303_, _05288_);
  nor (_05305_, _05304_, _05283_);
  and (_05306_, _05305_, _05166_);
  nor (_05307_, \oc8051_symbolic_cxrom1.regarray[2] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05308_, _10011_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05309_, _05308_, _05307_);
  and (_05310_, _05309_, _04586_);
  nor (_05311_, \oc8051_symbolic_cxrom1.regarray[4] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05312_, _10233_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05313_, _05312_, _05311_);
  and (_05314_, _05313_, _04585_);
  nor (_05315_, \oc8051_symbolic_cxrom1.regarray[6] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05316_, _10443_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05317_, _05316_, _05315_);
  and (_05318_, _05317_, _04235_);
  nor (_05319_, \oc8051_symbolic_cxrom1.regarray[0] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05320_, _09761_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05321_, _05320_, _05319_);
  and (_05322_, _05321_, _05057_);
  or (_05323_, _05322_, _05318_);
  or (_05324_, _05323_, _05314_);
  or (_05325_, _05324_, _05310_);
  and (_05326_, _05325_, _01279_);
  nor (_05327_, \oc8051_symbolic_cxrom1.regarray[10] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05328_, _11292_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05329_, _05328_, _05327_);
  and (_05330_, _05329_, _04586_);
  nor (_05331_, \oc8051_symbolic_cxrom1.regarray[12] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05332_, _12403_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05333_, _05332_, _05331_);
  and (_05334_, _05333_, _04585_);
  nor (_05335_, \oc8051_symbolic_cxrom1.regarray[14] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05336_, _12766_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05337_, _05336_, _05335_);
  and (_05338_, _05337_, _04235_);
  nor (_05339_, \oc8051_symbolic_cxrom1.regarray[8] [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05340_, _10660_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05341_, _05340_, _05339_);
  and (_05342_, _05341_, _05057_);
  or (_05343_, _05342_, _05338_);
  or (_05344_, _05343_, _05334_);
  or (_05345_, _05344_, _05330_);
  and (_05346_, _05345_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_05347_, _05346_, _05326_);
  and (_05348_, _05347_, _05166_);
  nor (_05349_, _05348_, _05306_);
  and (_05350_, _05349_, _05262_);
  nor (_05351_, \oc8051_symbolic_cxrom1.regarray[2] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05352_, _09985_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05353_, _05352_, _05351_);
  and (_05354_, _05353_, _04586_);
  nor (_05355_, \oc8051_symbolic_cxrom1.regarray[4] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05356_, _10209_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05357_, _05356_, _05355_);
  and (_05358_, _05357_, _04585_);
  nor (_05359_, \oc8051_symbolic_cxrom1.regarray[0] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05360_, _09734_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05361_, _05360_, _05359_);
  and (_05362_, _05361_, _05057_);
  nor (_05363_, \oc8051_symbolic_cxrom1.regarray[6] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05364_, _10420_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05365_, _05364_, _05363_);
  and (_05366_, _05365_, _04235_);
  or (_05367_, _05366_, _05362_);
  or (_05368_, _05367_, _05358_);
  or (_05369_, _05368_, _05354_);
  and (_05370_, _05369_, _01279_);
  nor (_05371_, \oc8051_symbolic_cxrom1.regarray[10] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05372_, _11267_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05373_, _05372_, _05371_);
  and (_05374_, _05373_, _04586_);
  nor (_05375_, \oc8051_symbolic_cxrom1.regarray[12] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05376_, _12378_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05377_, _05376_, _05375_);
  and (_05378_, _05377_, _04585_);
  nor (_05379_, \oc8051_symbolic_cxrom1.regarray[8] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05380_, _10636_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05381_, _05380_, _05379_);
  and (_05382_, _05381_, _05057_);
  nor (_05383_, \oc8051_symbolic_cxrom1.regarray[14] [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05384_, _12741_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05385_, _05384_, _05383_);
  and (_05386_, _05385_, _04235_);
  or (_05387_, _05386_, _05382_);
  or (_05388_, _05387_, _05378_);
  or (_05389_, _05388_, _05374_);
  and (_05390_, _05389_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_05391_, _05390_, _05370_);
  and (_05392_, _05391_, _05166_);
  nor (_05393_, \oc8051_symbolic_cxrom1.regarray[2] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05394_, _09998_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05395_, _05394_, _05393_);
  and (_05396_, _05395_, _04586_);
  nor (_05397_, \oc8051_symbolic_cxrom1.regarray[4] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05398_, _10221_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05399_, _05398_, _05397_);
  and (_05400_, _05399_, _04585_);
  nor (_05401_, \oc8051_symbolic_cxrom1.regarray[0] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05402_, _09749_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05403_, _05402_, _05401_);
  and (_05404_, _05403_, _05057_);
  nor (_05405_, \oc8051_symbolic_cxrom1.regarray[6] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05406_, _10431_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05407_, _05406_, _05405_);
  and (_05408_, _05407_, _04235_);
  or (_05409_, _05408_, _05404_);
  or (_05410_, _05409_, _05400_);
  or (_05411_, _05410_, _05396_);
  and (_05412_, _05411_, _01279_);
  nor (_05413_, \oc8051_symbolic_cxrom1.regarray[10] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05414_, _11279_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05415_, _05414_, _05413_);
  and (_05416_, _05415_, _04586_);
  nor (_05417_, \oc8051_symbolic_cxrom1.regarray[12] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05418_, _12391_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05419_, _05418_, _05417_);
  and (_05420_, _05419_, _04585_);
  nor (_05421_, \oc8051_symbolic_cxrom1.regarray[8] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05422_, _10649_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05423_, _05422_, _05421_);
  and (_05424_, _05423_, _05057_);
  nor (_05425_, \oc8051_symbolic_cxrom1.regarray[14] [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05426_, _12754_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05427_, _05426_, _05425_);
  and (_05428_, _05427_, _04235_);
  or (_05429_, _05428_, _05424_);
  or (_05430_, _05429_, _05420_);
  or (_05431_, _05430_, _05416_);
  and (_05432_, _05431_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_05433_, _05432_, _05412_);
  and (_05434_, _05433_, _05166_);
  nor (_05435_, _05434_, _05392_);
  nor (_05436_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[0] [7]);
  and (_05437_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08600_);
  nor (_05438_, _05437_, _05436_);
  and (_05439_, _05438_, _05057_);
  nor (_05440_, _05439_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  nor (_05441_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[4] [7]);
  and (_05442_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08595_);
  nor (_05443_, _05442_, _05441_);
  and (_05444_, _05443_, _04585_);
  not (_05445_, _05444_);
  nor (_05446_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[2] [7]);
  and (_05447_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08584_);
  nor (_05448_, _05447_, _05446_);
  and (_05449_, _05448_, _04586_);
  nor (_05450_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[6] [7]);
  and (_05451_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08590_);
  nor (_05452_, _05451_, _05450_);
  and (_05453_, _05452_, _04235_);
  nor (_05454_, _05453_, _05449_);
  and (_05455_, _05454_, _05445_);
  and (_05456_, _05455_, _05440_);
  nor (_05457_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[8] [7]);
  and (_05458_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08576_);
  nor (_05459_, _05458_, _05457_);
  and (_05460_, _05459_, _05057_);
  nor (_05461_, _05460_, _01279_);
  nor (_05462_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[12] [7]);
  and (_05463_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08571_);
  nor (_05464_, _05463_, _05462_);
  and (_05465_, _05464_, _04585_);
  not (_05466_, _05465_);
  nor (_05467_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[10] [7]);
  and (_05468_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08565_);
  nor (_05469_, _05468_, _05467_);
  and (_05470_, _05469_, _04586_);
  nor (_05471_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], \oc8051_symbolic_cxrom1.regarray[14] [7]);
  and (_05472_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _08560_);
  nor (_05473_, _05472_, _05471_);
  and (_05474_, _05473_, _04235_);
  nor (_05475_, _05474_, _05470_);
  and (_05476_, _05475_, _05466_);
  and (_05477_, _05476_, _05461_);
  nor (_05478_, _05477_, _05456_);
  and (_05479_, _05478_, _05166_);
  nor (_05480_, \oc8051_symbolic_cxrom1.regarray[2] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05481_, _10042_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05482_, _05481_, _05480_);
  and (_05483_, _05482_, _04586_);
  nor (_05484_, \oc8051_symbolic_cxrom1.regarray[4] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05485_, _10258_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05486_, _05485_, _05484_);
  and (_05487_, _05486_, _04585_);
  nor (_05488_, \oc8051_symbolic_cxrom1.regarray[6] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05489_, _10469_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05490_, _05489_, _05488_);
  and (_05491_, _05490_, _04235_);
  nor (_05492_, \oc8051_symbolic_cxrom1.regarray[0] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05493_, _09792_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05494_, _05493_, _05492_);
  and (_05495_, _05494_, _05057_);
  or (_05496_, _05495_, _05491_);
  or (_05497_, _05496_, _05487_);
  or (_05498_, _05497_, _05483_);
  and (_05499_, _05498_, _01279_);
  nor (_05500_, \oc8051_symbolic_cxrom1.regarray[10] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05501_, _11318_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05502_, _05501_, _05500_);
  and (_05503_, _05502_, _04586_);
  nor (_05504_, \oc8051_symbolic_cxrom1.regarray[12] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05505_, _12429_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05506_, _05505_, _05504_);
  and (_05507_, _05506_, _04585_);
  nor (_05508_, \oc8051_symbolic_cxrom1.regarray[14] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05509_, _12794_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05510_, _05509_, _05508_);
  and (_05511_, _05510_, _04235_);
  nor (_05512_, \oc8051_symbolic_cxrom1.regarray[8] [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05513_, _10685_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05514_, _05513_, _05512_);
  and (_05515_, _05514_, _05057_);
  or (_05516_, _05515_, _05511_);
  or (_05517_, _05516_, _05507_);
  or (_05518_, _05517_, _05503_);
  and (_05519_, _05518_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  or (_05520_, _05519_, _05499_);
  and (_05521_, _05520_, _05166_);
  not (_05522_, _05521_);
  and (_05523_, _05522_, _05479_);
  and (_05524_, _05523_, _05435_);
  and (_05525_, _05524_, _05350_);
  and (_05526_, _05525_, _05173_);
  and (_05527_, _05526_, _04881_);
  not (_05528_, _05479_);
  nand (_05529_, _05348_, _05305_);
  and (_05530_, _05392_, _05217_);
  nor (_05531_, _05530_, _05433_);
  nor (_05532_, _05531_, _05529_);
  not (_05533_, _05261_);
  and (_05534_, _05435_, _05533_);
  and (_05535_, _05534_, _05217_);
  not (_05536_, _05260_);
  not (_05537_, _05216_);
  not (_05538_, _05433_);
  and (_05539_, _05538_, _05392_);
  and (_05540_, _05539_, _05537_);
  and (_05541_, _05540_, _05536_);
  or (_05542_, _05541_, _05535_);
  or (_05543_, _05542_, _05532_);
  and (_05544_, _05543_, _05521_);
  not (_05545_, _05306_);
  nor (_05546_, _05520_, _05545_);
  and (_05547_, _05546_, _05540_);
  and (_05548_, _05540_, _05261_);
  and (_05549_, _05548_, _05545_);
  or (_05550_, _05549_, _05547_);
  or (_05551_, _05550_, _05544_);
  and (_05552_, _05551_, _05528_);
  and (_05553_, _05535_, _05545_);
  not (_05554_, _05305_);
  and (_05555_, _05521_, _05554_);
  and (_05556_, _05555_, _05534_);
  and (_05557_, _05521_, _05305_);
  and (_05558_, _05557_, _05548_);
  or (_05559_, _05558_, _05556_);
  or (_05560_, _05559_, _05553_);
  and (_05561_, _05560_, _05479_);
  and (_05562_, _05348_, _05554_);
  and (_05563_, _05562_, _05540_);
  not (_05564_, _05348_);
  and (_05565_, _05434_, _05564_);
  and (_05566_, _05530_, _05564_);
  or (_05567_, _05566_, _05565_);
  or (_05568_, _05567_, _05563_);
  and (_05569_, _05568_, _05523_);
  and (_05570_, _05534_, _05306_);
  and (_05571_, _05570_, _05523_);
  and (_05572_, _05548_, _05564_);
  and (_05573_, _05572_, _05521_);
  or (_05574_, _05573_, _05571_);
  or (_05575_, _05574_, _05569_);
  or (_05576_, _05575_, _05561_);
  or (_05577_, _05576_, _05552_);
  nor (_05578_, _04359_, _00664_);
  and (_05579_, _04359_, _00664_);
  or (_05580_, _05579_, _05578_);
  or (_05581_, _05580_, _04863_);
  and (_05582_, _04249_, _01580_);
  nor (_05583_, _04249_, _01580_);
  or (_05584_, _05583_, _05582_);
  or (_05585_, _05584_, _04757_);
  or (_05586_, _05585_, _05581_);
  nor (_05587_, _04363_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_05588_, _04363_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nor (_05589_, _05588_, _05587_);
  nor (_05590_, _04368_, _01142_);
  and (_05591_, _04368_, _01142_);
  or (_05592_, _05591_, _05590_);
  nor (_05593_, _04438_, _01128_);
  and (_05594_, _04438_, _01128_);
  or (_05595_, _05594_, _05593_);
  nor (_05596_, _04393_, _01106_);
  and (_05597_, _04393_, _01106_);
  or (_05598_, _05597_, _05596_);
  or (_05599_, _05598_, _05595_);
  and (_05600_, _04525_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_05601_, _04525_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_05602_, _05601_, _05600_);
  and (_05603_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_05604_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  nor (_05605_, _05604_, _05603_);
  nand (_05606_, _05605_, _04819_);
  and (_05607_, _04588_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  nor (_05608_, _04588_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05609_, _05608_, _05607_);
  or (_05610_, _05609_, _05606_);
  or (_05611_, _05610_, _05602_);
  nor (_05612_, _04482_, _01275_);
  and (_05613_, _04482_, _01275_);
  or (_05614_, _05613_, _05612_);
  or (_05615_, _05614_, _05611_);
  nor (_05616_, _04384_, _01872_);
  or (_05617_, _05616_, _05615_);
  or (_05618_, _05617_, _05599_);
  or (_05619_, _05618_, _05592_);
  and (_05620_, _04389_, _01076_);
  and (_05621_, _04384_, _01872_);
  nor (_05622_, _04389_, _01076_);
  or (_05623_, _05622_, _05621_);
  or (_05624_, _05623_, _05620_);
  or (_05625_, _05624_, _04774_);
  or (_05626_, _05625_, _05619_);
  or (_05627_, _05626_, _05589_);
  or (_05628_, _05627_, _05586_);
  and (_05629_, _05628_, _05577_);
  and (_05630_, _05261_, _05217_);
  and (_05631_, _05630_, _05435_);
  and (_05632_, _05541_, _05349_);
  or (_05633_, _05632_, _05631_);
  nor (_05634_, _05305_, _05260_);
  and (_05635_, _05634_, _05392_);
  nor (_05636_, _05635_, _05350_);
  nor (_05637_, _05636_, _05479_);
  or (_05638_, _05637_, _05633_);
  and (_05639_, _05638_, _05522_);
  and (_05640_, _05547_, _05564_);
  or (_05641_, _05539_, _05306_);
  or (_05642_, _05433_, _05536_);
  and (_05643_, _05642_, _05521_);
  and (_05644_, _05643_, _05641_);
  or (_05645_, _05644_, _05640_);
  and (_05646_, _05645_, _05479_);
  nand (_05647_, _05478_, _05217_);
  nor (_05648_, _05647_, _05642_);
  or (_05649_, _05648_, _05566_);
  and (_05650_, _05649_, _05521_);
  nor (_05651_, _05521_, _05479_);
  nand (_05652_, _05347_, _05545_);
  nor (_05653_, _05652_, _05434_);
  or (_05654_, _05653_, _05651_);
  and (_05655_, _05654_, _05530_);
  and (_05656_, _05522_, _05434_);
  not (_05657_, _05478_);
  or (_05658_, _05562_, _05657_);
  and (_05659_, _05658_, _05656_);
  nor (_05660_, _05478_, _05305_);
  and (_05661_, _05660_, _05434_);
  and (_05662_, _05565_, _05521_);
  or (_05663_, _05662_, _05661_);
  or (_05664_, _05663_, _05659_);
  or (_05665_, _05664_, _05655_);
  or (_05666_, _05665_, _05650_);
  or (_05667_, _05666_, _05646_);
  or (_05668_, _05667_, _05639_);
  nor (_05669_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05670_, _04368_, _13796_);
  nor (_05671_, _05670_, _05669_);
  and (_05672_, _05671_, _01142_);
  and (_05673_, _04247_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05674_, _05673_, _00601_);
  nor (_05675_, _05673_, _00601_);
  or (_05676_, _05675_, _05674_);
  nor (_05677_, _05676_, _00584_);
  or (_05678_, _05677_, _05672_);
  and (_05679_, _04244_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05680_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  and (_05681_, \oc8051_top_1.oc8051_memory_interface1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_05682_, _05681_, _05680_);
  nand (_05683_, _05682_, _05679_);
  or (_05684_, _05682_, _05679_);
  and (_05685_, _05684_, _05683_);
  and (_05686_, _05676_, _00584_);
  or (_05687_, _05686_, _05685_);
  or (_05688_, _05687_, _05678_);
  nor (_05689_, _05671_, _01142_);
  and (_05690_, _04387_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05691_, _05690_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  and (_05692_, _05690_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_05693_, _05692_, _05691_);
  nor (_05694_, _05693_, _01076_);
  and (_05695_, _04259_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nor (_05696_, _04259_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  or (_05697_, _05696_, _05695_);
  or (_05698_, _05697_, _05694_);
  and (_05699_, _04236_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05700_, _05699_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_05701_, _05699_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_05702_, _05701_, _05700_);
  nor (_05703_, _05702_, _01275_);
  and (_05704_, _05702_, _01275_);
  or (_05705_, _05704_, _05703_);
  and (_05706_, _04386_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05707_, _05706_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_05708_, _05707_, _05690_);
  nor (_05709_, _05708_, _01106_);
  and (_05710_, _05700_, _01110_);
  nor (_05711_, _05700_, _01110_);
  nor (_05712_, _05711_, _05710_);
  nor (_05713_, _05712_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_05714_, _05712_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_05715_, _05605_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  or (_05716_, _05605_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05717_, _05716_, _05715_);
  or (_05718_, _05717_, _04819_);
  nor (_05719_, _04255_, _04811_);
  and (_05720_, _04255_, _04811_);
  or (_05721_, _05720_, _05719_);
  or (_05722_, _05721_, _05718_);
  or (_05723_, _05722_, _05714_);
  or (_05724_, _05723_, _05713_);
  or (_05725_, _05724_, _05709_);
  or (_05726_, _05725_, _05705_);
  or (_05727_, _05726_, _05698_);
  and (_05728_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _13796_);
  and (_05729_, _04378_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nor (_05730_, _05729_, _05728_);
  nor (_05731_, _05730_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_05732_, _05693_, _01076_);
  and (_05733_, _05730_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  or (_05734_, _05733_, _05732_);
  or (_05735_, _05734_, _05731_);
  or (_05736_, _05735_, _05727_);
  or (_05737_, _05736_, _05689_);
  and (_05738_, _05708_, _01106_);
  or (_05739_, _04355_, _13796_);
  or (_05740_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05741_, _05740_, _05739_);
  nor (_05742_, _05741_, _01591_);
  or (_05743_, _08066_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  nand (_05744_, _04363_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05745_, _05744_, _05743_);
  nor (_05746_, _05745_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or (_05747_, _05746_, _05742_);
  or (_05748_, _05747_, _05738_);
  or (_05749_, _05748_, _05737_);
  nand (_05750_, _04246_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  and (_05751_, _05750_, _00621_);
  nor (_05752_, _05751_, _05673_);
  nor (_05753_, _05752_, _01580_);
  and (_05754_, _05752_, _01580_);
  or (_05755_, _05754_, _05753_);
  and (_05756_, _05741_, _01591_);
  or (_05757_, _05756_, _05755_);
  and (_05758_, _05699_, _04239_);
  and (_05759_, _05758_, _01066_);
  nor (_05760_, _05758_, _01066_);
  or (_05761_, _05760_, _05759_);
  nor (_05762_, _05761_, _01872_);
  and (_05763_, _05761_, _01872_);
  or (_05764_, _05763_, _05762_);
  and (_05765_, _05745_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  or (_05766_, _05765_, _05764_);
  or (_05767_, _05766_, _05757_);
  or (_05768_, _05767_, _05749_);
  or (_05769_, _05768_, _05688_);
  and (_05770_, _05769_, _05668_);
  and (_05771_, _05558_, _05348_);
  and (_05772_, _05529_, _05521_);
  and (_05773_, _05772_, _05631_);
  or (_05774_, _05773_, _05771_);
  and (_05775_, _05774_, _05528_);
  and (_05776_, _05435_, _05262_);
  and (_05777_, _05776_, _05562_);
  and (_05778_, _05572_, _05545_);
  or (_05779_, _05778_, _05777_);
  and (_05780_, _05779_, _05523_);
  or (_05781_, _05780_, _05775_);
  and (_05782_, _05053_, _04239_);
  and (_05783_, _05782_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  and (_05784_, _05783_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_05785_, _05784_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  and (_05786_, _05785_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_05787_, _05785_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  nor (_05788_, _05787_, _05786_);
  nor (_05789_, _05788_, _01602_);
  and (_05790_, _05788_, _01602_);
  or (_05791_, _05790_, _05789_);
  nor (_05792_, _05784_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  nor (_05793_, _05792_, _05785_);
  nor (_05794_, _05793_, _01142_);
  not (_05795_, _05786_);
  nor (_05796_, _05795_, _05682_);
  or (_05797_, _05796_, _05794_);
  and (_05798_, _05793_, _01142_);
  and (_05799_, _05795_, _05682_);
  or (_05800_, _05799_, _05798_);
  or (_05801_, _05800_, _05797_);
  nor (_05802_, _05782_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  nor (_05803_, _05802_, _05783_);
  nor (_05804_, _05803_, _01872_);
  or (_05805_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  nand (_05806_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  and (_05807_, _05806_, _05805_);
  nand (_05808_, _05807_, _05783_);
  or (_05809_, _05807_, _05783_);
  and (_05810_, _05809_, _05808_);
  or (_05811_, _05810_, _05804_);
  and (_05812_, _05803_, _01872_);
  and (_05813_, _05053_, _04237_);
  and (_05814_, _05813_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_05815_, _05814_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  nor (_05816_, _05815_, _05782_);
  and (_05817_, _05816_, _01076_);
  or (_05818_, _05817_, _05812_);
  or (_05819_, _05818_, _05811_);
  nor (_05820_, _05813_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  nor (_05821_, _05820_, _05814_);
  nor (_05822_, _05821_, _01106_);
  and (_05823_, _05821_, _01106_);
  nor (_05824_, _05055_, _04802_);
  and (_05825_, _05055_, _04802_);
  or (_05826_, _05825_, _05824_);
  nand (_05827_, _05717_, _04820_);
  and (_05828_, _05059_, _04811_);
  nor (_05829_, _05059_, _04811_);
  or (_05830_, _05829_, _05828_);
  or (_05831_, _05830_, _05827_);
  or (_05832_, _05831_, _05826_);
  or (_05833_, _05832_, _05823_);
  or (_05834_, _05833_, _05822_);
  nor (_05835_, _05816_, _01076_);
  or (_05836_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_05837_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_05838_, _05837_, _05836_);
  and (_05839_, _05053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  or (_05840_, _05839_, _05838_);
  nand (_05841_, _05839_, _05838_);
  and (_05842_, _05841_, _05840_);
  nor (_05843_, _05053_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  nor (_05844_, _05843_, _05839_);
  and (_05845_, _05844_, _01275_);
  nor (_05846_, _05844_, _01275_);
  or (_05847_, _05846_, _05845_);
  or (_05848_, _05847_, _05842_);
  or (_05849_, _05848_, _05835_);
  or (_05850_, _05849_, _05834_);
  or (_05851_, _05850_, _05819_);
  or (_05852_, _05851_, _05801_);
  or (_05853_, _05852_, _05791_);
  and (_05854_, _05786_, _04245_);
  and (_05855_, _05786_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  nor (_05856_, _05855_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  nor (_05857_, _05856_, _05854_);
  and (_05858_, _05857_, _01591_);
  nor (_05859_, _05857_, _01591_);
  or (_05860_, _05859_, _05858_);
  or (_05861_, _05860_, _05853_);
  and (_05862_, _05854_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_05863_, _05854_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  nor (_05864_, _05863_, _05862_);
  nor (_05865_, _05864_, _01580_);
  and (_05866_, _05864_, _01580_);
  or (_05867_, _05866_, _05865_);
  or (_05868_, _05867_, _05861_);
  nor (_05869_, _05862_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  and (_05870_, _05862_, \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  nor (_05871_, _05870_, _05869_);
  nor (_05872_, _05871_, _00584_);
  and (_05873_, _05871_, _00584_);
  or (_05874_, _05873_, _05872_);
  or (_05875_, _05874_, _05868_);
  and (_05876_, _05875_, _05781_);
  or (_05877_, _05876_, _05770_);
  or (_05878_, _05877_, _05629_);
  and (_05879_, _05878_, _05173_);
  or (_05880_, _04670_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  nand (_05881_, _04670_, \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  and (_05882_, _05881_, _05880_);
  and (_05883_, _04709_, _04977_);
  nor (_05884_, _04709_, _04977_);
  or (_05885_, _05884_, _05883_);
  or (_05886_, _05885_, _05882_);
  or (_05887_, _04578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  nand (_05888_, _04578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  and (_05889_, _05888_, _05887_);
  and (_05890_, _04631_, _04811_);
  nor (_05891_, _04631_, _04811_);
  or (_05892_, _05891_, _05890_);
  or (_05893_, _05892_, _05889_);
  or (_05894_, _05893_, _05886_);
  or (_05895_, _04476_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  nand (_05896_, _04476_, \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  and (_05897_, _05896_, _05895_);
  nor (_05898_, _04521_, _01275_);
  and (_05899_, _04521_, _01275_);
  or (_05900_, _05899_, _05898_);
  or (_05901_, _05900_, _05897_);
  and (_05902_, _04349_, _01076_);
  nor (_05903_, _04349_, _01076_);
  or (_05904_, _05903_, _05902_);
  nor (_05905_, _04431_, _01106_);
  and (_05906_, _04431_, _01106_);
  or (_05907_, _05906_, _05905_);
  or (_05908_, _05907_, _05904_);
  or (_05909_, _05908_, _05901_);
  or (_05910_, _05909_, _05894_);
  or (_05911_, _05479_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  nand (_05912_, _05479_, \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  and (_05913_, _05912_, _05911_);
  or (_05914_, _05913_, _05589_);
  or (_05915_, _05306_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  nand (_05916_, _05306_, \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  and (_05917_, _05916_, _05915_);
  nor (_05918_, _05521_, _01150_);
  and (_05919_, _05521_, _01150_);
  or (_05920_, _05919_, _05918_);
  or (_05921_, _05920_, _05917_);
  or (_05922_, _05921_, _05914_);
  or (_05923_, _05922_, _05586_);
  or (_05924_, _05923_, _05910_);
  and (_05925_, _05261_, _05537_);
  and (_05926_, _05925_, _05435_);
  and (_05927_, _05926_, _05173_);
  and (_05928_, _05927_, _05924_);
  and (_05929_, _05357_, _04586_);
  and (_05930_, _05365_, _04585_);
  and (_05931_, _05361_, _04235_);
  or (_05932_, _05931_, _05930_);
  or (_05933_, _05932_, _05929_);
  and (_05934_, _05353_, _05057_);
  or (_05935_, _05934_, _04526_);
  or (_05936_, _05935_, _05933_);
  and (_05937_, _05377_, _04586_);
  or (_05938_, _05937_, _04525_);
  and (_05939_, _05381_, _04235_);
  and (_05940_, _05373_, _05057_);
  and (_05941_, _05385_, _04585_);
  or (_05942_, _05941_, _05940_);
  or (_05943_, _05942_, _05939_);
  or (_05944_, _05943_, _05938_);
  nand (_05945_, _05944_, _05936_);
  nor (_05946_, _05945_, _05147_);
  nand (_05947_, _05946_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  or (_05948_, _05946_, \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  and (_05949_, _05948_, _05947_);
  and (_05950_, _05399_, _04586_);
  or (_05951_, _05950_, _04526_);
  and (_05952_, _05403_, _04235_);
  and (_05953_, _05395_, _05057_);
  and (_05954_, _05407_, _04585_);
  or (_05955_, _05954_, _05953_);
  or (_05956_, _05955_, _05952_);
  or (_05957_, _05956_, _05951_);
  and (_05958_, _05419_, _04586_);
  or (_05959_, _05958_, _04525_);
  and (_05960_, _05423_, _04235_);
  and (_05961_, _05415_, _05057_);
  and (_05962_, _05427_, _04585_);
  or (_05963_, _05962_, _05961_);
  or (_05964_, _05963_, _05960_);
  or (_05965_, _05964_, _05959_);
  nand (_05966_, _05965_, _05957_);
  nor (_05967_, _05966_, _05147_);
  nor (_05968_, _05967_, _04802_);
  and (_05969_, _05967_, _04802_);
  or (_05970_, _05969_, _05968_);
  or (_05971_, _05970_, _05949_);
  and (_05972_, _05181_, _04586_);
  or (_05973_, _05972_, _04526_);
  and (_05974_, _05176_, _04235_);
  and (_05975_, _05186_, _05057_);
  and (_05976_, _05190_, _04585_);
  or (_05977_, _05976_, _05975_);
  or (_05978_, _05977_, _05974_);
  or (_05979_, _05978_, _05973_);
  and (_05980_, _05202_, _04586_);
  or (_05981_, _05980_, _04525_);
  and (_05982_, _05197_, _04235_);
  and (_05983_, _05207_, _05057_);
  and (_05984_, _05211_, _04585_);
  or (_05985_, _05984_, _05983_);
  or (_05986_, _05985_, _05982_);
  or (_05987_, _05986_, _05981_);
  nand (_05988_, _05987_, _05979_);
  nor (_05989_, _05988_, _05147_);
  and (_05990_, _05989_, _04827_);
  nor (_05991_, _05989_, _04827_);
  or (_05992_, _05991_, _05990_);
  and (_05993_, _05225_, _04586_);
  or (_05994_, _05993_, _04526_);
  and (_05995_, _05220_, _04235_);
  and (_05996_, _05230_, _05057_);
  and (_05997_, _05234_, _04585_);
  or (_05998_, _05997_, _05996_);
  or (_05999_, _05998_, _05995_);
  or (_06000_, _05999_, _05994_);
  and (_06001_, _05246_, _04586_);
  or (_06002_, _06001_, _04525_);
  and (_06003_, _05241_, _04235_);
  and (_06004_, _05251_, _05057_);
  and (_06005_, _05255_, _04585_);
  or (_06006_, _06005_, _06004_);
  or (_06007_, _06006_, _06003_);
  or (_06008_, _06007_, _06002_);
  nand (_06009_, _06008_, _06000_);
  nor (_06010_, _06009_, _05147_);
  nor (_06011_, _06010_, _04977_);
  and (_06012_, _06010_, _04977_);
  or (_06013_, _06012_, _06011_);
  or (_06014_, _06013_, _05992_);
  or (_06015_, _06014_, _05971_);
  not (_06016_, _05147_);
  and (_06017_, _05313_, _04586_);
  nor (_06018_, _06017_, _04526_);
  and (_06019_, _05321_, _04235_);
  not (_06020_, _06019_);
  and (_06021_, _05309_, _05057_);
  and (_06022_, _05317_, _04585_);
  nor (_06023_, _06022_, _06021_);
  and (_06024_, _06023_, _06020_);
  and (_06025_, _06024_, _06018_);
  and (_06026_, _05337_, _04585_);
  and (_06027_, _05333_, _04586_);
  and (_06028_, _05341_, _04235_);
  or (_06029_, _06028_, _06027_);
  nor (_06030_, _06029_, _06026_);
  and (_06031_, _05329_, _05057_);
  nor (_06032_, _06031_, _04525_);
  and (_06033_, _06032_, _06030_);
  nor (_06034_, _06033_, _06025_);
  and (_06035_, _06034_, _06016_);
  nand (_06036_, _06035_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  or (_06037_, _06035_, \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  and (_06038_, _06037_, _06036_);
  and (_06039_, _05296_, _05057_);
  and (_06040_, _05300_, _04585_);
  and (_06041_, _05286_, _04235_);
  and (_06042_, _05291_, _04586_);
  or (_06043_, _06042_, _06041_);
  or (_06044_, _06043_, _06040_);
  or (_06045_, _06044_, _06039_);
  and (_06046_, _06045_, _04526_);
  and (_06047_, _05275_, _05057_);
  and (_06048_, _05279_, _04585_);
  and (_06049_, _05265_, _04235_);
  and (_06050_, _05270_, _04586_);
  or (_06051_, _06050_, _06049_);
  or (_06052_, _06051_, _06048_);
  or (_06053_, _06052_, _06047_);
  and (_06054_, _06053_, _04525_);
  or (_06055_, _06054_, _06046_);
  and (_06056_, _06055_, _06016_);
  and (_06057_, _06056_, _01128_);
  nor (_06058_, _06056_, _01128_);
  or (_06059_, _06058_, _06057_);
  or (_06060_, _06059_, _06038_);
  and (_06061_, _05510_, _04585_);
  and (_06062_, _05506_, _04586_);
  nor (_06063_, _06062_, _06061_);
  and (_06064_, _05502_, _05057_);
  and (_06065_, _05514_, _01279_);
  nor (_06066_, _06065_, _06064_);
  and (_06067_, _06066_, _06063_);
  nor (_06068_, _06067_, _04525_);
  and (_06069_, _05490_, _04585_);
  and (_06070_, _05486_, _04586_);
  nor (_06071_, _06070_, _06069_);
  and (_06072_, _05482_, _05057_);
  and (_06073_, _05494_, _04235_);
  nor (_06074_, _06073_, _06072_);
  and (_06075_, _06074_, _06071_);
  nor (_06076_, _06075_, _04526_);
  nor (_06077_, _06076_, _06068_);
  nor (_06078_, _06077_, _05147_);
  and (_06079_, _06078_, _01106_);
  nor (_06080_, _06078_, _01106_);
  or (_06081_, _06080_, _06079_);
  and (_06082_, _05459_, _01279_);
  and (_06083_, _05469_, _05057_);
  and (_06084_, _05464_, _04586_);
  and (_06085_, _05473_, _04585_);
  or (_06086_, _06085_, _06084_);
  or (_06087_, _06086_, _06083_);
  or (_06088_, _06087_, _06082_);
  and (_06089_, _06088_, _04526_);
  and (_06090_, _05438_, _04235_);
  and (_06091_, _05443_, _04586_);
  and (_06092_, _05448_, _05057_);
  and (_06093_, _05452_, _04585_);
  or (_06094_, _06093_, _06092_);
  or (_06095_, _06094_, _06091_);
  or (_06096_, _06095_, _06090_);
  and (_06097_, _06096_, _04525_);
  or (_06098_, _06097_, _06089_);
  and (_06099_, _06098_, _06016_);
  nand (_06100_, _06099_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  or (_06101_, _06099_, \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  and (_06102_, _06101_, _06100_);
  or (_06103_, _06102_, _06081_);
  or (_06104_, _06103_, _06060_);
  or (_06105_, _06104_, _06015_);
  or (_06106_, _04670_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  nand (_06107_, _04670_, \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  and (_06108_, _06107_, _06106_);
  nor (_06109_, _04709_, _01872_);
  and (_06110_, _04709_, _01872_);
  or (_06111_, _06110_, _06109_);
  or (_06112_, _06111_, _06108_);
  or (_06113_, _04578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  nand (_06114_, _04578_, \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  and (_06115_, _06114_, _06113_);
  and (_06116_, _04631_, _01142_);
  nor (_06117_, _04631_, _01142_);
  or (_06118_, _06117_, _06116_);
  or (_06119_, _06118_, _06115_);
  or (_06120_, _06119_, _06112_);
  or (_06121_, _04476_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  nand (_06122_, _04476_, \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  and (_06123_, _06122_, _06121_);
  nor (_06124_, _04521_, _00664_);
  and (_06125_, _04521_, _00664_);
  or (_06126_, _06125_, _06124_);
  or (_06127_, _06126_, _06123_);
  and (_06128_, _04349_, _00584_);
  nor (_06129_, _04349_, _00584_);
  or (_06130_, _06129_, _06128_);
  and (_06131_, _04431_, _01580_);
  nor (_06132_, _04431_, _01580_);
  or (_06133_, _06132_, _06131_);
  or (_06134_, _06133_, _06130_);
  or (_06135_, _06134_, _06127_);
  or (_06136_, _06135_, _06120_);
  or (_06137_, _06136_, _06105_);
  and (_06138_, _05651_, _05553_);
  and (_06139_, _06138_, _05173_);
  and (_06140_, _06139_, _06137_);
  or (_06141_, _06140_, _05928_);
  or (_06142_, _06141_, _05879_);
  or (property_invalid, _06142_, _05527_);
  and (_06143_, _05167_, first_instr);
  or (_00000_, _06143_, rst);
  and (_06144_, _07046_, \oc8051_top_1.oc8051_indi_addr1.buff[5] [6]);
  nor (_06145_, _10494_, _07046_);
  or (_06146_, _06145_, _06144_);
  and (_04894_, _06146_, _06444_);
  and (_06147_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  and (_06148_, _06147_, _07026_);
  and (_06149_, _07011_, _06996_);
  nor (_06150_, _06149_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  nor (_06151_, _06150_, _09507_);
  or (_06152_, _06151_, _07017_);
  or (_06153_, _06152_, _06148_);
  nor (_06154_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  nor (_06155_, _06154_, _06985_);
  and (_06156_, _06155_, _06153_);
  nor (_06157_, _10494_, _02538_);
  or (_06158_, _06157_, _06156_);
  or (_06159_, _06158_, _06989_);
  or (_06160_, _09503_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  and (_06161_, _06160_, _06444_);
  and (_04910_, _06161_, _06159_);
  and (_06162_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_06163_, _06162_, _07026_);
  and (_06164_, _02515_, _03116_);
  nor (_06165_, _06164_, _06149_);
  or (_06166_, _06165_, _07017_);
  or (_06167_, _06166_, _06163_);
  or (_06168_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  and (_06169_, _06168_, _02538_);
  and (_06170_, _06169_, _06167_);
  nor (_06171_, _02538_, _06666_);
  or (_06172_, _06171_, _06989_);
  or (_06173_, _06172_, _06170_);
  nand (_06174_, _06989_, _03116_);
  and (_06175_, _06174_, _06444_);
  and (_04916_, _06175_, _06173_);
  and (_06176_, _07011_, _07002_);
  or (_06177_, _06176_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_06178_, _06177_, _04189_);
  and (_06179_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  and (_06180_, _06179_, _07026_);
  or (_06181_, _06180_, _06178_);
  and (_06182_, _06181_, _07035_);
  and (_06183_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  or (_06184_, _06183_, _06985_);
  or (_06185_, _06184_, _06182_);
  or (_06186_, _02538_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  and (_06187_, _06186_, _09503_);
  and (_06188_, _06187_, _06185_);
  nor (_06189_, _07188_, _09503_);
  or (_06190_, _06189_, _06188_);
  and (_04926_, _06190_, _06444_);
  not (_06191_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  nand (_06192_, _07011_, _07001_);
  and (_06193_, _06192_, _06191_);
  or (_06194_, _06193_, _06176_);
  nor (_06195_, _07028_, _02903_);
  nand (_06196_, _06195_, _07026_);
  and (_06197_, _06196_, _06194_);
  nor (_06198_, _06197_, _07017_);
  and (_06199_, _07017_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  or (_06200_, _06199_, _06985_);
  or (_06201_, _06200_, _06198_);
  nand (_06202_, _06985_, _06191_);
  and (_06203_, _06202_, _09503_);
  and (_06204_, _06203_, _06201_);
  nor (_06205_, _07300_, _09503_);
  or (_06206_, _06205_, _06204_);
  and (_04935_, _06206_, _06444_);
  and (_06207_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  and (_06208_, _06207_, _07026_);
  and (_06209_, _07011_, _07000_);
  or (_06210_, _06209_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  and (_06211_, _06210_, _06192_);
  or (_06212_, _06211_, _07017_);
  or (_06213_, _06212_, _06208_);
  nor (_06214_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  nor (_06215_, _06214_, _06985_);
  and (_06216_, _06215_, _06213_);
  and (_06217_, _06985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  or (_06218_, _06217_, _06989_);
  or (_06219_, _06218_, _06216_);
  nand (_06220_, _11589_, _06989_);
  and (_06221_, _06220_, _06444_);
  and (_04937_, _06221_, _06219_);
  and (_06222_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  nor (_06223_, _08064_, _01275_);
  or (_06224_, _06223_, _06222_);
  and (_04943_, _06224_, _06444_);
  and (_06225_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  and (_06226_, _06225_, _07026_);
  and (_06227_, _07011_, _06999_);
  nor (_06228_, _06227_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  nor (_06229_, _06228_, _06209_);
  or (_06230_, _06229_, _07017_);
  or (_06231_, _06230_, _06226_);
  nor (_06232_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  nor (_06233_, _06232_, _06985_);
  and (_06234_, _06233_, _06231_);
  and (_06235_, _06985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  or (_06236_, _06235_, _06989_);
  or (_06237_, _06236_, _06234_);
  nand (_06238_, _07069_, _06989_);
  and (_06239_, _06238_, _06444_);
  and (_04945_, _06239_, _06237_);
  and (_06240_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  nor (_06241_, _08064_, _04802_);
  or (_06242_, _06241_, _06240_);
  and (_04950_, _06242_, _06444_);
  or (_06243_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3]);
  or (_06244_, _03404_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  nand (_06245_, _06244_, _06243_);
  nor (_06246_, _06245_, _06442_);
  and (_06247_, _03410_, _07070_);
  or (_06248_, _06247_, _06246_);
  and (_06249_, _04154_, _11882_);
  or (_06250_, _06249_, _06248_);
  and (_04960_, _06250_, _06444_);
  and (_06251_, _07029_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  and (_06252_, _06251_, _07026_);
  and (_06253_, _07011_, _06998_);
  nor (_06254_, _06253_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  nor (_06255_, _06254_, _06227_);
  or (_06256_, _06255_, _07017_);
  or (_06257_, _06256_, _06252_);
  nor (_06258_, _07035_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  nor (_06259_, _06258_, _06985_);
  and (_06260_, _06259_, _06257_);
  and (_06261_, _06985_, \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  or (_06262_, _06261_, _06989_);
  or (_06263_, _06262_, _06260_);
  nand (_06264_, _09526_, _06989_);
  and (_06265_, _06264_, _06444_);
  and (_04966_, _06265_, _06263_);
  or (_06266_, _00936_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2]);
  not (_06267_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  nand (_06268_, _00936_, _06267_);
  nand (_06269_, _06268_, _06266_);
  nor (_06270_, _06269_, _06442_);
  and (_06271_, _03410_, _09527_);
  or (_06272_, _06271_, _06270_);
  and (_06273_, _04154_, _07070_);
  or (_06274_, _06273_, _06272_);
  and (_04984_, _06274_, _06444_);
  or (_06275_, _00935_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  nand (_06276_, _00935_, _06267_);
  and (_06277_, _06276_, _06275_);
  and (_06278_, _06277_, _13849_);
  and (_06279_, _13847_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0]);
  or (_06280_, _06279_, \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1]);
  and (_06281_, _06280_, _13836_);
  nor (_06282_, _06281_, _06278_);
  nor (_06283_, _06282_, _06442_);
  and (_06284_, _03977_, _09527_);
  or (_06285_, _06284_, _06283_);
  and (_04986_, _06285_, _06444_);
  and (_06286_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  nor (_06287_, _08064_, _04811_);
  or (_06288_, _06287_, _06286_);
  and (_04990_, _06288_, _06444_);
  and (_06289_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  nor (_06290_, _08064_, _04827_);
  or (_06291_, _06290_, _06289_);
  and (_05020_, _06291_, _06444_);
  and (_06292_, _08064_, \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  nor (_06293_, _08064_, _04977_);
  or (_06294_, _06293_, _06292_);
  and (_05031_, _06294_, _06444_);
  dff (first_instr, _00000_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [0], _14555_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [1], _14556_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [2], _14557_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [3], _14558_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [4], _14559_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [5], _14560_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [6], _14561_);
  dff (\oc8051_symbolic_cxrom1.regarray[10] [7], _14562_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [0], _14600_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [1], _14601_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [2], _14602_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [3], _14603_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [4], _14604_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [5], _14605_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [6], _14606_);
  dff (\oc8051_symbolic_cxrom1.regarray[9] [7], _14607_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [0], _09446_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [1], _09449_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [2], _14594_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [3], _14595_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [4], _14596_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [5], _14597_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [6], _14598_);
  dff (\oc8051_symbolic_cxrom1.regarray[8] [7], _14599_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [0], _14586_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [1], _14587_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [2], _14588_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [3], _14589_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [4], _14590_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [5], _14591_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [6], _14592_);
  dff (\oc8051_symbolic_cxrom1.regarray[7] [7], _14593_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [0], _14563_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [1], _14564_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [2], _14565_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [3], _14566_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [4], _14567_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [5], _14568_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [6], _14569_);
  dff (\oc8051_symbolic_cxrom1.regarray[11] [7], _14570_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [0], _09240_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [1], _09245_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [2], _09248_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [3], _09253_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [4], _09258_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [5], _09261_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [6], _09265_);
  dff (\oc8051_symbolic_cxrom1.regarray[6] [7], _09270_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [0], _09148_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [1], _09150_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [2], _09153_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [3], _09156_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [4], _09159_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [5], _09162_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [6], _09166_);
  dff (\oc8051_symbolic_cxrom1.regarray[5] [7], _09170_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [0], _08741_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [1], _08743_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [2], _08745_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [3], _08750_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [4], _08755_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [5], _08757_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [6], _08762_);
  dff (\oc8051_symbolic_cxrom1.regarray[1] [7], _08767_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [0], _08621_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [1], _08625_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [2], _08629_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [3], _08633_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [4], _08637_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [5], _08641_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [6], _08647_);
  dff (\oc8051_symbolic_cxrom1.regarray[0] [7], _08650_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [0], _14581_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [1], _08943_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [2], _08945_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [3], _08948_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [4], _08951_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [5], _08954_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [6], _08957_);
  dff (\oc8051_symbolic_cxrom1.regarray[3] [7], _08960_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [0], _08851_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [1], _08854_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [2], _08858_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [3], _08861_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [4], _08864_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [5], _14580_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [6], _08873_);
  dff (\oc8051_symbolic_cxrom1.regarray[2] [7], _08876_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [0], _09044_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [1], _09047_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [2], _14582_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [3], _14583_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [4], _14584_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [5], _14585_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [6], _09058_);
  dff (\oc8051_symbolic_cxrom1.regarray[4] [7], _09061_);
  dff (\oc8051_symbolic_cxrom1.regvalid [0], _07097_);
  dff (\oc8051_symbolic_cxrom1.regvalid [1], _07129_);
  dff (\oc8051_symbolic_cxrom1.regvalid [2], _07165_);
  dff (\oc8051_symbolic_cxrom1.regvalid [3], _07212_);
  dff (\oc8051_symbolic_cxrom1.regvalid [4], _07279_);
  dff (\oc8051_symbolic_cxrom1.regvalid [5], _07337_);
  dff (\oc8051_symbolic_cxrom1.regvalid [6], _07395_);
  dff (\oc8051_symbolic_cxrom1.regvalid [7], _07485_);
  dff (\oc8051_symbolic_cxrom1.regvalid [8], _07563_);
  dff (\oc8051_symbolic_cxrom1.regvalid [9], _07663_);
  dff (\oc8051_symbolic_cxrom1.regvalid [10], _07759_);
  dff (\oc8051_symbolic_cxrom1.regvalid [11], _07867_);
  dff (\oc8051_symbolic_cxrom1.regvalid [12], _07977_);
  dff (\oc8051_symbolic_cxrom1.regvalid [13], _08118_);
  dff (\oc8051_symbolic_cxrom1.regvalid [14], _08240_);
  dff (\oc8051_symbolic_cxrom1.regvalid [15], _07051_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [0], _14572_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [1], _14573_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [2], _14574_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [3], _14575_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [4], _14576_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [5], _14577_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [6], _14578_);
  dff (\oc8051_symbolic_cxrom1.regarray[15] [7], _14579_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [0], _09955_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [1], _09960_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [2], _09964_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [3], _09969_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [4], _09974_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [5], _09976_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [6], _09981_);
  dff (\oc8051_symbolic_cxrom1.regarray[14] [7], _09983_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [0], _14571_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [1], _09872_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [2], _09877_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [3], _09880_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [4], _09884_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [5], _09887_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [6], _09890_);
  dff (\oc8051_symbolic_cxrom1.regarray[13] [7], _09894_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [0], _09784_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [1], _09786_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [2], _09789_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [3], _09791_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [4], _09793_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [5], _09796_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [6], _09799_);
  dff (\oc8051_symbolic_cxrom1.regarray[12] [7], _09801_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0], _13422_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1], _13050_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2], _13046_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3], _12889_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4], _04074_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5], _04203_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [0], _04088_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.cycle [1], _04192_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [0], _03293_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [1], _11898_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [2], _11916_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [3], _11913_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [4], _04094_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [5], _12057_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [6], _12317_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_rem [7], _04195_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [0], _11176_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.cycle [1], _12304_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [0], _11252_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [1], _11248_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [2], _11222_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [3], _11308_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [4], _11304_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [5], _11298_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [6], _11219_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [7], _07878_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [8], _11141_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [9], _11159_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [10], _11154_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [11], _11239_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [12], _11214_);
  dff (\oc8051_top_1.oc8051_alu1.oc8051_mul1.tmp_mul [13], _11198_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [0], _06713_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [1], _06715_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [2], _06717_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [3], _06719_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [4], _06721_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [5], _06724_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [6], _06726_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op1_r [7], _06566_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [2], _04491_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op2_r [7], _06569_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [0], _08694_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [6], _03747_);
  dff (\oc8051_top_1.oc8051_alu_src_sel1.op3_r [7], _00282_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [0], _03794_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [1], _03758_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_rd_sel_r [2], _03623_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [0], _03688_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [1], _03715_);
  dff (\oc8051_top_1.oc8051_decoder1.mem_act [2], _03625_);
  dff (\oc8051_top_1.oc8051_decoder1.state [0], _03718_);
  dff (\oc8051_top_1.oc8051_decoder1.state [1], _03627_);
  dff (\oc8051_top_1.oc8051_decoder1.op [0], _03831_);
  dff (\oc8051_top_1.oc8051_decoder1.op [1], _03833_);
  dff (\oc8051_top_1.oc8051_decoder1.op [2], _03835_);
  dff (\oc8051_top_1.oc8051_decoder1.op [3], _03837_);
  dff (\oc8051_top_1.oc8051_decoder1.op [4], _03839_);
  dff (\oc8051_top_1.oc8051_decoder1.op [5], _03840_);
  dff (\oc8051_top_1.oc8051_decoder1.op [6], _03851_);
  dff (\oc8051_top_1.oc8051_decoder1.op [7], _03630_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel3 , _03632_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [0], _03537_);
  dff (\oc8051_top_1.oc8051_decoder1.wr_sfr [1], _03634_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [0], _03545_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel2 [1], _03637_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [0], _03554_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [1], _03573_);
  dff (\oc8051_top_1.oc8051_decoder1.ram_wr_sel [2], _03646_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [0], _03710_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [1], _03743_);
  dff (\oc8051_top_1.oc8051_decoder1.src_sel1 [2], _03648_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [0], _03816_);
  dff (\oc8051_top_1.oc8051_decoder1.cy_sel [1], _03653_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [0], _03981_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [1], _03989_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [2], _03994_);
  dff (\oc8051_top_1.oc8051_decoder1.alu_op [3], _03656_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [0], _04011_);
  dff (\oc8051_top_1.oc8051_decoder1.psw_set [1], _03658_);
  dff (\oc8051_top_1.oc8051_decoder1.wr , _03660_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [0], _03765_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [1], _14515_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [2], _11806_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [3], _09234_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [4], _13300_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [5], _09050_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [6], _04105_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[0] [7], _14356_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [0], _01247_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [1], _04204_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [2], _13148_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [3], _04208_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [4], _02269_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [5], _07623_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [6], _04210_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[1] [7], _04025_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [0], _03036_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [1], _00471_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [2], _10727_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [3], _00509_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [4], _03325_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [5], _12642_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [6], _12351_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[2] [7], _02763_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [0], _03321_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [1], _03357_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [2], _13161_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [3], _01641_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [4], _00504_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [5], _03429_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [6], _01734_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[3] [7], _03986_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [0], _08409_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [1], _07824_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [2], _04095_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [3], _01560_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [4], _12259_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [5], _12465_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [6], _03425_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[4] [7], _02146_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [0], _10802_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [1], _11722_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [2], _03944_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [3], _12752_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [4], _03344_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [5], _03996_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [6], _04894_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[5] [7], _04587_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [0], _02645_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [1], _13387_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [2], _01183_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [3], _08690_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [4], _13150_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [5], _11956_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [6], _09410_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[6] [7], _12599_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [0], _01218_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [1], _12864_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [2], _10905_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [3], _13551_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [4], _07954_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [5], _06471_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [6], _02266_);
  dff (\oc8051_top_1.oc8051_indi_addr1.buff[7] [7], _01157_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [0], _08075_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [1], _07992_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [2], _07809_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [3], _07964_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rn_r [4], _03532_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [0], _05031_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [1], _05020_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [2], _04990_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [3], _04950_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [4], _04943_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [5], _00650_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [6], _04566_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [7], _02945_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [8], _02908_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [9], _02898_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [10], _00676_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [11], _02090_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [12], _01790_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [13], _02042_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [14], _01974_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log [15], _14073_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0], _11397_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1], _10809_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2], _00691_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3], _01394_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4], _01378_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5], _00572_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6], _00569_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7], _00475_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8], _00447_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9], _00688_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10], _00671_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11], _06473_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12], _14524_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13], _14522_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14], _14348_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15], _14207_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [0], _04313_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [1], _04533_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [2], _04362_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [3], _09949_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [4], _09624_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [5], _09742_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [6], _03700_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [7], _03692_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [8], _09962_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [9], _04057_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [10], _04052_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [11], _04050_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [12], _09958_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [13], _03147_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [14], _00724_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [15], _02566_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [16], _01803_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [17], _01708_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [18], _09972_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [19], _03460_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [20], _03502_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [21], _03495_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [22], _09967_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [23], _09619_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [24], _13974_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [25], _13783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [26], _13897_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [27], _13805_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [28], _09979_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [29], _00434_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [30], _00088_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_cur [31], _13965_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_addr_r , _14177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [0], _09996_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [1], _09610_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [2], _09730_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [3], _14055_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [4], _14295_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [5], _01145_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [6], _09849_);
  dff (\oc8051_top_1.oc8051_memory_interface1.ri_r [7], _03523_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [0], _09852_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [1], _09673_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [3], _00608_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [4], _09859_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [5], _10040_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm_r [6], _09590_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [1], _09863_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [2], _09668_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [3], _04000_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [4], _03812_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imm2_r [5], _03802_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r , _00272_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_wr_r2 , _03752_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [0], _10012_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [1], _04582_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [2], _04576_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [3], _04564_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [4], _04562_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [5], _10009_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [6], _09725_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [7], _04131_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [8], _04126_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [9], _04123_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [10], _04113_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [11], _04109_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [12], _10017_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [13], _04226_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [14], _04222_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc_buf [15], _03733_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [0], _03385_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [1], _03360_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [2], _03355_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [3], _10029_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [4], _03842_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [5], _03712_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [6], _03669_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [7], _03621_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [8], _10025_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [9], _09598_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [10], _02046_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [11], _01846_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [12], _02013_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [13], _01854_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [14], _01849_);
  dff (\oc8051_top_1.oc8051_memory_interface1.pc [15], _03720_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack , _13966_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_t , _03309_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_ack_buff , _03331_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [0], _00999_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [1], _00976_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [2], _10037_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [3], _01716_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [4], _01684_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [5], _01679_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [6], _01676_);
  dff (\oc8051_top_1.oc8051_memory_interface1.int_vec_buff [7], _03304_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [0], _09594_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [1], _00655_);
  dff (\oc8051_top_1.oc8051_memory_interface1.op_pos [2], _03295_);
  dff (\oc8051_top_1.oc8051_memory_interface1.reti , _03428_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [0], _10053_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [1], _00189_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [2], _00151_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [3], _00177_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [4], _00166_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [5], _00164_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [6], _00162_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdata [7], _03414_);
  dff (\oc8051_top_1.oc8051_memory_interface1.cdone , _03406_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst , _03398_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [0], _14197_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [1], _14182_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [2], _14180_);
  dff (\oc8051_top_1.oc8051_memory_interface1.out_of_rst_cycles [3], _00278_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [0], _13138_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [1], _13108_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [2], _13078_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [3], _13038_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [4], _10345_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [5], _09571_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [6], _12049_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [7], _12027_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [8], _11988_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [9], _10357_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [10], _12409_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [11], _12334_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [12], _12407_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [13], _12380_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [14], _12375_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [15], _12356_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [16], _12341_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [17], _10354_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [18], _09566_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [19], _09708_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [20], _11506_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [21], _11462_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [22], _10364_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [23], _11748_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [24], _11783_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [25], _11768_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [26], _11752_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [27], _10362_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [28], _09561_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [29], _10922_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [30], _01936_);
  dff (\oc8051_top_1.oc8051_memory_interface1.idat_old [31], _02583_);
  dff (\oc8051_top_1.oc8051_memory_interface1.dmem_wait , _03150_);
  dff (\oc8051_top_1.oc8051_memory_interface1.istb_t , _03144_);
  dff (\oc8051_top_1.oc8051_memory_interface1.imem_wait , _03132_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [0], _01786_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [1], _01752_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [2], _01697_);
  dff (\oc8051_top_1.oc8051_memory_interface1.iadr_t [3], _01650_);
  dff (\oc8051_top_1.oc8051_memory_interface1.rd_ind , _00287_);
  dff (\oc8051_top_1.oc8051_rom1.data_o [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  dff (\oc8051_top_1.oc8051_rom1.data_o [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  dff (\oc8051_top_1.oc8051_sfr1.pres_ow , _04220_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [0], _01806_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [1], _14012_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [2], _14009_);
  dff (\oc8051_top_1.oc8051_sfr1.prescaler [3], _04218_);
  dff (\oc8051_top_1.oc8051_sfr1.bit_out , _04214_);
  dff (\oc8051_top_1.oc8051_sfr1.wait_data , _04557_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [0], _01810_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [1], _13548_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [2], _13525_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [3], _13519_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [4], _01808_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [5], _01164_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [6], _13364_);
  dff (\oc8051_top_1.oc8051_sfr1.dat0 [7], _04366_);
  dff (\oc8051_top_1.oc8051_sfr1.wr_bit_r , _04364_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0], _06433_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1], _06429_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2], _03350_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3], _06536_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4], _06533_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5], _06517_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6], _03307_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7], _09630_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0], _03705_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1], _03804_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2], _03824_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3], _03807_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4], _03678_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5], _03708_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6], _03737_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7], _04377_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0], _07710_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1], _07705_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2], _07702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3], _07678_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4], _07658_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5], _07648_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6], _07645_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7], _13596_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0], _07449_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1], _07514_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2], _07498_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3], _07494_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4], _07469_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5], _07455_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6], _07452_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7], _13589_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0_buff , _02560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0], _00371_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1], _00368_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2], _00350_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3], _00345_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4], _00342_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5], _00339_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6], _00331_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7], _12487_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [0], _00326_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_dept [1], _12749_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_proc , _12769_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [0], _00299_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [1], _00295_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[0] [2], _03515_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [0], _00276_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [1], _00274_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.isrc[1] [2], _13339_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[0] [0], _00256_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_lev[1] [0], _00252_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 , _04592_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 , _04803_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 , _04826_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 , _01342_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0], _00211_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1], _00205_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2], _00191_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3], _04530_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0], _00172_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1], _00169_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2], _00153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3], _00143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4], _00149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5], _00147_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6], _00145_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7], _04535_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0], _00085_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1], _00082_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2], _00066_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3], _00064_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4], _00061_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5], _00056_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6], _00038_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7], _04538_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0], _02924_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1], _02893_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2], _03074_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3], _02926_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4], _03072_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5], _02890_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6], _03070_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7], _14416_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0], _02921_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1], _03080_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2], _02888_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3], _03076_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4], _03042_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5], _03040_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6], _02919_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7], _14346_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0], _03084_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1], _02883_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2], _03081_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3], _03046_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4], _03044_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5], _02886_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6], _03078_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7], _07328_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0], _02914_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1], _02879_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2], _03091_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3], _02916_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4], _03088_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5], _02881_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6], _03086_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7], _00501_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1], _03869_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2], _03860_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3], _03828_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4], _03784_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5], _03640_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6], _03547_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7], _02905_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.pop , _03196_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [0], _04806_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [1], _04808_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [2], _04810_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [3], _04812_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [4], _04814_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [5], _04822_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [6], _04824_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_sp1.sp [7], _03300_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0_buff , _02670_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1_buff , _02679_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0], _14392_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1], _14040_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2], _14032_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3], _14037_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4], _14026_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5], _14021_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6], _14023_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7], _02676_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0], _14047_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1], _13996_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2], _14000_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3], _13988_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4], _13991_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5], _13981_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6], _13978_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7], _02673_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_1 , _02666_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 , _02664_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0], _13925_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1], _13928_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2], _13834_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3], _13829_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4], _13831_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5], _13727_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6], _13721_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7], _02661_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0], _13714_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1], _13747_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2], _13739_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3], _13745_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4], _13742_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5], _13690_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6], _13693_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7], _02652_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf1_0 , _02658_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0], _13675_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1], _13637_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2], _13634_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3], _13661_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4], _13665_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5], _13844_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6], _13839_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7], _02649_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2_r , _10560_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tc2_event , _08140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.neg_trans , _08189_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex_r , _08204_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0], _03962_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1], _03958_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2], _03935_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3], _03911_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4], _03923_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5], _03917_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6], _03914_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7], _08719_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0], _03864_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1], _03787_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2], _03821_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3], _03800_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4], _03797_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5], _03791_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6], _03756_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7], _08068_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 , _08149_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0], _03685_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1], _03667_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2], _03663_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3], _03651_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4], _03644_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5], _04916_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6], _04910_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7], _08219_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0], _04966_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1], _04945_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2], _04937_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3], _04935_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4], _04926_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5], _04597_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6], _04595_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7], _11388_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2_set , _09435_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0], _04555_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1], _04551_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2], _04548_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3], _04545_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4], _03606_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5], _03599_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6], _03597_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7], _09333_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [0], _07970_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [1], _07876_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [2], _07849_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [3], _07863_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [4], _07860_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [5], _07855_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [6], _07852_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [7], _07909_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [8], _07934_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [9], _07983_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [10], _07973_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd_tmp [11], _13023_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf , _12089_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_re , _12083_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_re , _00247_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.receive , _12133_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_done , _12159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd_r , _12153_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [0], _02250_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rx_sam [1], _12143_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [0], _02236_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [1], _08701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [2], _03483_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.re_count [3], _12140_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0], _00550_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1], _00544_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2], _14544_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3], _14365_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4], _13011_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5], _12870_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6], _11894_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7], _00239_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.shift_tr , _12010_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod_clk_tr , _12007_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.trans , _12000_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tx_done , _11992_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [0], _14257_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [1], _10468_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [2], _06950_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tr_count [3], _11985_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [0], _04986_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [1], _04984_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [2], _04960_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [3], _04590_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [4], _04580_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [5], _04573_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [6], _04383_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [7], _04379_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [8], _04369_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [9], _04206_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_txd [10], _00280_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0], _03118_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1], _03061_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2], _03049_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3], _02632_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4], _02313_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5], _02191_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6], _02204_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7], _12036_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0], _01702_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1], _01700_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2], _00629_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3], _01159_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4], _00701_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5], _00695_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6], _13754_);
  dff (\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7], _12053_);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_for_ajmp [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [0], \oc8051_top_1.oc8051_memory_interface1.pc_buf [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.pc_out [1], \oc8051_top_1.oc8051_memory_interface1.pc_buf [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [1], \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [2], \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [5], \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op3_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [0], \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [1], \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [4], \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [5], \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.op2_buff [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.oc8051_memory_interface1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.int_v [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [0], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [6], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm2_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op3_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [2], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.imm_r [7], \oc8051_top_1.oc8051_alu_src_sel1.op2_r [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [0], ABINPUT[1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [1], ABINPUT[2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [2], ABINPUT[3]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [3], ABINPUT[4]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [4], ABINPUT[5]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [5], ABINPUT[6]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [6], ABINPUT[7]);
  buf(\oc8051_top_1.oc8051_memory_interface1.in_ram [7], ABINPUT[8]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.oc8051_memory_interface1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.oc8051_memory_interface1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.oc8051_memory_interface1.bit_in , ABINPUT[0]);
  buf(\oc8051_top_1.oc8051_memory_interface1.rst , rst);
  buf(\oc8051_top_1.oc8051_memory_interface1.clk , clk);
  buf(\oc8051_top_1.oc8051_indi_addr1.wr_bit_r , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_indi_addr1.rst , rst);
  buf(\oc8051_top_1.oc8051_indi_addr1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.oc8051_rom1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_rom1.clk , clk);
  buf(\oc8051_top_1.oc8051_rom1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.cprl2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.ct2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tr2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exen2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.exf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tf2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_tc21.clk , clk);
  buf(\oc8051_top_1.oc8051_decoder1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.oc8051_decoder1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.oc8051_decoder1.rst , rst);
  buf(\oc8051_top_1.oc8051_decoder1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.smod , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ri , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tb8 , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.ren , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pres_ow , \oc8051_top_1.oc8051_sfr1.pres_ow );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_uatr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.ip [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ip [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.ie [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [0]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [1]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [2]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [3]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [4]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [5]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [6]);
  buf(\oc8051_top_1.oc8051_sfr1.ie [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ie [7]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [0]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [1]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [2]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [3]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [4]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [5]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [6]);
  buf(\oc8051_top_1.oc8051_sfr1.sbuf [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.sbuf_rxd [7]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.pcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.pcon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [0], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [0]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [1], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [1]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [2], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [2]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [3], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [3]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [4], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [4]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [5], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [5]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [6], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [6]);
  buf(\oc8051_top_1.oc8051_sfr1.scon [7], \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.scon [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl1 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl1 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.th0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl0 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tl0 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tmod [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tmod [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2h [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2h [7]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [0]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [1]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [2]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [3]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [5]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [6]);
  buf(\oc8051_top_1.oc8051_sfr1.rcap2l [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.rcap2l [7]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.th2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.th2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [0]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [1]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [4]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [6]);
  buf(\oc8051_top_1.oc8051_sfr1.tl2 [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.tl2 [7]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [0], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [0]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [1], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [1]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [2], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [2]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [3], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [3]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [4], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [5], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [6], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [6]);
  buf(\oc8051_top_1.oc8051_sfr1.t2con [7], \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [7]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [0], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [1], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [2], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [3], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [4], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [5], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [6], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.b_reg [7], \oc8051_top_1.oc8051_sfr1.oc8051_b_register.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.brate2 , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.brate2 );
  buf(\oc8051_top_1.oc8051_sfr1.tclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [4]);
  buf(\oc8051_top_1.oc8051_sfr1.rclk , \oc8051_top_1.oc8051_sfr1.oc8051_tc21.t2con [5]);
  buf(\oc8051_top_1.oc8051_sfr1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.t2ex , t2ex_i);
  buf(\oc8051_top_1.oc8051_sfr1.t2 , t2_i);
  buf(\oc8051_top_1.oc8051_sfr1.t1 , t1_i);
  buf(\oc8051_top_1.oc8051_sfr1.t0 , t0_i);
  buf(\oc8051_top_1.oc8051_sfr1.rxd , rxd_i);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_sfr1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_sfr1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.oc8051_sfr1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.oc8051_sfr1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [8], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [9], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [10], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [11], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [12], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [13], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [14], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.dptr [15], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [0], \oc8051_top_1.oc8051_memory_interface1.imm_r [0]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [1], \oc8051_top_1.oc8051_memory_interface1.imm_r [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [3], \oc8051_top_1.oc8051_memory_interface1.imm_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [4], \oc8051_top_1.oc8051_memory_interface1.imm_r [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [5], \oc8051_top_1.oc8051_memory_interface1.imm_r [5]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op2_r [6], \oc8051_top_1.oc8051_memory_interface1.imm_r [6]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [1], \oc8051_top_1.oc8051_memory_interface1.imm2_r [1]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [2], \oc8051_top_1.oc8051_memory_interface1.imm2_r [2]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [3], \oc8051_top_1.oc8051_memory_interface1.imm2_r [3]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [4], \oc8051_top_1.oc8051_memory_interface1.imm2_r [4]);
  buf(\oc8051_top_1.oc8051_alu_src_sel1.op3_r [5], \oc8051_top_1.oc8051_memory_interface1.imm2_r [5]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.oc8051_cy_select1.cy_in , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_symbolic_cxrom1.clk , clk);
  buf(\oc8051_symbolic_cxrom1.rst , rst);
  buf(\oc8051_symbolic_cxrom1.word_in [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.word_in [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.word_in [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.word_in [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.word_in [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.word_in [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.word_in [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.word_in [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.word_in [8], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.word_in [9], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.word_in [10], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.word_in [11], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.word_in [12], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.word_in [13], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.word_in [14], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.word_in [15], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.word_in [16], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.word_in [17], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.word_in [18], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.word_in [19], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.word_in [20], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.word_in [21], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.word_in [22], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.word_in [23], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.word_in [24], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.word_in [25], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.word_in [26], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.word_in [27], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.word_in [28], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.word_in [29], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.word_in [30], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.word_in [31], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.pc1 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc1 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc1 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc1 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc1 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_symbolic_cxrom1.pc1 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_symbolic_cxrom1.pc1 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_symbolic_cxrom1.pc1 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_symbolic_cxrom1.pc1 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_symbolic_cxrom1.pc1 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_symbolic_cxrom1.pc1 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_symbolic_cxrom1.pc1 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_symbolic_cxrom1.pc1 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_symbolic_cxrom1.pc1 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_symbolic_cxrom1.pc1 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_symbolic_cxrom1.pc1 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_symbolic_cxrom1.pc2 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc2 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc2 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc2 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc2 [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_symbolic_cxrom1.pc2 [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_symbolic_cxrom1.pc2 [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_symbolic_cxrom1.pc2 [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_symbolic_cxrom1.pc2 [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_symbolic_cxrom1.pc2 [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_symbolic_cxrom1.pc2 [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_symbolic_cxrom1.pc2 [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_symbolic_cxrom1.pc2 [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_symbolic_cxrom1.pc2 [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_symbolic_cxrom1.pc2 [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_symbolic_cxrom1.pc2 [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [0], word_in[0]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [1], word_in[1]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [2], word_in[2]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [3], word_in[3]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [4], word_in[4]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [5], word_in[5]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [6], word_in[6]);
  buf(\oc8051_symbolic_cxrom1.bytein0 [7], word_in[7]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [0], word_in[8]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [1], word_in[9]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [2], word_in[10]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [3], word_in[11]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [4], word_in[12]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [5], word_in[13]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [6], word_in[14]);
  buf(\oc8051_symbolic_cxrom1.bytein1 [7], word_in[15]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [0], word_in[16]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [1], word_in[17]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [2], word_in[18]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [3], word_in[19]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [4], word_in[20]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [5], word_in[21]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [6], word_in[22]);
  buf(\oc8051_symbolic_cxrom1.bytein2 [7], word_in[23]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [0], word_in[24]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [1], word_in[25]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [2], word_in[26]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [3], word_in[27]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [4], word_in[28]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [5], word_in[29]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [6], word_in[30]);
  buf(\oc8051_symbolic_cxrom1.bytein3 [7], word_in[31]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_symbolic_cxrom1.byteout0 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_symbolic_cxrom1.byteout1 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_symbolic_cxrom1.byteout2 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [0], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [1], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [2], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [3], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [4], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [5], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [6], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_symbolic_cxrom1.byteout3 [7], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_symbolic_cxrom1.pc10 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc10 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_symbolic_cxrom1.pc10 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_symbolic_cxrom1.pc10 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_symbolic_cxrom1.pc12 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_symbolic_cxrom1.pc12 [1], pc1_plus_2[1]);
  buf(\oc8051_symbolic_cxrom1.pc12 [2], pc1_plus_2[2]);
  buf(\oc8051_symbolic_cxrom1.pc12 [3], pc1_plus_2[3]);
  buf(\oc8051_symbolic_cxrom1.pc20 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_symbolic_cxrom1.pc20 [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_symbolic_cxrom1.pc20 [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_symbolic_cxrom1.pc20 [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_symbolic_cxrom1.pc22 [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.oc8051_comp1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_comp1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.oc8051_comp1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.oc8051_comp1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.oc8051_comp1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.oc8051_comp1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.oc8051_comp1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.oc8051_comp1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.oc8051_comp1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div_out [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_alu1.clk , clk);
  buf(\oc8051_top_1.oc8051_alu1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.divsrc2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div1 , \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.div0 , \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [0], \oc8051_top_1.oc8051_alu1.divsrc2 [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [1], \oc8051_top_1.oc8051_alu1.divsrc2 [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [2], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [0]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [3], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [1]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [4], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [2]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [5], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [3]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [6], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [4]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.des2 [7], \oc8051_top_1.oc8051_alu1.oc8051_div1.tmp_div [5]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_div1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [0], p3_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [1], p3_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [2], p3_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [3], p3_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [4], p3_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [5], p3_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [6], p3_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_in [7], p3_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [0], p2_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [1], p2_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [2], p2_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [3], p2_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [4], p2_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [5], p2_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [6], p2_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_in [7], p2_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [0], p1_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [1], p1_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [2], p1_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [3], p1_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [4], p1_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [5], p1_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [6], p1_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_in [7], p1_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [0], p0_in[0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [1], p0_in[1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [2], p0_in[2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [3], p0_in[3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [4], p0_in[4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [5], p0_in[5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [6], p0_in[6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_in [7], p0_in[7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_ports1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_acc1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf1_buff , \oc8051_top_1.oc8051_sfr1.oc8051_uatr1.t1_ow_buf );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [4], \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.int_src [5], \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ip_l1 [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.ip [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_ie1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_tf1 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr1 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tr0 , \oc8051_top_1.oc8051_sfr1.oc8051_int1.tcon_s [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.uart_int , \oc8051_top_1.oc8051_sfr1.uart_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.t2_int , \oc8051_top_1.oc8051_sfr1.tc2_int );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_int1.tf0 , \oc8051_top_1.oc8051_sfr1.oc8051_tc1.tf0 );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [0], \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [1], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [2], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [2]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [3], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [3]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [4], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [4]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [5], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [5]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [6], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.data_out [7], \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.p , \oc8051_top_1.oc8051_sfr1.psw [0]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_psw1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_dptr1.clk , clk);
  buf(\oc8051_top_1.ABINPUT [0], ABINPUT[0]);
  buf(\oc8051_top_1.ABINPUT [1], ABINPUT[1]);
  buf(\oc8051_top_1.ABINPUT [2], ABINPUT[2]);
  buf(\oc8051_top_1.ABINPUT [3], ABINPUT[3]);
  buf(\oc8051_top_1.ABINPUT [4], ABINPUT[4]);
  buf(\oc8051_top_1.ABINPUT [5], ABINPUT[5]);
  buf(\oc8051_top_1.ABINPUT [6], ABINPUT[6]);
  buf(\oc8051_top_1.ABINPUT [7], ABINPUT[7]);
  buf(\oc8051_top_1.ABINPUT [8], ABINPUT[8]);
  buf(\oc8051_top_1.wb_rst_i , rst);
  buf(\oc8051_top_1.wb_clk_i , clk);
  buf(\oc8051_top_1.wait_data , \oc8051_top_1.oc8051_sfr1.wait_data );
  buf(\oc8051_top_1.bit_data , ABINPUT[0]);
  buf(\oc8051_top_1.rd_ind , \oc8051_top_1.oc8051_memory_interface1.rd_ind );
  buf(\oc8051_top_1.cy , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [7]);
  buf(\oc8051_top_1.srcAc , \oc8051_top_1.oc8051_sfr1.oc8051_psw1.data [6]);
  buf(\oc8051_top_1.irom_out_of_rst , \oc8051_top_1.oc8051_memory_interface1.out_of_rst );
  buf(\oc8051_top_1.psw_set [0], \oc8051_top_1.oc8051_decoder1.psw_set [0]);
  buf(\oc8051_top_1.psw_set [1], \oc8051_top_1.oc8051_decoder1.psw_set [1]);
  buf(\oc8051_top_1.mem_act [0], \oc8051_top_1.oc8051_decoder1.mem_act [0]);
  buf(\oc8051_top_1.mem_act [1], \oc8051_top_1.oc8051_decoder1.mem_act [1]);
  buf(\oc8051_top_1.mem_act [2], \oc8051_top_1.oc8051_decoder1.mem_act [2]);
  buf(\oc8051_top_1.int_src [0], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [0]);
  buf(\oc8051_top_1.int_src [1], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [1]);
  buf(\oc8051_top_1.int_src [2], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [2]);
  buf(\oc8051_top_1.int_src [3], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [3]);
  buf(\oc8051_top_1.int_src [4], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [4]);
  buf(\oc8051_top_1.int_src [5], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [5]);
  buf(\oc8051_top_1.int_src [6], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [6]);
  buf(\oc8051_top_1.int_src [7], \oc8051_top_1.oc8051_sfr1.oc8051_int1.int_vec [7]);
  buf(\oc8051_top_1.int_ack , \oc8051_top_1.oc8051_memory_interface1.int_ack );
  buf(\oc8051_top_1.reti , \oc8051_top_1.oc8051_memory_interface1.reti );
  buf(\oc8051_top_1.cy_sel [0], \oc8051_top_1.oc8051_decoder1.cy_sel [0]);
  buf(\oc8051_top_1.cy_sel [1], \oc8051_top_1.oc8051_decoder1.cy_sel [1]);
  buf(\oc8051_top_1.sfr_bit , \oc8051_top_1.oc8051_sfr1.bit_out );
  buf(\oc8051_top_1.sfr_out [0], \oc8051_top_1.oc8051_sfr1.dat0 [0]);
  buf(\oc8051_top_1.sfr_out [1], \oc8051_top_1.oc8051_sfr1.dat0 [1]);
  buf(\oc8051_top_1.sfr_out [2], \oc8051_top_1.oc8051_sfr1.dat0 [2]);
  buf(\oc8051_top_1.sfr_out [3], \oc8051_top_1.oc8051_sfr1.dat0 [3]);
  buf(\oc8051_top_1.sfr_out [4], \oc8051_top_1.oc8051_sfr1.dat0 [4]);
  buf(\oc8051_top_1.sfr_out [5], \oc8051_top_1.oc8051_sfr1.dat0 [5]);
  buf(\oc8051_top_1.sfr_out [6], \oc8051_top_1.oc8051_sfr1.dat0 [6]);
  buf(\oc8051_top_1.sfr_out [7], \oc8051_top_1.oc8051_sfr1.dat0 [7]);
  buf(\oc8051_top_1.ram_data [0], ABINPUT[1]);
  buf(\oc8051_top_1.ram_data [1], ABINPUT[2]);
  buf(\oc8051_top_1.ram_data [2], ABINPUT[3]);
  buf(\oc8051_top_1.ram_data [3], ABINPUT[4]);
  buf(\oc8051_top_1.ram_data [4], ABINPUT[5]);
  buf(\oc8051_top_1.ram_data [5], ABINPUT[6]);
  buf(\oc8051_top_1.ram_data [6], ABINPUT[7]);
  buf(\oc8051_top_1.ram_data [7], ABINPUT[8]);
  buf(\oc8051_top_1.src_sel1 [0], \oc8051_top_1.oc8051_decoder1.src_sel1 [0]);
  buf(\oc8051_top_1.src_sel1 [1], \oc8051_top_1.oc8051_decoder1.src_sel1 [1]);
  buf(\oc8051_top_1.src_sel1 [2], \oc8051_top_1.oc8051_decoder1.src_sel1 [2]);
  buf(\oc8051_top_1.src_sel2 [0], \oc8051_top_1.oc8051_decoder1.src_sel2 [0]);
  buf(\oc8051_top_1.src_sel2 [1], \oc8051_top_1.oc8051_decoder1.src_sel2 [1]);
  buf(\oc8051_top_1.src_sel3 , \oc8051_top_1.oc8051_decoder1.src_sel3 );
  buf(\oc8051_top_1.pc [0], \oc8051_top_1.oc8051_memory_interface1.pc [0]);
  buf(\oc8051_top_1.pc [1], \oc8051_top_1.oc8051_memory_interface1.pc [1]);
  buf(\oc8051_top_1.pc [2], \oc8051_top_1.oc8051_memory_interface1.pc [2]);
  buf(\oc8051_top_1.pc [3], \oc8051_top_1.oc8051_memory_interface1.pc [3]);
  buf(\oc8051_top_1.pc [4], \oc8051_top_1.oc8051_memory_interface1.pc [4]);
  buf(\oc8051_top_1.pc [5], \oc8051_top_1.oc8051_memory_interface1.pc [5]);
  buf(\oc8051_top_1.pc [6], \oc8051_top_1.oc8051_memory_interface1.pc [6]);
  buf(\oc8051_top_1.pc [7], \oc8051_top_1.oc8051_memory_interface1.pc [7]);
  buf(\oc8051_top_1.pc [8], \oc8051_top_1.oc8051_memory_interface1.pc [8]);
  buf(\oc8051_top_1.pc [9], \oc8051_top_1.oc8051_memory_interface1.pc [9]);
  buf(\oc8051_top_1.pc [10], \oc8051_top_1.oc8051_memory_interface1.pc [10]);
  buf(\oc8051_top_1.pc [11], \oc8051_top_1.oc8051_memory_interface1.pc [11]);
  buf(\oc8051_top_1.pc [12], \oc8051_top_1.oc8051_memory_interface1.pc [12]);
  buf(\oc8051_top_1.pc [13], \oc8051_top_1.oc8051_memory_interface1.pc [13]);
  buf(\oc8051_top_1.pc [14], \oc8051_top_1.oc8051_memory_interface1.pc [14]);
  buf(\oc8051_top_1.pc [15], \oc8051_top_1.oc8051_memory_interface1.pc [15]);
  buf(\oc8051_top_1.idat_onchip [0], \oc8051_top_1.oc8051_rom1.data_o [0]);
  buf(\oc8051_top_1.idat_onchip [1], \oc8051_top_1.oc8051_rom1.data_o [1]);
  buf(\oc8051_top_1.idat_onchip [2], \oc8051_top_1.oc8051_rom1.data_o [2]);
  buf(\oc8051_top_1.idat_onchip [3], \oc8051_top_1.oc8051_rom1.data_o [3]);
  buf(\oc8051_top_1.idat_onchip [4], \oc8051_top_1.oc8051_rom1.data_o [4]);
  buf(\oc8051_top_1.idat_onchip [5], \oc8051_top_1.oc8051_rom1.data_o [5]);
  buf(\oc8051_top_1.idat_onchip [6], \oc8051_top_1.oc8051_rom1.data_o [6]);
  buf(\oc8051_top_1.idat_onchip [7], \oc8051_top_1.oc8051_rom1.data_o [7]);
  buf(\oc8051_top_1.idat_onchip [8], \oc8051_top_1.oc8051_rom1.data_o [8]);
  buf(\oc8051_top_1.idat_onchip [9], \oc8051_top_1.oc8051_rom1.data_o [9]);
  buf(\oc8051_top_1.idat_onchip [10], \oc8051_top_1.oc8051_rom1.data_o [10]);
  buf(\oc8051_top_1.idat_onchip [11], \oc8051_top_1.oc8051_rom1.data_o [11]);
  buf(\oc8051_top_1.idat_onchip [12], \oc8051_top_1.oc8051_rom1.data_o [12]);
  buf(\oc8051_top_1.idat_onchip [13], \oc8051_top_1.oc8051_rom1.data_o [13]);
  buf(\oc8051_top_1.idat_onchip [14], \oc8051_top_1.oc8051_rom1.data_o [14]);
  buf(\oc8051_top_1.idat_onchip [15], \oc8051_top_1.oc8051_rom1.data_o [15]);
  buf(\oc8051_top_1.idat_onchip [16], \oc8051_top_1.oc8051_rom1.data_o [16]);
  buf(\oc8051_top_1.idat_onchip [17], \oc8051_top_1.oc8051_rom1.data_o [17]);
  buf(\oc8051_top_1.idat_onchip [18], \oc8051_top_1.oc8051_rom1.data_o [18]);
  buf(\oc8051_top_1.idat_onchip [19], \oc8051_top_1.oc8051_rom1.data_o [19]);
  buf(\oc8051_top_1.idat_onchip [20], \oc8051_top_1.oc8051_rom1.data_o [20]);
  buf(\oc8051_top_1.idat_onchip [21], \oc8051_top_1.oc8051_rom1.data_o [21]);
  buf(\oc8051_top_1.idat_onchip [22], \oc8051_top_1.oc8051_rom1.data_o [22]);
  buf(\oc8051_top_1.idat_onchip [23], \oc8051_top_1.oc8051_rom1.data_o [23]);
  buf(\oc8051_top_1.idat_onchip [24], \oc8051_top_1.oc8051_rom1.data_o [24]);
  buf(\oc8051_top_1.idat_onchip [25], \oc8051_top_1.oc8051_rom1.data_o [25]);
  buf(\oc8051_top_1.idat_onchip [26], \oc8051_top_1.oc8051_rom1.data_o [26]);
  buf(\oc8051_top_1.idat_onchip [27], \oc8051_top_1.oc8051_rom1.data_o [27]);
  buf(\oc8051_top_1.idat_onchip [28], \oc8051_top_1.oc8051_rom1.data_o [28]);
  buf(\oc8051_top_1.idat_onchip [29], \oc8051_top_1.oc8051_rom1.data_o [29]);
  buf(\oc8051_top_1.idat_onchip [30], \oc8051_top_1.oc8051_rom1.data_o [30]);
  buf(\oc8051_top_1.idat_onchip [31], \oc8051_top_1.oc8051_rom1.data_o [31]);
  buf(\oc8051_top_1.acc [0], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [0]);
  buf(\oc8051_top_1.acc [1], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [1]);
  buf(\oc8051_top_1.acc [2], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [2]);
  buf(\oc8051_top_1.acc [3], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [3]);
  buf(\oc8051_top_1.acc [4], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [4]);
  buf(\oc8051_top_1.acc [5], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [5]);
  buf(\oc8051_top_1.acc [6], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [6]);
  buf(\oc8051_top_1.acc [7], \oc8051_top_1.oc8051_sfr1.oc8051_acc1.data_out [7]);
  buf(\oc8051_top_1.pc_log [0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(\oc8051_top_1.pc_log [1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(\oc8051_top_1.pc_log [2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(\oc8051_top_1.pc_log [3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(\oc8051_top_1.pc_log [4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(\oc8051_top_1.pc_log [5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(\oc8051_top_1.pc_log [6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(\oc8051_top_1.pc_log [7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(\oc8051_top_1.pc_log [8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(\oc8051_top_1.pc_log [9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(\oc8051_top_1.pc_log [10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(\oc8051_top_1.pc_log [11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(\oc8051_top_1.pc_log [12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(\oc8051_top_1.pc_log [13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(\oc8051_top_1.pc_log [14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(\oc8051_top_1.pc_log [15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(\oc8051_top_1.pc_log_prev [0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(\oc8051_top_1.pc_log_prev [1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(\oc8051_top_1.pc_log_prev [2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(\oc8051_top_1.pc_log_prev [3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(\oc8051_top_1.pc_log_prev [4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(\oc8051_top_1.pc_log_prev [5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(\oc8051_top_1.pc_log_prev [6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(\oc8051_top_1.pc_log_prev [7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(\oc8051_top_1.pc_log_prev [8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(\oc8051_top_1.pc_log_prev [9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(\oc8051_top_1.pc_log_prev [10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(\oc8051_top_1.pc_log_prev [11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(\oc8051_top_1.pc_log_prev [12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(\oc8051_top_1.pc_log_prev [13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(\oc8051_top_1.pc_log_prev [14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(\oc8051_top_1.pc_log_prev [15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(\oc8051_top_1.dptr_lo [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [0]);
  buf(\oc8051_top_1.dptr_lo [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [1]);
  buf(\oc8051_top_1.dptr_lo [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [2]);
  buf(\oc8051_top_1.dptr_lo [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [3]);
  buf(\oc8051_top_1.dptr_lo [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [4]);
  buf(\oc8051_top_1.dptr_lo [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [5]);
  buf(\oc8051_top_1.dptr_lo [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [6]);
  buf(\oc8051_top_1.dptr_lo [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_lo [7]);
  buf(\oc8051_top_1.dptr_hi [0], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [0]);
  buf(\oc8051_top_1.dptr_hi [1], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [1]);
  buf(\oc8051_top_1.dptr_hi [2], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [2]);
  buf(\oc8051_top_1.dptr_hi [3], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [3]);
  buf(\oc8051_top_1.dptr_hi [4], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [4]);
  buf(\oc8051_top_1.dptr_hi [5], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [5]);
  buf(\oc8051_top_1.dptr_hi [6], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [6]);
  buf(\oc8051_top_1.dptr_hi [7], \oc8051_top_1.oc8051_sfr1.oc8051_dptr1.data_hi [7]);
  buf(\oc8051_top_1.t2ex_i , t2ex_i);
  buf(\oc8051_top_1.t2_i , t2_i);
  buf(\oc8051_top_1.t1_i , t1_i);
  buf(\oc8051_top_1.t0_i , t0_i);
  buf(\oc8051_top_1.rxd_i , rxd_i);
  buf(\oc8051_top_1.p3_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(\oc8051_top_1.p3_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(\oc8051_top_1.p3_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(\oc8051_top_1.p3_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(\oc8051_top_1.p3_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(\oc8051_top_1.p3_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(\oc8051_top_1.p3_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(\oc8051_top_1.p3_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(\oc8051_top_1.p3_i [0], p3_in[0]);
  buf(\oc8051_top_1.p3_i [1], p3_in[1]);
  buf(\oc8051_top_1.p3_i [2], p3_in[2]);
  buf(\oc8051_top_1.p3_i [3], p3_in[3]);
  buf(\oc8051_top_1.p3_i [4], p3_in[4]);
  buf(\oc8051_top_1.p3_i [5], p3_in[5]);
  buf(\oc8051_top_1.p3_i [6], p3_in[6]);
  buf(\oc8051_top_1.p3_i [7], p3_in[7]);
  buf(\oc8051_top_1.p2_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(\oc8051_top_1.p2_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(\oc8051_top_1.p2_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(\oc8051_top_1.p2_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(\oc8051_top_1.p2_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(\oc8051_top_1.p2_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(\oc8051_top_1.p2_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(\oc8051_top_1.p2_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(\oc8051_top_1.p2_i [0], p2_in[0]);
  buf(\oc8051_top_1.p2_i [1], p2_in[1]);
  buf(\oc8051_top_1.p2_i [2], p2_in[2]);
  buf(\oc8051_top_1.p2_i [3], p2_in[3]);
  buf(\oc8051_top_1.p2_i [4], p2_in[4]);
  buf(\oc8051_top_1.p2_i [5], p2_in[5]);
  buf(\oc8051_top_1.p2_i [6], p2_in[6]);
  buf(\oc8051_top_1.p2_i [7], p2_in[7]);
  buf(\oc8051_top_1.p1_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(\oc8051_top_1.p1_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(\oc8051_top_1.p1_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(\oc8051_top_1.p1_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(\oc8051_top_1.p1_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(\oc8051_top_1.p1_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(\oc8051_top_1.p1_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(\oc8051_top_1.p1_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(\oc8051_top_1.p1_i [0], p1_in[0]);
  buf(\oc8051_top_1.p1_i [1], p1_in[1]);
  buf(\oc8051_top_1.p1_i [2], p1_in[2]);
  buf(\oc8051_top_1.p1_i [3], p1_in[3]);
  buf(\oc8051_top_1.p1_i [4], p1_in[4]);
  buf(\oc8051_top_1.p1_i [5], p1_in[5]);
  buf(\oc8051_top_1.p1_i [6], p1_in[6]);
  buf(\oc8051_top_1.p1_i [7], p1_in[7]);
  buf(\oc8051_top_1.p0_o [0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(\oc8051_top_1.p0_o [1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(\oc8051_top_1.p0_o [2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(\oc8051_top_1.p0_o [3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(\oc8051_top_1.p0_o [4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(\oc8051_top_1.p0_o [5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(\oc8051_top_1.p0_o [6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(\oc8051_top_1.p0_o [7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
  buf(\oc8051_top_1.p0_i [0], p0_in[0]);
  buf(\oc8051_top_1.p0_i [1], p0_in[1]);
  buf(\oc8051_top_1.p0_i [2], p0_in[2]);
  buf(\oc8051_top_1.p0_i [3], p0_in[3]);
  buf(\oc8051_top_1.p0_i [4], p0_in[4]);
  buf(\oc8051_top_1.p0_i [5], p0_in[5]);
  buf(\oc8051_top_1.p0_i [6], p0_in[6]);
  buf(\oc8051_top_1.p0_i [7], p0_in[7]);
  buf(\oc8051_top_1.cxrom_data_out [0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(\oc8051_top_1.cxrom_data_out [1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(\oc8051_top_1.cxrom_data_out [2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(\oc8051_top_1.cxrom_data_out [3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(\oc8051_top_1.cxrom_data_out [4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(\oc8051_top_1.cxrom_data_out [5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(\oc8051_top_1.cxrom_data_out [6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(\oc8051_top_1.cxrom_data_out [7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(\oc8051_top_1.cxrom_data_out [8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(\oc8051_top_1.cxrom_data_out [9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(\oc8051_top_1.cxrom_data_out [10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(\oc8051_top_1.cxrom_data_out [11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(\oc8051_top_1.cxrom_data_out [12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(\oc8051_top_1.cxrom_data_out [13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(\oc8051_top_1.cxrom_data_out [14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(\oc8051_top_1.cxrom_data_out [15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(\oc8051_top_1.cxrom_data_out [16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(\oc8051_top_1.cxrom_data_out [17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(\oc8051_top_1.cxrom_data_out [18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(\oc8051_top_1.cxrom_data_out [19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(\oc8051_top_1.cxrom_data_out [20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(\oc8051_top_1.cxrom_data_out [21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(\oc8051_top_1.cxrom_data_out [22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(\oc8051_top_1.cxrom_data_out [23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(\oc8051_top_1.cxrom_data_out [24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(\oc8051_top_1.cxrom_data_out [25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(\oc8051_top_1.cxrom_data_out [26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(\oc8051_top_1.cxrom_data_out [27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(\oc8051_top_1.cxrom_data_out [28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(\oc8051_top_1.cxrom_data_out [29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(\oc8051_top_1.cxrom_data_out [30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(\oc8051_top_1.cxrom_data_out [31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.rst , rst);
  buf(\oc8051_top_1.oc8051_alu1.oc8051_mul1.clk , clk);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_sp1.clk , clk);
  buf(pc1_plus_2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[0], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [0]);
  buf(pc1[1], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [1]);
  buf(pc1[2], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [2]);
  buf(pc1[3], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [3]);
  buf(pc1[4], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [4]);
  buf(pc1[5], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [5]);
  buf(pc1[6], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [6]);
  buf(pc1[7], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [7]);
  buf(pc1[8], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [8]);
  buf(pc1[9], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [9]);
  buf(pc1[10], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [10]);
  buf(pc1[11], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [11]);
  buf(pc1[12], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [12]);
  buf(pc1[13], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [13]);
  buf(pc1[14], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [14]);
  buf(pc1[15], \oc8051_top_1.oc8051_memory_interface1.pc_log_prev [15]);
  buf(pc2[0], \oc8051_top_1.oc8051_memory_interface1.pc_log [0]);
  buf(pc2[1], \oc8051_top_1.oc8051_memory_interface1.pc_log [1]);
  buf(pc2[2], \oc8051_top_1.oc8051_memory_interface1.pc_log [2]);
  buf(pc2[3], \oc8051_top_1.oc8051_memory_interface1.pc_log [3]);
  buf(pc2[4], \oc8051_top_1.oc8051_memory_interface1.pc_log [4]);
  buf(pc2[5], \oc8051_top_1.oc8051_memory_interface1.pc_log [5]);
  buf(pc2[6], \oc8051_top_1.oc8051_memory_interface1.pc_log [6]);
  buf(pc2[7], \oc8051_top_1.oc8051_memory_interface1.pc_log [7]);
  buf(pc2[8], \oc8051_top_1.oc8051_memory_interface1.pc_log [8]);
  buf(pc2[9], \oc8051_top_1.oc8051_memory_interface1.pc_log [9]);
  buf(pc2[10], \oc8051_top_1.oc8051_memory_interface1.pc_log [10]);
  buf(pc2[11], \oc8051_top_1.oc8051_memory_interface1.pc_log [11]);
  buf(pc2[12], \oc8051_top_1.oc8051_memory_interface1.pc_log [12]);
  buf(pc2[13], \oc8051_top_1.oc8051_memory_interface1.pc_log [13]);
  buf(pc2[14], \oc8051_top_1.oc8051_memory_interface1.pc_log [14]);
  buf(pc2[15], \oc8051_top_1.oc8051_memory_interface1.pc_log [15]);
  buf(cxrom_data_out[0], \oc8051_symbolic_cxrom1.cxrom_data_out [0]);
  buf(cxrom_data_out[1], \oc8051_symbolic_cxrom1.cxrom_data_out [1]);
  buf(cxrom_data_out[2], \oc8051_symbolic_cxrom1.cxrom_data_out [2]);
  buf(cxrom_data_out[3], \oc8051_symbolic_cxrom1.cxrom_data_out [3]);
  buf(cxrom_data_out[4], \oc8051_symbolic_cxrom1.cxrom_data_out [4]);
  buf(cxrom_data_out[5], \oc8051_symbolic_cxrom1.cxrom_data_out [5]);
  buf(cxrom_data_out[6], \oc8051_symbolic_cxrom1.cxrom_data_out [6]);
  buf(cxrom_data_out[7], \oc8051_symbolic_cxrom1.cxrom_data_out [7]);
  buf(cxrom_data_out[8], \oc8051_symbolic_cxrom1.cxrom_data_out [8]);
  buf(cxrom_data_out[9], \oc8051_symbolic_cxrom1.cxrom_data_out [9]);
  buf(cxrom_data_out[10], \oc8051_symbolic_cxrom1.cxrom_data_out [10]);
  buf(cxrom_data_out[11], \oc8051_symbolic_cxrom1.cxrom_data_out [11]);
  buf(cxrom_data_out[12], \oc8051_symbolic_cxrom1.cxrom_data_out [12]);
  buf(cxrom_data_out[13], \oc8051_symbolic_cxrom1.cxrom_data_out [13]);
  buf(cxrom_data_out[14], \oc8051_symbolic_cxrom1.cxrom_data_out [14]);
  buf(cxrom_data_out[15], \oc8051_symbolic_cxrom1.cxrom_data_out [15]);
  buf(cxrom_data_out[16], \oc8051_symbolic_cxrom1.cxrom_data_out [16]);
  buf(cxrom_data_out[17], \oc8051_symbolic_cxrom1.cxrom_data_out [17]);
  buf(cxrom_data_out[18], \oc8051_symbolic_cxrom1.cxrom_data_out [18]);
  buf(cxrom_data_out[19], \oc8051_symbolic_cxrom1.cxrom_data_out [19]);
  buf(cxrom_data_out[20], \oc8051_symbolic_cxrom1.cxrom_data_out [20]);
  buf(cxrom_data_out[21], \oc8051_symbolic_cxrom1.cxrom_data_out [21]);
  buf(cxrom_data_out[22], \oc8051_symbolic_cxrom1.cxrom_data_out [22]);
  buf(cxrom_data_out[23], \oc8051_symbolic_cxrom1.cxrom_data_out [23]);
  buf(cxrom_data_out[24], \oc8051_symbolic_cxrom1.cxrom_data_out [24]);
  buf(cxrom_data_out[25], \oc8051_symbolic_cxrom1.cxrom_data_out [25]);
  buf(cxrom_data_out[26], \oc8051_symbolic_cxrom1.cxrom_data_out [26]);
  buf(cxrom_data_out[27], \oc8051_symbolic_cxrom1.cxrom_data_out [27]);
  buf(cxrom_data_out[28], \oc8051_symbolic_cxrom1.cxrom_data_out [28]);
  buf(cxrom_data_out[29], \oc8051_symbolic_cxrom1.cxrom_data_out [29]);
  buf(cxrom_data_out[30], \oc8051_symbolic_cxrom1.cxrom_data_out [30]);
  buf(cxrom_data_out[31], \oc8051_symbolic_cxrom1.cxrom_data_out [31]);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.wr_bit , \oc8051_top_1.oc8051_sfr1.wr_bit_r );
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.rst , rst);
  buf(\oc8051_top_1.oc8051_sfr1.oc8051_b_register.clk , clk);
  buf(p3_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [0]);
  buf(p3_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [1]);
  buf(p3_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [2]);
  buf(p3_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [3]);
  buf(p3_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [4]);
  buf(p3_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [5]);
  buf(p3_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [6]);
  buf(p3_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p3_out [7]);
  buf(p2_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [0]);
  buf(p2_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [1]);
  buf(p2_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [2]);
  buf(p2_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [3]);
  buf(p2_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [4]);
  buf(p2_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [5]);
  buf(p2_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [6]);
  buf(p2_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p2_out [7]);
  buf(p1_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [0]);
  buf(p1_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [1]);
  buf(p1_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [2]);
  buf(p1_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [3]);
  buf(p1_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [4]);
  buf(p1_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [5]);
  buf(p1_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [6]);
  buf(p1_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p1_out [7]);
  buf(p0_out[0], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [0]);
  buf(p0_out[1], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [1]);
  buf(p0_out[2], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [2]);
  buf(p0_out[3], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [3]);
  buf(p0_out[4], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [4]);
  buf(p0_out[5], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [5]);
  buf(p0_out[6], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [6]);
  buf(p0_out[7], \oc8051_top_1.oc8051_sfr1.oc8051_ports1.p0_out [7]);
endmodule
